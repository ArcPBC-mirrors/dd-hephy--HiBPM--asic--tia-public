magic
tech sky130A
magscale 1 2
timestamp 1683544843
<< metal3 >>
rect -2186 1512 2186 1540
rect -2186 -1512 2102 1512
rect 2166 -1512 2186 1512
rect -2186 -1540 2186 -1512
<< via3 >>
rect 2102 -1512 2166 1512
<< mimcap >>
rect -2146 1460 1854 1500
rect -2146 -1460 -2106 1460
rect 1814 -1460 1854 1460
rect -2146 -1500 1854 -1460
<< mimcapcontact >>
rect -2106 -1460 1814 1460
<< metal4 >>
rect 2086 1512 2182 1528
rect -2107 1460 1815 1461
rect -2107 -1460 -2106 1460
rect 1814 -1460 1815 1460
rect -2107 -1461 1815 -1460
rect 2086 -1512 2102 1512
rect 2166 -1512 2182 1512
rect 2086 -1528 2182 -1512
<< properties >>
string FIXED_BBOX -2186 -1540 1894 1540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20 l 15 val 613.3 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
