magic
tech sky130A
magscale 1 2
timestamp 1683558843
<< pwell >>
rect -307 -998 307 998
<< psubdiff >>
rect -271 928 -175 962
rect 175 928 271 962
rect -271 866 -237 928
rect 237 866 271 928
rect -271 -928 -237 -866
rect 237 -928 271 -866
rect -271 -962 -175 -928
rect 175 -962 271 -928
<< psubdiffcont >>
rect -175 928 175 962
rect -271 -866 -237 866
rect 237 -866 271 866
rect -175 -962 175 -928
<< xpolycontact >>
rect -141 400 141 832
rect -141 -832 141 -400
<< xpolyres >>
rect -141 -400 141 400
<< locali >>
rect -271 928 -175 962
rect 175 928 271 962
rect -271 866 -237 928
rect 237 866 271 928
rect -271 -928 -237 -866
rect 237 -928 271 -866
rect -271 -962 -175 -928
rect 175 -962 271 -928
<< viali >>
rect -125 417 125 814
rect -125 -814 125 -417
<< metal1 >>
rect -131 814 131 826
rect -131 417 -125 814
rect 125 417 131 814
rect -131 405 131 417
rect -131 -417 131 -405
rect -131 -814 -125 -417
rect 125 -814 131 -417
rect -131 -826 131 -814
<< res1p41 >>
rect -143 -402 143 402
<< properties >>
string FIXED_BBOX -254 -945 254 945
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.0 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 5.94k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
