magic
tech sky130A
magscale 1 2
timestamp 1683561438
<< nwell >>
rect -4913 1381 -2647 1963
rect -2393 1381 -127 1963
rect 127 1381 2393 1963
rect 2647 1381 4913 1963
rect -4913 545 -2647 1127
rect -2393 545 -127 1127
rect 127 545 2393 1127
rect 2647 545 4913 1127
rect -4913 -291 -2647 291
rect -2393 -291 -127 291
rect 127 -291 2393 291
rect 2647 -291 4913 291
rect -4913 -1127 -2647 -545
rect -2393 -1127 -127 -545
rect 127 -1127 2393 -545
rect 2647 -1127 4913 -545
rect -4913 -1963 -2647 -1381
rect -2393 -1963 -127 -1381
rect 127 -1963 2393 -1381
rect 2647 -1963 4913 -1381
<< pwell >>
rect -5023 1963 5023 2073
rect -5023 1381 -4913 1963
rect -2647 1381 -2393 1963
rect -127 1381 127 1963
rect 2393 1381 2647 1963
rect 4913 1381 5023 1963
rect -5023 1127 5023 1381
rect -5023 545 -4913 1127
rect -2647 545 -2393 1127
rect -127 545 127 1127
rect 2393 545 2647 1127
rect 4913 545 5023 1127
rect -5023 291 5023 545
rect -5023 -291 -4913 291
rect -2647 -291 -2393 291
rect -127 -291 127 291
rect 2393 -291 2647 291
rect 4913 -291 5023 291
rect -5023 -545 5023 -291
rect -5023 -1127 -4913 -545
rect -2647 -1127 -2393 -545
rect -127 -1127 127 -545
rect 2393 -1127 2647 -545
rect 4913 -1127 5023 -545
rect -5023 -1381 5023 -1127
rect -5023 -1963 -4913 -1381
rect -2647 -1963 -2393 -1381
rect -127 -1963 127 -1381
rect 2393 -1963 2647 -1381
rect 4913 -1963 5023 -1381
rect -5023 -2073 5023 -1963
<< varactor >>
rect -4780 1472 -2780 1872
rect -2260 1472 -260 1872
rect 260 1472 2260 1872
rect 2780 1472 4780 1872
rect -4780 636 -2780 1036
rect -2260 636 -260 1036
rect 260 636 2260 1036
rect 2780 636 4780 1036
rect -4780 -200 -2780 200
rect -2260 -200 -260 200
rect 260 -200 2260 200
rect 2780 -200 4780 200
rect -4780 -1036 -2780 -636
rect -2260 -1036 -260 -636
rect 260 -1036 2260 -636
rect 2780 -1036 4780 -636
rect -4780 -1872 -2780 -1472
rect -2260 -1872 -260 -1472
rect 260 -1872 2260 -1472
rect 2780 -1872 4780 -1472
<< psubdiff >>
rect -4987 2003 -4891 2037
rect 4891 2003 4987 2037
rect -4987 1941 -4953 2003
rect 4953 1941 4987 2003
rect -4987 -2003 -4953 -1941
rect 4953 -2003 4987 -1941
rect -4987 -2037 -4891 -2003
rect 4891 -2037 4987 -2003
<< nsubdiff >>
rect -4877 1848 -4780 1872
rect -4877 1496 -4865 1848
rect -4831 1496 -4780 1848
rect -4877 1472 -4780 1496
rect -2780 1848 -2683 1872
rect -2780 1496 -2729 1848
rect -2695 1496 -2683 1848
rect -2780 1472 -2683 1496
rect -2357 1848 -2260 1872
rect -2357 1496 -2345 1848
rect -2311 1496 -2260 1848
rect -2357 1472 -2260 1496
rect -260 1848 -163 1872
rect -260 1496 -209 1848
rect -175 1496 -163 1848
rect -260 1472 -163 1496
rect 163 1848 260 1872
rect 163 1496 175 1848
rect 209 1496 260 1848
rect 163 1472 260 1496
rect 2260 1848 2357 1872
rect 2260 1496 2311 1848
rect 2345 1496 2357 1848
rect 2260 1472 2357 1496
rect 2683 1848 2780 1872
rect 2683 1496 2695 1848
rect 2729 1496 2780 1848
rect 2683 1472 2780 1496
rect 4780 1848 4877 1872
rect 4780 1496 4831 1848
rect 4865 1496 4877 1848
rect 4780 1472 4877 1496
rect -4877 1012 -4780 1036
rect -4877 660 -4865 1012
rect -4831 660 -4780 1012
rect -4877 636 -4780 660
rect -2780 1012 -2683 1036
rect -2780 660 -2729 1012
rect -2695 660 -2683 1012
rect -2780 636 -2683 660
rect -2357 1012 -2260 1036
rect -2357 660 -2345 1012
rect -2311 660 -2260 1012
rect -2357 636 -2260 660
rect -260 1012 -163 1036
rect -260 660 -209 1012
rect -175 660 -163 1012
rect -260 636 -163 660
rect 163 1012 260 1036
rect 163 660 175 1012
rect 209 660 260 1012
rect 163 636 260 660
rect 2260 1012 2357 1036
rect 2260 660 2311 1012
rect 2345 660 2357 1012
rect 2260 636 2357 660
rect 2683 1012 2780 1036
rect 2683 660 2695 1012
rect 2729 660 2780 1012
rect 2683 636 2780 660
rect 4780 1012 4877 1036
rect 4780 660 4831 1012
rect 4865 660 4877 1012
rect 4780 636 4877 660
rect -4877 176 -4780 200
rect -4877 -176 -4865 176
rect -4831 -176 -4780 176
rect -4877 -200 -4780 -176
rect -2780 176 -2683 200
rect -2780 -176 -2729 176
rect -2695 -176 -2683 176
rect -2780 -200 -2683 -176
rect -2357 176 -2260 200
rect -2357 -176 -2345 176
rect -2311 -176 -2260 176
rect -2357 -200 -2260 -176
rect -260 176 -163 200
rect -260 -176 -209 176
rect -175 -176 -163 176
rect -260 -200 -163 -176
rect 163 176 260 200
rect 163 -176 175 176
rect 209 -176 260 176
rect 163 -200 260 -176
rect 2260 176 2357 200
rect 2260 -176 2311 176
rect 2345 -176 2357 176
rect 2260 -200 2357 -176
rect 2683 176 2780 200
rect 2683 -176 2695 176
rect 2729 -176 2780 176
rect 2683 -200 2780 -176
rect 4780 176 4877 200
rect 4780 -176 4831 176
rect 4865 -176 4877 176
rect 4780 -200 4877 -176
rect -4877 -660 -4780 -636
rect -4877 -1012 -4865 -660
rect -4831 -1012 -4780 -660
rect -4877 -1036 -4780 -1012
rect -2780 -660 -2683 -636
rect -2780 -1012 -2729 -660
rect -2695 -1012 -2683 -660
rect -2780 -1036 -2683 -1012
rect -2357 -660 -2260 -636
rect -2357 -1012 -2345 -660
rect -2311 -1012 -2260 -660
rect -2357 -1036 -2260 -1012
rect -260 -660 -163 -636
rect -260 -1012 -209 -660
rect -175 -1012 -163 -660
rect -260 -1036 -163 -1012
rect 163 -660 260 -636
rect 163 -1012 175 -660
rect 209 -1012 260 -660
rect 163 -1036 260 -1012
rect 2260 -660 2357 -636
rect 2260 -1012 2311 -660
rect 2345 -1012 2357 -660
rect 2260 -1036 2357 -1012
rect 2683 -660 2780 -636
rect 2683 -1012 2695 -660
rect 2729 -1012 2780 -660
rect 2683 -1036 2780 -1012
rect 4780 -660 4877 -636
rect 4780 -1012 4831 -660
rect 4865 -1012 4877 -660
rect 4780 -1036 4877 -1012
rect -4877 -1496 -4780 -1472
rect -4877 -1848 -4865 -1496
rect -4831 -1848 -4780 -1496
rect -4877 -1872 -4780 -1848
rect -2780 -1496 -2683 -1472
rect -2780 -1848 -2729 -1496
rect -2695 -1848 -2683 -1496
rect -2780 -1872 -2683 -1848
rect -2357 -1496 -2260 -1472
rect -2357 -1848 -2345 -1496
rect -2311 -1848 -2260 -1496
rect -2357 -1872 -2260 -1848
rect -260 -1496 -163 -1472
rect -260 -1848 -209 -1496
rect -175 -1848 -163 -1496
rect -260 -1872 -163 -1848
rect 163 -1496 260 -1472
rect 163 -1848 175 -1496
rect 209 -1848 260 -1496
rect 163 -1872 260 -1848
rect 2260 -1496 2357 -1472
rect 2260 -1848 2311 -1496
rect 2345 -1848 2357 -1496
rect 2260 -1872 2357 -1848
rect 2683 -1496 2780 -1472
rect 2683 -1848 2695 -1496
rect 2729 -1848 2780 -1496
rect 2683 -1872 2780 -1848
rect 4780 -1496 4877 -1472
rect 4780 -1848 4831 -1496
rect 4865 -1848 4877 -1496
rect 4780 -1872 4877 -1848
<< psubdiffcont >>
rect -4891 2003 4891 2037
rect -4987 -1941 -4953 1941
rect 4953 -1941 4987 1941
rect -4891 -2037 4891 -2003
<< nsubdiffcont >>
rect -4865 1496 -4831 1848
rect -2729 1496 -2695 1848
rect -2345 1496 -2311 1848
rect -209 1496 -175 1848
rect 175 1496 209 1848
rect 2311 1496 2345 1848
rect 2695 1496 2729 1848
rect 4831 1496 4865 1848
rect -4865 660 -4831 1012
rect -2729 660 -2695 1012
rect -2345 660 -2311 1012
rect -209 660 -175 1012
rect 175 660 209 1012
rect 2311 660 2345 1012
rect 2695 660 2729 1012
rect 4831 660 4865 1012
rect -4865 -176 -4831 176
rect -2729 -176 -2695 176
rect -2345 -176 -2311 176
rect -209 -176 -175 176
rect 175 -176 209 176
rect 2311 -176 2345 176
rect 2695 -176 2729 176
rect 4831 -176 4865 176
rect -4865 -1012 -4831 -660
rect -2729 -1012 -2695 -660
rect -2345 -1012 -2311 -660
rect -209 -1012 -175 -660
rect 175 -1012 209 -660
rect 2311 -1012 2345 -660
rect 2695 -1012 2729 -660
rect 4831 -1012 4865 -660
rect -4865 -1848 -4831 -1496
rect -2729 -1848 -2695 -1496
rect -2345 -1848 -2311 -1496
rect -209 -1848 -175 -1496
rect 175 -1848 209 -1496
rect 2311 -1848 2345 -1496
rect 2695 -1848 2729 -1496
rect 4831 -1848 4865 -1496
<< poly >>
rect -4780 1944 -2780 1960
rect -4780 1910 -4764 1944
rect -2796 1910 -2780 1944
rect -4780 1872 -2780 1910
rect -2260 1944 -260 1960
rect -2260 1910 -2244 1944
rect -276 1910 -260 1944
rect -2260 1872 -260 1910
rect 260 1944 2260 1960
rect 260 1910 276 1944
rect 2244 1910 2260 1944
rect 260 1872 2260 1910
rect 2780 1944 4780 1960
rect 2780 1910 2796 1944
rect 4764 1910 4780 1944
rect 2780 1872 4780 1910
rect -4780 1434 -2780 1472
rect -4780 1400 -4764 1434
rect -2796 1400 -2780 1434
rect -4780 1384 -2780 1400
rect -2260 1434 -260 1472
rect -2260 1400 -2244 1434
rect -276 1400 -260 1434
rect -2260 1384 -260 1400
rect 260 1434 2260 1472
rect 260 1400 276 1434
rect 2244 1400 2260 1434
rect 260 1384 2260 1400
rect 2780 1434 4780 1472
rect 2780 1400 2796 1434
rect 4764 1400 4780 1434
rect 2780 1384 4780 1400
rect -4780 1108 -2780 1124
rect -4780 1074 -4764 1108
rect -2796 1074 -2780 1108
rect -4780 1036 -2780 1074
rect -2260 1108 -260 1124
rect -2260 1074 -2244 1108
rect -276 1074 -260 1108
rect -2260 1036 -260 1074
rect 260 1108 2260 1124
rect 260 1074 276 1108
rect 2244 1074 2260 1108
rect 260 1036 2260 1074
rect 2780 1108 4780 1124
rect 2780 1074 2796 1108
rect 4764 1074 4780 1108
rect 2780 1036 4780 1074
rect -4780 598 -2780 636
rect -4780 564 -4764 598
rect -2796 564 -2780 598
rect -4780 548 -2780 564
rect -2260 598 -260 636
rect -2260 564 -2244 598
rect -276 564 -260 598
rect -2260 548 -260 564
rect 260 598 2260 636
rect 260 564 276 598
rect 2244 564 2260 598
rect 260 548 2260 564
rect 2780 598 4780 636
rect 2780 564 2796 598
rect 4764 564 4780 598
rect 2780 548 4780 564
rect -4780 272 -2780 288
rect -4780 238 -4764 272
rect -2796 238 -2780 272
rect -4780 200 -2780 238
rect -2260 272 -260 288
rect -2260 238 -2244 272
rect -276 238 -260 272
rect -2260 200 -260 238
rect 260 272 2260 288
rect 260 238 276 272
rect 2244 238 2260 272
rect 260 200 2260 238
rect 2780 272 4780 288
rect 2780 238 2796 272
rect 4764 238 4780 272
rect 2780 200 4780 238
rect -4780 -238 -2780 -200
rect -4780 -272 -4764 -238
rect -2796 -272 -2780 -238
rect -4780 -288 -2780 -272
rect -2260 -238 -260 -200
rect -2260 -272 -2244 -238
rect -276 -272 -260 -238
rect -2260 -288 -260 -272
rect 260 -238 2260 -200
rect 260 -272 276 -238
rect 2244 -272 2260 -238
rect 260 -288 2260 -272
rect 2780 -238 4780 -200
rect 2780 -272 2796 -238
rect 4764 -272 4780 -238
rect 2780 -288 4780 -272
rect -4780 -564 -2780 -548
rect -4780 -598 -4764 -564
rect -2796 -598 -2780 -564
rect -4780 -636 -2780 -598
rect -2260 -564 -260 -548
rect -2260 -598 -2244 -564
rect -276 -598 -260 -564
rect -2260 -636 -260 -598
rect 260 -564 2260 -548
rect 260 -598 276 -564
rect 2244 -598 2260 -564
rect 260 -636 2260 -598
rect 2780 -564 4780 -548
rect 2780 -598 2796 -564
rect 4764 -598 4780 -564
rect 2780 -636 4780 -598
rect -4780 -1074 -2780 -1036
rect -4780 -1108 -4764 -1074
rect -2796 -1108 -2780 -1074
rect -4780 -1124 -2780 -1108
rect -2260 -1074 -260 -1036
rect -2260 -1108 -2244 -1074
rect -276 -1108 -260 -1074
rect -2260 -1124 -260 -1108
rect 260 -1074 2260 -1036
rect 260 -1108 276 -1074
rect 2244 -1108 2260 -1074
rect 260 -1124 2260 -1108
rect 2780 -1074 4780 -1036
rect 2780 -1108 2796 -1074
rect 4764 -1108 4780 -1074
rect 2780 -1124 4780 -1108
rect -4780 -1400 -2780 -1384
rect -4780 -1434 -4764 -1400
rect -2796 -1434 -2780 -1400
rect -4780 -1472 -2780 -1434
rect -2260 -1400 -260 -1384
rect -2260 -1434 -2244 -1400
rect -276 -1434 -260 -1400
rect -2260 -1472 -260 -1434
rect 260 -1400 2260 -1384
rect 260 -1434 276 -1400
rect 2244 -1434 2260 -1400
rect 260 -1472 2260 -1434
rect 2780 -1400 4780 -1384
rect 2780 -1434 2796 -1400
rect 4764 -1434 4780 -1400
rect 2780 -1472 4780 -1434
rect -4780 -1910 -2780 -1872
rect -4780 -1944 -4764 -1910
rect -2796 -1944 -2780 -1910
rect -4780 -1960 -2780 -1944
rect -2260 -1910 -260 -1872
rect -2260 -1944 -2244 -1910
rect -276 -1944 -260 -1910
rect -2260 -1960 -260 -1944
rect 260 -1910 2260 -1872
rect 260 -1944 276 -1910
rect 2244 -1944 2260 -1910
rect 260 -1960 2260 -1944
rect 2780 -1910 4780 -1872
rect 2780 -1944 2796 -1910
rect 4764 -1944 4780 -1910
rect 2780 -1960 4780 -1944
<< polycont >>
rect -4764 1910 -2796 1944
rect -2244 1910 -276 1944
rect 276 1910 2244 1944
rect 2796 1910 4764 1944
rect -4764 1400 -2796 1434
rect -2244 1400 -276 1434
rect 276 1400 2244 1434
rect 2796 1400 4764 1434
rect -4764 1074 -2796 1108
rect -2244 1074 -276 1108
rect 276 1074 2244 1108
rect 2796 1074 4764 1108
rect -4764 564 -2796 598
rect -2244 564 -276 598
rect 276 564 2244 598
rect 2796 564 4764 598
rect -4764 238 -2796 272
rect -2244 238 -276 272
rect 276 238 2244 272
rect 2796 238 4764 272
rect -4764 -272 -2796 -238
rect -2244 -272 -276 -238
rect 276 -272 2244 -238
rect 2796 -272 4764 -238
rect -4764 -598 -2796 -564
rect -2244 -598 -276 -564
rect 276 -598 2244 -564
rect 2796 -598 4764 -564
rect -4764 -1108 -2796 -1074
rect -2244 -1108 -276 -1074
rect 276 -1108 2244 -1074
rect 2796 -1108 4764 -1074
rect -4764 -1434 -2796 -1400
rect -2244 -1434 -276 -1400
rect 276 -1434 2244 -1400
rect 2796 -1434 4764 -1400
rect -4764 -1944 -2796 -1910
rect -2244 -1944 -276 -1910
rect 276 -1944 2244 -1910
rect 2796 -1944 4764 -1910
<< locali >>
rect -4987 2003 -4891 2037
rect 4891 2003 4987 2037
rect -4987 1941 -4953 2003
rect -4780 1910 -4764 1944
rect -2796 1910 -2780 1944
rect -2260 1910 -2244 1944
rect -276 1910 -260 1944
rect 260 1910 276 1944
rect 2244 1910 2260 1944
rect 2780 1910 2796 1944
rect 4764 1910 4780 1944
rect 4953 1941 4987 2003
rect -4865 1848 -4831 1864
rect -4865 1480 -4831 1496
rect -2729 1848 -2695 1864
rect -2729 1480 -2695 1496
rect -2345 1848 -2311 1864
rect -2345 1480 -2311 1496
rect -209 1848 -175 1864
rect -209 1480 -175 1496
rect 175 1848 209 1864
rect 175 1480 209 1496
rect 2311 1848 2345 1864
rect 2311 1480 2345 1496
rect 2695 1848 2729 1864
rect 2695 1480 2729 1496
rect 4831 1848 4865 1864
rect 4831 1480 4865 1496
rect -4780 1400 -4764 1434
rect -2796 1400 -2780 1434
rect -2260 1400 -2244 1434
rect -276 1400 -260 1434
rect 260 1400 276 1434
rect 2244 1400 2260 1434
rect 2780 1400 2796 1434
rect 4764 1400 4780 1434
rect -4780 1074 -4764 1108
rect -2796 1074 -2780 1108
rect -2260 1074 -2244 1108
rect -276 1074 -260 1108
rect 260 1074 276 1108
rect 2244 1074 2260 1108
rect 2780 1074 2796 1108
rect 4764 1074 4780 1108
rect -4865 1012 -4831 1028
rect -4865 644 -4831 660
rect -2729 1012 -2695 1028
rect -2729 644 -2695 660
rect -2345 1012 -2311 1028
rect -2345 644 -2311 660
rect -209 1012 -175 1028
rect -209 644 -175 660
rect 175 1012 209 1028
rect 175 644 209 660
rect 2311 1012 2345 1028
rect 2311 644 2345 660
rect 2695 1012 2729 1028
rect 2695 644 2729 660
rect 4831 1012 4865 1028
rect 4831 644 4865 660
rect -4780 564 -4764 598
rect -2796 564 -2780 598
rect -2260 564 -2244 598
rect -276 564 -260 598
rect 260 564 276 598
rect 2244 564 2260 598
rect 2780 564 2796 598
rect 4764 564 4780 598
rect -4780 238 -4764 272
rect -2796 238 -2780 272
rect -2260 238 -2244 272
rect -276 238 -260 272
rect 260 238 276 272
rect 2244 238 2260 272
rect 2780 238 2796 272
rect 4764 238 4780 272
rect -4865 176 -4831 192
rect -4865 -192 -4831 -176
rect -2729 176 -2695 192
rect -2729 -192 -2695 -176
rect -2345 176 -2311 192
rect -2345 -192 -2311 -176
rect -209 176 -175 192
rect -209 -192 -175 -176
rect 175 176 209 192
rect 175 -192 209 -176
rect 2311 176 2345 192
rect 2311 -192 2345 -176
rect 2695 176 2729 192
rect 2695 -192 2729 -176
rect 4831 176 4865 192
rect 4831 -192 4865 -176
rect -4780 -272 -4764 -238
rect -2796 -272 -2780 -238
rect -2260 -272 -2244 -238
rect -276 -272 -260 -238
rect 260 -272 276 -238
rect 2244 -272 2260 -238
rect 2780 -272 2796 -238
rect 4764 -272 4780 -238
rect -4780 -598 -4764 -564
rect -2796 -598 -2780 -564
rect -2260 -598 -2244 -564
rect -276 -598 -260 -564
rect 260 -598 276 -564
rect 2244 -598 2260 -564
rect 2780 -598 2796 -564
rect 4764 -598 4780 -564
rect -4865 -660 -4831 -644
rect -4865 -1028 -4831 -1012
rect -2729 -660 -2695 -644
rect -2729 -1028 -2695 -1012
rect -2345 -660 -2311 -644
rect -2345 -1028 -2311 -1012
rect -209 -660 -175 -644
rect -209 -1028 -175 -1012
rect 175 -660 209 -644
rect 175 -1028 209 -1012
rect 2311 -660 2345 -644
rect 2311 -1028 2345 -1012
rect 2695 -660 2729 -644
rect 2695 -1028 2729 -1012
rect 4831 -660 4865 -644
rect 4831 -1028 4865 -1012
rect -4780 -1108 -4764 -1074
rect -2796 -1108 -2780 -1074
rect -2260 -1108 -2244 -1074
rect -276 -1108 -260 -1074
rect 260 -1108 276 -1074
rect 2244 -1108 2260 -1074
rect 2780 -1108 2796 -1074
rect 4764 -1108 4780 -1074
rect -4780 -1434 -4764 -1400
rect -2796 -1434 -2780 -1400
rect -2260 -1434 -2244 -1400
rect -276 -1434 -260 -1400
rect 260 -1434 276 -1400
rect 2244 -1434 2260 -1400
rect 2780 -1434 2796 -1400
rect 4764 -1434 4780 -1400
rect -4865 -1496 -4831 -1480
rect -4865 -1864 -4831 -1848
rect -2729 -1496 -2695 -1480
rect -2729 -1864 -2695 -1848
rect -2345 -1496 -2311 -1480
rect -2345 -1864 -2311 -1848
rect -209 -1496 -175 -1480
rect -209 -1864 -175 -1848
rect 175 -1496 209 -1480
rect 175 -1864 209 -1848
rect 2311 -1496 2345 -1480
rect 2311 -1864 2345 -1848
rect 2695 -1496 2729 -1480
rect 2695 -1864 2729 -1848
rect 4831 -1496 4865 -1480
rect 4831 -1864 4865 -1848
rect -4987 -2003 -4953 -1941
rect -4780 -1944 -4764 -1910
rect -2796 -1944 -2780 -1910
rect -2260 -1944 -2244 -1910
rect -276 -1944 -260 -1910
rect 260 -1944 276 -1910
rect 2244 -1944 2260 -1910
rect 2780 -1944 2796 -1910
rect 4764 -1944 4780 -1910
rect 4953 -2003 4987 -1941
rect -4987 -2037 -4891 -2003
rect 4891 -2037 4987 -2003
<< viali >>
rect -4764 1910 -2796 1944
rect -2244 1910 -276 1944
rect 276 1910 2244 1944
rect 2796 1910 4764 1944
rect -4865 1496 -4831 1848
rect -2729 1496 -2695 1848
rect -2345 1496 -2311 1848
rect -209 1496 -175 1848
rect 175 1496 209 1848
rect 2311 1496 2345 1848
rect 2695 1496 2729 1848
rect 4831 1496 4865 1848
rect -4764 1400 -2796 1434
rect -2244 1400 -276 1434
rect 276 1400 2244 1434
rect 2796 1400 4764 1434
rect -4764 1074 -2796 1108
rect -2244 1074 -276 1108
rect 276 1074 2244 1108
rect 2796 1074 4764 1108
rect -4865 660 -4831 1012
rect -2729 660 -2695 1012
rect -2345 660 -2311 1012
rect -209 660 -175 1012
rect 175 660 209 1012
rect 2311 660 2345 1012
rect 2695 660 2729 1012
rect 4831 660 4865 1012
rect -4764 564 -2796 598
rect -2244 564 -276 598
rect 276 564 2244 598
rect 2796 564 4764 598
rect -4764 238 -2796 272
rect -2244 238 -276 272
rect 276 238 2244 272
rect 2796 238 4764 272
rect -4865 -176 -4831 176
rect -2729 -176 -2695 176
rect -2345 -176 -2311 176
rect -209 -176 -175 176
rect 175 -176 209 176
rect 2311 -176 2345 176
rect 2695 -176 2729 176
rect 4831 -176 4865 176
rect -4764 -272 -2796 -238
rect -2244 -272 -276 -238
rect 276 -272 2244 -238
rect 2796 -272 4764 -238
rect -4764 -598 -2796 -564
rect -2244 -598 -276 -564
rect 276 -598 2244 -564
rect 2796 -598 4764 -564
rect -4865 -1012 -4831 -660
rect -2729 -1012 -2695 -660
rect -2345 -1012 -2311 -660
rect -209 -1012 -175 -660
rect 175 -1012 209 -660
rect 2311 -1012 2345 -660
rect 2695 -1012 2729 -660
rect 4831 -1012 4865 -660
rect -4764 -1108 -2796 -1074
rect -2244 -1108 -276 -1074
rect 276 -1108 2244 -1074
rect 2796 -1108 4764 -1074
rect -4764 -1434 -2796 -1400
rect -2244 -1434 -276 -1400
rect 276 -1434 2244 -1400
rect 2796 -1434 4764 -1400
rect -4865 -1848 -4831 -1496
rect -2729 -1848 -2695 -1496
rect -2345 -1848 -2311 -1496
rect -209 -1848 -175 -1496
rect 175 -1848 209 -1496
rect 2311 -1848 2345 -1496
rect 2695 -1848 2729 -1496
rect 4831 -1848 4865 -1496
rect -4764 -1944 -2796 -1910
rect -2244 -1944 -276 -1910
rect 276 -1944 2244 -1910
rect 2796 -1944 4764 -1910
<< metal1 >>
rect -4776 1944 -2784 1950
rect -4776 1910 -4764 1944
rect -2796 1910 -2784 1944
rect -4776 1904 -2784 1910
rect -2256 1944 -264 1950
rect -2256 1910 -2244 1944
rect -276 1910 -264 1944
rect -2256 1904 -264 1910
rect 264 1944 2256 1950
rect 264 1910 276 1944
rect 2244 1910 2256 1944
rect 264 1904 2256 1910
rect 2784 1944 4776 1950
rect 2784 1910 2796 1944
rect 4764 1910 4776 1944
rect 2784 1904 4776 1910
rect -4871 1848 -4825 1860
rect -2735 1848 -2689 1860
rect -4871 1496 -4865 1848
rect -4831 1496 -2729 1848
rect -2695 1496 -2689 1848
rect -4871 1484 -4825 1496
rect -2735 1484 -2689 1496
rect -2351 1848 -2305 1860
rect -215 1848 -169 1860
rect -2351 1496 -2345 1848
rect -2311 1496 -209 1848
rect -175 1496 -169 1848
rect -2351 1484 -2305 1496
rect -215 1484 -169 1496
rect 169 1848 215 1860
rect 2305 1848 2351 1860
rect 169 1496 175 1848
rect 209 1496 2311 1848
rect 2345 1496 2351 1848
rect 169 1484 215 1496
rect 2305 1484 2351 1496
rect 2689 1848 2735 1860
rect 4825 1848 4871 1860
rect 2689 1496 2695 1848
rect 2729 1496 4831 1848
rect 4865 1496 4871 1848
rect 2689 1484 2735 1496
rect 4825 1484 4871 1496
rect -4776 1434 -2784 1440
rect -4776 1400 -4764 1434
rect -2796 1400 -2784 1434
rect -4776 1394 -2784 1400
rect -2256 1434 -264 1440
rect -2256 1400 -2244 1434
rect -276 1400 -264 1434
rect -2256 1394 -264 1400
rect 264 1434 2256 1440
rect 264 1400 276 1434
rect 2244 1400 2256 1434
rect 264 1394 2256 1400
rect 2784 1434 4776 1440
rect 2784 1400 2796 1434
rect 4764 1400 4776 1434
rect 2784 1394 4776 1400
rect -4776 1108 -2784 1114
rect -4776 1074 -4764 1108
rect -2796 1074 -2784 1108
rect -4776 1068 -2784 1074
rect -2256 1108 -264 1114
rect -2256 1074 -2244 1108
rect -276 1074 -264 1108
rect -2256 1068 -264 1074
rect 264 1108 2256 1114
rect 264 1074 276 1108
rect 2244 1074 2256 1108
rect 264 1068 2256 1074
rect 2784 1108 4776 1114
rect 2784 1074 2796 1108
rect 4764 1074 4776 1108
rect 2784 1068 4776 1074
rect -4871 1012 -4825 1024
rect -2735 1012 -2689 1024
rect -4871 660 -4865 1012
rect -4831 660 -2729 1012
rect -2695 660 -2689 1012
rect -4871 648 -4825 660
rect -2735 648 -2689 660
rect -2351 1012 -2305 1024
rect -215 1012 -169 1024
rect -2351 660 -2345 1012
rect -2311 660 -209 1012
rect -175 660 -169 1012
rect -2351 648 -2305 660
rect -215 648 -169 660
rect 169 1012 215 1024
rect 2305 1012 2351 1024
rect 169 660 175 1012
rect 209 660 2311 1012
rect 2345 660 2351 1012
rect 169 648 215 660
rect 2305 648 2351 660
rect 2689 1012 2735 1024
rect 4825 1012 4871 1024
rect 2689 660 2695 1012
rect 2729 660 4831 1012
rect 4865 660 4871 1012
rect 2689 648 2735 660
rect 4825 648 4871 660
rect -4776 598 -2784 604
rect -4776 564 -4764 598
rect -2796 564 -2784 598
rect -4776 558 -2784 564
rect -2256 598 -264 604
rect -2256 564 -2244 598
rect -276 564 -264 598
rect -2256 558 -264 564
rect 264 598 2256 604
rect 264 564 276 598
rect 2244 564 2256 598
rect 264 558 2256 564
rect 2784 598 4776 604
rect 2784 564 2796 598
rect 4764 564 4776 598
rect 2784 558 4776 564
rect -4776 272 -2784 278
rect -4776 238 -4764 272
rect -2796 238 -2784 272
rect -4776 232 -2784 238
rect -2256 272 -264 278
rect -2256 238 -2244 272
rect -276 238 -264 272
rect -2256 232 -264 238
rect 264 272 2256 278
rect 264 238 276 272
rect 2244 238 2256 272
rect 264 232 2256 238
rect 2784 272 4776 278
rect 2784 238 2796 272
rect 4764 238 4776 272
rect 2784 232 4776 238
rect -4871 176 -4825 188
rect -2735 176 -2689 188
rect -4871 -176 -4865 176
rect -4831 -176 -2729 176
rect -2695 -176 -2689 176
rect -4871 -188 -4825 -176
rect -2735 -188 -2689 -176
rect -2351 176 -2305 188
rect -215 176 -169 188
rect -2351 -176 -2345 176
rect -2311 -176 -209 176
rect -175 -176 -169 176
rect -2351 -188 -2305 -176
rect -215 -188 -169 -176
rect 169 176 215 188
rect 2305 176 2351 188
rect 169 -176 175 176
rect 209 -176 2311 176
rect 2345 -176 2351 176
rect 169 -188 215 -176
rect 2305 -188 2351 -176
rect 2689 176 2735 188
rect 4825 176 4871 188
rect 2689 -176 2695 176
rect 2729 -176 4831 176
rect 4865 -176 4871 176
rect 2689 -188 2735 -176
rect 4825 -188 4871 -176
rect -4776 -238 -2784 -232
rect -4776 -272 -4764 -238
rect -2796 -272 -2784 -238
rect -4776 -278 -2784 -272
rect -2256 -238 -264 -232
rect -2256 -272 -2244 -238
rect -276 -272 -264 -238
rect -2256 -278 -264 -272
rect 264 -238 2256 -232
rect 264 -272 276 -238
rect 2244 -272 2256 -238
rect 264 -278 2256 -272
rect 2784 -238 4776 -232
rect 2784 -272 2796 -238
rect 4764 -272 4776 -238
rect 2784 -278 4776 -272
rect -4776 -564 -2784 -558
rect -4776 -598 -4764 -564
rect -2796 -598 -2784 -564
rect -4776 -604 -2784 -598
rect -2256 -564 -264 -558
rect -2256 -598 -2244 -564
rect -276 -598 -264 -564
rect -2256 -604 -264 -598
rect 264 -564 2256 -558
rect 264 -598 276 -564
rect 2244 -598 2256 -564
rect 264 -604 2256 -598
rect 2784 -564 4776 -558
rect 2784 -598 2796 -564
rect 4764 -598 4776 -564
rect 2784 -604 4776 -598
rect -4871 -660 -4825 -648
rect -2735 -660 -2689 -648
rect -4871 -1012 -4865 -660
rect -4831 -1012 -2729 -660
rect -2695 -1012 -2689 -660
rect -4871 -1024 -4825 -1012
rect -2735 -1024 -2689 -1012
rect -2351 -660 -2305 -648
rect -215 -660 -169 -648
rect -2351 -1012 -2345 -660
rect -2311 -1012 -209 -660
rect -175 -1012 -169 -660
rect -2351 -1024 -2305 -1012
rect -215 -1024 -169 -1012
rect 169 -660 215 -648
rect 2305 -660 2351 -648
rect 169 -1012 175 -660
rect 209 -1012 2311 -660
rect 2345 -1012 2351 -660
rect 169 -1024 215 -1012
rect 2305 -1024 2351 -1012
rect 2689 -660 2735 -648
rect 4825 -660 4871 -648
rect 2689 -1012 2695 -660
rect 2729 -1012 4831 -660
rect 4865 -1012 4871 -660
rect 2689 -1024 2735 -1012
rect 4825 -1024 4871 -1012
rect -4776 -1074 -2784 -1068
rect -4776 -1108 -4764 -1074
rect -2796 -1108 -2784 -1074
rect -4776 -1114 -2784 -1108
rect -2256 -1074 -264 -1068
rect -2256 -1108 -2244 -1074
rect -276 -1108 -264 -1074
rect -2256 -1114 -264 -1108
rect 264 -1074 2256 -1068
rect 264 -1108 276 -1074
rect 2244 -1108 2256 -1074
rect 264 -1114 2256 -1108
rect 2784 -1074 4776 -1068
rect 2784 -1108 2796 -1074
rect 4764 -1108 4776 -1074
rect 2784 -1114 4776 -1108
rect -4776 -1400 -2784 -1394
rect -4776 -1434 -4764 -1400
rect -2796 -1434 -2784 -1400
rect -4776 -1440 -2784 -1434
rect -2256 -1400 -264 -1394
rect -2256 -1434 -2244 -1400
rect -276 -1434 -264 -1400
rect -2256 -1440 -264 -1434
rect 264 -1400 2256 -1394
rect 264 -1434 276 -1400
rect 2244 -1434 2256 -1400
rect 264 -1440 2256 -1434
rect 2784 -1400 4776 -1394
rect 2784 -1434 2796 -1400
rect 4764 -1434 4776 -1400
rect 2784 -1440 4776 -1434
rect -4871 -1496 -4825 -1484
rect -2735 -1496 -2689 -1484
rect -4871 -1848 -4865 -1496
rect -4831 -1848 -2729 -1496
rect -2695 -1848 -2689 -1496
rect -4871 -1860 -4825 -1848
rect -2735 -1860 -2689 -1848
rect -2351 -1496 -2305 -1484
rect -215 -1496 -169 -1484
rect -2351 -1848 -2345 -1496
rect -2311 -1848 -209 -1496
rect -175 -1848 -169 -1496
rect -2351 -1860 -2305 -1848
rect -215 -1860 -169 -1848
rect 169 -1496 215 -1484
rect 2305 -1496 2351 -1484
rect 169 -1848 175 -1496
rect 209 -1848 2311 -1496
rect 2345 -1848 2351 -1496
rect 169 -1860 215 -1848
rect 2305 -1860 2351 -1848
rect 2689 -1496 2735 -1484
rect 4825 -1496 4871 -1484
rect 2689 -1848 2695 -1496
rect 2729 -1848 4831 -1496
rect 4865 -1848 4871 -1496
rect 2689 -1860 2735 -1848
rect 4825 -1860 4871 -1848
rect -4776 -1910 -2784 -1904
rect -4776 -1944 -4764 -1910
rect -2796 -1944 -2784 -1910
rect -4776 -1950 -2784 -1944
rect -2256 -1910 -264 -1904
rect -2256 -1944 -2244 -1910
rect -276 -1944 -264 -1910
rect -2256 -1950 -264 -1944
rect 264 -1910 2256 -1904
rect 264 -1944 276 -1910
rect 2244 -1944 2256 -1910
rect 264 -1950 2256 -1944
rect 2784 -1910 4776 -1904
rect 2784 -1944 2796 -1910
rect 4764 -1944 4776 -1910
rect 2784 -1950 4776 -1944
<< properties >>
string FIXED_BBOX -4970 -2020 4970 2020
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 10 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
