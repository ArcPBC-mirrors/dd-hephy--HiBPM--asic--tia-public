magic
tech sky130A
timestamp 1689778598
<< metal3 >>
rect 16500 19100 17000 21400
rect 55800 19100 56250 21450
rect 16500 14100 17000 16400
rect 55800 14050 56250 16400
rect 16800 6600 17100 8900
rect 55900 6600 56200 8900
rect 16800 -3400 17100 -1100
rect 55900 -3400 56200 -1100
rect 16800 -13400 17100 -11100
rect 55900 -13400 56200 -11100
rect 16800 -23400 17100 -21100
rect 55900 -23400 56200 -21100
<< end >>
