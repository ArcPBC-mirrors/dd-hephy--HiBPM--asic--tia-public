magic
tech sky130A
magscale 1 2
timestamp 1683806952
<< error_p >>
rect -147 581 -89 587
rect -29 581 29 587
rect 89 581 147 587
rect -147 547 -135 581
rect -29 547 -17 581
rect 89 547 101 581
rect -147 541 -89 547
rect -29 541 29 547
rect 89 541 147 547
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect -147 -37 -89 -31
rect -29 -37 29 -31
rect 89 -37 147 -31
rect -147 -71 -135 -37
rect -29 -71 -17 -37
rect 89 -71 101 -37
rect -147 -77 -89 -71
rect -29 -77 29 -71
rect 89 -77 147 -71
rect -147 -547 -89 -541
rect -29 -547 29 -541
rect 89 -547 147 -541
rect -147 -581 -135 -547
rect -29 -581 -17 -547
rect 89 -581 101 -547
rect -147 -587 -89 -581
rect -29 -587 29 -581
rect 89 -587 147 -581
<< pwell >>
rect -344 -719 344 719
<< nmoslvt >>
rect -148 109 -88 509
rect -30 109 30 509
rect 88 109 148 509
rect -148 -509 -88 -109
rect -30 -509 30 -109
rect 88 -509 148 -109
<< ndiff >>
rect -206 497 -148 509
rect -206 121 -194 497
rect -160 121 -148 497
rect -206 109 -148 121
rect -88 497 -30 509
rect -88 121 -76 497
rect -42 121 -30 497
rect -88 109 -30 121
rect 30 497 88 509
rect 30 121 42 497
rect 76 121 88 497
rect 30 109 88 121
rect 148 497 206 509
rect 148 121 160 497
rect 194 121 206 497
rect 148 109 206 121
rect -206 -121 -148 -109
rect -206 -497 -194 -121
rect -160 -497 -148 -121
rect -206 -509 -148 -497
rect -88 -121 -30 -109
rect -88 -497 -76 -121
rect -42 -497 -30 -121
rect -88 -509 -30 -497
rect 30 -121 88 -109
rect 30 -497 42 -121
rect 76 -497 88 -121
rect 30 -509 88 -497
rect 148 -121 206 -109
rect 148 -497 160 -121
rect 194 -497 206 -121
rect 148 -509 206 -497
<< ndiffc >>
rect -194 121 -160 497
rect -76 121 -42 497
rect 42 121 76 497
rect 160 121 194 497
rect -194 -497 -160 -121
rect -76 -497 -42 -121
rect 42 -497 76 -121
rect 160 -497 194 -121
<< psubdiff >>
rect -308 649 -212 683
rect 212 649 308 683
rect -308 587 -274 649
rect 274 587 308 649
rect -308 -649 -274 -587
rect 274 -649 308 -587
rect -308 -683 -212 -649
rect 212 -683 308 -649
<< psubdiffcont >>
rect -212 649 212 683
rect -308 -587 -274 587
rect 274 -587 308 587
rect -212 -683 212 -649
<< poly >>
rect -151 581 -85 597
rect -151 547 -135 581
rect -101 547 -85 581
rect -151 531 -85 547
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect 85 581 151 597
rect 85 547 101 581
rect 135 547 151 581
rect 85 531 151 547
rect -148 509 -88 531
rect -30 509 30 531
rect 88 509 148 531
rect -148 87 -88 109
rect -30 87 30 109
rect 88 87 148 109
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect -151 -37 -85 -21
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -151 -87 -85 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 85 -37 151 -21
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 85 -87 151 -71
rect -148 -109 -88 -87
rect -30 -109 30 -87
rect 88 -109 148 -87
rect -148 -531 -88 -509
rect -30 -531 30 -509
rect 88 -531 148 -509
rect -151 -547 -85 -531
rect -151 -581 -135 -547
rect -101 -581 -85 -547
rect -151 -597 -85 -581
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect 85 -547 151 -531
rect 85 -581 101 -547
rect 135 -581 151 -547
rect 85 -597 151 -581
<< polycont >>
rect -135 547 -101 581
rect -17 547 17 581
rect 101 547 135 581
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect -135 -581 -101 -547
rect -17 -581 17 -547
rect 101 -581 135 -547
<< locali >>
rect -308 649 -212 683
rect 212 649 308 683
rect -308 587 -274 649
rect 274 587 308 649
rect -151 547 -135 581
rect -101 547 -85 581
rect -33 547 -17 581
rect 17 547 33 581
rect 85 547 101 581
rect 135 547 151 581
rect -194 497 -160 513
rect -194 105 -160 121
rect -76 497 -42 513
rect -76 105 -42 121
rect 42 497 76 513
rect 42 105 76 121
rect 160 497 194 513
rect 160 105 194 121
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 85 -71 101 -37
rect 135 -71 151 -37
rect -194 -121 -160 -105
rect -194 -513 -160 -497
rect -76 -121 -42 -105
rect -76 -513 -42 -497
rect 42 -121 76 -105
rect 42 -513 76 -497
rect 160 -121 194 -105
rect 160 -513 194 -497
rect -151 -581 -135 -547
rect -101 -581 -85 -547
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect 85 -581 101 -547
rect 135 -581 151 -547
rect -308 -649 -274 -587
rect 274 -649 308 -587
rect -308 -683 -212 -649
rect 212 -683 308 -649
<< viali >>
rect -135 547 -101 581
rect -17 547 17 581
rect 101 547 135 581
rect -194 121 -160 497
rect -76 121 -42 497
rect 42 121 76 497
rect 160 121 194 497
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect -194 -497 -160 -121
rect -76 -497 -42 -121
rect 42 -497 76 -121
rect 160 -497 194 -121
rect -135 -581 -101 -547
rect -17 -581 17 -547
rect 101 -581 135 -547
<< metal1 >>
rect -147 581 -89 587
rect -147 547 -135 581
rect -101 547 -89 581
rect -147 541 -89 547
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect 89 581 147 587
rect 89 547 101 581
rect 135 547 147 581
rect 89 541 147 547
rect -200 497 -154 509
rect -200 121 -194 497
rect -160 121 -154 497
rect -200 109 -154 121
rect -82 497 -36 509
rect -82 121 -76 497
rect -42 121 -36 497
rect -82 109 -36 121
rect 36 497 82 509
rect 36 121 42 497
rect 76 121 82 497
rect 36 109 82 121
rect 154 497 200 509
rect 154 121 160 497
rect 194 121 200 497
rect 154 109 200 121
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect -147 -37 -89 -31
rect -147 -71 -135 -37
rect -101 -71 -89 -37
rect -147 -77 -89 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 89 -37 147 -31
rect 89 -71 101 -37
rect 135 -71 147 -37
rect 89 -77 147 -71
rect -200 -121 -154 -109
rect -200 -497 -194 -121
rect -160 -497 -154 -121
rect -200 -509 -154 -497
rect -82 -121 -36 -109
rect -82 -497 -76 -121
rect -42 -497 -36 -121
rect -82 -509 -36 -497
rect 36 -121 82 -109
rect 36 -497 42 -121
rect 76 -497 82 -121
rect 36 -509 82 -497
rect 154 -121 200 -109
rect 154 -497 160 -121
rect 194 -497 200 -121
rect 154 -509 200 -497
rect -147 -547 -89 -541
rect -147 -581 -135 -547
rect -101 -581 -89 -547
rect -147 -587 -89 -581
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect 89 -547 147 -541
rect 89 -581 101 -547
rect 135 -581 147 -547
rect 89 -587 147 -581
<< properties >>
string FIXED_BBOX -291 -666 291 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 2 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
