magic
tech sky130A
magscale 1 2
timestamp 1683553776
<< error_p >>
rect -461 599 -403 605
rect -269 599 -211 605
rect -77 599 -19 605
rect 115 599 173 605
rect 307 599 365 605
rect -461 565 -449 599
rect -269 565 -257 599
rect -77 565 -65 599
rect 115 565 127 599
rect 307 565 319 599
rect -461 559 -403 565
rect -269 559 -211 565
rect -77 559 -19 565
rect 115 559 173 565
rect 307 559 365 565
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect -461 -565 -403 -559
rect -269 -565 -211 -559
rect -77 -565 -19 -559
rect 115 -565 173 -559
rect 307 -565 365 -559
rect -461 -599 -449 -565
rect -269 -599 -257 -565
rect -77 -599 -65 -565
rect 115 -599 127 -565
rect 307 -599 319 -565
rect -461 -605 -403 -599
rect -269 -605 -211 -599
rect -77 -605 -19 -599
rect 115 -605 173 -599
rect 307 -605 365 -599
<< nwell >>
rect -647 -737 647 737
<< pmos >>
rect -447 118 -417 518
rect -351 118 -321 518
rect -255 118 -225 518
rect -159 118 -129 518
rect -63 118 -33 518
rect 33 118 63 518
rect 129 118 159 518
rect 225 118 255 518
rect 321 118 351 518
rect 417 118 447 518
rect -447 -518 -417 -118
rect -351 -518 -321 -118
rect -255 -518 -225 -118
rect -159 -518 -129 -118
rect -63 -518 -33 -118
rect 33 -518 63 -118
rect 129 -518 159 -118
rect 225 -518 255 -118
rect 321 -518 351 -118
rect 417 -518 447 -118
<< pdiff >>
rect -509 506 -447 518
rect -509 130 -497 506
rect -463 130 -447 506
rect -509 118 -447 130
rect -417 506 -351 518
rect -417 130 -401 506
rect -367 130 -351 506
rect -417 118 -351 130
rect -321 506 -255 518
rect -321 130 -305 506
rect -271 130 -255 506
rect -321 118 -255 130
rect -225 506 -159 518
rect -225 130 -209 506
rect -175 130 -159 506
rect -225 118 -159 130
rect -129 506 -63 518
rect -129 130 -113 506
rect -79 130 -63 506
rect -129 118 -63 130
rect -33 506 33 518
rect -33 130 -17 506
rect 17 130 33 506
rect -33 118 33 130
rect 63 506 129 518
rect 63 130 79 506
rect 113 130 129 506
rect 63 118 129 130
rect 159 506 225 518
rect 159 130 175 506
rect 209 130 225 506
rect 159 118 225 130
rect 255 506 321 518
rect 255 130 271 506
rect 305 130 321 506
rect 255 118 321 130
rect 351 506 417 518
rect 351 130 367 506
rect 401 130 417 506
rect 351 118 417 130
rect 447 506 509 518
rect 447 130 463 506
rect 497 130 509 506
rect 447 118 509 130
rect -509 -130 -447 -118
rect -509 -506 -497 -130
rect -463 -506 -447 -130
rect -509 -518 -447 -506
rect -417 -130 -351 -118
rect -417 -506 -401 -130
rect -367 -506 -351 -130
rect -417 -518 -351 -506
rect -321 -130 -255 -118
rect -321 -506 -305 -130
rect -271 -506 -255 -130
rect -321 -518 -255 -506
rect -225 -130 -159 -118
rect -225 -506 -209 -130
rect -175 -506 -159 -130
rect -225 -518 -159 -506
rect -129 -130 -63 -118
rect -129 -506 -113 -130
rect -79 -506 -63 -130
rect -129 -518 -63 -506
rect -33 -130 33 -118
rect -33 -506 -17 -130
rect 17 -506 33 -130
rect -33 -518 33 -506
rect 63 -130 129 -118
rect 63 -506 79 -130
rect 113 -506 129 -130
rect 63 -518 129 -506
rect 159 -130 225 -118
rect 159 -506 175 -130
rect 209 -506 225 -130
rect 159 -518 225 -506
rect 255 -130 321 -118
rect 255 -506 271 -130
rect 305 -506 321 -130
rect 255 -518 321 -506
rect 351 -130 417 -118
rect 351 -506 367 -130
rect 401 -506 417 -130
rect 351 -518 417 -506
rect 447 -130 509 -118
rect 447 -506 463 -130
rect 497 -506 509 -130
rect 447 -518 509 -506
<< pdiffc >>
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
<< nsubdiff >>
rect -611 667 -515 701
rect 515 667 611 701
rect -611 605 -577 667
rect 577 605 611 667
rect -611 -667 -577 -605
rect 577 -667 611 -605
rect -611 -701 -515 -667
rect 515 -701 611 -667
<< nsubdiffcont >>
rect -515 667 515 701
rect -611 -605 -577 605
rect 577 -605 611 605
rect -515 -701 515 -667
<< poly >>
rect -465 599 -399 615
rect -465 565 -449 599
rect -415 565 -399 599
rect -465 549 -399 565
rect -273 599 -207 615
rect -273 565 -257 599
rect -223 565 -207 599
rect -273 549 -207 565
rect -81 599 -15 615
rect -81 565 -65 599
rect -31 565 -15 599
rect -81 549 -15 565
rect 111 599 177 615
rect 111 565 127 599
rect 161 565 177 599
rect 111 549 177 565
rect 303 599 369 615
rect 303 565 319 599
rect 353 565 369 599
rect 303 549 369 565
rect -447 518 -417 549
rect -351 518 -321 544
rect -255 518 -225 549
rect -159 518 -129 544
rect -63 518 -33 549
rect 33 518 63 544
rect 129 518 159 549
rect 225 518 255 544
rect 321 518 351 549
rect 417 518 447 544
rect -447 92 -417 118
rect -351 87 -321 118
rect -255 92 -225 118
rect -159 87 -129 118
rect -63 92 -33 118
rect 33 87 63 118
rect 129 92 159 118
rect 225 87 255 118
rect 321 92 351 118
rect 417 87 447 118
rect -369 71 -303 87
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 399 -87 465 -71
rect -447 -118 -417 -92
rect -351 -118 -321 -87
rect -255 -118 -225 -92
rect -159 -118 -129 -87
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect 129 -118 159 -92
rect 225 -118 255 -87
rect 321 -118 351 -92
rect 417 -118 447 -87
rect -447 -549 -417 -518
rect -351 -544 -321 -518
rect -255 -549 -225 -518
rect -159 -544 -129 -518
rect -63 -549 -33 -518
rect 33 -544 63 -518
rect 129 -549 159 -518
rect 225 -544 255 -518
rect 321 -549 351 -518
rect 417 -544 447 -518
rect -465 -565 -399 -549
rect -465 -599 -449 -565
rect -415 -599 -399 -565
rect -465 -615 -399 -599
rect -273 -565 -207 -549
rect -273 -599 -257 -565
rect -223 -599 -207 -565
rect -273 -615 -207 -599
rect -81 -565 -15 -549
rect -81 -599 -65 -565
rect -31 -599 -15 -565
rect -81 -615 -15 -599
rect 111 -565 177 -549
rect 111 -599 127 -565
rect 161 -599 177 -565
rect 111 -615 177 -599
rect 303 -565 369 -549
rect 303 -599 319 -565
rect 353 -599 369 -565
rect 303 -615 369 -599
<< polycont >>
rect -449 565 -415 599
rect -257 565 -223 599
rect -65 565 -31 599
rect 127 565 161 599
rect 319 565 353 599
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -449 -599 -415 -565
rect -257 -599 -223 -565
rect -65 -599 -31 -565
rect 127 -599 161 -565
rect 319 -599 353 -565
<< locali >>
rect -611 667 -515 701
rect 515 667 611 701
rect -611 605 -577 667
rect 577 605 611 667
rect -465 565 -449 599
rect -415 565 -399 599
rect -273 565 -257 599
rect -223 565 -207 599
rect -81 565 -65 599
rect -31 565 -15 599
rect 111 565 127 599
rect 161 565 177 599
rect 303 565 319 599
rect 353 565 369 599
rect -497 506 -463 522
rect -497 114 -463 130
rect -401 506 -367 522
rect -401 114 -367 130
rect -305 506 -271 522
rect -305 114 -271 130
rect -209 506 -175 522
rect -209 114 -175 130
rect -113 506 -79 522
rect -113 114 -79 130
rect -17 506 17 522
rect -17 114 17 130
rect 79 506 113 522
rect 79 114 113 130
rect 175 506 209 522
rect 175 114 209 130
rect 271 506 305 522
rect 271 114 305 130
rect 367 506 401 522
rect 367 114 401 130
rect 463 506 497 522
rect 463 114 497 130
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect -497 -130 -463 -114
rect -497 -522 -463 -506
rect -401 -130 -367 -114
rect -401 -522 -367 -506
rect -305 -130 -271 -114
rect -305 -522 -271 -506
rect -209 -130 -175 -114
rect -209 -522 -175 -506
rect -113 -130 -79 -114
rect -113 -522 -79 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 79 -130 113 -114
rect 79 -522 113 -506
rect 175 -130 209 -114
rect 175 -522 209 -506
rect 271 -130 305 -114
rect 271 -522 305 -506
rect 367 -130 401 -114
rect 367 -522 401 -506
rect 463 -130 497 -114
rect 463 -522 497 -506
rect -465 -599 -449 -565
rect -415 -599 -399 -565
rect -273 -599 -257 -565
rect -223 -599 -207 -565
rect -81 -599 -65 -565
rect -31 -599 -15 -565
rect 111 -599 127 -565
rect 161 -599 177 -565
rect 303 -599 319 -565
rect 353 -599 369 -565
rect -611 -667 -577 -605
rect 577 -667 611 -605
rect -611 -701 -515 -667
rect 515 -701 611 -667
<< viali >>
rect -449 565 -415 599
rect -257 565 -223 599
rect -65 565 -31 599
rect 127 565 161 599
rect 319 565 353 599
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect -449 -599 -415 -565
rect -257 -599 -223 -565
rect -65 -599 -31 -565
rect 127 -599 161 -565
rect 319 -599 353 -565
<< metal1 >>
rect -461 599 -403 605
rect -461 565 -449 599
rect -415 565 -403 599
rect -461 559 -403 565
rect -269 599 -211 605
rect -269 565 -257 599
rect -223 565 -211 599
rect -269 559 -211 565
rect -77 599 -19 605
rect -77 565 -65 599
rect -31 565 -19 599
rect -77 559 -19 565
rect 115 599 173 605
rect 115 565 127 599
rect 161 565 173 599
rect 115 559 173 565
rect 307 599 365 605
rect 307 565 319 599
rect 353 565 365 599
rect 307 559 365 565
rect -503 506 -457 518
rect -503 130 -497 506
rect -463 130 -457 506
rect -503 118 -457 130
rect -407 506 -361 518
rect -407 130 -401 506
rect -367 130 -361 506
rect -407 118 -361 130
rect -311 506 -265 518
rect -311 130 -305 506
rect -271 130 -265 506
rect -311 118 -265 130
rect -215 506 -169 518
rect -215 130 -209 506
rect -175 130 -169 506
rect -215 118 -169 130
rect -119 506 -73 518
rect -119 130 -113 506
rect -79 130 -73 506
rect -119 118 -73 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 73 506 119 518
rect 73 130 79 506
rect 113 130 119 506
rect 73 118 119 130
rect 169 506 215 518
rect 169 130 175 506
rect 209 130 215 506
rect 169 118 215 130
rect 265 506 311 518
rect 265 130 271 506
rect 305 130 311 506
rect 265 118 311 130
rect 361 506 407 518
rect 361 130 367 506
rect 401 130 407 506
rect 361 118 407 130
rect 457 506 503 518
rect 457 130 463 506
rect 497 130 503 506
rect 457 118 503 130
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect -503 -130 -457 -118
rect -503 -506 -497 -130
rect -463 -506 -457 -130
rect -503 -518 -457 -506
rect -407 -130 -361 -118
rect -407 -506 -401 -130
rect -367 -506 -361 -130
rect -407 -518 -361 -506
rect -311 -130 -265 -118
rect -311 -506 -305 -130
rect -271 -506 -265 -130
rect -311 -518 -265 -506
rect -215 -130 -169 -118
rect -215 -506 -209 -130
rect -175 -506 -169 -130
rect -215 -518 -169 -506
rect -119 -130 -73 -118
rect -119 -506 -113 -130
rect -79 -506 -73 -130
rect -119 -518 -73 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 73 -130 119 -118
rect 73 -506 79 -130
rect 113 -506 119 -130
rect 73 -518 119 -506
rect 169 -130 215 -118
rect 169 -506 175 -130
rect 209 -506 215 -130
rect 169 -518 215 -506
rect 265 -130 311 -118
rect 265 -506 271 -130
rect 305 -506 311 -130
rect 265 -518 311 -506
rect 361 -130 407 -118
rect 361 -506 367 -130
rect 401 -506 407 -130
rect 361 -518 407 -506
rect 457 -130 503 -118
rect 457 -506 463 -130
rect 497 -506 503 -130
rect 457 -518 503 -506
rect -461 -565 -403 -559
rect -461 -599 -449 -565
rect -415 -599 -403 -565
rect -461 -605 -403 -599
rect -269 -565 -211 -559
rect -269 -599 -257 -565
rect -223 -599 -211 -565
rect -269 -605 -211 -599
rect -77 -565 -19 -559
rect -77 -599 -65 -565
rect -31 -599 -19 -565
rect -77 -605 -19 -599
rect 115 -565 173 -559
rect 115 -599 127 -565
rect 161 -599 173 -565
rect 115 -605 173 -599
rect 307 -565 365 -559
rect 307 -599 319 -565
rect 353 -599 365 -565
rect 307 -605 365 -599
<< properties >>
string FIXED_BBOX -594 -684 594 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
