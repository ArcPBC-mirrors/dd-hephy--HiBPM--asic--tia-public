magic
tech sky130A
magscale 1 2
timestamp 1683887376
<< error_p >>
rect -324 272 -266 278
rect -206 272 -148 278
rect -88 272 -30 278
rect 30 272 88 278
rect 148 272 206 278
rect 266 272 324 278
rect -324 238 -312 272
rect -206 238 -194 272
rect -88 238 -76 272
rect 30 238 42 272
rect 148 238 160 272
rect 266 238 278 272
rect -324 232 -266 238
rect -206 232 -148 238
rect -88 232 -30 238
rect 30 232 88 238
rect 148 232 206 238
rect 266 232 324 238
rect -324 -238 -266 -232
rect -206 -238 -148 -232
rect -88 -238 -30 -232
rect 30 -238 88 -232
rect 148 -238 206 -232
rect 266 -238 324 -232
rect -324 -272 -312 -238
rect -206 -272 -194 -238
rect -88 -272 -76 -238
rect 30 -272 42 -238
rect 148 -272 160 -238
rect 266 -272 278 -238
rect -324 -278 -266 -272
rect -206 -278 -148 -272
rect -88 -278 -30 -272
rect 30 -278 88 -272
rect 148 -278 206 -272
rect 266 -278 324 -272
<< pwell >>
rect -521 -410 521 410
<< nmoslvt >>
rect -325 -200 -265 200
rect -207 -200 -147 200
rect -89 -200 -29 200
rect 29 -200 89 200
rect 147 -200 207 200
rect 265 -200 325 200
<< ndiff >>
rect -383 188 -325 200
rect -383 -188 -371 188
rect -337 -188 -325 188
rect -383 -200 -325 -188
rect -265 188 -207 200
rect -265 -188 -253 188
rect -219 -188 -207 188
rect -265 -200 -207 -188
rect -147 188 -89 200
rect -147 -188 -135 188
rect -101 -188 -89 188
rect -147 -200 -89 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 89 188 147 200
rect 89 -188 101 188
rect 135 -188 147 188
rect 89 -200 147 -188
rect 207 188 265 200
rect 207 -188 219 188
rect 253 -188 265 188
rect 207 -200 265 -188
rect 325 188 383 200
rect 325 -188 337 188
rect 371 -188 383 188
rect 325 -200 383 -188
<< ndiffc >>
rect -371 -188 -337 188
rect -253 -188 -219 188
rect -135 -188 -101 188
rect -17 -188 17 188
rect 101 -188 135 188
rect 219 -188 253 188
rect 337 -188 371 188
<< psubdiff >>
rect -485 340 -389 374
rect 389 340 485 374
rect -485 278 -451 340
rect 451 278 485 340
rect -485 -340 -451 -278
rect 451 -340 485 -278
rect -485 -374 -389 -340
rect 389 -374 485 -340
<< psubdiffcont >>
rect -389 340 389 374
rect -485 -278 -451 278
rect 451 -278 485 278
rect -389 -374 389 -340
<< poly >>
rect -328 272 -262 288
rect -328 238 -312 272
rect -278 238 -262 272
rect -328 222 -262 238
rect -210 272 -144 288
rect -210 238 -194 272
rect -160 238 -144 272
rect -210 222 -144 238
rect -92 272 -26 288
rect -92 238 -76 272
rect -42 238 -26 272
rect -92 222 -26 238
rect 26 272 92 288
rect 26 238 42 272
rect 76 238 92 272
rect 26 222 92 238
rect 144 272 210 288
rect 144 238 160 272
rect 194 238 210 272
rect 144 222 210 238
rect 262 272 328 288
rect 262 238 278 272
rect 312 238 328 272
rect 262 222 328 238
rect -325 200 -265 222
rect -207 200 -147 222
rect -89 200 -29 222
rect 29 200 89 222
rect 147 200 207 222
rect 265 200 325 222
rect -325 -222 -265 -200
rect -207 -222 -147 -200
rect -89 -222 -29 -200
rect 29 -222 89 -200
rect 147 -222 207 -200
rect 265 -222 325 -200
rect -328 -238 -262 -222
rect -328 -272 -312 -238
rect -278 -272 -262 -238
rect -328 -288 -262 -272
rect -210 -238 -144 -222
rect -210 -272 -194 -238
rect -160 -272 -144 -238
rect -210 -288 -144 -272
rect -92 -238 -26 -222
rect -92 -272 -76 -238
rect -42 -272 -26 -238
rect -92 -288 -26 -272
rect 26 -238 92 -222
rect 26 -272 42 -238
rect 76 -272 92 -238
rect 26 -288 92 -272
rect 144 -238 210 -222
rect 144 -272 160 -238
rect 194 -272 210 -238
rect 144 -288 210 -272
rect 262 -238 328 -222
rect 262 -272 278 -238
rect 312 -272 328 -238
rect 262 -288 328 -272
<< polycont >>
rect -312 238 -278 272
rect -194 238 -160 272
rect -76 238 -42 272
rect 42 238 76 272
rect 160 238 194 272
rect 278 238 312 272
rect -312 -272 -278 -238
rect -194 -272 -160 -238
rect -76 -272 -42 -238
rect 42 -272 76 -238
rect 160 -272 194 -238
rect 278 -272 312 -238
<< locali >>
rect -485 340 -389 374
rect 389 340 485 374
rect -485 278 -451 340
rect 451 278 485 340
rect -328 238 -312 272
rect -278 238 -262 272
rect -210 238 -194 272
rect -160 238 -144 272
rect -92 238 -76 272
rect -42 238 -26 272
rect 26 238 42 272
rect 76 238 92 272
rect 144 238 160 272
rect 194 238 210 272
rect 262 238 278 272
rect 312 238 328 272
rect -371 188 -337 204
rect -371 -204 -337 -188
rect -253 188 -219 204
rect -253 -204 -219 -188
rect -135 188 -101 204
rect -135 -204 -101 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 101 188 135 204
rect 101 -204 135 -188
rect 219 188 253 204
rect 219 -204 253 -188
rect 337 188 371 204
rect 337 -204 371 -188
rect -328 -272 -312 -238
rect -278 -272 -262 -238
rect -210 -272 -194 -238
rect -160 -272 -144 -238
rect -92 -272 -76 -238
rect -42 -272 -26 -238
rect 26 -272 42 -238
rect 76 -272 92 -238
rect 144 -272 160 -238
rect 194 -272 210 -238
rect 262 -272 278 -238
rect 312 -272 328 -238
rect -485 -340 -451 -278
rect 451 -340 485 -278
rect -485 -374 -389 -340
rect 389 -374 485 -340
<< viali >>
rect -312 238 -278 272
rect -194 238 -160 272
rect -76 238 -42 272
rect 42 238 76 272
rect 160 238 194 272
rect 278 238 312 272
rect -371 -188 -337 188
rect -253 -188 -219 188
rect -135 -188 -101 188
rect -17 -188 17 188
rect 101 -188 135 188
rect 219 -188 253 188
rect 337 -188 371 188
rect -312 -272 -278 -238
rect -194 -272 -160 -238
rect -76 -272 -42 -238
rect 42 -272 76 -238
rect 160 -272 194 -238
rect 278 -272 312 -238
<< metal1 >>
rect -324 272 -266 278
rect -324 238 -312 272
rect -278 238 -266 272
rect -324 232 -266 238
rect -206 272 -148 278
rect -206 238 -194 272
rect -160 238 -148 272
rect -206 232 -148 238
rect -88 272 -30 278
rect -88 238 -76 272
rect -42 238 -30 272
rect -88 232 -30 238
rect 30 272 88 278
rect 30 238 42 272
rect 76 238 88 272
rect 30 232 88 238
rect 148 272 206 278
rect 148 238 160 272
rect 194 238 206 272
rect 148 232 206 238
rect 266 272 324 278
rect 266 238 278 272
rect 312 238 324 272
rect 266 232 324 238
rect -377 188 -331 200
rect -377 -188 -371 188
rect -337 -188 -331 188
rect -377 -200 -331 -188
rect -259 188 -213 200
rect -259 -188 -253 188
rect -219 -188 -213 188
rect -259 -200 -213 -188
rect -141 188 -95 200
rect -141 -188 -135 188
rect -101 -188 -95 188
rect -141 -200 -95 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 95 188 141 200
rect 95 -188 101 188
rect 135 -188 141 188
rect 95 -200 141 -188
rect 213 188 259 200
rect 213 -188 219 188
rect 253 -188 259 188
rect 213 -200 259 -188
rect 331 188 377 200
rect 331 -188 337 188
rect 371 -188 377 188
rect 331 -200 377 -188
rect -324 -238 -266 -232
rect -324 -272 -312 -238
rect -278 -272 -266 -238
rect -324 -278 -266 -272
rect -206 -238 -148 -232
rect -206 -272 -194 -238
rect -160 -272 -148 -238
rect -206 -278 -148 -272
rect -88 -238 -30 -232
rect -88 -272 -76 -238
rect -42 -272 -30 -238
rect -88 -278 -30 -272
rect 30 -238 88 -232
rect 30 -272 42 -238
rect 76 -272 88 -238
rect 30 -278 88 -272
rect 148 -238 206 -232
rect 148 -272 160 -238
rect 194 -272 206 -238
rect 148 -278 206 -272
rect 266 -238 324 -232
rect 266 -272 278 -238
rect 312 -272 324 -238
rect 266 -278 324 -272
<< properties >>
string FIXED_BBOX -468 -357 468 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
