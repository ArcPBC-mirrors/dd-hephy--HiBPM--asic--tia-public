magic
tech sky130A
magscale 1 2
timestamp 1687116508
<< locali >>
rect 100 -40 4080 60
<< metal1 >>
rect 230 3160 240 3600
rect 3940 3160 3950 3600
rect 230 1920 240 2360
rect 3940 1920 3950 2360
rect 230 1400 240 1840
rect 3940 1400 3950 1840
rect 230 160 240 600
rect 3940 160 3950 600
rect 276 -180 4028 -88
rect 226 -392 236 -212
rect 288 -392 298 -212
rect 418 -396 428 -216
rect 480 -396 490 -216
rect 610 -392 620 -212
rect 672 -392 682 -212
rect 802 -392 812 -212
rect 864 -392 874 -212
rect 994 -392 1004 -212
rect 1056 -392 1066 -212
rect 1186 -392 1196 -212
rect 1248 -392 1258 -212
rect 1378 -392 1388 -212
rect 1440 -392 1450 -212
rect 1570 -392 1580 -212
rect 1632 -392 1642 -212
rect 1762 -388 1772 -208
rect 1824 -388 1834 -208
rect 1954 -388 1964 -208
rect 2016 -388 2026 -208
rect 2146 -388 2156 -208
rect 2208 -388 2218 -208
rect 2338 -388 2348 -208
rect 2400 -388 2410 -208
rect 2530 -388 2540 -208
rect 2592 -388 2602 -208
rect 2722 -388 2732 -208
rect 2784 -388 2794 -208
rect 2914 -388 2924 -208
rect 2976 -388 2986 -208
rect 3106 -388 3116 -208
rect 3168 -388 3178 -208
rect 3298 -388 3308 -208
rect 3360 -388 3370 -208
rect 3490 -388 3500 -208
rect 3552 -388 3562 -208
rect 3682 -388 3692 -208
rect 3744 -388 3754 -208
rect 3874 -388 3884 -208
rect 3936 -388 3946 -208
rect 130 -608 140 -428
rect 192 -608 202 -428
rect 322 -608 332 -428
rect 384 -608 394 -428
rect 514 -608 524 -428
rect 576 -608 586 -428
rect 706 -608 716 -428
rect 768 -608 778 -428
rect 898 -608 908 -428
rect 960 -608 970 -428
rect 1090 -608 1100 -428
rect 1152 -608 1162 -428
rect 1282 -608 1292 -428
rect 1344 -608 1354 -428
rect 1474 -608 1484 -428
rect 1536 -608 1546 -428
rect 1666 -608 1676 -428
rect 1728 -608 1738 -428
rect 1858 -608 1868 -428
rect 1920 -608 1930 -428
rect 2050 -608 2060 -428
rect 2112 -608 2122 -428
rect 2242 -608 2252 -428
rect 2304 -608 2314 -428
rect 2434 -608 2444 -428
rect 2496 -608 2506 -428
rect 2626 -608 2636 -428
rect 2688 -608 2698 -428
rect 2818 -608 2828 -428
rect 2880 -608 2890 -428
rect 3010 -608 3020 -428
rect 3072 -608 3082 -428
rect 3202 -608 3212 -428
rect 3264 -608 3274 -428
rect 3394 -608 3404 -428
rect 3456 -608 3466 -428
rect 3586 -608 3596 -428
rect 3648 -608 3658 -428
rect 3778 -608 3788 -428
rect 3840 -608 3850 -428
rect 3970 -608 3980 -428
rect 4032 -608 4042 -428
rect 144 -732 3896 -640
<< via1 >>
rect 240 3160 3940 3600
rect 240 1920 3940 2360
rect 240 1400 3940 1840
rect 240 160 3940 600
rect 236 -392 288 -212
rect 428 -396 480 -216
rect 620 -392 672 -212
rect 812 -392 864 -212
rect 1004 -392 1056 -212
rect 1196 -392 1248 -212
rect 1388 -392 1440 -212
rect 1580 -392 1632 -212
rect 1772 -388 1824 -208
rect 1964 -388 2016 -208
rect 2156 -388 2208 -208
rect 2348 -388 2400 -208
rect 2540 -388 2592 -208
rect 2732 -388 2784 -208
rect 2924 -388 2976 -208
rect 3116 -388 3168 -208
rect 3308 -388 3360 -208
rect 3500 -388 3552 -208
rect 3692 -388 3744 -208
rect 3884 -388 3936 -208
rect 140 -608 192 -428
rect 332 -608 384 -428
rect 524 -608 576 -428
rect 716 -608 768 -428
rect 908 -608 960 -428
rect 1100 -608 1152 -428
rect 1292 -608 1344 -428
rect 1484 -608 1536 -428
rect 1676 -608 1728 -428
rect 1868 -608 1920 -428
rect 2060 -608 2112 -428
rect 2252 -608 2304 -428
rect 2444 -608 2496 -428
rect 2636 -608 2688 -428
rect 2828 -608 2880 -428
rect 3020 -608 3072 -428
rect 3212 -608 3264 -428
rect 3404 -608 3456 -428
rect 3596 -608 3648 -428
rect 3788 -608 3840 -428
rect 3980 -608 4032 -428
<< metal2 >>
rect 240 3600 3940 3610
rect 240 3150 3940 3160
rect 240 2360 3940 2370
rect 240 1910 3940 1920
rect 240 1840 3940 1850
rect 240 1390 3940 1400
rect 208 600 3940 620
rect 208 160 240 600
rect 208 -4 3940 160
rect 232 -76 3940 -4
rect 232 -144 3964 -76
rect 208 -208 3964 -144
rect 208 -212 1772 -208
rect 208 -372 236 -212
rect 288 -216 620 -212
rect 288 -340 428 -216
rect 288 -372 316 -340
rect 400 -372 428 -340
rect 236 -402 288 -392
rect 480 -340 620 -216
rect 480 -372 508 -340
rect 592 -372 620 -340
rect 428 -406 480 -396
rect 672 -340 812 -212
rect 672 -372 700 -340
rect 784 -372 812 -340
rect 620 -402 672 -392
rect 864 -340 1004 -212
rect 864 -372 892 -340
rect 976 -372 1004 -340
rect 812 -402 864 -392
rect 1056 -340 1196 -212
rect 1056 -372 1084 -340
rect 1168 -372 1196 -340
rect 1004 -402 1056 -392
rect 1248 -340 1388 -212
rect 1248 -372 1276 -340
rect 1360 -372 1388 -340
rect 1196 -402 1248 -392
rect 1440 -340 1580 -212
rect 1440 -372 1468 -340
rect 1552 -372 1580 -340
rect 1388 -402 1440 -392
rect 1632 -340 1772 -212
rect 1632 -372 1660 -340
rect 1744 -372 1772 -340
rect 1580 -402 1632 -392
rect 1824 -340 1964 -208
rect 1824 -372 1852 -340
rect 1936 -372 1964 -340
rect 1772 -398 1824 -388
rect 2016 -340 2156 -208
rect 2016 -372 2044 -340
rect 2128 -372 2156 -340
rect 1964 -398 2016 -388
rect 2208 -340 2348 -208
rect 2208 -372 2236 -340
rect 2320 -372 2348 -340
rect 2156 -398 2208 -388
rect 2400 -340 2540 -208
rect 2400 -372 2428 -340
rect 2512 -372 2540 -340
rect 2348 -398 2400 -388
rect 2592 -340 2732 -208
rect 2592 -372 2620 -340
rect 2704 -372 2732 -340
rect 2540 -398 2592 -388
rect 2784 -340 2924 -208
rect 2784 -372 2812 -340
rect 2896 -372 2924 -340
rect 2732 -398 2784 -388
rect 2976 -340 3116 -208
rect 2976 -372 3004 -340
rect 3088 -372 3116 -340
rect 2924 -398 2976 -388
rect 3168 -340 3308 -208
rect 3168 -372 3196 -340
rect 3280 -372 3308 -340
rect 3116 -398 3168 -388
rect 3360 -340 3500 -208
rect 3360 -372 3388 -340
rect 3472 -372 3500 -340
rect 3308 -398 3360 -388
rect 3552 -340 3692 -208
rect 3552 -372 3580 -340
rect 3664 -372 3692 -340
rect 3500 -398 3552 -388
rect 3744 -340 3884 -208
rect 3744 -372 3772 -340
rect 3856 -372 3884 -340
rect 3692 -398 3744 -388
rect 3936 -372 3964 -208
rect 3884 -398 3936 -388
rect 140 -428 192 -418
rect 112 -472 140 -440
rect 84 -608 140 -472
rect 332 -428 384 -418
rect 192 -472 220 -440
rect 304 -472 332 -440
rect 192 -608 332 -472
rect 524 -428 576 -418
rect 384 -472 412 -440
rect 496 -472 524 -440
rect 384 -608 524 -472
rect 716 -428 768 -418
rect 576 -472 604 -440
rect 688 -472 716 -440
rect 576 -608 716 -472
rect 908 -428 960 -418
rect 768 -472 796 -440
rect 880 -472 908 -440
rect 768 -608 908 -472
rect 1100 -428 1152 -418
rect 960 -472 988 -440
rect 1072 -472 1100 -440
rect 960 -608 1100 -472
rect 1292 -428 1344 -418
rect 1152 -472 1180 -440
rect 1264 -472 1292 -440
rect 1152 -608 1292 -472
rect 1484 -428 1536 -418
rect 1344 -472 1372 -440
rect 1456 -472 1484 -440
rect 1344 -608 1484 -472
rect 1676 -428 1728 -418
rect 1536 -472 1564 -440
rect 1648 -472 1676 -440
rect 1536 -608 1676 -472
rect 1868 -428 1920 -418
rect 1728 -472 1756 -440
rect 1840 -472 1868 -440
rect 1728 -608 1868 -472
rect 2060 -428 2112 -418
rect 1920 -472 1948 -440
rect 2032 -472 2060 -440
rect 1920 -608 2060 -472
rect 2252 -428 2304 -418
rect 2112 -472 2140 -440
rect 2224 -472 2252 -440
rect 2112 -608 2252 -472
rect 2444 -428 2496 -418
rect 2304 -472 2332 -440
rect 2416 -472 2444 -440
rect 2304 -608 2444 -472
rect 2636 -428 2688 -418
rect 2496 -472 2524 -440
rect 2608 -472 2636 -440
rect 2496 -608 2636 -472
rect 2828 -428 2880 -418
rect 2688 -472 2716 -440
rect 2800 -472 2828 -440
rect 2688 -608 2828 -472
rect 3020 -428 3072 -418
rect 2880 -472 2908 -440
rect 2992 -472 3020 -440
rect 2880 -608 3020 -472
rect 3212 -428 3264 -418
rect 3072 -472 3100 -440
rect 3184 -472 3212 -440
rect 3072 -608 3212 -472
rect 3404 -428 3456 -418
rect 3264 -472 3292 -440
rect 3376 -472 3404 -440
rect 3264 -608 3404 -472
rect 3596 -428 3648 -418
rect 3456 -472 3484 -440
rect 3568 -472 3596 -440
rect 3456 -608 3596 -472
rect 3788 -428 3840 -418
rect 3648 -472 3676 -440
rect 3760 -472 3788 -440
rect 3648 -608 3788 -472
rect 3980 -428 4032 -418
rect 3840 -472 3868 -440
rect 3952 -472 3980 -440
rect 3840 -608 3980 -472
rect 4032 -472 4060 -440
rect 4032 -608 4136 -472
rect 84 -816 4136 -608
<< via2 >>
rect 240 3160 520 3600
rect 1000 3160 1280 3600
rect 1760 3160 2040 3600
rect 2520 3160 2800 3600
rect 3280 3160 3560 3600
rect 620 1940 900 2360
rect 1380 1940 1660 2360
rect 2140 1940 2420 2360
rect 2900 1940 3180 2360
rect 3660 1940 3940 2360
rect 240 1400 520 1840
rect 1000 1400 1280 1840
rect 1760 1400 2040 1840
rect 2520 1400 2800 1840
rect 3280 1400 3560 1840
rect 620 160 900 600
rect 1380 160 1660 600
rect 2140 160 2420 600
rect 2900 160 3180 600
rect 3640 160 3920 600
<< metal3 >>
rect 80 3720 4100 4040
rect 220 3600 540 3720
rect 220 3160 240 3600
rect 520 3160 540 3600
rect 220 1840 540 3160
rect 980 3600 1300 3720
rect 980 3160 1000 3600
rect 1280 3160 1300 3600
rect 620 2365 920 2380
rect 610 2360 920 2365
rect 610 1940 620 2360
rect 900 1940 920 2360
rect 610 1935 920 1940
rect 220 1400 240 1840
rect 520 1400 540 1840
rect 220 1380 540 1400
rect 620 605 920 1935
rect 980 1840 1300 3160
rect 1740 3600 2060 3720
rect 1740 3160 1760 3600
rect 2040 3160 2060 3600
rect 980 1400 1000 1840
rect 1280 1400 1300 1840
rect 980 1380 1300 1400
rect 1360 2365 1660 2380
rect 1360 2360 1670 2365
rect 1360 1940 1380 2360
rect 1660 1940 1670 2360
rect 1360 1935 1670 1940
rect 610 600 920 605
rect 610 160 620 600
rect 900 160 920 600
rect 1360 605 1660 1935
rect 1740 1840 2060 3160
rect 2500 3600 2820 3720
rect 2500 3160 2520 3600
rect 2800 3160 2820 3600
rect 1740 1400 1760 1840
rect 2040 1400 2060 1840
rect 1740 1380 2060 1400
rect 2120 2365 2420 2380
rect 2120 2360 2430 2365
rect 2120 1940 2140 2360
rect 2420 1940 2430 2360
rect 2120 1935 2430 1940
rect 2120 605 2420 1935
rect 2500 1840 2820 3160
rect 3260 3600 3580 3720
rect 3260 3160 3280 3600
rect 3560 3160 3580 3600
rect 2500 1400 2520 1840
rect 2800 1400 2820 1840
rect 2500 1380 2820 1400
rect 2880 2365 3180 2380
rect 2880 2360 3190 2365
rect 2880 1940 2900 2360
rect 3180 1940 3190 2360
rect 2880 1935 3190 1940
rect 2880 605 3180 1935
rect 3260 1840 3580 3160
rect 3260 1400 3280 1840
rect 3560 1400 3580 1840
rect 3260 1380 3580 1400
rect 3640 2365 3940 2380
rect 3640 2360 3950 2365
rect 3640 1940 3660 2360
rect 3940 1940 3950 2360
rect 3640 1935 3950 1940
rect 3640 605 3940 1935
rect 1360 600 1670 605
rect 1360 160 1380 600
rect 1660 160 1670 600
rect 2120 600 2430 605
rect 2120 160 2140 600
rect 2420 160 2430 600
rect 2880 600 3190 605
rect 2880 160 2900 600
rect 3180 160 3190 600
rect 610 155 910 160
rect 1370 155 1670 160
rect 2130 155 2430 160
rect 2890 155 3190 160
rect 3630 600 3940 605
rect 3630 160 3640 600
rect 3920 160 3940 600
rect 3630 155 3930 160
use sky130_fd_pr__nfet_01v8_lvt_U9F2PH  sky130_fd_pr__nfet_01v8_lvt_U9F2PH_0
timestamp 1685105324
transform 1 0 2087 0 1 -410
box -2087 -410 2087 410
use sky130_fd_pr__res_high_po_1p41_YU66GB  sky130_fd_pr__res_high_po_1p41_YU66GB_0
timestamp 1685105324
transform 1 0 2088 0 1 1882
box -2008 -1882 2008 1882
<< end >>
