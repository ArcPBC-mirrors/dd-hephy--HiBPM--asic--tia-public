magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< error_p >>
rect -365 281 -307 287
rect -173 281 -115 287
rect 19 281 77 287
rect 211 281 269 287
rect 403 281 461 287
rect -365 247 -353 281
rect -173 247 -161 281
rect 19 247 31 281
rect 211 247 223 281
rect 403 247 415 281
rect -365 241 -307 247
rect -173 241 -115 247
rect 19 241 77 247
rect 211 241 269 247
rect 403 241 461 247
rect -461 -247 -403 -241
rect -269 -247 -211 -241
rect -77 -247 -19 -241
rect 115 -247 173 -241
rect 307 -247 365 -241
rect -461 -281 -449 -247
rect -269 -281 -257 -247
rect -77 -281 -65 -247
rect 115 -281 127 -247
rect 307 -281 319 -247
rect -461 -287 -403 -281
rect -269 -287 -211 -281
rect -77 -287 -19 -281
rect 115 -287 173 -281
rect 307 -287 365 -281
<< nwell >>
rect -647 -419 647 419
<< pmos >>
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
<< pdiff >>
rect -509 188 -447 200
rect -509 -188 -497 188
rect -463 -188 -447 188
rect -509 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 509 200
rect 447 -188 463 188
rect 497 -188 509 188
rect 447 -200 509 -188
<< pdiffc >>
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
<< nsubdiff >>
rect -611 349 -515 383
rect 515 349 611 383
rect -611 287 -577 349
rect 577 287 611 349
rect -611 -349 -577 -287
rect 577 -349 611 -287
rect -611 -383 -515 -349
rect 515 -383 611 -349
<< nsubdiffcont >>
rect -515 349 515 383
rect -611 -287 -577 287
rect 577 -287 611 287
rect -515 -383 515 -349
<< poly >>
rect -369 281 -303 297
rect -369 247 -353 281
rect -319 247 -303 281
rect -369 231 -303 247
rect -177 281 -111 297
rect -177 247 -161 281
rect -127 247 -111 281
rect -177 231 -111 247
rect 15 281 81 297
rect 15 247 31 281
rect 65 247 81 281
rect 15 231 81 247
rect 207 281 273 297
rect 207 247 223 281
rect 257 247 273 281
rect 207 231 273 247
rect 399 281 465 297
rect 399 247 415 281
rect 449 247 465 281
rect 399 231 465 247
rect -447 200 -417 226
rect -351 200 -321 231
rect -255 200 -225 226
rect -159 200 -129 231
rect -63 200 -33 226
rect 33 200 63 231
rect 129 200 159 226
rect 225 200 255 231
rect 321 200 351 226
rect 417 200 447 231
rect -447 -231 -417 -200
rect -351 -226 -321 -200
rect -255 -231 -225 -200
rect -159 -226 -129 -200
rect -63 -231 -33 -200
rect 33 -226 63 -200
rect 129 -231 159 -200
rect 225 -226 255 -200
rect 321 -231 351 -200
rect 417 -226 447 -200
rect -465 -247 -399 -231
rect -465 -281 -449 -247
rect -415 -281 -399 -247
rect -465 -297 -399 -281
rect -273 -247 -207 -231
rect -273 -281 -257 -247
rect -223 -281 -207 -247
rect -273 -297 -207 -281
rect -81 -247 -15 -231
rect -81 -281 -65 -247
rect -31 -281 -15 -247
rect -81 -297 -15 -281
rect 111 -247 177 -231
rect 111 -281 127 -247
rect 161 -281 177 -247
rect 111 -297 177 -281
rect 303 -247 369 -231
rect 303 -281 319 -247
rect 353 -281 369 -247
rect 303 -297 369 -281
<< polycont >>
rect -353 247 -319 281
rect -161 247 -127 281
rect 31 247 65 281
rect 223 247 257 281
rect 415 247 449 281
rect -449 -281 -415 -247
rect -257 -281 -223 -247
rect -65 -281 -31 -247
rect 127 -281 161 -247
rect 319 -281 353 -247
<< locali >>
rect -611 349 -515 383
rect 515 349 611 383
rect -611 287 -577 349
rect 577 287 611 349
rect -369 247 -353 281
rect -319 247 -303 281
rect -177 247 -161 281
rect -127 247 -111 281
rect 15 247 31 281
rect 65 247 81 281
rect 207 247 223 281
rect 257 247 273 281
rect 399 247 415 281
rect 449 247 465 281
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect -465 -281 -449 -247
rect -415 -281 -399 -247
rect -273 -281 -257 -247
rect -223 -281 -207 -247
rect -81 -281 -65 -247
rect -31 -281 -15 -247
rect 111 -281 127 -247
rect 161 -281 177 -247
rect 303 -281 319 -247
rect 353 -281 369 -247
rect -611 -349 -577 -287
rect 577 -349 611 -287
rect -611 -383 -515 -349
rect 515 -383 611 -349
<< viali >>
rect -353 247 -319 281
rect -161 247 -127 281
rect 31 247 65 281
rect 223 247 257 281
rect 415 247 449 281
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -449 -281 -415 -247
rect -257 -281 -223 -247
rect -65 -281 -31 -247
rect 127 -281 161 -247
rect 319 -281 353 -247
<< metal1 >>
rect -365 281 -307 287
rect -365 247 -353 281
rect -319 247 -307 281
rect -365 241 -307 247
rect -173 281 -115 287
rect -173 247 -161 281
rect -127 247 -115 281
rect -173 241 -115 247
rect 19 281 77 287
rect 19 247 31 281
rect 65 247 77 281
rect 19 241 77 247
rect 211 281 269 287
rect 211 247 223 281
rect 257 247 269 281
rect 211 241 269 247
rect 403 281 461 287
rect 403 247 415 281
rect 449 247 461 281
rect 403 241 461 247
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect -461 -247 -403 -241
rect -461 -281 -449 -247
rect -415 -281 -403 -247
rect -461 -287 -403 -281
rect -269 -247 -211 -241
rect -269 -281 -257 -247
rect -223 -281 -211 -247
rect -269 -287 -211 -281
rect -77 -247 -19 -241
rect -77 -281 -65 -247
rect -31 -281 -19 -247
rect -77 -287 -19 -281
rect 115 -247 173 -241
rect 115 -281 127 -247
rect 161 -281 173 -247
rect 115 -287 173 -281
rect 307 -247 365 -241
rect 307 -281 319 -247
rect 353 -281 365 -247
rect 307 -287 365 -281
<< properties >>
string FIXED_BBOX -594 -366 594 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
