magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< error_p >>
rect -365 890 -307 896
rect -173 890 -115 896
rect 19 890 77 896
rect 211 890 269 896
rect 403 890 461 896
rect -365 856 -353 890
rect -173 856 -161 890
rect 19 856 31 890
rect 211 856 223 890
rect 403 856 415 890
rect -365 850 -307 856
rect -173 850 -115 856
rect 19 850 77 856
rect 211 850 269 856
rect 403 850 461 856
rect -461 380 -403 386
rect -269 380 -211 386
rect -77 380 -19 386
rect 115 380 173 386
rect 307 380 365 386
rect -461 346 -449 380
rect -269 346 -257 380
rect -77 346 -65 380
rect 115 346 127 380
rect 307 346 319 380
rect -461 340 -403 346
rect -269 340 -211 346
rect -77 340 -19 346
rect 115 340 173 346
rect 307 340 365 346
rect -461 272 -403 278
rect -269 272 -211 278
rect -77 272 -19 278
rect 115 272 173 278
rect 307 272 365 278
rect -461 238 -449 272
rect -269 238 -257 272
rect -77 238 -65 272
rect 115 238 127 272
rect 307 238 319 272
rect -461 232 -403 238
rect -269 232 -211 238
rect -77 232 -19 238
rect 115 232 173 238
rect 307 232 365 238
rect -365 -238 -307 -232
rect -173 -238 -115 -232
rect 19 -238 77 -232
rect 211 -238 269 -232
rect 403 -238 461 -232
rect -365 -272 -353 -238
rect -173 -272 -161 -238
rect 19 -272 31 -238
rect 211 -272 223 -238
rect 403 -272 415 -238
rect -365 -278 -307 -272
rect -173 -278 -115 -272
rect 19 -278 77 -272
rect 211 -278 269 -272
rect 403 -278 461 -272
rect -365 -346 -307 -340
rect -173 -346 -115 -340
rect 19 -346 77 -340
rect 211 -346 269 -340
rect 403 -346 461 -340
rect -365 -380 -353 -346
rect -173 -380 -161 -346
rect 19 -380 31 -346
rect 211 -380 223 -346
rect 403 -380 415 -346
rect -365 -386 -307 -380
rect -173 -386 -115 -380
rect 19 -386 77 -380
rect 211 -386 269 -380
rect 403 -386 461 -380
rect -461 -856 -403 -850
rect -269 -856 -211 -850
rect -77 -856 -19 -850
rect 115 -856 173 -850
rect 307 -856 365 -850
rect -461 -890 -449 -856
rect -269 -890 -257 -856
rect -77 -890 -65 -856
rect 115 -890 127 -856
rect 307 -890 319 -856
rect -461 -896 -403 -890
rect -269 -896 -211 -890
rect -77 -896 -19 -890
rect 115 -896 173 -890
rect 307 -896 365 -890
<< pwell >>
rect -647 -1028 647 1028
<< nmoslvt >>
rect -447 418 -417 818
rect -351 418 -321 818
rect -255 418 -225 818
rect -159 418 -129 818
rect -63 418 -33 818
rect 33 418 63 818
rect 129 418 159 818
rect 225 418 255 818
rect 321 418 351 818
rect 417 418 447 818
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect -447 -818 -417 -418
rect -351 -818 -321 -418
rect -255 -818 -225 -418
rect -159 -818 -129 -418
rect -63 -818 -33 -418
rect 33 -818 63 -418
rect 129 -818 159 -418
rect 225 -818 255 -418
rect 321 -818 351 -418
rect 417 -818 447 -418
<< ndiff >>
rect -509 806 -447 818
rect -509 430 -497 806
rect -463 430 -447 806
rect -509 418 -447 430
rect -417 806 -351 818
rect -417 430 -401 806
rect -367 430 -351 806
rect -417 418 -351 430
rect -321 806 -255 818
rect -321 430 -305 806
rect -271 430 -255 806
rect -321 418 -255 430
rect -225 806 -159 818
rect -225 430 -209 806
rect -175 430 -159 806
rect -225 418 -159 430
rect -129 806 -63 818
rect -129 430 -113 806
rect -79 430 -63 806
rect -129 418 -63 430
rect -33 806 33 818
rect -33 430 -17 806
rect 17 430 33 806
rect -33 418 33 430
rect 63 806 129 818
rect 63 430 79 806
rect 113 430 129 806
rect 63 418 129 430
rect 159 806 225 818
rect 159 430 175 806
rect 209 430 225 806
rect 159 418 225 430
rect 255 806 321 818
rect 255 430 271 806
rect 305 430 321 806
rect 255 418 321 430
rect 351 806 417 818
rect 351 430 367 806
rect 401 430 417 806
rect 351 418 417 430
rect 447 806 509 818
rect 447 430 463 806
rect 497 430 509 806
rect 447 418 509 430
rect -509 188 -447 200
rect -509 -188 -497 188
rect -463 -188 -447 188
rect -509 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 509 200
rect 447 -188 463 188
rect 497 -188 509 188
rect 447 -200 509 -188
rect -509 -430 -447 -418
rect -509 -806 -497 -430
rect -463 -806 -447 -430
rect -509 -818 -447 -806
rect -417 -430 -351 -418
rect -417 -806 -401 -430
rect -367 -806 -351 -430
rect -417 -818 -351 -806
rect -321 -430 -255 -418
rect -321 -806 -305 -430
rect -271 -806 -255 -430
rect -321 -818 -255 -806
rect -225 -430 -159 -418
rect -225 -806 -209 -430
rect -175 -806 -159 -430
rect -225 -818 -159 -806
rect -129 -430 -63 -418
rect -129 -806 -113 -430
rect -79 -806 -63 -430
rect -129 -818 -63 -806
rect -33 -430 33 -418
rect -33 -806 -17 -430
rect 17 -806 33 -430
rect -33 -818 33 -806
rect 63 -430 129 -418
rect 63 -806 79 -430
rect 113 -806 129 -430
rect 63 -818 129 -806
rect 159 -430 225 -418
rect 159 -806 175 -430
rect 209 -806 225 -430
rect 159 -818 225 -806
rect 255 -430 321 -418
rect 255 -806 271 -430
rect 305 -806 321 -430
rect 255 -818 321 -806
rect 351 -430 417 -418
rect 351 -806 367 -430
rect 401 -806 417 -430
rect 351 -818 417 -806
rect 447 -430 509 -418
rect 447 -806 463 -430
rect 497 -806 509 -430
rect 447 -818 509 -806
<< ndiffc >>
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
<< psubdiff >>
rect -611 958 -515 992
rect 515 958 611 992
rect -611 896 -577 958
rect 577 896 611 958
rect -611 -958 -577 -896
rect 577 -958 611 -896
rect -611 -992 -515 -958
rect 515 -992 611 -958
<< psubdiffcont >>
rect -515 958 515 992
rect -611 -896 -577 896
rect 577 -896 611 896
rect -515 -992 515 -958
<< poly >>
rect -369 890 -303 906
rect -369 856 -353 890
rect -319 856 -303 890
rect -447 818 -417 844
rect -369 840 -303 856
rect -177 890 -111 906
rect -177 856 -161 890
rect -127 856 -111 890
rect -351 818 -321 840
rect -255 818 -225 844
rect -177 840 -111 856
rect 15 890 81 906
rect 15 856 31 890
rect 65 856 81 890
rect -159 818 -129 840
rect -63 818 -33 844
rect 15 840 81 856
rect 207 890 273 906
rect 207 856 223 890
rect 257 856 273 890
rect 33 818 63 840
rect 129 818 159 844
rect 207 840 273 856
rect 399 890 465 906
rect 399 856 415 890
rect 449 856 465 890
rect 225 818 255 840
rect 321 818 351 844
rect 399 840 465 856
rect 417 818 447 840
rect -447 396 -417 418
rect -465 380 -399 396
rect -351 392 -321 418
rect -255 396 -225 418
rect -465 346 -449 380
rect -415 346 -399 380
rect -465 330 -399 346
rect -273 380 -207 396
rect -159 392 -129 418
rect -63 396 -33 418
rect -273 346 -257 380
rect -223 346 -207 380
rect -273 330 -207 346
rect -81 380 -15 396
rect 33 392 63 418
rect 129 396 159 418
rect -81 346 -65 380
rect -31 346 -15 380
rect -81 330 -15 346
rect 111 380 177 396
rect 225 392 255 418
rect 321 396 351 418
rect 111 346 127 380
rect 161 346 177 380
rect 111 330 177 346
rect 303 380 369 396
rect 417 392 447 418
rect 303 346 319 380
rect 353 346 369 380
rect 303 330 369 346
rect -465 272 -399 288
rect -465 238 -449 272
rect -415 238 -399 272
rect -465 222 -399 238
rect -273 272 -207 288
rect -273 238 -257 272
rect -223 238 -207 272
rect -447 200 -417 222
rect -351 200 -321 226
rect -273 222 -207 238
rect -81 272 -15 288
rect -81 238 -65 272
rect -31 238 -15 272
rect -255 200 -225 222
rect -159 200 -129 226
rect -81 222 -15 238
rect 111 272 177 288
rect 111 238 127 272
rect 161 238 177 272
rect -63 200 -33 222
rect 33 200 63 226
rect 111 222 177 238
rect 303 272 369 288
rect 303 238 319 272
rect 353 238 369 272
rect 129 200 159 222
rect 225 200 255 226
rect 303 222 369 238
rect 321 200 351 222
rect 417 200 447 226
rect -447 -226 -417 -200
rect -351 -222 -321 -200
rect -369 -238 -303 -222
rect -255 -226 -225 -200
rect -159 -222 -129 -200
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -369 -288 -303 -272
rect -177 -238 -111 -222
rect -63 -226 -33 -200
rect 33 -222 63 -200
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect -177 -288 -111 -272
rect 15 -238 81 -222
rect 129 -226 159 -200
rect 225 -222 255 -200
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 15 -288 81 -272
rect 207 -238 273 -222
rect 321 -226 351 -200
rect 417 -222 447 -200
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 207 -288 273 -272
rect 399 -238 465 -222
rect 399 -272 415 -238
rect 449 -272 465 -238
rect 399 -288 465 -272
rect -369 -346 -303 -330
rect -369 -380 -353 -346
rect -319 -380 -303 -346
rect -447 -418 -417 -392
rect -369 -396 -303 -380
rect -177 -346 -111 -330
rect -177 -380 -161 -346
rect -127 -380 -111 -346
rect -351 -418 -321 -396
rect -255 -418 -225 -392
rect -177 -396 -111 -380
rect 15 -346 81 -330
rect 15 -380 31 -346
rect 65 -380 81 -346
rect -159 -418 -129 -396
rect -63 -418 -33 -392
rect 15 -396 81 -380
rect 207 -346 273 -330
rect 207 -380 223 -346
rect 257 -380 273 -346
rect 33 -418 63 -396
rect 129 -418 159 -392
rect 207 -396 273 -380
rect 399 -346 465 -330
rect 399 -380 415 -346
rect 449 -380 465 -346
rect 225 -418 255 -396
rect 321 -418 351 -392
rect 399 -396 465 -380
rect 417 -418 447 -396
rect -447 -840 -417 -818
rect -465 -856 -399 -840
rect -351 -844 -321 -818
rect -255 -840 -225 -818
rect -465 -890 -449 -856
rect -415 -890 -399 -856
rect -465 -906 -399 -890
rect -273 -856 -207 -840
rect -159 -844 -129 -818
rect -63 -840 -33 -818
rect -273 -890 -257 -856
rect -223 -890 -207 -856
rect -273 -906 -207 -890
rect -81 -856 -15 -840
rect 33 -844 63 -818
rect 129 -840 159 -818
rect -81 -890 -65 -856
rect -31 -890 -15 -856
rect -81 -906 -15 -890
rect 111 -856 177 -840
rect 225 -844 255 -818
rect 321 -840 351 -818
rect 111 -890 127 -856
rect 161 -890 177 -856
rect 111 -906 177 -890
rect 303 -856 369 -840
rect 417 -844 447 -818
rect 303 -890 319 -856
rect 353 -890 369 -856
rect 303 -906 369 -890
<< polycont >>
rect -353 856 -319 890
rect -161 856 -127 890
rect 31 856 65 890
rect 223 856 257 890
rect 415 856 449 890
rect -449 346 -415 380
rect -257 346 -223 380
rect -65 346 -31 380
rect 127 346 161 380
rect 319 346 353 380
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
rect -353 -380 -319 -346
rect -161 -380 -127 -346
rect 31 -380 65 -346
rect 223 -380 257 -346
rect 415 -380 449 -346
rect -449 -890 -415 -856
rect -257 -890 -223 -856
rect -65 -890 -31 -856
rect 127 -890 161 -856
rect 319 -890 353 -856
<< locali >>
rect -611 958 -515 992
rect 515 958 611 992
rect -611 896 -577 958
rect 577 896 611 958
rect -369 856 -353 890
rect -319 856 -303 890
rect -177 856 -161 890
rect -127 856 -111 890
rect 15 856 31 890
rect 65 856 81 890
rect 207 856 223 890
rect 257 856 273 890
rect 399 856 415 890
rect 449 856 465 890
rect -497 806 -463 822
rect -497 414 -463 430
rect -401 806 -367 822
rect -401 414 -367 430
rect -305 806 -271 822
rect -305 414 -271 430
rect -209 806 -175 822
rect -209 414 -175 430
rect -113 806 -79 822
rect -113 414 -79 430
rect -17 806 17 822
rect -17 414 17 430
rect 79 806 113 822
rect 79 414 113 430
rect 175 806 209 822
rect 175 414 209 430
rect 271 806 305 822
rect 271 414 305 430
rect 367 806 401 822
rect 367 414 401 430
rect 463 806 497 822
rect 463 414 497 430
rect -465 346 -449 380
rect -415 346 -399 380
rect -273 346 -257 380
rect -223 346 -207 380
rect -81 346 -65 380
rect -31 346 -15 380
rect 111 346 127 380
rect 161 346 177 380
rect 303 346 319 380
rect 353 346 369 380
rect -465 238 -449 272
rect -415 238 -399 272
rect -273 238 -257 272
rect -223 238 -207 272
rect -81 238 -65 272
rect -31 238 -15 272
rect 111 238 127 272
rect 161 238 177 272
rect 303 238 319 272
rect 353 238 369 272
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 399 -272 415 -238
rect 449 -272 465 -238
rect -369 -380 -353 -346
rect -319 -380 -303 -346
rect -177 -380 -161 -346
rect -127 -380 -111 -346
rect 15 -380 31 -346
rect 65 -380 81 -346
rect 207 -380 223 -346
rect 257 -380 273 -346
rect 399 -380 415 -346
rect 449 -380 465 -346
rect -497 -430 -463 -414
rect -497 -822 -463 -806
rect -401 -430 -367 -414
rect -401 -822 -367 -806
rect -305 -430 -271 -414
rect -305 -822 -271 -806
rect -209 -430 -175 -414
rect -209 -822 -175 -806
rect -113 -430 -79 -414
rect -113 -822 -79 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 79 -430 113 -414
rect 79 -822 113 -806
rect 175 -430 209 -414
rect 175 -822 209 -806
rect 271 -430 305 -414
rect 271 -822 305 -806
rect 367 -430 401 -414
rect 367 -822 401 -806
rect 463 -430 497 -414
rect 463 -822 497 -806
rect -465 -890 -449 -856
rect -415 -890 -399 -856
rect -273 -890 -257 -856
rect -223 -890 -207 -856
rect -81 -890 -65 -856
rect -31 -890 -15 -856
rect 111 -890 127 -856
rect 161 -890 177 -856
rect 303 -890 319 -856
rect 353 -890 369 -856
rect -611 -958 -577 -896
rect 577 -958 611 -896
rect -611 -992 -515 -958
rect 515 -992 611 -958
<< viali >>
rect -353 856 -319 890
rect -161 856 -127 890
rect 31 856 65 890
rect 223 856 257 890
rect 415 856 449 890
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect -449 346 -415 380
rect -257 346 -223 380
rect -65 346 -31 380
rect 127 346 161 380
rect 319 346 353 380
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
rect -353 -380 -319 -346
rect -161 -380 -127 -346
rect 31 -380 65 -346
rect 223 -380 257 -346
rect 415 -380 449 -346
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect -449 -890 -415 -856
rect -257 -890 -223 -856
rect -65 -890 -31 -856
rect 127 -890 161 -856
rect 319 -890 353 -856
<< metal1 >>
rect -365 890 -307 896
rect -365 856 -353 890
rect -319 856 -307 890
rect -365 850 -307 856
rect -173 890 -115 896
rect -173 856 -161 890
rect -127 856 -115 890
rect -173 850 -115 856
rect 19 890 77 896
rect 19 856 31 890
rect 65 856 77 890
rect 19 850 77 856
rect 211 890 269 896
rect 211 856 223 890
rect 257 856 269 890
rect 211 850 269 856
rect 403 890 461 896
rect 403 856 415 890
rect 449 856 461 890
rect 403 850 461 856
rect -503 806 -457 818
rect -503 430 -497 806
rect -463 430 -457 806
rect -503 418 -457 430
rect -407 806 -361 818
rect -407 430 -401 806
rect -367 430 -361 806
rect -407 418 -361 430
rect -311 806 -265 818
rect -311 430 -305 806
rect -271 430 -265 806
rect -311 418 -265 430
rect -215 806 -169 818
rect -215 430 -209 806
rect -175 430 -169 806
rect -215 418 -169 430
rect -119 806 -73 818
rect -119 430 -113 806
rect -79 430 -73 806
rect -119 418 -73 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 73 806 119 818
rect 73 430 79 806
rect 113 430 119 806
rect 73 418 119 430
rect 169 806 215 818
rect 169 430 175 806
rect 209 430 215 806
rect 169 418 215 430
rect 265 806 311 818
rect 265 430 271 806
rect 305 430 311 806
rect 265 418 311 430
rect 361 806 407 818
rect 361 430 367 806
rect 401 430 407 806
rect 361 418 407 430
rect 457 806 503 818
rect 457 430 463 806
rect 497 430 503 806
rect 457 418 503 430
rect -461 380 -403 386
rect -461 346 -449 380
rect -415 346 -403 380
rect -461 340 -403 346
rect -269 380 -211 386
rect -269 346 -257 380
rect -223 346 -211 380
rect -269 340 -211 346
rect -77 380 -19 386
rect -77 346 -65 380
rect -31 346 -19 380
rect -77 340 -19 346
rect 115 380 173 386
rect 115 346 127 380
rect 161 346 173 380
rect 115 340 173 346
rect 307 380 365 386
rect 307 346 319 380
rect 353 346 365 380
rect 307 340 365 346
rect -461 272 -403 278
rect -461 238 -449 272
rect -415 238 -403 272
rect -461 232 -403 238
rect -269 272 -211 278
rect -269 238 -257 272
rect -223 238 -211 272
rect -269 232 -211 238
rect -77 272 -19 278
rect -77 238 -65 272
rect -31 238 -19 272
rect -77 232 -19 238
rect 115 272 173 278
rect 115 238 127 272
rect 161 238 173 272
rect 115 232 173 238
rect 307 272 365 278
rect 307 238 319 272
rect 353 238 365 272
rect 307 232 365 238
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect -365 -238 -307 -232
rect -365 -272 -353 -238
rect -319 -272 -307 -238
rect -365 -278 -307 -272
rect -173 -238 -115 -232
rect -173 -272 -161 -238
rect -127 -272 -115 -238
rect -173 -278 -115 -272
rect 19 -238 77 -232
rect 19 -272 31 -238
rect 65 -272 77 -238
rect 19 -278 77 -272
rect 211 -238 269 -232
rect 211 -272 223 -238
rect 257 -272 269 -238
rect 211 -278 269 -272
rect 403 -238 461 -232
rect 403 -272 415 -238
rect 449 -272 461 -238
rect 403 -278 461 -272
rect -365 -346 -307 -340
rect -365 -380 -353 -346
rect -319 -380 -307 -346
rect -365 -386 -307 -380
rect -173 -346 -115 -340
rect -173 -380 -161 -346
rect -127 -380 -115 -346
rect -173 -386 -115 -380
rect 19 -346 77 -340
rect 19 -380 31 -346
rect 65 -380 77 -346
rect 19 -386 77 -380
rect 211 -346 269 -340
rect 211 -380 223 -346
rect 257 -380 269 -346
rect 211 -386 269 -380
rect 403 -346 461 -340
rect 403 -380 415 -346
rect 449 -380 461 -346
rect 403 -386 461 -380
rect -503 -430 -457 -418
rect -503 -806 -497 -430
rect -463 -806 -457 -430
rect -503 -818 -457 -806
rect -407 -430 -361 -418
rect -407 -806 -401 -430
rect -367 -806 -361 -430
rect -407 -818 -361 -806
rect -311 -430 -265 -418
rect -311 -806 -305 -430
rect -271 -806 -265 -430
rect -311 -818 -265 -806
rect -215 -430 -169 -418
rect -215 -806 -209 -430
rect -175 -806 -169 -430
rect -215 -818 -169 -806
rect -119 -430 -73 -418
rect -119 -806 -113 -430
rect -79 -806 -73 -430
rect -119 -818 -73 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 73 -430 119 -418
rect 73 -806 79 -430
rect 113 -806 119 -430
rect 73 -818 119 -806
rect 169 -430 215 -418
rect 169 -806 175 -430
rect 209 -806 215 -430
rect 169 -818 215 -806
rect 265 -430 311 -418
rect 265 -806 271 -430
rect 305 -806 311 -430
rect 265 -818 311 -806
rect 361 -430 407 -418
rect 361 -806 367 -430
rect 401 -806 407 -430
rect 361 -818 407 -806
rect 457 -430 503 -418
rect 457 -806 463 -430
rect 497 -806 503 -430
rect 457 -818 503 -806
rect -461 -856 -403 -850
rect -461 -890 -449 -856
rect -415 -890 -403 -856
rect -461 -896 -403 -890
rect -269 -856 -211 -850
rect -269 -890 -257 -856
rect -223 -890 -211 -856
rect -269 -896 -211 -890
rect -77 -856 -19 -850
rect -77 -890 -65 -856
rect -31 -890 -19 -856
rect -77 -896 -19 -890
rect 115 -856 173 -850
rect 115 -890 127 -856
rect 161 -890 173 -856
rect 115 -896 173 -890
rect 307 -856 365 -850
rect 307 -890 319 -856
rect 353 -890 365 -856
rect 307 -896 365 -890
<< properties >>
string FIXED_BBOX -594 -975 594 975
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 3 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
