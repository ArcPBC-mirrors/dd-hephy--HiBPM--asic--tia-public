magic
tech sky130A
magscale 1 2
timestamp 1685028972
<< metal3 >>
rect -2686 212 2686 240
rect -2686 -212 2602 212
rect 2666 -212 2686 212
rect -2686 -240 2686 -212
<< via3 >>
rect 2602 -212 2666 212
<< mimcap >>
rect -2646 160 2354 200
rect -2646 -160 -2606 160
rect 2314 -160 2354 160
rect -2646 -200 2354 -160
<< mimcapcontact >>
rect -2606 -160 2314 160
<< metal4 >>
rect 2586 212 2682 228
rect -2607 160 2315 161
rect -2607 -160 -2606 160
rect 2314 -160 2315 160
rect -2607 -161 2315 -160
rect 2586 -212 2602 212
rect 2666 -212 2682 212
rect 2586 -228 2682 -212
<< properties >>
string FIXED_BBOX -2686 -240 2394 240
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25 l 2.00 val 110.26 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
