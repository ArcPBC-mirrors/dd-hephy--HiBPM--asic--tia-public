magic
tech sky130A
magscale 1 2
timestamp 1684166381
<< pwell >>
rect 14566 13206 17674 15634
rect 14566 9082 17674 11510
rect 16400 5066 17718 7334
<< psubdiff >>
rect 8476 13900 8500 15280
rect 10040 13900 10064 15280
<< psubdiffcont >>
rect 8500 13900 10040 15280
<< locali >>
rect 8484 14040 8500 15280
rect -40 14020 8500 14040
rect -280 13900 8500 14020
rect 10040 14620 10056 15280
rect 10420 13900 11080 14620
rect -280 13760 11080 13900
rect 12442 13858 12652 13938
rect 12296 13760 12652 13858
rect -280 13460 12652 13760
rect -280 -2300 80 13460
rect 9900 13448 12652 13460
rect 9900 13440 12534 13448
rect 11060 13420 12440 13440
rect 12920 13380 13200 13440
rect 12900 8480 13220 13380
rect 18900 9790 19320 9800
rect 18900 9700 21010 9790
rect 12920 7330 13200 8480
rect 18900 7440 21010 7530
rect 12920 7320 13250 7330
rect 12920 7220 13340 7320
rect 12930 6180 13340 7220
rect 12930 6170 13260 6180
rect 12980 5000 13260 6170
rect 18880 5290 18930 5340
rect 18880 5200 20360 5290
rect 12910 4810 13280 5000
rect 12940 1720 13280 4810
rect 12910 1540 13280 1720
rect 18880 3010 18930 5200
rect 18880 2920 20360 3010
rect 12910 1340 18620 1540
rect 12880 1310 18620 1340
rect 12880 -860 13440 1310
rect 16580 -840 16820 1310
rect 18020 -1180 18620 1310
rect 13060 -2140 13220 -1360
rect 18260 -2140 18420 -1360
rect 18530 -1560 18620 -1180
rect 18880 760 18930 2920
rect 18880 670 20360 760
rect 18880 -1560 18930 670
rect -280 -2540 18540 -2300
rect 40 -2560 18540 -2540
rect 20760 -4780 21220 -4120
<< viali >>
rect 9300 14620 9800 15280
rect 9300 13900 10040 14620
rect 10040 13900 10420 14620
rect 17920 6300 18040 6480
rect 16446 5046 16624 5142
<< metal1 >>
rect 17670 15580 17680 15780
rect 17790 15580 17800 15780
rect 9294 15280 9806 15292
rect 9290 13900 9300 15280
rect 9800 14626 9810 15280
rect 9800 14620 10432 14626
rect 10420 13900 10432 14620
rect 12990 14600 13000 14720
rect 13080 14600 13090 14720
rect 17420 14360 17840 14480
rect 18000 14360 18010 14480
rect 12970 14080 12980 14200
rect 13060 14080 13070 14200
rect 13970 13980 13980 14100
rect 14100 14098 14140 14100
rect 14200 14098 14360 14100
rect 14100 13980 14360 14098
rect 14132 13976 14228 13980
rect 9294 13894 10432 13900
rect 9294 13888 9806 13894
rect 12320 13740 12400 13800
rect 12320 13620 12520 13740
rect 12620 13620 12630 13740
rect 14900 11260 15040 13440
rect 17670 12400 17680 12580
rect 17980 12400 17990 12580
rect 17680 11480 17980 12400
rect 18800 11840 19020 11920
rect 18800 10980 18960 11840
rect 17420 10230 17540 10360
rect 14030 9840 14040 9980
rect 14180 9840 14360 9980
rect 18800 9920 18980 10980
rect 18800 9840 19040 9920
rect 18800 9660 18980 9840
rect 18800 9580 19040 9660
rect 18610 8500 18620 8760
rect 18800 7660 18980 9580
rect 12930 7180 13390 7240
rect 13430 7200 13610 7480
rect 17610 7400 17620 7660
rect 17800 7400 17810 7660
rect 18800 7580 19000 7660
rect 17620 7100 17800 7400
rect 18800 7310 18980 7580
rect 17914 6480 18046 6492
rect 12920 6250 13380 6310
rect 17910 6300 17920 6480
rect 18040 6300 18050 6480
rect 17914 6288 18046 6300
rect 16434 5142 16636 5148
rect 16434 5046 16446 5142
rect 16624 5046 16636 5142
rect 16434 5040 16636 5046
rect 14040 1340 14340 1800
rect 18190 1600 18200 2120
rect 18560 1600 18570 2120
rect 14040 -1310 14330 1340
rect 16290 580 16760 810
rect 18800 620 18980 5090
rect 18800 520 19020 620
rect 18800 490 18980 520
<< via1 >>
rect 17680 15580 17790 15780
rect 9300 14620 9800 15280
rect 9300 13900 10420 14620
rect 13000 14600 13080 14720
rect 17840 14360 18000 14480
rect 12980 14080 13060 14200
rect 13980 13980 14100 14100
rect 12520 13620 12620 13740
rect 17680 12400 17980 12580
rect 14040 9840 14180 9980
rect 18620 8500 18800 8760
rect 17620 7400 17800 7660
rect 17920 6300 18040 6480
rect 16446 5046 16624 5142
rect 18200 1600 18560 2120
<< metal2 >>
rect 13060 15780 13500 15790
rect 17680 15780 17790 15790
rect 13500 15580 17680 15780
rect 17790 15580 21200 15780
rect 17680 15570 17790 15580
rect 18880 15560 19080 15580
rect 13060 15310 13500 15320
rect 9300 15280 9800 15290
rect 13060 14730 13320 15310
rect 13000 14720 13320 14730
rect 9800 14620 10420 14630
rect 13080 14600 13320 14720
rect 13760 15040 13880 15050
rect 13000 14590 13080 14600
rect 12980 14200 13060 14210
rect 13760 14200 13880 14900
rect 20920 15000 21200 15580
rect 18500 14520 18680 14536
rect 17640 14480 19080 14520
rect 17640 14360 17840 14480
rect 18000 14360 19080 14480
rect 17640 14320 19080 14360
rect 10420 13940 11260 14140
rect 13060 14080 13880 14200
rect 13980 14160 14520 14300
rect 13980 14100 14100 14160
rect 12980 14070 13060 14080
rect 9300 13890 10420 13900
rect 13980 13932 14100 13980
rect 13980 13790 14102 13932
rect 12520 13740 12620 13750
rect 13980 13720 14100 13790
rect 12520 13610 12620 13620
rect 13040 13500 14100 13720
rect 13040 9480 13720 13500
rect 17680 12580 17980 12590
rect 17680 12390 17980 12400
rect 13260 9240 13720 9480
rect 13860 11140 14060 11150
rect 14060 10900 14234 11140
rect 13860 10180 14234 10900
rect 18880 10560 19080 14320
rect 20920 12950 21180 15000
rect 20800 12940 21300 12950
rect 20800 12460 21300 12500
rect 20800 12220 21440 12460
rect 13860 10020 14380 10180
rect 13860 9980 14234 10020
rect 13860 9840 14040 9980
rect 14180 9840 14234 9980
rect 13040 9230 13260 9240
rect 13860 8306 14234 9840
rect 16800 8760 17020 8770
rect 17660 8760 18000 10380
rect 18620 8760 18800 8770
rect 18880 8760 19080 8940
rect 17020 8500 18620 8760
rect 18800 8500 19080 8760
rect 16800 8490 17020 8500
rect 17660 8480 18000 8500
rect 18620 8490 18800 8500
rect 13860 8120 14320 8306
rect 18880 8300 19080 8500
rect 12140 7760 12340 7770
rect 13220 7760 14320 8120
rect 12340 7560 12720 7760
rect 13140 7560 14320 7760
rect 20920 7780 21440 12220
rect 21140 7700 21440 7780
rect 17620 7660 17800 7670
rect 12140 7550 12340 7560
rect 18240 7400 18520 7660
rect 17620 7390 17800 7400
rect 21360 7560 21440 7700
rect 21360 7340 23100 7560
rect 20920 7320 23100 7340
rect 12720 6920 13360 7120
rect 18360 7080 18680 7090
rect 18180 6800 18360 7080
rect 18180 6790 18680 6800
rect 17920 6480 18040 6490
rect 18180 6480 18660 6790
rect 17720 6300 17920 6480
rect 18040 6300 18660 6480
rect 17920 6290 18040 6300
rect 15840 5760 16380 6100
rect 16200 5140 16380 5760
rect 16446 5142 16624 5152
rect 16200 5046 16446 5140
rect 16200 5036 16624 5046
rect 16200 5020 16620 5036
rect 18200 2120 18560 2130
rect 18200 1590 18560 1600
rect 19160 1520 19300 6680
rect 20820 5600 21280 5610
rect 20820 4830 21280 4840
rect 20820 3340 21360 3350
rect 20720 2580 20820 2740
rect 21360 2580 21780 2740
rect 20720 2540 21780 2580
rect 22900 700 23100 7320
rect 20800 660 23100 700
rect 20800 380 20840 660
rect 21360 540 23100 660
rect 20800 370 21360 380
rect 18040 160 18200 170
rect 18040 -50 18200 -40
rect 20800 -1360 21040 370
rect 16950 -1640 17820 -1400
rect 17600 -3020 18440 -3010
rect 17600 -3830 18440 -3820
rect 20760 -4240 21060 -4230
rect 20760 -4670 21060 -4660
<< via2 >>
rect 13060 15320 13500 15780
rect 9300 14620 9800 15280
rect 9300 13900 10420 14620
rect 13760 14900 13880 15040
rect 12520 13620 12620 13740
rect 17680 12400 17980 12580
rect 13040 9240 13260 9480
rect 13860 10900 14060 11140
rect 20800 12500 21300 12940
rect 16800 8500 17020 8760
rect 12140 7560 12340 7760
rect 20920 7700 21140 7780
rect 20920 7340 21360 7700
rect 18360 6800 18680 7080
rect 18200 1600 18560 2120
rect 20820 4840 21280 5600
rect 20820 2580 21360 3340
rect 20840 380 21360 660
rect 18040 -40 18200 160
rect 17600 -3820 18440 -3020
rect 20760 -4660 21060 -4240
<< metal3 >>
rect 13050 15780 13510 15785
rect 13050 15320 13060 15780
rect 13500 15320 13510 15780
rect 13050 15315 13510 15320
rect 9290 15280 9810 15285
rect 9290 13900 9300 15280
rect 9800 14625 9810 15280
rect 13750 15040 13890 15045
rect 13750 14900 13760 15040
rect 13880 14900 17000 15040
rect 13750 14895 13890 14900
rect 9800 14620 10430 14625
rect 10420 13900 10430 14620
rect 9290 13895 10430 13900
rect 12510 13740 12630 13745
rect 12510 13620 12520 13740
rect 12620 13620 14100 13740
rect 12510 13615 12630 13620
rect 12818 13500 14100 13620
rect 11850 11840 11860 11940
rect 12060 11840 12070 11940
rect 11380 7260 11680 7440
rect 11870 1540 11880 11840
rect 12040 1540 12050 11840
rect 13860 11145 14060 13500
rect 13850 11140 14070 11145
rect 13850 10900 13860 11140
rect 14060 10900 14070 11140
rect 13850 10895 14070 10900
rect 13030 9480 13270 9485
rect 12480 9250 13040 9480
rect 12680 9240 13040 9250
rect 13260 9240 13270 9480
rect 13030 9235 13270 9240
rect 16820 8765 17000 14900
rect 17660 12940 21380 12960
rect 17660 12580 20800 12940
rect 17660 12400 17680 12580
rect 17980 12500 20800 12580
rect 21300 12500 21380 12940
rect 17980 12400 21380 12500
rect 17670 12395 17990 12400
rect 18880 11840 19080 12140
rect 16790 8760 17030 8765
rect 16790 8500 16800 8760
rect 17020 8500 17520 8760
rect 16790 8495 17030 8500
rect 20910 7780 21150 7785
rect 12130 7760 12350 7765
rect 12130 7560 12140 7760
rect 12340 7560 12350 7760
rect 12130 7555 12350 7560
rect 20910 7340 20920 7780
rect 21140 7705 21150 7780
rect 21140 7700 21370 7705
rect 21360 7340 21370 7700
rect 20910 7335 21370 7340
rect 18350 7080 18690 7085
rect 18350 6800 18360 7080
rect 18680 6800 18690 7080
rect 18350 6795 18690 6800
rect 20810 5600 21290 5605
rect 20810 4840 20820 5600
rect 21280 4840 21290 5600
rect 20810 4835 21290 4840
rect 20810 3340 21370 3345
rect 20810 2580 20820 3340
rect 21360 2580 21370 3340
rect 20810 2575 21370 2580
rect 18190 2120 18570 2125
rect 18190 1600 18200 2120
rect 18560 1600 18570 2120
rect 18190 1595 18570 1600
rect 20830 660 21370 665
rect 20830 380 20840 660
rect 21360 380 21370 660
rect 20830 375 21370 380
rect 18030 160 18210 165
rect 14900 -40 18040 160
rect 18200 -40 18210 160
rect 14900 -2994 15080 -40
rect 18030 -45 18210 -40
rect 17590 -3020 18450 -3015
rect 17590 -3820 17600 -3020
rect 18440 -3820 18450 -3020
rect 17590 -3825 18450 -3820
rect 20750 -4240 21070 -4235
rect 20750 -4660 20760 -4240
rect 21060 -4660 21070 -4240
rect 20750 -4665 21070 -4660
<< via3 >>
rect 13060 15320 13500 15780
rect 9300 14620 9800 15280
rect 9300 13900 10420 14620
rect 11860 11840 12060 11940
rect 11880 1540 12040 11840
rect 20800 12500 21300 12940
rect 20920 7700 21140 7780
rect 20920 7340 21360 7700
rect 20820 4840 21280 5600
rect 20820 2580 21360 3340
rect 18200 1600 18560 2120
rect 20840 380 21360 660
rect 17600 -3820 18440 -3020
rect 20760 -4660 21060 -4240
<< metal4 >>
rect -308 15780 21640 17576
rect -308 15564 13060 15780
rect 4720 4540 5500 15564
rect 13059 15320 13060 15564
rect 13500 15564 21640 15780
rect 13500 15320 13501 15564
rect 13059 15319 13501 15320
rect 9299 15280 9801 15281
rect 9299 13900 9300 15280
rect 9800 14800 9801 15280
rect 9800 14621 10420 14800
rect 9800 14620 10421 14621
rect 10420 13900 10421 14620
rect 9299 13899 10421 13900
rect 9620 -2880 10420 13899
rect 20802 12941 21382 15564
rect 20799 12940 21382 12941
rect 20799 12500 20800 12940
rect 21300 12500 21382 12940
rect 20799 12499 21382 12500
rect 20800 12380 21382 12499
rect 20802 12220 21382 12380
rect 11480 11940 12320 12020
rect 11480 11840 11860 11940
rect 12060 11840 12320 11940
rect 11480 1540 11880 11840
rect 12040 1540 12320 11840
rect 20800 11820 21382 12220
rect 20802 8280 21382 11820
rect 20802 7780 21400 8280
rect 20802 7340 20920 7780
rect 21140 7700 21400 7780
rect 21360 7340 21400 7700
rect 20802 7320 21400 7340
rect 20802 5600 21382 7320
rect 20802 4840 20820 5600
rect 21280 4840 21382 5600
rect 20802 3340 21382 4840
rect 20802 2580 20820 3340
rect 21360 2580 21382 3340
rect 11480 -2880 12320 1540
rect 17600 2120 18720 2340
rect 17600 1600 18200 2120
rect 18560 1600 18720 2120
rect 17600 -2880 18720 1600
rect 20802 660 21382 2580
rect 20802 538 20840 660
rect 20839 380 20840 538
rect 21360 538 21382 660
rect 21360 380 21361 538
rect 20839 379 21361 380
rect -220 -3020 23140 -2880
rect -220 -3820 17600 -3020
rect 18440 -3820 23140 -3020
rect -220 -4240 23140 -3820
rect -220 -4660 20760 -4240
rect 21060 -4660 23140 -4240
rect -220 -5900 23140 -4660
use isource_cmirror#0  isource_cmirror_2
timestamp 1654768133
transform 1 0 18900 0 1 9740
box 0 0 2044 2280
use isource_cmirror#0  isource_cmirror_3
timestamp 1654768133
transform 1 0 18900 0 1 7480
box 0 0 2044 2280
use isource_conv  isource_conv_0
timestamp 1654768133
transform 1 0 9200 0 1 -6200
box 3980 6900 13920 13860
use isource_conv_tsmal_nwell  isource_conv_tsmal_nwell_0
timestamp 1654768133
transform 1 0 12044 0 1 -1430
box 4070 6210 5960 9050
use isource_diffamp  isource_diffamp_0
timestamp 1654768133
transform 1 0 -280 0 1 16996
box 14560 -8200 18240 -5200
use isource_diffamp  isource_diffamp_1
timestamp 1654768133
transform 1 0 -280 0 1 21120
box 14560 -8200 18240 -5200
use isource_out  isource_out_0
timestamp 1654768133
transform 1 0 -4300 0 1 -13810
box 4320 8980 25514 15188
use isource_ref  isource_ref_0
timestamp 1654768133
transform 1 0 20 0 1 40
box -30 -40 13220 13420
use isource_startup  isource_startup_0
timestamp 1654768133
transform 1 0 10820 0 1 13700
box 200 0 2352 1238
use sky130_fd_pr__cap_mim_m3_1_SJ85NT  sky130_fd_pr__cap_mim_m3_1_SJ85NT_0
timestamp 1684165924
transform 1 0 7026 0 1 5280
box -2686 -6200 2686 6200
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ#0  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0
timestamp 1654768133
transform 1 0 19490 0 1 10040
box -2150 -2100 2149 2100
<< labels >>
rlabel metal1 14040 730 14330 920 1 VM3G
rlabel metal2 17660 -1630 17810 -1400 3 VM3D
rlabel metal1 16290 580 16490 800 3 VM22D
rlabel metal3 11380 7260 11680 7440 1 VM12D
rlabel metal1 13440 7380 13580 7460 1 VM12G
rlabel metal2 13720 7620 14040 8060 1 VM11D
rlabel metal2 18260 7400 18480 7660 1 VM14D
rlabel metal1 14908 12062 15034 12202 1 VM9D
rlabel metal2 17100 8540 17460 8740 1 VM8D
rlabel metal2 13280 12860 13440 13080 1 VM2D
rlabel metal3 14920 -2860 15060 -2600 1 I_ref
port 1 n
rlabel metal4 160 -5460 980 -4140 1 VN
port 2 n
rlabel metal4 -20 15880 1220 17200 1 VP
port 3 n
<< end >>
