magic
tech sky130A
magscale 1 2
timestamp 1683737876
<< error_p >>
rect -3725 890 -3667 896
rect -3533 890 -3475 896
rect -3341 890 -3283 896
rect -3149 890 -3091 896
rect -2957 890 -2899 896
rect -2765 890 -2707 896
rect -2573 890 -2515 896
rect -2381 890 -2323 896
rect -2189 890 -2131 896
rect -1997 890 -1939 896
rect -1805 890 -1747 896
rect -1613 890 -1555 896
rect -1421 890 -1363 896
rect -1229 890 -1171 896
rect -1037 890 -979 896
rect -845 890 -787 896
rect -653 890 -595 896
rect -461 890 -403 896
rect -269 890 -211 896
rect -77 890 -19 896
rect 115 890 173 896
rect 307 890 365 896
rect 499 890 557 896
rect 691 890 749 896
rect 883 890 941 896
rect 1075 890 1133 896
rect 1267 890 1325 896
rect 1459 890 1517 896
rect 1651 890 1709 896
rect 1843 890 1901 896
rect 2035 890 2093 896
rect 2227 890 2285 896
rect 2419 890 2477 896
rect 2611 890 2669 896
rect 2803 890 2861 896
rect 2995 890 3053 896
rect 3187 890 3245 896
rect 3379 890 3437 896
rect 3571 890 3629 896
rect 3763 890 3821 896
rect -3725 856 -3713 890
rect -3533 856 -3521 890
rect -3341 856 -3329 890
rect -3149 856 -3137 890
rect -2957 856 -2945 890
rect -2765 856 -2753 890
rect -2573 856 -2561 890
rect -2381 856 -2369 890
rect -2189 856 -2177 890
rect -1997 856 -1985 890
rect -1805 856 -1793 890
rect -1613 856 -1601 890
rect -1421 856 -1409 890
rect -1229 856 -1217 890
rect -1037 856 -1025 890
rect -845 856 -833 890
rect -653 856 -641 890
rect -461 856 -449 890
rect -269 856 -257 890
rect -77 856 -65 890
rect 115 856 127 890
rect 307 856 319 890
rect 499 856 511 890
rect 691 856 703 890
rect 883 856 895 890
rect 1075 856 1087 890
rect 1267 856 1279 890
rect 1459 856 1471 890
rect 1651 856 1663 890
rect 1843 856 1855 890
rect 2035 856 2047 890
rect 2227 856 2239 890
rect 2419 856 2431 890
rect 2611 856 2623 890
rect 2803 856 2815 890
rect 2995 856 3007 890
rect 3187 856 3199 890
rect 3379 856 3391 890
rect 3571 856 3583 890
rect 3763 856 3775 890
rect -3725 850 -3667 856
rect -3533 850 -3475 856
rect -3341 850 -3283 856
rect -3149 850 -3091 856
rect -2957 850 -2899 856
rect -2765 850 -2707 856
rect -2573 850 -2515 856
rect -2381 850 -2323 856
rect -2189 850 -2131 856
rect -1997 850 -1939 856
rect -1805 850 -1747 856
rect -1613 850 -1555 856
rect -1421 850 -1363 856
rect -1229 850 -1171 856
rect -1037 850 -979 856
rect -845 850 -787 856
rect -653 850 -595 856
rect -461 850 -403 856
rect -269 850 -211 856
rect -77 850 -19 856
rect 115 850 173 856
rect 307 850 365 856
rect 499 850 557 856
rect 691 850 749 856
rect 883 850 941 856
rect 1075 850 1133 856
rect 1267 850 1325 856
rect 1459 850 1517 856
rect 1651 850 1709 856
rect 1843 850 1901 856
rect 2035 850 2093 856
rect 2227 850 2285 856
rect 2419 850 2477 856
rect 2611 850 2669 856
rect 2803 850 2861 856
rect 2995 850 3053 856
rect 3187 850 3245 856
rect 3379 850 3437 856
rect 3571 850 3629 856
rect 3763 850 3821 856
rect -3821 380 -3763 386
rect -3629 380 -3571 386
rect -3437 380 -3379 386
rect -3245 380 -3187 386
rect -3053 380 -2995 386
rect -2861 380 -2803 386
rect -2669 380 -2611 386
rect -2477 380 -2419 386
rect -2285 380 -2227 386
rect -2093 380 -2035 386
rect -1901 380 -1843 386
rect -1709 380 -1651 386
rect -1517 380 -1459 386
rect -1325 380 -1267 386
rect -1133 380 -1075 386
rect -941 380 -883 386
rect -749 380 -691 386
rect -557 380 -499 386
rect -365 380 -307 386
rect -173 380 -115 386
rect 19 380 77 386
rect 211 380 269 386
rect 403 380 461 386
rect 595 380 653 386
rect 787 380 845 386
rect 979 380 1037 386
rect 1171 380 1229 386
rect 1363 380 1421 386
rect 1555 380 1613 386
rect 1747 380 1805 386
rect 1939 380 1997 386
rect 2131 380 2189 386
rect 2323 380 2381 386
rect 2515 380 2573 386
rect 2707 380 2765 386
rect 2899 380 2957 386
rect 3091 380 3149 386
rect 3283 380 3341 386
rect 3475 380 3533 386
rect 3667 380 3725 386
rect -3821 346 -3809 380
rect -3629 346 -3617 380
rect -3437 346 -3425 380
rect -3245 346 -3233 380
rect -3053 346 -3041 380
rect -2861 346 -2849 380
rect -2669 346 -2657 380
rect -2477 346 -2465 380
rect -2285 346 -2273 380
rect -2093 346 -2081 380
rect -1901 346 -1889 380
rect -1709 346 -1697 380
rect -1517 346 -1505 380
rect -1325 346 -1313 380
rect -1133 346 -1121 380
rect -941 346 -929 380
rect -749 346 -737 380
rect -557 346 -545 380
rect -365 346 -353 380
rect -173 346 -161 380
rect 19 346 31 380
rect 211 346 223 380
rect 403 346 415 380
rect 595 346 607 380
rect 787 346 799 380
rect 979 346 991 380
rect 1171 346 1183 380
rect 1363 346 1375 380
rect 1555 346 1567 380
rect 1747 346 1759 380
rect 1939 346 1951 380
rect 2131 346 2143 380
rect 2323 346 2335 380
rect 2515 346 2527 380
rect 2707 346 2719 380
rect 2899 346 2911 380
rect 3091 346 3103 380
rect 3283 346 3295 380
rect 3475 346 3487 380
rect 3667 346 3679 380
rect -3821 340 -3763 346
rect -3629 340 -3571 346
rect -3437 340 -3379 346
rect -3245 340 -3187 346
rect -3053 340 -2995 346
rect -2861 340 -2803 346
rect -2669 340 -2611 346
rect -2477 340 -2419 346
rect -2285 340 -2227 346
rect -2093 340 -2035 346
rect -1901 340 -1843 346
rect -1709 340 -1651 346
rect -1517 340 -1459 346
rect -1325 340 -1267 346
rect -1133 340 -1075 346
rect -941 340 -883 346
rect -749 340 -691 346
rect -557 340 -499 346
rect -365 340 -307 346
rect -173 340 -115 346
rect 19 340 77 346
rect 211 340 269 346
rect 403 340 461 346
rect 595 340 653 346
rect 787 340 845 346
rect 979 340 1037 346
rect 1171 340 1229 346
rect 1363 340 1421 346
rect 1555 340 1613 346
rect 1747 340 1805 346
rect 1939 340 1997 346
rect 2131 340 2189 346
rect 2323 340 2381 346
rect 2515 340 2573 346
rect 2707 340 2765 346
rect 2899 340 2957 346
rect 3091 340 3149 346
rect 3283 340 3341 346
rect 3475 340 3533 346
rect 3667 340 3725 346
rect -3821 272 -3763 278
rect -3629 272 -3571 278
rect -3437 272 -3379 278
rect -3245 272 -3187 278
rect -3053 272 -2995 278
rect -2861 272 -2803 278
rect -2669 272 -2611 278
rect -2477 272 -2419 278
rect -2285 272 -2227 278
rect -2093 272 -2035 278
rect -1901 272 -1843 278
rect -1709 272 -1651 278
rect -1517 272 -1459 278
rect -1325 272 -1267 278
rect -1133 272 -1075 278
rect -941 272 -883 278
rect -749 272 -691 278
rect -557 272 -499 278
rect -365 272 -307 278
rect -173 272 -115 278
rect 19 272 77 278
rect 211 272 269 278
rect 403 272 461 278
rect 595 272 653 278
rect 787 272 845 278
rect 979 272 1037 278
rect 1171 272 1229 278
rect 1363 272 1421 278
rect 1555 272 1613 278
rect 1747 272 1805 278
rect 1939 272 1997 278
rect 2131 272 2189 278
rect 2323 272 2381 278
rect 2515 272 2573 278
rect 2707 272 2765 278
rect 2899 272 2957 278
rect 3091 272 3149 278
rect 3283 272 3341 278
rect 3475 272 3533 278
rect 3667 272 3725 278
rect -3821 238 -3809 272
rect -3629 238 -3617 272
rect -3437 238 -3425 272
rect -3245 238 -3233 272
rect -3053 238 -3041 272
rect -2861 238 -2849 272
rect -2669 238 -2657 272
rect -2477 238 -2465 272
rect -2285 238 -2273 272
rect -2093 238 -2081 272
rect -1901 238 -1889 272
rect -1709 238 -1697 272
rect -1517 238 -1505 272
rect -1325 238 -1313 272
rect -1133 238 -1121 272
rect -941 238 -929 272
rect -749 238 -737 272
rect -557 238 -545 272
rect -365 238 -353 272
rect -173 238 -161 272
rect 19 238 31 272
rect 211 238 223 272
rect 403 238 415 272
rect 595 238 607 272
rect 787 238 799 272
rect 979 238 991 272
rect 1171 238 1183 272
rect 1363 238 1375 272
rect 1555 238 1567 272
rect 1747 238 1759 272
rect 1939 238 1951 272
rect 2131 238 2143 272
rect 2323 238 2335 272
rect 2515 238 2527 272
rect 2707 238 2719 272
rect 2899 238 2911 272
rect 3091 238 3103 272
rect 3283 238 3295 272
rect 3475 238 3487 272
rect 3667 238 3679 272
rect -3821 232 -3763 238
rect -3629 232 -3571 238
rect -3437 232 -3379 238
rect -3245 232 -3187 238
rect -3053 232 -2995 238
rect -2861 232 -2803 238
rect -2669 232 -2611 238
rect -2477 232 -2419 238
rect -2285 232 -2227 238
rect -2093 232 -2035 238
rect -1901 232 -1843 238
rect -1709 232 -1651 238
rect -1517 232 -1459 238
rect -1325 232 -1267 238
rect -1133 232 -1075 238
rect -941 232 -883 238
rect -749 232 -691 238
rect -557 232 -499 238
rect -365 232 -307 238
rect -173 232 -115 238
rect 19 232 77 238
rect 211 232 269 238
rect 403 232 461 238
rect 595 232 653 238
rect 787 232 845 238
rect 979 232 1037 238
rect 1171 232 1229 238
rect 1363 232 1421 238
rect 1555 232 1613 238
rect 1747 232 1805 238
rect 1939 232 1997 238
rect 2131 232 2189 238
rect 2323 232 2381 238
rect 2515 232 2573 238
rect 2707 232 2765 238
rect 2899 232 2957 238
rect 3091 232 3149 238
rect 3283 232 3341 238
rect 3475 232 3533 238
rect 3667 232 3725 238
rect -3725 -238 -3667 -232
rect -3533 -238 -3475 -232
rect -3341 -238 -3283 -232
rect -3149 -238 -3091 -232
rect -2957 -238 -2899 -232
rect -2765 -238 -2707 -232
rect -2573 -238 -2515 -232
rect -2381 -238 -2323 -232
rect -2189 -238 -2131 -232
rect -1997 -238 -1939 -232
rect -1805 -238 -1747 -232
rect -1613 -238 -1555 -232
rect -1421 -238 -1363 -232
rect -1229 -238 -1171 -232
rect -1037 -238 -979 -232
rect -845 -238 -787 -232
rect -653 -238 -595 -232
rect -461 -238 -403 -232
rect -269 -238 -211 -232
rect -77 -238 -19 -232
rect 115 -238 173 -232
rect 307 -238 365 -232
rect 499 -238 557 -232
rect 691 -238 749 -232
rect 883 -238 941 -232
rect 1075 -238 1133 -232
rect 1267 -238 1325 -232
rect 1459 -238 1517 -232
rect 1651 -238 1709 -232
rect 1843 -238 1901 -232
rect 2035 -238 2093 -232
rect 2227 -238 2285 -232
rect 2419 -238 2477 -232
rect 2611 -238 2669 -232
rect 2803 -238 2861 -232
rect 2995 -238 3053 -232
rect 3187 -238 3245 -232
rect 3379 -238 3437 -232
rect 3571 -238 3629 -232
rect 3763 -238 3821 -232
rect -3725 -272 -3713 -238
rect -3533 -272 -3521 -238
rect -3341 -272 -3329 -238
rect -3149 -272 -3137 -238
rect -2957 -272 -2945 -238
rect -2765 -272 -2753 -238
rect -2573 -272 -2561 -238
rect -2381 -272 -2369 -238
rect -2189 -272 -2177 -238
rect -1997 -272 -1985 -238
rect -1805 -272 -1793 -238
rect -1613 -272 -1601 -238
rect -1421 -272 -1409 -238
rect -1229 -272 -1217 -238
rect -1037 -272 -1025 -238
rect -845 -272 -833 -238
rect -653 -272 -641 -238
rect -461 -272 -449 -238
rect -269 -272 -257 -238
rect -77 -272 -65 -238
rect 115 -272 127 -238
rect 307 -272 319 -238
rect 499 -272 511 -238
rect 691 -272 703 -238
rect 883 -272 895 -238
rect 1075 -272 1087 -238
rect 1267 -272 1279 -238
rect 1459 -272 1471 -238
rect 1651 -272 1663 -238
rect 1843 -272 1855 -238
rect 2035 -272 2047 -238
rect 2227 -272 2239 -238
rect 2419 -272 2431 -238
rect 2611 -272 2623 -238
rect 2803 -272 2815 -238
rect 2995 -272 3007 -238
rect 3187 -272 3199 -238
rect 3379 -272 3391 -238
rect 3571 -272 3583 -238
rect 3763 -272 3775 -238
rect -3725 -278 -3667 -272
rect -3533 -278 -3475 -272
rect -3341 -278 -3283 -272
rect -3149 -278 -3091 -272
rect -2957 -278 -2899 -272
rect -2765 -278 -2707 -272
rect -2573 -278 -2515 -272
rect -2381 -278 -2323 -272
rect -2189 -278 -2131 -272
rect -1997 -278 -1939 -272
rect -1805 -278 -1747 -272
rect -1613 -278 -1555 -272
rect -1421 -278 -1363 -272
rect -1229 -278 -1171 -272
rect -1037 -278 -979 -272
rect -845 -278 -787 -272
rect -653 -278 -595 -272
rect -461 -278 -403 -272
rect -269 -278 -211 -272
rect -77 -278 -19 -272
rect 115 -278 173 -272
rect 307 -278 365 -272
rect 499 -278 557 -272
rect 691 -278 749 -272
rect 883 -278 941 -272
rect 1075 -278 1133 -272
rect 1267 -278 1325 -272
rect 1459 -278 1517 -272
rect 1651 -278 1709 -272
rect 1843 -278 1901 -272
rect 2035 -278 2093 -272
rect 2227 -278 2285 -272
rect 2419 -278 2477 -272
rect 2611 -278 2669 -272
rect 2803 -278 2861 -272
rect 2995 -278 3053 -272
rect 3187 -278 3245 -272
rect 3379 -278 3437 -272
rect 3571 -278 3629 -272
rect 3763 -278 3821 -272
rect -3725 -346 -3667 -340
rect -3533 -346 -3475 -340
rect -3341 -346 -3283 -340
rect -3149 -346 -3091 -340
rect -2957 -346 -2899 -340
rect -2765 -346 -2707 -340
rect -2573 -346 -2515 -340
rect -2381 -346 -2323 -340
rect -2189 -346 -2131 -340
rect -1997 -346 -1939 -340
rect -1805 -346 -1747 -340
rect -1613 -346 -1555 -340
rect -1421 -346 -1363 -340
rect -1229 -346 -1171 -340
rect -1037 -346 -979 -340
rect -845 -346 -787 -340
rect -653 -346 -595 -340
rect -461 -346 -403 -340
rect -269 -346 -211 -340
rect -77 -346 -19 -340
rect 115 -346 173 -340
rect 307 -346 365 -340
rect 499 -346 557 -340
rect 691 -346 749 -340
rect 883 -346 941 -340
rect 1075 -346 1133 -340
rect 1267 -346 1325 -340
rect 1459 -346 1517 -340
rect 1651 -346 1709 -340
rect 1843 -346 1901 -340
rect 2035 -346 2093 -340
rect 2227 -346 2285 -340
rect 2419 -346 2477 -340
rect 2611 -346 2669 -340
rect 2803 -346 2861 -340
rect 2995 -346 3053 -340
rect 3187 -346 3245 -340
rect 3379 -346 3437 -340
rect 3571 -346 3629 -340
rect 3763 -346 3821 -340
rect -3725 -380 -3713 -346
rect -3533 -380 -3521 -346
rect -3341 -380 -3329 -346
rect -3149 -380 -3137 -346
rect -2957 -380 -2945 -346
rect -2765 -380 -2753 -346
rect -2573 -380 -2561 -346
rect -2381 -380 -2369 -346
rect -2189 -380 -2177 -346
rect -1997 -380 -1985 -346
rect -1805 -380 -1793 -346
rect -1613 -380 -1601 -346
rect -1421 -380 -1409 -346
rect -1229 -380 -1217 -346
rect -1037 -380 -1025 -346
rect -845 -380 -833 -346
rect -653 -380 -641 -346
rect -461 -380 -449 -346
rect -269 -380 -257 -346
rect -77 -380 -65 -346
rect 115 -380 127 -346
rect 307 -380 319 -346
rect 499 -380 511 -346
rect 691 -380 703 -346
rect 883 -380 895 -346
rect 1075 -380 1087 -346
rect 1267 -380 1279 -346
rect 1459 -380 1471 -346
rect 1651 -380 1663 -346
rect 1843 -380 1855 -346
rect 2035 -380 2047 -346
rect 2227 -380 2239 -346
rect 2419 -380 2431 -346
rect 2611 -380 2623 -346
rect 2803 -380 2815 -346
rect 2995 -380 3007 -346
rect 3187 -380 3199 -346
rect 3379 -380 3391 -346
rect 3571 -380 3583 -346
rect 3763 -380 3775 -346
rect -3725 -386 -3667 -380
rect -3533 -386 -3475 -380
rect -3341 -386 -3283 -380
rect -3149 -386 -3091 -380
rect -2957 -386 -2899 -380
rect -2765 -386 -2707 -380
rect -2573 -386 -2515 -380
rect -2381 -386 -2323 -380
rect -2189 -386 -2131 -380
rect -1997 -386 -1939 -380
rect -1805 -386 -1747 -380
rect -1613 -386 -1555 -380
rect -1421 -386 -1363 -380
rect -1229 -386 -1171 -380
rect -1037 -386 -979 -380
rect -845 -386 -787 -380
rect -653 -386 -595 -380
rect -461 -386 -403 -380
rect -269 -386 -211 -380
rect -77 -386 -19 -380
rect 115 -386 173 -380
rect 307 -386 365 -380
rect 499 -386 557 -380
rect 691 -386 749 -380
rect 883 -386 941 -380
rect 1075 -386 1133 -380
rect 1267 -386 1325 -380
rect 1459 -386 1517 -380
rect 1651 -386 1709 -380
rect 1843 -386 1901 -380
rect 2035 -386 2093 -380
rect 2227 -386 2285 -380
rect 2419 -386 2477 -380
rect 2611 -386 2669 -380
rect 2803 -386 2861 -380
rect 2995 -386 3053 -380
rect 3187 -386 3245 -380
rect 3379 -386 3437 -380
rect 3571 -386 3629 -380
rect 3763 -386 3821 -380
rect -3821 -856 -3763 -850
rect -3629 -856 -3571 -850
rect -3437 -856 -3379 -850
rect -3245 -856 -3187 -850
rect -3053 -856 -2995 -850
rect -2861 -856 -2803 -850
rect -2669 -856 -2611 -850
rect -2477 -856 -2419 -850
rect -2285 -856 -2227 -850
rect -2093 -856 -2035 -850
rect -1901 -856 -1843 -850
rect -1709 -856 -1651 -850
rect -1517 -856 -1459 -850
rect -1325 -856 -1267 -850
rect -1133 -856 -1075 -850
rect -941 -856 -883 -850
rect -749 -856 -691 -850
rect -557 -856 -499 -850
rect -365 -856 -307 -850
rect -173 -856 -115 -850
rect 19 -856 77 -850
rect 211 -856 269 -850
rect 403 -856 461 -850
rect 595 -856 653 -850
rect 787 -856 845 -850
rect 979 -856 1037 -850
rect 1171 -856 1229 -850
rect 1363 -856 1421 -850
rect 1555 -856 1613 -850
rect 1747 -856 1805 -850
rect 1939 -856 1997 -850
rect 2131 -856 2189 -850
rect 2323 -856 2381 -850
rect 2515 -856 2573 -850
rect 2707 -856 2765 -850
rect 2899 -856 2957 -850
rect 3091 -856 3149 -850
rect 3283 -856 3341 -850
rect 3475 -856 3533 -850
rect 3667 -856 3725 -850
rect -3821 -890 -3809 -856
rect -3629 -890 -3617 -856
rect -3437 -890 -3425 -856
rect -3245 -890 -3233 -856
rect -3053 -890 -3041 -856
rect -2861 -890 -2849 -856
rect -2669 -890 -2657 -856
rect -2477 -890 -2465 -856
rect -2285 -890 -2273 -856
rect -2093 -890 -2081 -856
rect -1901 -890 -1889 -856
rect -1709 -890 -1697 -856
rect -1517 -890 -1505 -856
rect -1325 -890 -1313 -856
rect -1133 -890 -1121 -856
rect -941 -890 -929 -856
rect -749 -890 -737 -856
rect -557 -890 -545 -856
rect -365 -890 -353 -856
rect -173 -890 -161 -856
rect 19 -890 31 -856
rect 211 -890 223 -856
rect 403 -890 415 -856
rect 595 -890 607 -856
rect 787 -890 799 -856
rect 979 -890 991 -856
rect 1171 -890 1183 -856
rect 1363 -890 1375 -856
rect 1555 -890 1567 -856
rect 1747 -890 1759 -856
rect 1939 -890 1951 -856
rect 2131 -890 2143 -856
rect 2323 -890 2335 -856
rect 2515 -890 2527 -856
rect 2707 -890 2719 -856
rect 2899 -890 2911 -856
rect 3091 -890 3103 -856
rect 3283 -890 3295 -856
rect 3475 -890 3487 -856
rect 3667 -890 3679 -856
rect -3821 -896 -3763 -890
rect -3629 -896 -3571 -890
rect -3437 -896 -3379 -890
rect -3245 -896 -3187 -890
rect -3053 -896 -2995 -890
rect -2861 -896 -2803 -890
rect -2669 -896 -2611 -890
rect -2477 -896 -2419 -890
rect -2285 -896 -2227 -890
rect -2093 -896 -2035 -890
rect -1901 -896 -1843 -890
rect -1709 -896 -1651 -890
rect -1517 -896 -1459 -890
rect -1325 -896 -1267 -890
rect -1133 -896 -1075 -890
rect -941 -896 -883 -890
rect -749 -896 -691 -890
rect -557 -896 -499 -890
rect -365 -896 -307 -890
rect -173 -896 -115 -890
rect 19 -896 77 -890
rect 211 -896 269 -890
rect 403 -896 461 -890
rect 595 -896 653 -890
rect 787 -896 845 -890
rect 979 -896 1037 -890
rect 1171 -896 1229 -890
rect 1363 -896 1421 -890
rect 1555 -896 1613 -890
rect 1747 -896 1805 -890
rect 1939 -896 1997 -890
rect 2131 -896 2189 -890
rect 2323 -896 2381 -890
rect 2515 -896 2573 -890
rect 2707 -896 2765 -890
rect 2899 -896 2957 -890
rect 3091 -896 3149 -890
rect 3283 -896 3341 -890
rect 3475 -896 3533 -890
rect 3667 -896 3725 -890
<< pwell >>
rect -4007 -1028 4007 1028
<< nmoslvt >>
rect -3807 418 -3777 818
rect -3711 418 -3681 818
rect -3615 418 -3585 818
rect -3519 418 -3489 818
rect -3423 418 -3393 818
rect -3327 418 -3297 818
rect -3231 418 -3201 818
rect -3135 418 -3105 818
rect -3039 418 -3009 818
rect -2943 418 -2913 818
rect -2847 418 -2817 818
rect -2751 418 -2721 818
rect -2655 418 -2625 818
rect -2559 418 -2529 818
rect -2463 418 -2433 818
rect -2367 418 -2337 818
rect -2271 418 -2241 818
rect -2175 418 -2145 818
rect -2079 418 -2049 818
rect -1983 418 -1953 818
rect -1887 418 -1857 818
rect -1791 418 -1761 818
rect -1695 418 -1665 818
rect -1599 418 -1569 818
rect -1503 418 -1473 818
rect -1407 418 -1377 818
rect -1311 418 -1281 818
rect -1215 418 -1185 818
rect -1119 418 -1089 818
rect -1023 418 -993 818
rect -927 418 -897 818
rect -831 418 -801 818
rect -735 418 -705 818
rect -639 418 -609 818
rect -543 418 -513 818
rect -447 418 -417 818
rect -351 418 -321 818
rect -255 418 -225 818
rect -159 418 -129 818
rect -63 418 -33 818
rect 33 418 63 818
rect 129 418 159 818
rect 225 418 255 818
rect 321 418 351 818
rect 417 418 447 818
rect 513 418 543 818
rect 609 418 639 818
rect 705 418 735 818
rect 801 418 831 818
rect 897 418 927 818
rect 993 418 1023 818
rect 1089 418 1119 818
rect 1185 418 1215 818
rect 1281 418 1311 818
rect 1377 418 1407 818
rect 1473 418 1503 818
rect 1569 418 1599 818
rect 1665 418 1695 818
rect 1761 418 1791 818
rect 1857 418 1887 818
rect 1953 418 1983 818
rect 2049 418 2079 818
rect 2145 418 2175 818
rect 2241 418 2271 818
rect 2337 418 2367 818
rect 2433 418 2463 818
rect 2529 418 2559 818
rect 2625 418 2655 818
rect 2721 418 2751 818
rect 2817 418 2847 818
rect 2913 418 2943 818
rect 3009 418 3039 818
rect 3105 418 3135 818
rect 3201 418 3231 818
rect 3297 418 3327 818
rect 3393 418 3423 818
rect 3489 418 3519 818
rect 3585 418 3615 818
rect 3681 418 3711 818
rect 3777 418 3807 818
rect -3807 -200 -3777 200
rect -3711 -200 -3681 200
rect -3615 -200 -3585 200
rect -3519 -200 -3489 200
rect -3423 -200 -3393 200
rect -3327 -200 -3297 200
rect -3231 -200 -3201 200
rect -3135 -200 -3105 200
rect -3039 -200 -3009 200
rect -2943 -200 -2913 200
rect -2847 -200 -2817 200
rect -2751 -200 -2721 200
rect -2655 -200 -2625 200
rect -2559 -200 -2529 200
rect -2463 -200 -2433 200
rect -2367 -200 -2337 200
rect -2271 -200 -2241 200
rect -2175 -200 -2145 200
rect -2079 -200 -2049 200
rect -1983 -200 -1953 200
rect -1887 -200 -1857 200
rect -1791 -200 -1761 200
rect -1695 -200 -1665 200
rect -1599 -200 -1569 200
rect -1503 -200 -1473 200
rect -1407 -200 -1377 200
rect -1311 -200 -1281 200
rect -1215 -200 -1185 200
rect -1119 -200 -1089 200
rect -1023 -200 -993 200
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
rect 993 -200 1023 200
rect 1089 -200 1119 200
rect 1185 -200 1215 200
rect 1281 -200 1311 200
rect 1377 -200 1407 200
rect 1473 -200 1503 200
rect 1569 -200 1599 200
rect 1665 -200 1695 200
rect 1761 -200 1791 200
rect 1857 -200 1887 200
rect 1953 -200 1983 200
rect 2049 -200 2079 200
rect 2145 -200 2175 200
rect 2241 -200 2271 200
rect 2337 -200 2367 200
rect 2433 -200 2463 200
rect 2529 -200 2559 200
rect 2625 -200 2655 200
rect 2721 -200 2751 200
rect 2817 -200 2847 200
rect 2913 -200 2943 200
rect 3009 -200 3039 200
rect 3105 -200 3135 200
rect 3201 -200 3231 200
rect 3297 -200 3327 200
rect 3393 -200 3423 200
rect 3489 -200 3519 200
rect 3585 -200 3615 200
rect 3681 -200 3711 200
rect 3777 -200 3807 200
rect -3807 -818 -3777 -418
rect -3711 -818 -3681 -418
rect -3615 -818 -3585 -418
rect -3519 -818 -3489 -418
rect -3423 -818 -3393 -418
rect -3327 -818 -3297 -418
rect -3231 -818 -3201 -418
rect -3135 -818 -3105 -418
rect -3039 -818 -3009 -418
rect -2943 -818 -2913 -418
rect -2847 -818 -2817 -418
rect -2751 -818 -2721 -418
rect -2655 -818 -2625 -418
rect -2559 -818 -2529 -418
rect -2463 -818 -2433 -418
rect -2367 -818 -2337 -418
rect -2271 -818 -2241 -418
rect -2175 -818 -2145 -418
rect -2079 -818 -2049 -418
rect -1983 -818 -1953 -418
rect -1887 -818 -1857 -418
rect -1791 -818 -1761 -418
rect -1695 -818 -1665 -418
rect -1599 -818 -1569 -418
rect -1503 -818 -1473 -418
rect -1407 -818 -1377 -418
rect -1311 -818 -1281 -418
rect -1215 -818 -1185 -418
rect -1119 -818 -1089 -418
rect -1023 -818 -993 -418
rect -927 -818 -897 -418
rect -831 -818 -801 -418
rect -735 -818 -705 -418
rect -639 -818 -609 -418
rect -543 -818 -513 -418
rect -447 -818 -417 -418
rect -351 -818 -321 -418
rect -255 -818 -225 -418
rect -159 -818 -129 -418
rect -63 -818 -33 -418
rect 33 -818 63 -418
rect 129 -818 159 -418
rect 225 -818 255 -418
rect 321 -818 351 -418
rect 417 -818 447 -418
rect 513 -818 543 -418
rect 609 -818 639 -418
rect 705 -818 735 -418
rect 801 -818 831 -418
rect 897 -818 927 -418
rect 993 -818 1023 -418
rect 1089 -818 1119 -418
rect 1185 -818 1215 -418
rect 1281 -818 1311 -418
rect 1377 -818 1407 -418
rect 1473 -818 1503 -418
rect 1569 -818 1599 -418
rect 1665 -818 1695 -418
rect 1761 -818 1791 -418
rect 1857 -818 1887 -418
rect 1953 -818 1983 -418
rect 2049 -818 2079 -418
rect 2145 -818 2175 -418
rect 2241 -818 2271 -418
rect 2337 -818 2367 -418
rect 2433 -818 2463 -418
rect 2529 -818 2559 -418
rect 2625 -818 2655 -418
rect 2721 -818 2751 -418
rect 2817 -818 2847 -418
rect 2913 -818 2943 -418
rect 3009 -818 3039 -418
rect 3105 -818 3135 -418
rect 3201 -818 3231 -418
rect 3297 -818 3327 -418
rect 3393 -818 3423 -418
rect 3489 -818 3519 -418
rect 3585 -818 3615 -418
rect 3681 -818 3711 -418
rect 3777 -818 3807 -418
<< ndiff >>
rect -3869 806 -3807 818
rect -3869 430 -3857 806
rect -3823 430 -3807 806
rect -3869 418 -3807 430
rect -3777 806 -3711 818
rect -3777 430 -3761 806
rect -3727 430 -3711 806
rect -3777 418 -3711 430
rect -3681 806 -3615 818
rect -3681 430 -3665 806
rect -3631 430 -3615 806
rect -3681 418 -3615 430
rect -3585 806 -3519 818
rect -3585 430 -3569 806
rect -3535 430 -3519 806
rect -3585 418 -3519 430
rect -3489 806 -3423 818
rect -3489 430 -3473 806
rect -3439 430 -3423 806
rect -3489 418 -3423 430
rect -3393 806 -3327 818
rect -3393 430 -3377 806
rect -3343 430 -3327 806
rect -3393 418 -3327 430
rect -3297 806 -3231 818
rect -3297 430 -3281 806
rect -3247 430 -3231 806
rect -3297 418 -3231 430
rect -3201 806 -3135 818
rect -3201 430 -3185 806
rect -3151 430 -3135 806
rect -3201 418 -3135 430
rect -3105 806 -3039 818
rect -3105 430 -3089 806
rect -3055 430 -3039 806
rect -3105 418 -3039 430
rect -3009 806 -2943 818
rect -3009 430 -2993 806
rect -2959 430 -2943 806
rect -3009 418 -2943 430
rect -2913 806 -2847 818
rect -2913 430 -2897 806
rect -2863 430 -2847 806
rect -2913 418 -2847 430
rect -2817 806 -2751 818
rect -2817 430 -2801 806
rect -2767 430 -2751 806
rect -2817 418 -2751 430
rect -2721 806 -2655 818
rect -2721 430 -2705 806
rect -2671 430 -2655 806
rect -2721 418 -2655 430
rect -2625 806 -2559 818
rect -2625 430 -2609 806
rect -2575 430 -2559 806
rect -2625 418 -2559 430
rect -2529 806 -2463 818
rect -2529 430 -2513 806
rect -2479 430 -2463 806
rect -2529 418 -2463 430
rect -2433 806 -2367 818
rect -2433 430 -2417 806
rect -2383 430 -2367 806
rect -2433 418 -2367 430
rect -2337 806 -2271 818
rect -2337 430 -2321 806
rect -2287 430 -2271 806
rect -2337 418 -2271 430
rect -2241 806 -2175 818
rect -2241 430 -2225 806
rect -2191 430 -2175 806
rect -2241 418 -2175 430
rect -2145 806 -2079 818
rect -2145 430 -2129 806
rect -2095 430 -2079 806
rect -2145 418 -2079 430
rect -2049 806 -1983 818
rect -2049 430 -2033 806
rect -1999 430 -1983 806
rect -2049 418 -1983 430
rect -1953 806 -1887 818
rect -1953 430 -1937 806
rect -1903 430 -1887 806
rect -1953 418 -1887 430
rect -1857 806 -1791 818
rect -1857 430 -1841 806
rect -1807 430 -1791 806
rect -1857 418 -1791 430
rect -1761 806 -1695 818
rect -1761 430 -1745 806
rect -1711 430 -1695 806
rect -1761 418 -1695 430
rect -1665 806 -1599 818
rect -1665 430 -1649 806
rect -1615 430 -1599 806
rect -1665 418 -1599 430
rect -1569 806 -1503 818
rect -1569 430 -1553 806
rect -1519 430 -1503 806
rect -1569 418 -1503 430
rect -1473 806 -1407 818
rect -1473 430 -1457 806
rect -1423 430 -1407 806
rect -1473 418 -1407 430
rect -1377 806 -1311 818
rect -1377 430 -1361 806
rect -1327 430 -1311 806
rect -1377 418 -1311 430
rect -1281 806 -1215 818
rect -1281 430 -1265 806
rect -1231 430 -1215 806
rect -1281 418 -1215 430
rect -1185 806 -1119 818
rect -1185 430 -1169 806
rect -1135 430 -1119 806
rect -1185 418 -1119 430
rect -1089 806 -1023 818
rect -1089 430 -1073 806
rect -1039 430 -1023 806
rect -1089 418 -1023 430
rect -993 806 -927 818
rect -993 430 -977 806
rect -943 430 -927 806
rect -993 418 -927 430
rect -897 806 -831 818
rect -897 430 -881 806
rect -847 430 -831 806
rect -897 418 -831 430
rect -801 806 -735 818
rect -801 430 -785 806
rect -751 430 -735 806
rect -801 418 -735 430
rect -705 806 -639 818
rect -705 430 -689 806
rect -655 430 -639 806
rect -705 418 -639 430
rect -609 806 -543 818
rect -609 430 -593 806
rect -559 430 -543 806
rect -609 418 -543 430
rect -513 806 -447 818
rect -513 430 -497 806
rect -463 430 -447 806
rect -513 418 -447 430
rect -417 806 -351 818
rect -417 430 -401 806
rect -367 430 -351 806
rect -417 418 -351 430
rect -321 806 -255 818
rect -321 430 -305 806
rect -271 430 -255 806
rect -321 418 -255 430
rect -225 806 -159 818
rect -225 430 -209 806
rect -175 430 -159 806
rect -225 418 -159 430
rect -129 806 -63 818
rect -129 430 -113 806
rect -79 430 -63 806
rect -129 418 -63 430
rect -33 806 33 818
rect -33 430 -17 806
rect 17 430 33 806
rect -33 418 33 430
rect 63 806 129 818
rect 63 430 79 806
rect 113 430 129 806
rect 63 418 129 430
rect 159 806 225 818
rect 159 430 175 806
rect 209 430 225 806
rect 159 418 225 430
rect 255 806 321 818
rect 255 430 271 806
rect 305 430 321 806
rect 255 418 321 430
rect 351 806 417 818
rect 351 430 367 806
rect 401 430 417 806
rect 351 418 417 430
rect 447 806 513 818
rect 447 430 463 806
rect 497 430 513 806
rect 447 418 513 430
rect 543 806 609 818
rect 543 430 559 806
rect 593 430 609 806
rect 543 418 609 430
rect 639 806 705 818
rect 639 430 655 806
rect 689 430 705 806
rect 639 418 705 430
rect 735 806 801 818
rect 735 430 751 806
rect 785 430 801 806
rect 735 418 801 430
rect 831 806 897 818
rect 831 430 847 806
rect 881 430 897 806
rect 831 418 897 430
rect 927 806 993 818
rect 927 430 943 806
rect 977 430 993 806
rect 927 418 993 430
rect 1023 806 1089 818
rect 1023 430 1039 806
rect 1073 430 1089 806
rect 1023 418 1089 430
rect 1119 806 1185 818
rect 1119 430 1135 806
rect 1169 430 1185 806
rect 1119 418 1185 430
rect 1215 806 1281 818
rect 1215 430 1231 806
rect 1265 430 1281 806
rect 1215 418 1281 430
rect 1311 806 1377 818
rect 1311 430 1327 806
rect 1361 430 1377 806
rect 1311 418 1377 430
rect 1407 806 1473 818
rect 1407 430 1423 806
rect 1457 430 1473 806
rect 1407 418 1473 430
rect 1503 806 1569 818
rect 1503 430 1519 806
rect 1553 430 1569 806
rect 1503 418 1569 430
rect 1599 806 1665 818
rect 1599 430 1615 806
rect 1649 430 1665 806
rect 1599 418 1665 430
rect 1695 806 1761 818
rect 1695 430 1711 806
rect 1745 430 1761 806
rect 1695 418 1761 430
rect 1791 806 1857 818
rect 1791 430 1807 806
rect 1841 430 1857 806
rect 1791 418 1857 430
rect 1887 806 1953 818
rect 1887 430 1903 806
rect 1937 430 1953 806
rect 1887 418 1953 430
rect 1983 806 2049 818
rect 1983 430 1999 806
rect 2033 430 2049 806
rect 1983 418 2049 430
rect 2079 806 2145 818
rect 2079 430 2095 806
rect 2129 430 2145 806
rect 2079 418 2145 430
rect 2175 806 2241 818
rect 2175 430 2191 806
rect 2225 430 2241 806
rect 2175 418 2241 430
rect 2271 806 2337 818
rect 2271 430 2287 806
rect 2321 430 2337 806
rect 2271 418 2337 430
rect 2367 806 2433 818
rect 2367 430 2383 806
rect 2417 430 2433 806
rect 2367 418 2433 430
rect 2463 806 2529 818
rect 2463 430 2479 806
rect 2513 430 2529 806
rect 2463 418 2529 430
rect 2559 806 2625 818
rect 2559 430 2575 806
rect 2609 430 2625 806
rect 2559 418 2625 430
rect 2655 806 2721 818
rect 2655 430 2671 806
rect 2705 430 2721 806
rect 2655 418 2721 430
rect 2751 806 2817 818
rect 2751 430 2767 806
rect 2801 430 2817 806
rect 2751 418 2817 430
rect 2847 806 2913 818
rect 2847 430 2863 806
rect 2897 430 2913 806
rect 2847 418 2913 430
rect 2943 806 3009 818
rect 2943 430 2959 806
rect 2993 430 3009 806
rect 2943 418 3009 430
rect 3039 806 3105 818
rect 3039 430 3055 806
rect 3089 430 3105 806
rect 3039 418 3105 430
rect 3135 806 3201 818
rect 3135 430 3151 806
rect 3185 430 3201 806
rect 3135 418 3201 430
rect 3231 806 3297 818
rect 3231 430 3247 806
rect 3281 430 3297 806
rect 3231 418 3297 430
rect 3327 806 3393 818
rect 3327 430 3343 806
rect 3377 430 3393 806
rect 3327 418 3393 430
rect 3423 806 3489 818
rect 3423 430 3439 806
rect 3473 430 3489 806
rect 3423 418 3489 430
rect 3519 806 3585 818
rect 3519 430 3535 806
rect 3569 430 3585 806
rect 3519 418 3585 430
rect 3615 806 3681 818
rect 3615 430 3631 806
rect 3665 430 3681 806
rect 3615 418 3681 430
rect 3711 806 3777 818
rect 3711 430 3727 806
rect 3761 430 3777 806
rect 3711 418 3777 430
rect 3807 806 3869 818
rect 3807 430 3823 806
rect 3857 430 3869 806
rect 3807 418 3869 430
rect -3869 188 -3807 200
rect -3869 -188 -3857 188
rect -3823 -188 -3807 188
rect -3869 -200 -3807 -188
rect -3777 188 -3711 200
rect -3777 -188 -3761 188
rect -3727 -188 -3711 188
rect -3777 -200 -3711 -188
rect -3681 188 -3615 200
rect -3681 -188 -3665 188
rect -3631 -188 -3615 188
rect -3681 -200 -3615 -188
rect -3585 188 -3519 200
rect -3585 -188 -3569 188
rect -3535 -188 -3519 188
rect -3585 -200 -3519 -188
rect -3489 188 -3423 200
rect -3489 -188 -3473 188
rect -3439 -188 -3423 188
rect -3489 -200 -3423 -188
rect -3393 188 -3327 200
rect -3393 -188 -3377 188
rect -3343 -188 -3327 188
rect -3393 -200 -3327 -188
rect -3297 188 -3231 200
rect -3297 -188 -3281 188
rect -3247 -188 -3231 188
rect -3297 -200 -3231 -188
rect -3201 188 -3135 200
rect -3201 -188 -3185 188
rect -3151 -188 -3135 188
rect -3201 -200 -3135 -188
rect -3105 188 -3039 200
rect -3105 -188 -3089 188
rect -3055 -188 -3039 188
rect -3105 -200 -3039 -188
rect -3009 188 -2943 200
rect -3009 -188 -2993 188
rect -2959 -188 -2943 188
rect -3009 -200 -2943 -188
rect -2913 188 -2847 200
rect -2913 -188 -2897 188
rect -2863 -188 -2847 188
rect -2913 -200 -2847 -188
rect -2817 188 -2751 200
rect -2817 -188 -2801 188
rect -2767 -188 -2751 188
rect -2817 -200 -2751 -188
rect -2721 188 -2655 200
rect -2721 -188 -2705 188
rect -2671 -188 -2655 188
rect -2721 -200 -2655 -188
rect -2625 188 -2559 200
rect -2625 -188 -2609 188
rect -2575 -188 -2559 188
rect -2625 -200 -2559 -188
rect -2529 188 -2463 200
rect -2529 -188 -2513 188
rect -2479 -188 -2463 188
rect -2529 -200 -2463 -188
rect -2433 188 -2367 200
rect -2433 -188 -2417 188
rect -2383 -188 -2367 188
rect -2433 -200 -2367 -188
rect -2337 188 -2271 200
rect -2337 -188 -2321 188
rect -2287 -188 -2271 188
rect -2337 -200 -2271 -188
rect -2241 188 -2175 200
rect -2241 -188 -2225 188
rect -2191 -188 -2175 188
rect -2241 -200 -2175 -188
rect -2145 188 -2079 200
rect -2145 -188 -2129 188
rect -2095 -188 -2079 188
rect -2145 -200 -2079 -188
rect -2049 188 -1983 200
rect -2049 -188 -2033 188
rect -1999 -188 -1983 188
rect -2049 -200 -1983 -188
rect -1953 188 -1887 200
rect -1953 -188 -1937 188
rect -1903 -188 -1887 188
rect -1953 -200 -1887 -188
rect -1857 188 -1791 200
rect -1857 -188 -1841 188
rect -1807 -188 -1791 188
rect -1857 -200 -1791 -188
rect -1761 188 -1695 200
rect -1761 -188 -1745 188
rect -1711 -188 -1695 188
rect -1761 -200 -1695 -188
rect -1665 188 -1599 200
rect -1665 -188 -1649 188
rect -1615 -188 -1599 188
rect -1665 -200 -1599 -188
rect -1569 188 -1503 200
rect -1569 -188 -1553 188
rect -1519 -188 -1503 188
rect -1569 -200 -1503 -188
rect -1473 188 -1407 200
rect -1473 -188 -1457 188
rect -1423 -188 -1407 188
rect -1473 -200 -1407 -188
rect -1377 188 -1311 200
rect -1377 -188 -1361 188
rect -1327 -188 -1311 188
rect -1377 -200 -1311 -188
rect -1281 188 -1215 200
rect -1281 -188 -1265 188
rect -1231 -188 -1215 188
rect -1281 -200 -1215 -188
rect -1185 188 -1119 200
rect -1185 -188 -1169 188
rect -1135 -188 -1119 188
rect -1185 -200 -1119 -188
rect -1089 188 -1023 200
rect -1089 -188 -1073 188
rect -1039 -188 -1023 188
rect -1089 -200 -1023 -188
rect -993 188 -927 200
rect -993 -188 -977 188
rect -943 -188 -927 188
rect -993 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 993 200
rect 927 -188 943 188
rect 977 -188 993 188
rect 927 -200 993 -188
rect 1023 188 1089 200
rect 1023 -188 1039 188
rect 1073 -188 1089 188
rect 1023 -200 1089 -188
rect 1119 188 1185 200
rect 1119 -188 1135 188
rect 1169 -188 1185 188
rect 1119 -200 1185 -188
rect 1215 188 1281 200
rect 1215 -188 1231 188
rect 1265 -188 1281 188
rect 1215 -200 1281 -188
rect 1311 188 1377 200
rect 1311 -188 1327 188
rect 1361 -188 1377 188
rect 1311 -200 1377 -188
rect 1407 188 1473 200
rect 1407 -188 1423 188
rect 1457 -188 1473 188
rect 1407 -200 1473 -188
rect 1503 188 1569 200
rect 1503 -188 1519 188
rect 1553 -188 1569 188
rect 1503 -200 1569 -188
rect 1599 188 1665 200
rect 1599 -188 1615 188
rect 1649 -188 1665 188
rect 1599 -200 1665 -188
rect 1695 188 1761 200
rect 1695 -188 1711 188
rect 1745 -188 1761 188
rect 1695 -200 1761 -188
rect 1791 188 1857 200
rect 1791 -188 1807 188
rect 1841 -188 1857 188
rect 1791 -200 1857 -188
rect 1887 188 1953 200
rect 1887 -188 1903 188
rect 1937 -188 1953 188
rect 1887 -200 1953 -188
rect 1983 188 2049 200
rect 1983 -188 1999 188
rect 2033 -188 2049 188
rect 1983 -200 2049 -188
rect 2079 188 2145 200
rect 2079 -188 2095 188
rect 2129 -188 2145 188
rect 2079 -200 2145 -188
rect 2175 188 2241 200
rect 2175 -188 2191 188
rect 2225 -188 2241 188
rect 2175 -200 2241 -188
rect 2271 188 2337 200
rect 2271 -188 2287 188
rect 2321 -188 2337 188
rect 2271 -200 2337 -188
rect 2367 188 2433 200
rect 2367 -188 2383 188
rect 2417 -188 2433 188
rect 2367 -200 2433 -188
rect 2463 188 2529 200
rect 2463 -188 2479 188
rect 2513 -188 2529 188
rect 2463 -200 2529 -188
rect 2559 188 2625 200
rect 2559 -188 2575 188
rect 2609 -188 2625 188
rect 2559 -200 2625 -188
rect 2655 188 2721 200
rect 2655 -188 2671 188
rect 2705 -188 2721 188
rect 2655 -200 2721 -188
rect 2751 188 2817 200
rect 2751 -188 2767 188
rect 2801 -188 2817 188
rect 2751 -200 2817 -188
rect 2847 188 2913 200
rect 2847 -188 2863 188
rect 2897 -188 2913 188
rect 2847 -200 2913 -188
rect 2943 188 3009 200
rect 2943 -188 2959 188
rect 2993 -188 3009 188
rect 2943 -200 3009 -188
rect 3039 188 3105 200
rect 3039 -188 3055 188
rect 3089 -188 3105 188
rect 3039 -200 3105 -188
rect 3135 188 3201 200
rect 3135 -188 3151 188
rect 3185 -188 3201 188
rect 3135 -200 3201 -188
rect 3231 188 3297 200
rect 3231 -188 3247 188
rect 3281 -188 3297 188
rect 3231 -200 3297 -188
rect 3327 188 3393 200
rect 3327 -188 3343 188
rect 3377 -188 3393 188
rect 3327 -200 3393 -188
rect 3423 188 3489 200
rect 3423 -188 3439 188
rect 3473 -188 3489 188
rect 3423 -200 3489 -188
rect 3519 188 3585 200
rect 3519 -188 3535 188
rect 3569 -188 3585 188
rect 3519 -200 3585 -188
rect 3615 188 3681 200
rect 3615 -188 3631 188
rect 3665 -188 3681 188
rect 3615 -200 3681 -188
rect 3711 188 3777 200
rect 3711 -188 3727 188
rect 3761 -188 3777 188
rect 3711 -200 3777 -188
rect 3807 188 3869 200
rect 3807 -188 3823 188
rect 3857 -188 3869 188
rect 3807 -200 3869 -188
rect -3869 -430 -3807 -418
rect -3869 -806 -3857 -430
rect -3823 -806 -3807 -430
rect -3869 -818 -3807 -806
rect -3777 -430 -3711 -418
rect -3777 -806 -3761 -430
rect -3727 -806 -3711 -430
rect -3777 -818 -3711 -806
rect -3681 -430 -3615 -418
rect -3681 -806 -3665 -430
rect -3631 -806 -3615 -430
rect -3681 -818 -3615 -806
rect -3585 -430 -3519 -418
rect -3585 -806 -3569 -430
rect -3535 -806 -3519 -430
rect -3585 -818 -3519 -806
rect -3489 -430 -3423 -418
rect -3489 -806 -3473 -430
rect -3439 -806 -3423 -430
rect -3489 -818 -3423 -806
rect -3393 -430 -3327 -418
rect -3393 -806 -3377 -430
rect -3343 -806 -3327 -430
rect -3393 -818 -3327 -806
rect -3297 -430 -3231 -418
rect -3297 -806 -3281 -430
rect -3247 -806 -3231 -430
rect -3297 -818 -3231 -806
rect -3201 -430 -3135 -418
rect -3201 -806 -3185 -430
rect -3151 -806 -3135 -430
rect -3201 -818 -3135 -806
rect -3105 -430 -3039 -418
rect -3105 -806 -3089 -430
rect -3055 -806 -3039 -430
rect -3105 -818 -3039 -806
rect -3009 -430 -2943 -418
rect -3009 -806 -2993 -430
rect -2959 -806 -2943 -430
rect -3009 -818 -2943 -806
rect -2913 -430 -2847 -418
rect -2913 -806 -2897 -430
rect -2863 -806 -2847 -430
rect -2913 -818 -2847 -806
rect -2817 -430 -2751 -418
rect -2817 -806 -2801 -430
rect -2767 -806 -2751 -430
rect -2817 -818 -2751 -806
rect -2721 -430 -2655 -418
rect -2721 -806 -2705 -430
rect -2671 -806 -2655 -430
rect -2721 -818 -2655 -806
rect -2625 -430 -2559 -418
rect -2625 -806 -2609 -430
rect -2575 -806 -2559 -430
rect -2625 -818 -2559 -806
rect -2529 -430 -2463 -418
rect -2529 -806 -2513 -430
rect -2479 -806 -2463 -430
rect -2529 -818 -2463 -806
rect -2433 -430 -2367 -418
rect -2433 -806 -2417 -430
rect -2383 -806 -2367 -430
rect -2433 -818 -2367 -806
rect -2337 -430 -2271 -418
rect -2337 -806 -2321 -430
rect -2287 -806 -2271 -430
rect -2337 -818 -2271 -806
rect -2241 -430 -2175 -418
rect -2241 -806 -2225 -430
rect -2191 -806 -2175 -430
rect -2241 -818 -2175 -806
rect -2145 -430 -2079 -418
rect -2145 -806 -2129 -430
rect -2095 -806 -2079 -430
rect -2145 -818 -2079 -806
rect -2049 -430 -1983 -418
rect -2049 -806 -2033 -430
rect -1999 -806 -1983 -430
rect -2049 -818 -1983 -806
rect -1953 -430 -1887 -418
rect -1953 -806 -1937 -430
rect -1903 -806 -1887 -430
rect -1953 -818 -1887 -806
rect -1857 -430 -1791 -418
rect -1857 -806 -1841 -430
rect -1807 -806 -1791 -430
rect -1857 -818 -1791 -806
rect -1761 -430 -1695 -418
rect -1761 -806 -1745 -430
rect -1711 -806 -1695 -430
rect -1761 -818 -1695 -806
rect -1665 -430 -1599 -418
rect -1665 -806 -1649 -430
rect -1615 -806 -1599 -430
rect -1665 -818 -1599 -806
rect -1569 -430 -1503 -418
rect -1569 -806 -1553 -430
rect -1519 -806 -1503 -430
rect -1569 -818 -1503 -806
rect -1473 -430 -1407 -418
rect -1473 -806 -1457 -430
rect -1423 -806 -1407 -430
rect -1473 -818 -1407 -806
rect -1377 -430 -1311 -418
rect -1377 -806 -1361 -430
rect -1327 -806 -1311 -430
rect -1377 -818 -1311 -806
rect -1281 -430 -1215 -418
rect -1281 -806 -1265 -430
rect -1231 -806 -1215 -430
rect -1281 -818 -1215 -806
rect -1185 -430 -1119 -418
rect -1185 -806 -1169 -430
rect -1135 -806 -1119 -430
rect -1185 -818 -1119 -806
rect -1089 -430 -1023 -418
rect -1089 -806 -1073 -430
rect -1039 -806 -1023 -430
rect -1089 -818 -1023 -806
rect -993 -430 -927 -418
rect -993 -806 -977 -430
rect -943 -806 -927 -430
rect -993 -818 -927 -806
rect -897 -430 -831 -418
rect -897 -806 -881 -430
rect -847 -806 -831 -430
rect -897 -818 -831 -806
rect -801 -430 -735 -418
rect -801 -806 -785 -430
rect -751 -806 -735 -430
rect -801 -818 -735 -806
rect -705 -430 -639 -418
rect -705 -806 -689 -430
rect -655 -806 -639 -430
rect -705 -818 -639 -806
rect -609 -430 -543 -418
rect -609 -806 -593 -430
rect -559 -806 -543 -430
rect -609 -818 -543 -806
rect -513 -430 -447 -418
rect -513 -806 -497 -430
rect -463 -806 -447 -430
rect -513 -818 -447 -806
rect -417 -430 -351 -418
rect -417 -806 -401 -430
rect -367 -806 -351 -430
rect -417 -818 -351 -806
rect -321 -430 -255 -418
rect -321 -806 -305 -430
rect -271 -806 -255 -430
rect -321 -818 -255 -806
rect -225 -430 -159 -418
rect -225 -806 -209 -430
rect -175 -806 -159 -430
rect -225 -818 -159 -806
rect -129 -430 -63 -418
rect -129 -806 -113 -430
rect -79 -806 -63 -430
rect -129 -818 -63 -806
rect -33 -430 33 -418
rect -33 -806 -17 -430
rect 17 -806 33 -430
rect -33 -818 33 -806
rect 63 -430 129 -418
rect 63 -806 79 -430
rect 113 -806 129 -430
rect 63 -818 129 -806
rect 159 -430 225 -418
rect 159 -806 175 -430
rect 209 -806 225 -430
rect 159 -818 225 -806
rect 255 -430 321 -418
rect 255 -806 271 -430
rect 305 -806 321 -430
rect 255 -818 321 -806
rect 351 -430 417 -418
rect 351 -806 367 -430
rect 401 -806 417 -430
rect 351 -818 417 -806
rect 447 -430 513 -418
rect 447 -806 463 -430
rect 497 -806 513 -430
rect 447 -818 513 -806
rect 543 -430 609 -418
rect 543 -806 559 -430
rect 593 -806 609 -430
rect 543 -818 609 -806
rect 639 -430 705 -418
rect 639 -806 655 -430
rect 689 -806 705 -430
rect 639 -818 705 -806
rect 735 -430 801 -418
rect 735 -806 751 -430
rect 785 -806 801 -430
rect 735 -818 801 -806
rect 831 -430 897 -418
rect 831 -806 847 -430
rect 881 -806 897 -430
rect 831 -818 897 -806
rect 927 -430 993 -418
rect 927 -806 943 -430
rect 977 -806 993 -430
rect 927 -818 993 -806
rect 1023 -430 1089 -418
rect 1023 -806 1039 -430
rect 1073 -806 1089 -430
rect 1023 -818 1089 -806
rect 1119 -430 1185 -418
rect 1119 -806 1135 -430
rect 1169 -806 1185 -430
rect 1119 -818 1185 -806
rect 1215 -430 1281 -418
rect 1215 -806 1231 -430
rect 1265 -806 1281 -430
rect 1215 -818 1281 -806
rect 1311 -430 1377 -418
rect 1311 -806 1327 -430
rect 1361 -806 1377 -430
rect 1311 -818 1377 -806
rect 1407 -430 1473 -418
rect 1407 -806 1423 -430
rect 1457 -806 1473 -430
rect 1407 -818 1473 -806
rect 1503 -430 1569 -418
rect 1503 -806 1519 -430
rect 1553 -806 1569 -430
rect 1503 -818 1569 -806
rect 1599 -430 1665 -418
rect 1599 -806 1615 -430
rect 1649 -806 1665 -430
rect 1599 -818 1665 -806
rect 1695 -430 1761 -418
rect 1695 -806 1711 -430
rect 1745 -806 1761 -430
rect 1695 -818 1761 -806
rect 1791 -430 1857 -418
rect 1791 -806 1807 -430
rect 1841 -806 1857 -430
rect 1791 -818 1857 -806
rect 1887 -430 1953 -418
rect 1887 -806 1903 -430
rect 1937 -806 1953 -430
rect 1887 -818 1953 -806
rect 1983 -430 2049 -418
rect 1983 -806 1999 -430
rect 2033 -806 2049 -430
rect 1983 -818 2049 -806
rect 2079 -430 2145 -418
rect 2079 -806 2095 -430
rect 2129 -806 2145 -430
rect 2079 -818 2145 -806
rect 2175 -430 2241 -418
rect 2175 -806 2191 -430
rect 2225 -806 2241 -430
rect 2175 -818 2241 -806
rect 2271 -430 2337 -418
rect 2271 -806 2287 -430
rect 2321 -806 2337 -430
rect 2271 -818 2337 -806
rect 2367 -430 2433 -418
rect 2367 -806 2383 -430
rect 2417 -806 2433 -430
rect 2367 -818 2433 -806
rect 2463 -430 2529 -418
rect 2463 -806 2479 -430
rect 2513 -806 2529 -430
rect 2463 -818 2529 -806
rect 2559 -430 2625 -418
rect 2559 -806 2575 -430
rect 2609 -806 2625 -430
rect 2559 -818 2625 -806
rect 2655 -430 2721 -418
rect 2655 -806 2671 -430
rect 2705 -806 2721 -430
rect 2655 -818 2721 -806
rect 2751 -430 2817 -418
rect 2751 -806 2767 -430
rect 2801 -806 2817 -430
rect 2751 -818 2817 -806
rect 2847 -430 2913 -418
rect 2847 -806 2863 -430
rect 2897 -806 2913 -430
rect 2847 -818 2913 -806
rect 2943 -430 3009 -418
rect 2943 -806 2959 -430
rect 2993 -806 3009 -430
rect 2943 -818 3009 -806
rect 3039 -430 3105 -418
rect 3039 -806 3055 -430
rect 3089 -806 3105 -430
rect 3039 -818 3105 -806
rect 3135 -430 3201 -418
rect 3135 -806 3151 -430
rect 3185 -806 3201 -430
rect 3135 -818 3201 -806
rect 3231 -430 3297 -418
rect 3231 -806 3247 -430
rect 3281 -806 3297 -430
rect 3231 -818 3297 -806
rect 3327 -430 3393 -418
rect 3327 -806 3343 -430
rect 3377 -806 3393 -430
rect 3327 -818 3393 -806
rect 3423 -430 3489 -418
rect 3423 -806 3439 -430
rect 3473 -806 3489 -430
rect 3423 -818 3489 -806
rect 3519 -430 3585 -418
rect 3519 -806 3535 -430
rect 3569 -806 3585 -430
rect 3519 -818 3585 -806
rect 3615 -430 3681 -418
rect 3615 -806 3631 -430
rect 3665 -806 3681 -430
rect 3615 -818 3681 -806
rect 3711 -430 3777 -418
rect 3711 -806 3727 -430
rect 3761 -806 3777 -430
rect 3711 -818 3777 -806
rect 3807 -430 3869 -418
rect 3807 -806 3823 -430
rect 3857 -806 3869 -430
rect 3807 -818 3869 -806
<< ndiffc >>
rect -3857 430 -3823 806
rect -3761 430 -3727 806
rect -3665 430 -3631 806
rect -3569 430 -3535 806
rect -3473 430 -3439 806
rect -3377 430 -3343 806
rect -3281 430 -3247 806
rect -3185 430 -3151 806
rect -3089 430 -3055 806
rect -2993 430 -2959 806
rect -2897 430 -2863 806
rect -2801 430 -2767 806
rect -2705 430 -2671 806
rect -2609 430 -2575 806
rect -2513 430 -2479 806
rect -2417 430 -2383 806
rect -2321 430 -2287 806
rect -2225 430 -2191 806
rect -2129 430 -2095 806
rect -2033 430 -1999 806
rect -1937 430 -1903 806
rect -1841 430 -1807 806
rect -1745 430 -1711 806
rect -1649 430 -1615 806
rect -1553 430 -1519 806
rect -1457 430 -1423 806
rect -1361 430 -1327 806
rect -1265 430 -1231 806
rect -1169 430 -1135 806
rect -1073 430 -1039 806
rect -977 430 -943 806
rect -881 430 -847 806
rect -785 430 -751 806
rect -689 430 -655 806
rect -593 430 -559 806
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect 559 430 593 806
rect 655 430 689 806
rect 751 430 785 806
rect 847 430 881 806
rect 943 430 977 806
rect 1039 430 1073 806
rect 1135 430 1169 806
rect 1231 430 1265 806
rect 1327 430 1361 806
rect 1423 430 1457 806
rect 1519 430 1553 806
rect 1615 430 1649 806
rect 1711 430 1745 806
rect 1807 430 1841 806
rect 1903 430 1937 806
rect 1999 430 2033 806
rect 2095 430 2129 806
rect 2191 430 2225 806
rect 2287 430 2321 806
rect 2383 430 2417 806
rect 2479 430 2513 806
rect 2575 430 2609 806
rect 2671 430 2705 806
rect 2767 430 2801 806
rect 2863 430 2897 806
rect 2959 430 2993 806
rect 3055 430 3089 806
rect 3151 430 3185 806
rect 3247 430 3281 806
rect 3343 430 3377 806
rect 3439 430 3473 806
rect 3535 430 3569 806
rect 3631 430 3665 806
rect 3727 430 3761 806
rect 3823 430 3857 806
rect -3857 -188 -3823 188
rect -3761 -188 -3727 188
rect -3665 -188 -3631 188
rect -3569 -188 -3535 188
rect -3473 -188 -3439 188
rect -3377 -188 -3343 188
rect -3281 -188 -3247 188
rect -3185 -188 -3151 188
rect -3089 -188 -3055 188
rect -2993 -188 -2959 188
rect -2897 -188 -2863 188
rect -2801 -188 -2767 188
rect -2705 -188 -2671 188
rect -2609 -188 -2575 188
rect -2513 -188 -2479 188
rect -2417 -188 -2383 188
rect -2321 -188 -2287 188
rect -2225 -188 -2191 188
rect -2129 -188 -2095 188
rect -2033 -188 -1999 188
rect -1937 -188 -1903 188
rect -1841 -188 -1807 188
rect -1745 -188 -1711 188
rect -1649 -188 -1615 188
rect -1553 -188 -1519 188
rect -1457 -188 -1423 188
rect -1361 -188 -1327 188
rect -1265 -188 -1231 188
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect 1231 -188 1265 188
rect 1327 -188 1361 188
rect 1423 -188 1457 188
rect 1519 -188 1553 188
rect 1615 -188 1649 188
rect 1711 -188 1745 188
rect 1807 -188 1841 188
rect 1903 -188 1937 188
rect 1999 -188 2033 188
rect 2095 -188 2129 188
rect 2191 -188 2225 188
rect 2287 -188 2321 188
rect 2383 -188 2417 188
rect 2479 -188 2513 188
rect 2575 -188 2609 188
rect 2671 -188 2705 188
rect 2767 -188 2801 188
rect 2863 -188 2897 188
rect 2959 -188 2993 188
rect 3055 -188 3089 188
rect 3151 -188 3185 188
rect 3247 -188 3281 188
rect 3343 -188 3377 188
rect 3439 -188 3473 188
rect 3535 -188 3569 188
rect 3631 -188 3665 188
rect 3727 -188 3761 188
rect 3823 -188 3857 188
rect -3857 -806 -3823 -430
rect -3761 -806 -3727 -430
rect -3665 -806 -3631 -430
rect -3569 -806 -3535 -430
rect -3473 -806 -3439 -430
rect -3377 -806 -3343 -430
rect -3281 -806 -3247 -430
rect -3185 -806 -3151 -430
rect -3089 -806 -3055 -430
rect -2993 -806 -2959 -430
rect -2897 -806 -2863 -430
rect -2801 -806 -2767 -430
rect -2705 -806 -2671 -430
rect -2609 -806 -2575 -430
rect -2513 -806 -2479 -430
rect -2417 -806 -2383 -430
rect -2321 -806 -2287 -430
rect -2225 -806 -2191 -430
rect -2129 -806 -2095 -430
rect -2033 -806 -1999 -430
rect -1937 -806 -1903 -430
rect -1841 -806 -1807 -430
rect -1745 -806 -1711 -430
rect -1649 -806 -1615 -430
rect -1553 -806 -1519 -430
rect -1457 -806 -1423 -430
rect -1361 -806 -1327 -430
rect -1265 -806 -1231 -430
rect -1169 -806 -1135 -430
rect -1073 -806 -1039 -430
rect -977 -806 -943 -430
rect -881 -806 -847 -430
rect -785 -806 -751 -430
rect -689 -806 -655 -430
rect -593 -806 -559 -430
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect 559 -806 593 -430
rect 655 -806 689 -430
rect 751 -806 785 -430
rect 847 -806 881 -430
rect 943 -806 977 -430
rect 1039 -806 1073 -430
rect 1135 -806 1169 -430
rect 1231 -806 1265 -430
rect 1327 -806 1361 -430
rect 1423 -806 1457 -430
rect 1519 -806 1553 -430
rect 1615 -806 1649 -430
rect 1711 -806 1745 -430
rect 1807 -806 1841 -430
rect 1903 -806 1937 -430
rect 1999 -806 2033 -430
rect 2095 -806 2129 -430
rect 2191 -806 2225 -430
rect 2287 -806 2321 -430
rect 2383 -806 2417 -430
rect 2479 -806 2513 -430
rect 2575 -806 2609 -430
rect 2671 -806 2705 -430
rect 2767 -806 2801 -430
rect 2863 -806 2897 -430
rect 2959 -806 2993 -430
rect 3055 -806 3089 -430
rect 3151 -806 3185 -430
rect 3247 -806 3281 -430
rect 3343 -806 3377 -430
rect 3439 -806 3473 -430
rect 3535 -806 3569 -430
rect 3631 -806 3665 -430
rect 3727 -806 3761 -430
rect 3823 -806 3857 -430
<< psubdiff >>
rect -3971 958 -3875 992
rect 3875 958 3971 992
rect -3971 896 -3937 958
rect 3937 896 3971 958
rect -3971 -958 -3937 -896
rect 3937 -958 3971 -896
rect -3971 -992 -3875 -958
rect 3875 -992 3971 -958
<< psubdiffcont >>
rect -3875 958 3875 992
rect -3971 -896 -3937 896
rect 3937 -896 3971 896
rect -3875 -992 3875 -958
<< poly >>
rect -3729 890 -3663 906
rect -3729 856 -3713 890
rect -3679 856 -3663 890
rect -3807 818 -3777 844
rect -3729 840 -3663 856
rect -3537 890 -3471 906
rect -3537 856 -3521 890
rect -3487 856 -3471 890
rect -3711 818 -3681 840
rect -3615 818 -3585 844
rect -3537 840 -3471 856
rect -3345 890 -3279 906
rect -3345 856 -3329 890
rect -3295 856 -3279 890
rect -3519 818 -3489 840
rect -3423 818 -3393 844
rect -3345 840 -3279 856
rect -3153 890 -3087 906
rect -3153 856 -3137 890
rect -3103 856 -3087 890
rect -3327 818 -3297 840
rect -3231 818 -3201 844
rect -3153 840 -3087 856
rect -2961 890 -2895 906
rect -2961 856 -2945 890
rect -2911 856 -2895 890
rect -3135 818 -3105 840
rect -3039 818 -3009 844
rect -2961 840 -2895 856
rect -2769 890 -2703 906
rect -2769 856 -2753 890
rect -2719 856 -2703 890
rect -2943 818 -2913 840
rect -2847 818 -2817 844
rect -2769 840 -2703 856
rect -2577 890 -2511 906
rect -2577 856 -2561 890
rect -2527 856 -2511 890
rect -2751 818 -2721 840
rect -2655 818 -2625 844
rect -2577 840 -2511 856
rect -2385 890 -2319 906
rect -2385 856 -2369 890
rect -2335 856 -2319 890
rect -2559 818 -2529 840
rect -2463 818 -2433 844
rect -2385 840 -2319 856
rect -2193 890 -2127 906
rect -2193 856 -2177 890
rect -2143 856 -2127 890
rect -2367 818 -2337 840
rect -2271 818 -2241 844
rect -2193 840 -2127 856
rect -2001 890 -1935 906
rect -2001 856 -1985 890
rect -1951 856 -1935 890
rect -2175 818 -2145 840
rect -2079 818 -2049 844
rect -2001 840 -1935 856
rect -1809 890 -1743 906
rect -1809 856 -1793 890
rect -1759 856 -1743 890
rect -1983 818 -1953 840
rect -1887 818 -1857 844
rect -1809 840 -1743 856
rect -1617 890 -1551 906
rect -1617 856 -1601 890
rect -1567 856 -1551 890
rect -1791 818 -1761 840
rect -1695 818 -1665 844
rect -1617 840 -1551 856
rect -1425 890 -1359 906
rect -1425 856 -1409 890
rect -1375 856 -1359 890
rect -1599 818 -1569 840
rect -1503 818 -1473 844
rect -1425 840 -1359 856
rect -1233 890 -1167 906
rect -1233 856 -1217 890
rect -1183 856 -1167 890
rect -1407 818 -1377 840
rect -1311 818 -1281 844
rect -1233 840 -1167 856
rect -1041 890 -975 906
rect -1041 856 -1025 890
rect -991 856 -975 890
rect -1215 818 -1185 840
rect -1119 818 -1089 844
rect -1041 840 -975 856
rect -849 890 -783 906
rect -849 856 -833 890
rect -799 856 -783 890
rect -1023 818 -993 840
rect -927 818 -897 844
rect -849 840 -783 856
rect -657 890 -591 906
rect -657 856 -641 890
rect -607 856 -591 890
rect -831 818 -801 840
rect -735 818 -705 844
rect -657 840 -591 856
rect -465 890 -399 906
rect -465 856 -449 890
rect -415 856 -399 890
rect -639 818 -609 840
rect -543 818 -513 844
rect -465 840 -399 856
rect -273 890 -207 906
rect -273 856 -257 890
rect -223 856 -207 890
rect -447 818 -417 840
rect -351 818 -321 844
rect -273 840 -207 856
rect -81 890 -15 906
rect -81 856 -65 890
rect -31 856 -15 890
rect -255 818 -225 840
rect -159 818 -129 844
rect -81 840 -15 856
rect 111 890 177 906
rect 111 856 127 890
rect 161 856 177 890
rect -63 818 -33 840
rect 33 818 63 844
rect 111 840 177 856
rect 303 890 369 906
rect 303 856 319 890
rect 353 856 369 890
rect 129 818 159 840
rect 225 818 255 844
rect 303 840 369 856
rect 495 890 561 906
rect 495 856 511 890
rect 545 856 561 890
rect 321 818 351 840
rect 417 818 447 844
rect 495 840 561 856
rect 687 890 753 906
rect 687 856 703 890
rect 737 856 753 890
rect 513 818 543 840
rect 609 818 639 844
rect 687 840 753 856
rect 879 890 945 906
rect 879 856 895 890
rect 929 856 945 890
rect 705 818 735 840
rect 801 818 831 844
rect 879 840 945 856
rect 1071 890 1137 906
rect 1071 856 1087 890
rect 1121 856 1137 890
rect 897 818 927 840
rect 993 818 1023 844
rect 1071 840 1137 856
rect 1263 890 1329 906
rect 1263 856 1279 890
rect 1313 856 1329 890
rect 1089 818 1119 840
rect 1185 818 1215 844
rect 1263 840 1329 856
rect 1455 890 1521 906
rect 1455 856 1471 890
rect 1505 856 1521 890
rect 1281 818 1311 840
rect 1377 818 1407 844
rect 1455 840 1521 856
rect 1647 890 1713 906
rect 1647 856 1663 890
rect 1697 856 1713 890
rect 1473 818 1503 840
rect 1569 818 1599 844
rect 1647 840 1713 856
rect 1839 890 1905 906
rect 1839 856 1855 890
rect 1889 856 1905 890
rect 1665 818 1695 840
rect 1761 818 1791 844
rect 1839 840 1905 856
rect 2031 890 2097 906
rect 2031 856 2047 890
rect 2081 856 2097 890
rect 1857 818 1887 840
rect 1953 818 1983 844
rect 2031 840 2097 856
rect 2223 890 2289 906
rect 2223 856 2239 890
rect 2273 856 2289 890
rect 2049 818 2079 840
rect 2145 818 2175 844
rect 2223 840 2289 856
rect 2415 890 2481 906
rect 2415 856 2431 890
rect 2465 856 2481 890
rect 2241 818 2271 840
rect 2337 818 2367 844
rect 2415 840 2481 856
rect 2607 890 2673 906
rect 2607 856 2623 890
rect 2657 856 2673 890
rect 2433 818 2463 840
rect 2529 818 2559 844
rect 2607 840 2673 856
rect 2799 890 2865 906
rect 2799 856 2815 890
rect 2849 856 2865 890
rect 2625 818 2655 840
rect 2721 818 2751 844
rect 2799 840 2865 856
rect 2991 890 3057 906
rect 2991 856 3007 890
rect 3041 856 3057 890
rect 2817 818 2847 840
rect 2913 818 2943 844
rect 2991 840 3057 856
rect 3183 890 3249 906
rect 3183 856 3199 890
rect 3233 856 3249 890
rect 3009 818 3039 840
rect 3105 818 3135 844
rect 3183 840 3249 856
rect 3375 890 3441 906
rect 3375 856 3391 890
rect 3425 856 3441 890
rect 3201 818 3231 840
rect 3297 818 3327 844
rect 3375 840 3441 856
rect 3567 890 3633 906
rect 3567 856 3583 890
rect 3617 856 3633 890
rect 3393 818 3423 840
rect 3489 818 3519 844
rect 3567 840 3633 856
rect 3759 890 3825 906
rect 3759 856 3775 890
rect 3809 856 3825 890
rect 3585 818 3615 840
rect 3681 818 3711 844
rect 3759 840 3825 856
rect 3777 818 3807 840
rect -3807 396 -3777 418
rect -3825 380 -3759 396
rect -3711 392 -3681 418
rect -3615 396 -3585 418
rect -3825 346 -3809 380
rect -3775 346 -3759 380
rect -3825 330 -3759 346
rect -3633 380 -3567 396
rect -3519 392 -3489 418
rect -3423 396 -3393 418
rect -3633 346 -3617 380
rect -3583 346 -3567 380
rect -3633 330 -3567 346
rect -3441 380 -3375 396
rect -3327 392 -3297 418
rect -3231 396 -3201 418
rect -3441 346 -3425 380
rect -3391 346 -3375 380
rect -3441 330 -3375 346
rect -3249 380 -3183 396
rect -3135 392 -3105 418
rect -3039 396 -3009 418
rect -3249 346 -3233 380
rect -3199 346 -3183 380
rect -3249 330 -3183 346
rect -3057 380 -2991 396
rect -2943 392 -2913 418
rect -2847 396 -2817 418
rect -3057 346 -3041 380
rect -3007 346 -2991 380
rect -3057 330 -2991 346
rect -2865 380 -2799 396
rect -2751 392 -2721 418
rect -2655 396 -2625 418
rect -2865 346 -2849 380
rect -2815 346 -2799 380
rect -2865 330 -2799 346
rect -2673 380 -2607 396
rect -2559 392 -2529 418
rect -2463 396 -2433 418
rect -2673 346 -2657 380
rect -2623 346 -2607 380
rect -2673 330 -2607 346
rect -2481 380 -2415 396
rect -2367 392 -2337 418
rect -2271 396 -2241 418
rect -2481 346 -2465 380
rect -2431 346 -2415 380
rect -2481 330 -2415 346
rect -2289 380 -2223 396
rect -2175 392 -2145 418
rect -2079 396 -2049 418
rect -2289 346 -2273 380
rect -2239 346 -2223 380
rect -2289 330 -2223 346
rect -2097 380 -2031 396
rect -1983 392 -1953 418
rect -1887 396 -1857 418
rect -2097 346 -2081 380
rect -2047 346 -2031 380
rect -2097 330 -2031 346
rect -1905 380 -1839 396
rect -1791 392 -1761 418
rect -1695 396 -1665 418
rect -1905 346 -1889 380
rect -1855 346 -1839 380
rect -1905 330 -1839 346
rect -1713 380 -1647 396
rect -1599 392 -1569 418
rect -1503 396 -1473 418
rect -1713 346 -1697 380
rect -1663 346 -1647 380
rect -1713 330 -1647 346
rect -1521 380 -1455 396
rect -1407 392 -1377 418
rect -1311 396 -1281 418
rect -1521 346 -1505 380
rect -1471 346 -1455 380
rect -1521 330 -1455 346
rect -1329 380 -1263 396
rect -1215 392 -1185 418
rect -1119 396 -1089 418
rect -1329 346 -1313 380
rect -1279 346 -1263 380
rect -1329 330 -1263 346
rect -1137 380 -1071 396
rect -1023 392 -993 418
rect -927 396 -897 418
rect -1137 346 -1121 380
rect -1087 346 -1071 380
rect -1137 330 -1071 346
rect -945 380 -879 396
rect -831 392 -801 418
rect -735 396 -705 418
rect -945 346 -929 380
rect -895 346 -879 380
rect -945 330 -879 346
rect -753 380 -687 396
rect -639 392 -609 418
rect -543 396 -513 418
rect -753 346 -737 380
rect -703 346 -687 380
rect -753 330 -687 346
rect -561 380 -495 396
rect -447 392 -417 418
rect -351 396 -321 418
rect -561 346 -545 380
rect -511 346 -495 380
rect -561 330 -495 346
rect -369 380 -303 396
rect -255 392 -225 418
rect -159 396 -129 418
rect -369 346 -353 380
rect -319 346 -303 380
rect -369 330 -303 346
rect -177 380 -111 396
rect -63 392 -33 418
rect 33 396 63 418
rect -177 346 -161 380
rect -127 346 -111 380
rect -177 330 -111 346
rect 15 380 81 396
rect 129 392 159 418
rect 225 396 255 418
rect 15 346 31 380
rect 65 346 81 380
rect 15 330 81 346
rect 207 380 273 396
rect 321 392 351 418
rect 417 396 447 418
rect 207 346 223 380
rect 257 346 273 380
rect 207 330 273 346
rect 399 380 465 396
rect 513 392 543 418
rect 609 396 639 418
rect 399 346 415 380
rect 449 346 465 380
rect 399 330 465 346
rect 591 380 657 396
rect 705 392 735 418
rect 801 396 831 418
rect 591 346 607 380
rect 641 346 657 380
rect 591 330 657 346
rect 783 380 849 396
rect 897 392 927 418
rect 993 396 1023 418
rect 783 346 799 380
rect 833 346 849 380
rect 783 330 849 346
rect 975 380 1041 396
rect 1089 392 1119 418
rect 1185 396 1215 418
rect 975 346 991 380
rect 1025 346 1041 380
rect 975 330 1041 346
rect 1167 380 1233 396
rect 1281 392 1311 418
rect 1377 396 1407 418
rect 1167 346 1183 380
rect 1217 346 1233 380
rect 1167 330 1233 346
rect 1359 380 1425 396
rect 1473 392 1503 418
rect 1569 396 1599 418
rect 1359 346 1375 380
rect 1409 346 1425 380
rect 1359 330 1425 346
rect 1551 380 1617 396
rect 1665 392 1695 418
rect 1761 396 1791 418
rect 1551 346 1567 380
rect 1601 346 1617 380
rect 1551 330 1617 346
rect 1743 380 1809 396
rect 1857 392 1887 418
rect 1953 396 1983 418
rect 1743 346 1759 380
rect 1793 346 1809 380
rect 1743 330 1809 346
rect 1935 380 2001 396
rect 2049 392 2079 418
rect 2145 396 2175 418
rect 1935 346 1951 380
rect 1985 346 2001 380
rect 1935 330 2001 346
rect 2127 380 2193 396
rect 2241 392 2271 418
rect 2337 396 2367 418
rect 2127 346 2143 380
rect 2177 346 2193 380
rect 2127 330 2193 346
rect 2319 380 2385 396
rect 2433 392 2463 418
rect 2529 396 2559 418
rect 2319 346 2335 380
rect 2369 346 2385 380
rect 2319 330 2385 346
rect 2511 380 2577 396
rect 2625 392 2655 418
rect 2721 396 2751 418
rect 2511 346 2527 380
rect 2561 346 2577 380
rect 2511 330 2577 346
rect 2703 380 2769 396
rect 2817 392 2847 418
rect 2913 396 2943 418
rect 2703 346 2719 380
rect 2753 346 2769 380
rect 2703 330 2769 346
rect 2895 380 2961 396
rect 3009 392 3039 418
rect 3105 396 3135 418
rect 2895 346 2911 380
rect 2945 346 2961 380
rect 2895 330 2961 346
rect 3087 380 3153 396
rect 3201 392 3231 418
rect 3297 396 3327 418
rect 3087 346 3103 380
rect 3137 346 3153 380
rect 3087 330 3153 346
rect 3279 380 3345 396
rect 3393 392 3423 418
rect 3489 396 3519 418
rect 3279 346 3295 380
rect 3329 346 3345 380
rect 3279 330 3345 346
rect 3471 380 3537 396
rect 3585 392 3615 418
rect 3681 396 3711 418
rect 3471 346 3487 380
rect 3521 346 3537 380
rect 3471 330 3537 346
rect 3663 380 3729 396
rect 3777 392 3807 418
rect 3663 346 3679 380
rect 3713 346 3729 380
rect 3663 330 3729 346
rect -3825 272 -3759 288
rect -3825 238 -3809 272
rect -3775 238 -3759 272
rect -3825 222 -3759 238
rect -3633 272 -3567 288
rect -3633 238 -3617 272
rect -3583 238 -3567 272
rect -3807 200 -3777 222
rect -3711 200 -3681 226
rect -3633 222 -3567 238
rect -3441 272 -3375 288
rect -3441 238 -3425 272
rect -3391 238 -3375 272
rect -3615 200 -3585 222
rect -3519 200 -3489 226
rect -3441 222 -3375 238
rect -3249 272 -3183 288
rect -3249 238 -3233 272
rect -3199 238 -3183 272
rect -3423 200 -3393 222
rect -3327 200 -3297 226
rect -3249 222 -3183 238
rect -3057 272 -2991 288
rect -3057 238 -3041 272
rect -3007 238 -2991 272
rect -3231 200 -3201 222
rect -3135 200 -3105 226
rect -3057 222 -2991 238
rect -2865 272 -2799 288
rect -2865 238 -2849 272
rect -2815 238 -2799 272
rect -3039 200 -3009 222
rect -2943 200 -2913 226
rect -2865 222 -2799 238
rect -2673 272 -2607 288
rect -2673 238 -2657 272
rect -2623 238 -2607 272
rect -2847 200 -2817 222
rect -2751 200 -2721 226
rect -2673 222 -2607 238
rect -2481 272 -2415 288
rect -2481 238 -2465 272
rect -2431 238 -2415 272
rect -2655 200 -2625 222
rect -2559 200 -2529 226
rect -2481 222 -2415 238
rect -2289 272 -2223 288
rect -2289 238 -2273 272
rect -2239 238 -2223 272
rect -2463 200 -2433 222
rect -2367 200 -2337 226
rect -2289 222 -2223 238
rect -2097 272 -2031 288
rect -2097 238 -2081 272
rect -2047 238 -2031 272
rect -2271 200 -2241 222
rect -2175 200 -2145 226
rect -2097 222 -2031 238
rect -1905 272 -1839 288
rect -1905 238 -1889 272
rect -1855 238 -1839 272
rect -2079 200 -2049 222
rect -1983 200 -1953 226
rect -1905 222 -1839 238
rect -1713 272 -1647 288
rect -1713 238 -1697 272
rect -1663 238 -1647 272
rect -1887 200 -1857 222
rect -1791 200 -1761 226
rect -1713 222 -1647 238
rect -1521 272 -1455 288
rect -1521 238 -1505 272
rect -1471 238 -1455 272
rect -1695 200 -1665 222
rect -1599 200 -1569 226
rect -1521 222 -1455 238
rect -1329 272 -1263 288
rect -1329 238 -1313 272
rect -1279 238 -1263 272
rect -1503 200 -1473 222
rect -1407 200 -1377 226
rect -1329 222 -1263 238
rect -1137 272 -1071 288
rect -1137 238 -1121 272
rect -1087 238 -1071 272
rect -1311 200 -1281 222
rect -1215 200 -1185 226
rect -1137 222 -1071 238
rect -945 272 -879 288
rect -945 238 -929 272
rect -895 238 -879 272
rect -1119 200 -1089 222
rect -1023 200 -993 226
rect -945 222 -879 238
rect -753 272 -687 288
rect -753 238 -737 272
rect -703 238 -687 272
rect -927 200 -897 222
rect -831 200 -801 226
rect -753 222 -687 238
rect -561 272 -495 288
rect -561 238 -545 272
rect -511 238 -495 272
rect -735 200 -705 222
rect -639 200 -609 226
rect -561 222 -495 238
rect -369 272 -303 288
rect -369 238 -353 272
rect -319 238 -303 272
rect -543 200 -513 222
rect -447 200 -417 226
rect -369 222 -303 238
rect -177 272 -111 288
rect -177 238 -161 272
rect -127 238 -111 272
rect -351 200 -321 222
rect -255 200 -225 226
rect -177 222 -111 238
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -159 200 -129 222
rect -63 200 -33 226
rect 15 222 81 238
rect 207 272 273 288
rect 207 238 223 272
rect 257 238 273 272
rect 33 200 63 222
rect 129 200 159 226
rect 207 222 273 238
rect 399 272 465 288
rect 399 238 415 272
rect 449 238 465 272
rect 225 200 255 222
rect 321 200 351 226
rect 399 222 465 238
rect 591 272 657 288
rect 591 238 607 272
rect 641 238 657 272
rect 417 200 447 222
rect 513 200 543 226
rect 591 222 657 238
rect 783 272 849 288
rect 783 238 799 272
rect 833 238 849 272
rect 609 200 639 222
rect 705 200 735 226
rect 783 222 849 238
rect 975 272 1041 288
rect 975 238 991 272
rect 1025 238 1041 272
rect 801 200 831 222
rect 897 200 927 226
rect 975 222 1041 238
rect 1167 272 1233 288
rect 1167 238 1183 272
rect 1217 238 1233 272
rect 993 200 1023 222
rect 1089 200 1119 226
rect 1167 222 1233 238
rect 1359 272 1425 288
rect 1359 238 1375 272
rect 1409 238 1425 272
rect 1185 200 1215 222
rect 1281 200 1311 226
rect 1359 222 1425 238
rect 1551 272 1617 288
rect 1551 238 1567 272
rect 1601 238 1617 272
rect 1377 200 1407 222
rect 1473 200 1503 226
rect 1551 222 1617 238
rect 1743 272 1809 288
rect 1743 238 1759 272
rect 1793 238 1809 272
rect 1569 200 1599 222
rect 1665 200 1695 226
rect 1743 222 1809 238
rect 1935 272 2001 288
rect 1935 238 1951 272
rect 1985 238 2001 272
rect 1761 200 1791 222
rect 1857 200 1887 226
rect 1935 222 2001 238
rect 2127 272 2193 288
rect 2127 238 2143 272
rect 2177 238 2193 272
rect 1953 200 1983 222
rect 2049 200 2079 226
rect 2127 222 2193 238
rect 2319 272 2385 288
rect 2319 238 2335 272
rect 2369 238 2385 272
rect 2145 200 2175 222
rect 2241 200 2271 226
rect 2319 222 2385 238
rect 2511 272 2577 288
rect 2511 238 2527 272
rect 2561 238 2577 272
rect 2337 200 2367 222
rect 2433 200 2463 226
rect 2511 222 2577 238
rect 2703 272 2769 288
rect 2703 238 2719 272
rect 2753 238 2769 272
rect 2529 200 2559 222
rect 2625 200 2655 226
rect 2703 222 2769 238
rect 2895 272 2961 288
rect 2895 238 2911 272
rect 2945 238 2961 272
rect 2721 200 2751 222
rect 2817 200 2847 226
rect 2895 222 2961 238
rect 3087 272 3153 288
rect 3087 238 3103 272
rect 3137 238 3153 272
rect 2913 200 2943 222
rect 3009 200 3039 226
rect 3087 222 3153 238
rect 3279 272 3345 288
rect 3279 238 3295 272
rect 3329 238 3345 272
rect 3105 200 3135 222
rect 3201 200 3231 226
rect 3279 222 3345 238
rect 3471 272 3537 288
rect 3471 238 3487 272
rect 3521 238 3537 272
rect 3297 200 3327 222
rect 3393 200 3423 226
rect 3471 222 3537 238
rect 3663 272 3729 288
rect 3663 238 3679 272
rect 3713 238 3729 272
rect 3489 200 3519 222
rect 3585 200 3615 226
rect 3663 222 3729 238
rect 3681 200 3711 222
rect 3777 200 3807 226
rect -3807 -226 -3777 -200
rect -3711 -222 -3681 -200
rect -3729 -238 -3663 -222
rect -3615 -226 -3585 -200
rect -3519 -222 -3489 -200
rect -3729 -272 -3713 -238
rect -3679 -272 -3663 -238
rect -3729 -288 -3663 -272
rect -3537 -238 -3471 -222
rect -3423 -226 -3393 -200
rect -3327 -222 -3297 -200
rect -3537 -272 -3521 -238
rect -3487 -272 -3471 -238
rect -3537 -288 -3471 -272
rect -3345 -238 -3279 -222
rect -3231 -226 -3201 -200
rect -3135 -222 -3105 -200
rect -3345 -272 -3329 -238
rect -3295 -272 -3279 -238
rect -3345 -288 -3279 -272
rect -3153 -238 -3087 -222
rect -3039 -226 -3009 -200
rect -2943 -222 -2913 -200
rect -3153 -272 -3137 -238
rect -3103 -272 -3087 -238
rect -3153 -288 -3087 -272
rect -2961 -238 -2895 -222
rect -2847 -226 -2817 -200
rect -2751 -222 -2721 -200
rect -2961 -272 -2945 -238
rect -2911 -272 -2895 -238
rect -2961 -288 -2895 -272
rect -2769 -238 -2703 -222
rect -2655 -226 -2625 -200
rect -2559 -222 -2529 -200
rect -2769 -272 -2753 -238
rect -2719 -272 -2703 -238
rect -2769 -288 -2703 -272
rect -2577 -238 -2511 -222
rect -2463 -226 -2433 -200
rect -2367 -222 -2337 -200
rect -2577 -272 -2561 -238
rect -2527 -272 -2511 -238
rect -2577 -288 -2511 -272
rect -2385 -238 -2319 -222
rect -2271 -226 -2241 -200
rect -2175 -222 -2145 -200
rect -2385 -272 -2369 -238
rect -2335 -272 -2319 -238
rect -2385 -288 -2319 -272
rect -2193 -238 -2127 -222
rect -2079 -226 -2049 -200
rect -1983 -222 -1953 -200
rect -2193 -272 -2177 -238
rect -2143 -272 -2127 -238
rect -2193 -288 -2127 -272
rect -2001 -238 -1935 -222
rect -1887 -226 -1857 -200
rect -1791 -222 -1761 -200
rect -2001 -272 -1985 -238
rect -1951 -272 -1935 -238
rect -2001 -288 -1935 -272
rect -1809 -238 -1743 -222
rect -1695 -226 -1665 -200
rect -1599 -222 -1569 -200
rect -1809 -272 -1793 -238
rect -1759 -272 -1743 -238
rect -1809 -288 -1743 -272
rect -1617 -238 -1551 -222
rect -1503 -226 -1473 -200
rect -1407 -222 -1377 -200
rect -1617 -272 -1601 -238
rect -1567 -272 -1551 -238
rect -1617 -288 -1551 -272
rect -1425 -238 -1359 -222
rect -1311 -226 -1281 -200
rect -1215 -222 -1185 -200
rect -1425 -272 -1409 -238
rect -1375 -272 -1359 -238
rect -1425 -288 -1359 -272
rect -1233 -238 -1167 -222
rect -1119 -226 -1089 -200
rect -1023 -222 -993 -200
rect -1233 -272 -1217 -238
rect -1183 -272 -1167 -238
rect -1233 -288 -1167 -272
rect -1041 -238 -975 -222
rect -927 -226 -897 -200
rect -831 -222 -801 -200
rect -1041 -272 -1025 -238
rect -991 -272 -975 -238
rect -1041 -288 -975 -272
rect -849 -238 -783 -222
rect -735 -226 -705 -200
rect -639 -222 -609 -200
rect -849 -272 -833 -238
rect -799 -272 -783 -238
rect -849 -288 -783 -272
rect -657 -238 -591 -222
rect -543 -226 -513 -200
rect -447 -222 -417 -200
rect -657 -272 -641 -238
rect -607 -272 -591 -238
rect -657 -288 -591 -272
rect -465 -238 -399 -222
rect -351 -226 -321 -200
rect -255 -222 -225 -200
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -465 -288 -399 -272
rect -273 -238 -207 -222
rect -159 -226 -129 -200
rect -63 -222 -33 -200
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -273 -288 -207 -272
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect 129 -222 159 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
rect 111 -238 177 -222
rect 225 -226 255 -200
rect 321 -222 351 -200
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 111 -288 177 -272
rect 303 -238 369 -222
rect 417 -226 447 -200
rect 513 -222 543 -200
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 303 -288 369 -272
rect 495 -238 561 -222
rect 609 -226 639 -200
rect 705 -222 735 -200
rect 495 -272 511 -238
rect 545 -272 561 -238
rect 495 -288 561 -272
rect 687 -238 753 -222
rect 801 -226 831 -200
rect 897 -222 927 -200
rect 687 -272 703 -238
rect 737 -272 753 -238
rect 687 -288 753 -272
rect 879 -238 945 -222
rect 993 -226 1023 -200
rect 1089 -222 1119 -200
rect 879 -272 895 -238
rect 929 -272 945 -238
rect 879 -288 945 -272
rect 1071 -238 1137 -222
rect 1185 -226 1215 -200
rect 1281 -222 1311 -200
rect 1071 -272 1087 -238
rect 1121 -272 1137 -238
rect 1071 -288 1137 -272
rect 1263 -238 1329 -222
rect 1377 -226 1407 -200
rect 1473 -222 1503 -200
rect 1263 -272 1279 -238
rect 1313 -272 1329 -238
rect 1263 -288 1329 -272
rect 1455 -238 1521 -222
rect 1569 -226 1599 -200
rect 1665 -222 1695 -200
rect 1455 -272 1471 -238
rect 1505 -272 1521 -238
rect 1455 -288 1521 -272
rect 1647 -238 1713 -222
rect 1761 -226 1791 -200
rect 1857 -222 1887 -200
rect 1647 -272 1663 -238
rect 1697 -272 1713 -238
rect 1647 -288 1713 -272
rect 1839 -238 1905 -222
rect 1953 -226 1983 -200
rect 2049 -222 2079 -200
rect 1839 -272 1855 -238
rect 1889 -272 1905 -238
rect 1839 -288 1905 -272
rect 2031 -238 2097 -222
rect 2145 -226 2175 -200
rect 2241 -222 2271 -200
rect 2031 -272 2047 -238
rect 2081 -272 2097 -238
rect 2031 -288 2097 -272
rect 2223 -238 2289 -222
rect 2337 -226 2367 -200
rect 2433 -222 2463 -200
rect 2223 -272 2239 -238
rect 2273 -272 2289 -238
rect 2223 -288 2289 -272
rect 2415 -238 2481 -222
rect 2529 -226 2559 -200
rect 2625 -222 2655 -200
rect 2415 -272 2431 -238
rect 2465 -272 2481 -238
rect 2415 -288 2481 -272
rect 2607 -238 2673 -222
rect 2721 -226 2751 -200
rect 2817 -222 2847 -200
rect 2607 -272 2623 -238
rect 2657 -272 2673 -238
rect 2607 -288 2673 -272
rect 2799 -238 2865 -222
rect 2913 -226 2943 -200
rect 3009 -222 3039 -200
rect 2799 -272 2815 -238
rect 2849 -272 2865 -238
rect 2799 -288 2865 -272
rect 2991 -238 3057 -222
rect 3105 -226 3135 -200
rect 3201 -222 3231 -200
rect 2991 -272 3007 -238
rect 3041 -272 3057 -238
rect 2991 -288 3057 -272
rect 3183 -238 3249 -222
rect 3297 -226 3327 -200
rect 3393 -222 3423 -200
rect 3183 -272 3199 -238
rect 3233 -272 3249 -238
rect 3183 -288 3249 -272
rect 3375 -238 3441 -222
rect 3489 -226 3519 -200
rect 3585 -222 3615 -200
rect 3375 -272 3391 -238
rect 3425 -272 3441 -238
rect 3375 -288 3441 -272
rect 3567 -238 3633 -222
rect 3681 -226 3711 -200
rect 3777 -222 3807 -200
rect 3567 -272 3583 -238
rect 3617 -272 3633 -238
rect 3567 -288 3633 -272
rect 3759 -238 3825 -222
rect 3759 -272 3775 -238
rect 3809 -272 3825 -238
rect 3759 -288 3825 -272
rect -3729 -346 -3663 -330
rect -3729 -380 -3713 -346
rect -3679 -380 -3663 -346
rect -3807 -418 -3777 -392
rect -3729 -396 -3663 -380
rect -3537 -346 -3471 -330
rect -3537 -380 -3521 -346
rect -3487 -380 -3471 -346
rect -3711 -418 -3681 -396
rect -3615 -418 -3585 -392
rect -3537 -396 -3471 -380
rect -3345 -346 -3279 -330
rect -3345 -380 -3329 -346
rect -3295 -380 -3279 -346
rect -3519 -418 -3489 -396
rect -3423 -418 -3393 -392
rect -3345 -396 -3279 -380
rect -3153 -346 -3087 -330
rect -3153 -380 -3137 -346
rect -3103 -380 -3087 -346
rect -3327 -418 -3297 -396
rect -3231 -418 -3201 -392
rect -3153 -396 -3087 -380
rect -2961 -346 -2895 -330
rect -2961 -380 -2945 -346
rect -2911 -380 -2895 -346
rect -3135 -418 -3105 -396
rect -3039 -418 -3009 -392
rect -2961 -396 -2895 -380
rect -2769 -346 -2703 -330
rect -2769 -380 -2753 -346
rect -2719 -380 -2703 -346
rect -2943 -418 -2913 -396
rect -2847 -418 -2817 -392
rect -2769 -396 -2703 -380
rect -2577 -346 -2511 -330
rect -2577 -380 -2561 -346
rect -2527 -380 -2511 -346
rect -2751 -418 -2721 -396
rect -2655 -418 -2625 -392
rect -2577 -396 -2511 -380
rect -2385 -346 -2319 -330
rect -2385 -380 -2369 -346
rect -2335 -380 -2319 -346
rect -2559 -418 -2529 -396
rect -2463 -418 -2433 -392
rect -2385 -396 -2319 -380
rect -2193 -346 -2127 -330
rect -2193 -380 -2177 -346
rect -2143 -380 -2127 -346
rect -2367 -418 -2337 -396
rect -2271 -418 -2241 -392
rect -2193 -396 -2127 -380
rect -2001 -346 -1935 -330
rect -2001 -380 -1985 -346
rect -1951 -380 -1935 -346
rect -2175 -418 -2145 -396
rect -2079 -418 -2049 -392
rect -2001 -396 -1935 -380
rect -1809 -346 -1743 -330
rect -1809 -380 -1793 -346
rect -1759 -380 -1743 -346
rect -1983 -418 -1953 -396
rect -1887 -418 -1857 -392
rect -1809 -396 -1743 -380
rect -1617 -346 -1551 -330
rect -1617 -380 -1601 -346
rect -1567 -380 -1551 -346
rect -1791 -418 -1761 -396
rect -1695 -418 -1665 -392
rect -1617 -396 -1551 -380
rect -1425 -346 -1359 -330
rect -1425 -380 -1409 -346
rect -1375 -380 -1359 -346
rect -1599 -418 -1569 -396
rect -1503 -418 -1473 -392
rect -1425 -396 -1359 -380
rect -1233 -346 -1167 -330
rect -1233 -380 -1217 -346
rect -1183 -380 -1167 -346
rect -1407 -418 -1377 -396
rect -1311 -418 -1281 -392
rect -1233 -396 -1167 -380
rect -1041 -346 -975 -330
rect -1041 -380 -1025 -346
rect -991 -380 -975 -346
rect -1215 -418 -1185 -396
rect -1119 -418 -1089 -392
rect -1041 -396 -975 -380
rect -849 -346 -783 -330
rect -849 -380 -833 -346
rect -799 -380 -783 -346
rect -1023 -418 -993 -396
rect -927 -418 -897 -392
rect -849 -396 -783 -380
rect -657 -346 -591 -330
rect -657 -380 -641 -346
rect -607 -380 -591 -346
rect -831 -418 -801 -396
rect -735 -418 -705 -392
rect -657 -396 -591 -380
rect -465 -346 -399 -330
rect -465 -380 -449 -346
rect -415 -380 -399 -346
rect -639 -418 -609 -396
rect -543 -418 -513 -392
rect -465 -396 -399 -380
rect -273 -346 -207 -330
rect -273 -380 -257 -346
rect -223 -380 -207 -346
rect -447 -418 -417 -396
rect -351 -418 -321 -392
rect -273 -396 -207 -380
rect -81 -346 -15 -330
rect -81 -380 -65 -346
rect -31 -380 -15 -346
rect -255 -418 -225 -396
rect -159 -418 -129 -392
rect -81 -396 -15 -380
rect 111 -346 177 -330
rect 111 -380 127 -346
rect 161 -380 177 -346
rect -63 -418 -33 -396
rect 33 -418 63 -392
rect 111 -396 177 -380
rect 303 -346 369 -330
rect 303 -380 319 -346
rect 353 -380 369 -346
rect 129 -418 159 -396
rect 225 -418 255 -392
rect 303 -396 369 -380
rect 495 -346 561 -330
rect 495 -380 511 -346
rect 545 -380 561 -346
rect 321 -418 351 -396
rect 417 -418 447 -392
rect 495 -396 561 -380
rect 687 -346 753 -330
rect 687 -380 703 -346
rect 737 -380 753 -346
rect 513 -418 543 -396
rect 609 -418 639 -392
rect 687 -396 753 -380
rect 879 -346 945 -330
rect 879 -380 895 -346
rect 929 -380 945 -346
rect 705 -418 735 -396
rect 801 -418 831 -392
rect 879 -396 945 -380
rect 1071 -346 1137 -330
rect 1071 -380 1087 -346
rect 1121 -380 1137 -346
rect 897 -418 927 -396
rect 993 -418 1023 -392
rect 1071 -396 1137 -380
rect 1263 -346 1329 -330
rect 1263 -380 1279 -346
rect 1313 -380 1329 -346
rect 1089 -418 1119 -396
rect 1185 -418 1215 -392
rect 1263 -396 1329 -380
rect 1455 -346 1521 -330
rect 1455 -380 1471 -346
rect 1505 -380 1521 -346
rect 1281 -418 1311 -396
rect 1377 -418 1407 -392
rect 1455 -396 1521 -380
rect 1647 -346 1713 -330
rect 1647 -380 1663 -346
rect 1697 -380 1713 -346
rect 1473 -418 1503 -396
rect 1569 -418 1599 -392
rect 1647 -396 1713 -380
rect 1839 -346 1905 -330
rect 1839 -380 1855 -346
rect 1889 -380 1905 -346
rect 1665 -418 1695 -396
rect 1761 -418 1791 -392
rect 1839 -396 1905 -380
rect 2031 -346 2097 -330
rect 2031 -380 2047 -346
rect 2081 -380 2097 -346
rect 1857 -418 1887 -396
rect 1953 -418 1983 -392
rect 2031 -396 2097 -380
rect 2223 -346 2289 -330
rect 2223 -380 2239 -346
rect 2273 -380 2289 -346
rect 2049 -418 2079 -396
rect 2145 -418 2175 -392
rect 2223 -396 2289 -380
rect 2415 -346 2481 -330
rect 2415 -380 2431 -346
rect 2465 -380 2481 -346
rect 2241 -418 2271 -396
rect 2337 -418 2367 -392
rect 2415 -396 2481 -380
rect 2607 -346 2673 -330
rect 2607 -380 2623 -346
rect 2657 -380 2673 -346
rect 2433 -418 2463 -396
rect 2529 -418 2559 -392
rect 2607 -396 2673 -380
rect 2799 -346 2865 -330
rect 2799 -380 2815 -346
rect 2849 -380 2865 -346
rect 2625 -418 2655 -396
rect 2721 -418 2751 -392
rect 2799 -396 2865 -380
rect 2991 -346 3057 -330
rect 2991 -380 3007 -346
rect 3041 -380 3057 -346
rect 2817 -418 2847 -396
rect 2913 -418 2943 -392
rect 2991 -396 3057 -380
rect 3183 -346 3249 -330
rect 3183 -380 3199 -346
rect 3233 -380 3249 -346
rect 3009 -418 3039 -396
rect 3105 -418 3135 -392
rect 3183 -396 3249 -380
rect 3375 -346 3441 -330
rect 3375 -380 3391 -346
rect 3425 -380 3441 -346
rect 3201 -418 3231 -396
rect 3297 -418 3327 -392
rect 3375 -396 3441 -380
rect 3567 -346 3633 -330
rect 3567 -380 3583 -346
rect 3617 -380 3633 -346
rect 3393 -418 3423 -396
rect 3489 -418 3519 -392
rect 3567 -396 3633 -380
rect 3759 -346 3825 -330
rect 3759 -380 3775 -346
rect 3809 -380 3825 -346
rect 3585 -418 3615 -396
rect 3681 -418 3711 -392
rect 3759 -396 3825 -380
rect 3777 -418 3807 -396
rect -3807 -840 -3777 -818
rect -3825 -856 -3759 -840
rect -3711 -844 -3681 -818
rect -3615 -840 -3585 -818
rect -3825 -890 -3809 -856
rect -3775 -890 -3759 -856
rect -3825 -906 -3759 -890
rect -3633 -856 -3567 -840
rect -3519 -844 -3489 -818
rect -3423 -840 -3393 -818
rect -3633 -890 -3617 -856
rect -3583 -890 -3567 -856
rect -3633 -906 -3567 -890
rect -3441 -856 -3375 -840
rect -3327 -844 -3297 -818
rect -3231 -840 -3201 -818
rect -3441 -890 -3425 -856
rect -3391 -890 -3375 -856
rect -3441 -906 -3375 -890
rect -3249 -856 -3183 -840
rect -3135 -844 -3105 -818
rect -3039 -840 -3009 -818
rect -3249 -890 -3233 -856
rect -3199 -890 -3183 -856
rect -3249 -906 -3183 -890
rect -3057 -856 -2991 -840
rect -2943 -844 -2913 -818
rect -2847 -840 -2817 -818
rect -3057 -890 -3041 -856
rect -3007 -890 -2991 -856
rect -3057 -906 -2991 -890
rect -2865 -856 -2799 -840
rect -2751 -844 -2721 -818
rect -2655 -840 -2625 -818
rect -2865 -890 -2849 -856
rect -2815 -890 -2799 -856
rect -2865 -906 -2799 -890
rect -2673 -856 -2607 -840
rect -2559 -844 -2529 -818
rect -2463 -840 -2433 -818
rect -2673 -890 -2657 -856
rect -2623 -890 -2607 -856
rect -2673 -906 -2607 -890
rect -2481 -856 -2415 -840
rect -2367 -844 -2337 -818
rect -2271 -840 -2241 -818
rect -2481 -890 -2465 -856
rect -2431 -890 -2415 -856
rect -2481 -906 -2415 -890
rect -2289 -856 -2223 -840
rect -2175 -844 -2145 -818
rect -2079 -840 -2049 -818
rect -2289 -890 -2273 -856
rect -2239 -890 -2223 -856
rect -2289 -906 -2223 -890
rect -2097 -856 -2031 -840
rect -1983 -844 -1953 -818
rect -1887 -840 -1857 -818
rect -2097 -890 -2081 -856
rect -2047 -890 -2031 -856
rect -2097 -906 -2031 -890
rect -1905 -856 -1839 -840
rect -1791 -844 -1761 -818
rect -1695 -840 -1665 -818
rect -1905 -890 -1889 -856
rect -1855 -890 -1839 -856
rect -1905 -906 -1839 -890
rect -1713 -856 -1647 -840
rect -1599 -844 -1569 -818
rect -1503 -840 -1473 -818
rect -1713 -890 -1697 -856
rect -1663 -890 -1647 -856
rect -1713 -906 -1647 -890
rect -1521 -856 -1455 -840
rect -1407 -844 -1377 -818
rect -1311 -840 -1281 -818
rect -1521 -890 -1505 -856
rect -1471 -890 -1455 -856
rect -1521 -906 -1455 -890
rect -1329 -856 -1263 -840
rect -1215 -844 -1185 -818
rect -1119 -840 -1089 -818
rect -1329 -890 -1313 -856
rect -1279 -890 -1263 -856
rect -1329 -906 -1263 -890
rect -1137 -856 -1071 -840
rect -1023 -844 -993 -818
rect -927 -840 -897 -818
rect -1137 -890 -1121 -856
rect -1087 -890 -1071 -856
rect -1137 -906 -1071 -890
rect -945 -856 -879 -840
rect -831 -844 -801 -818
rect -735 -840 -705 -818
rect -945 -890 -929 -856
rect -895 -890 -879 -856
rect -945 -906 -879 -890
rect -753 -856 -687 -840
rect -639 -844 -609 -818
rect -543 -840 -513 -818
rect -753 -890 -737 -856
rect -703 -890 -687 -856
rect -753 -906 -687 -890
rect -561 -856 -495 -840
rect -447 -844 -417 -818
rect -351 -840 -321 -818
rect -561 -890 -545 -856
rect -511 -890 -495 -856
rect -561 -906 -495 -890
rect -369 -856 -303 -840
rect -255 -844 -225 -818
rect -159 -840 -129 -818
rect -369 -890 -353 -856
rect -319 -890 -303 -856
rect -369 -906 -303 -890
rect -177 -856 -111 -840
rect -63 -844 -33 -818
rect 33 -840 63 -818
rect -177 -890 -161 -856
rect -127 -890 -111 -856
rect -177 -906 -111 -890
rect 15 -856 81 -840
rect 129 -844 159 -818
rect 225 -840 255 -818
rect 15 -890 31 -856
rect 65 -890 81 -856
rect 15 -906 81 -890
rect 207 -856 273 -840
rect 321 -844 351 -818
rect 417 -840 447 -818
rect 207 -890 223 -856
rect 257 -890 273 -856
rect 207 -906 273 -890
rect 399 -856 465 -840
rect 513 -844 543 -818
rect 609 -840 639 -818
rect 399 -890 415 -856
rect 449 -890 465 -856
rect 399 -906 465 -890
rect 591 -856 657 -840
rect 705 -844 735 -818
rect 801 -840 831 -818
rect 591 -890 607 -856
rect 641 -890 657 -856
rect 591 -906 657 -890
rect 783 -856 849 -840
rect 897 -844 927 -818
rect 993 -840 1023 -818
rect 783 -890 799 -856
rect 833 -890 849 -856
rect 783 -906 849 -890
rect 975 -856 1041 -840
rect 1089 -844 1119 -818
rect 1185 -840 1215 -818
rect 975 -890 991 -856
rect 1025 -890 1041 -856
rect 975 -906 1041 -890
rect 1167 -856 1233 -840
rect 1281 -844 1311 -818
rect 1377 -840 1407 -818
rect 1167 -890 1183 -856
rect 1217 -890 1233 -856
rect 1167 -906 1233 -890
rect 1359 -856 1425 -840
rect 1473 -844 1503 -818
rect 1569 -840 1599 -818
rect 1359 -890 1375 -856
rect 1409 -890 1425 -856
rect 1359 -906 1425 -890
rect 1551 -856 1617 -840
rect 1665 -844 1695 -818
rect 1761 -840 1791 -818
rect 1551 -890 1567 -856
rect 1601 -890 1617 -856
rect 1551 -906 1617 -890
rect 1743 -856 1809 -840
rect 1857 -844 1887 -818
rect 1953 -840 1983 -818
rect 1743 -890 1759 -856
rect 1793 -890 1809 -856
rect 1743 -906 1809 -890
rect 1935 -856 2001 -840
rect 2049 -844 2079 -818
rect 2145 -840 2175 -818
rect 1935 -890 1951 -856
rect 1985 -890 2001 -856
rect 1935 -906 2001 -890
rect 2127 -856 2193 -840
rect 2241 -844 2271 -818
rect 2337 -840 2367 -818
rect 2127 -890 2143 -856
rect 2177 -890 2193 -856
rect 2127 -906 2193 -890
rect 2319 -856 2385 -840
rect 2433 -844 2463 -818
rect 2529 -840 2559 -818
rect 2319 -890 2335 -856
rect 2369 -890 2385 -856
rect 2319 -906 2385 -890
rect 2511 -856 2577 -840
rect 2625 -844 2655 -818
rect 2721 -840 2751 -818
rect 2511 -890 2527 -856
rect 2561 -890 2577 -856
rect 2511 -906 2577 -890
rect 2703 -856 2769 -840
rect 2817 -844 2847 -818
rect 2913 -840 2943 -818
rect 2703 -890 2719 -856
rect 2753 -890 2769 -856
rect 2703 -906 2769 -890
rect 2895 -856 2961 -840
rect 3009 -844 3039 -818
rect 3105 -840 3135 -818
rect 2895 -890 2911 -856
rect 2945 -890 2961 -856
rect 2895 -906 2961 -890
rect 3087 -856 3153 -840
rect 3201 -844 3231 -818
rect 3297 -840 3327 -818
rect 3087 -890 3103 -856
rect 3137 -890 3153 -856
rect 3087 -906 3153 -890
rect 3279 -856 3345 -840
rect 3393 -844 3423 -818
rect 3489 -840 3519 -818
rect 3279 -890 3295 -856
rect 3329 -890 3345 -856
rect 3279 -906 3345 -890
rect 3471 -856 3537 -840
rect 3585 -844 3615 -818
rect 3681 -840 3711 -818
rect 3471 -890 3487 -856
rect 3521 -890 3537 -856
rect 3471 -906 3537 -890
rect 3663 -856 3729 -840
rect 3777 -844 3807 -818
rect 3663 -890 3679 -856
rect 3713 -890 3729 -856
rect 3663 -906 3729 -890
<< polycont >>
rect -3713 856 -3679 890
rect -3521 856 -3487 890
rect -3329 856 -3295 890
rect -3137 856 -3103 890
rect -2945 856 -2911 890
rect -2753 856 -2719 890
rect -2561 856 -2527 890
rect -2369 856 -2335 890
rect -2177 856 -2143 890
rect -1985 856 -1951 890
rect -1793 856 -1759 890
rect -1601 856 -1567 890
rect -1409 856 -1375 890
rect -1217 856 -1183 890
rect -1025 856 -991 890
rect -833 856 -799 890
rect -641 856 -607 890
rect -449 856 -415 890
rect -257 856 -223 890
rect -65 856 -31 890
rect 127 856 161 890
rect 319 856 353 890
rect 511 856 545 890
rect 703 856 737 890
rect 895 856 929 890
rect 1087 856 1121 890
rect 1279 856 1313 890
rect 1471 856 1505 890
rect 1663 856 1697 890
rect 1855 856 1889 890
rect 2047 856 2081 890
rect 2239 856 2273 890
rect 2431 856 2465 890
rect 2623 856 2657 890
rect 2815 856 2849 890
rect 3007 856 3041 890
rect 3199 856 3233 890
rect 3391 856 3425 890
rect 3583 856 3617 890
rect 3775 856 3809 890
rect -3809 346 -3775 380
rect -3617 346 -3583 380
rect -3425 346 -3391 380
rect -3233 346 -3199 380
rect -3041 346 -3007 380
rect -2849 346 -2815 380
rect -2657 346 -2623 380
rect -2465 346 -2431 380
rect -2273 346 -2239 380
rect -2081 346 -2047 380
rect -1889 346 -1855 380
rect -1697 346 -1663 380
rect -1505 346 -1471 380
rect -1313 346 -1279 380
rect -1121 346 -1087 380
rect -929 346 -895 380
rect -737 346 -703 380
rect -545 346 -511 380
rect -353 346 -319 380
rect -161 346 -127 380
rect 31 346 65 380
rect 223 346 257 380
rect 415 346 449 380
rect 607 346 641 380
rect 799 346 833 380
rect 991 346 1025 380
rect 1183 346 1217 380
rect 1375 346 1409 380
rect 1567 346 1601 380
rect 1759 346 1793 380
rect 1951 346 1985 380
rect 2143 346 2177 380
rect 2335 346 2369 380
rect 2527 346 2561 380
rect 2719 346 2753 380
rect 2911 346 2945 380
rect 3103 346 3137 380
rect 3295 346 3329 380
rect 3487 346 3521 380
rect 3679 346 3713 380
rect -3809 238 -3775 272
rect -3617 238 -3583 272
rect -3425 238 -3391 272
rect -3233 238 -3199 272
rect -3041 238 -3007 272
rect -2849 238 -2815 272
rect -2657 238 -2623 272
rect -2465 238 -2431 272
rect -2273 238 -2239 272
rect -2081 238 -2047 272
rect -1889 238 -1855 272
rect -1697 238 -1663 272
rect -1505 238 -1471 272
rect -1313 238 -1279 272
rect -1121 238 -1087 272
rect -929 238 -895 272
rect -737 238 -703 272
rect -545 238 -511 272
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect 607 238 641 272
rect 799 238 833 272
rect 991 238 1025 272
rect 1183 238 1217 272
rect 1375 238 1409 272
rect 1567 238 1601 272
rect 1759 238 1793 272
rect 1951 238 1985 272
rect 2143 238 2177 272
rect 2335 238 2369 272
rect 2527 238 2561 272
rect 2719 238 2753 272
rect 2911 238 2945 272
rect 3103 238 3137 272
rect 3295 238 3329 272
rect 3487 238 3521 272
rect 3679 238 3713 272
rect -3713 -272 -3679 -238
rect -3521 -272 -3487 -238
rect -3329 -272 -3295 -238
rect -3137 -272 -3103 -238
rect -2945 -272 -2911 -238
rect -2753 -272 -2719 -238
rect -2561 -272 -2527 -238
rect -2369 -272 -2335 -238
rect -2177 -272 -2143 -238
rect -1985 -272 -1951 -238
rect -1793 -272 -1759 -238
rect -1601 -272 -1567 -238
rect -1409 -272 -1375 -238
rect -1217 -272 -1183 -238
rect -1025 -272 -991 -238
rect -833 -272 -799 -238
rect -641 -272 -607 -238
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect 511 -272 545 -238
rect 703 -272 737 -238
rect 895 -272 929 -238
rect 1087 -272 1121 -238
rect 1279 -272 1313 -238
rect 1471 -272 1505 -238
rect 1663 -272 1697 -238
rect 1855 -272 1889 -238
rect 2047 -272 2081 -238
rect 2239 -272 2273 -238
rect 2431 -272 2465 -238
rect 2623 -272 2657 -238
rect 2815 -272 2849 -238
rect 3007 -272 3041 -238
rect 3199 -272 3233 -238
rect 3391 -272 3425 -238
rect 3583 -272 3617 -238
rect 3775 -272 3809 -238
rect -3713 -380 -3679 -346
rect -3521 -380 -3487 -346
rect -3329 -380 -3295 -346
rect -3137 -380 -3103 -346
rect -2945 -380 -2911 -346
rect -2753 -380 -2719 -346
rect -2561 -380 -2527 -346
rect -2369 -380 -2335 -346
rect -2177 -380 -2143 -346
rect -1985 -380 -1951 -346
rect -1793 -380 -1759 -346
rect -1601 -380 -1567 -346
rect -1409 -380 -1375 -346
rect -1217 -380 -1183 -346
rect -1025 -380 -991 -346
rect -833 -380 -799 -346
rect -641 -380 -607 -346
rect -449 -380 -415 -346
rect -257 -380 -223 -346
rect -65 -380 -31 -346
rect 127 -380 161 -346
rect 319 -380 353 -346
rect 511 -380 545 -346
rect 703 -380 737 -346
rect 895 -380 929 -346
rect 1087 -380 1121 -346
rect 1279 -380 1313 -346
rect 1471 -380 1505 -346
rect 1663 -380 1697 -346
rect 1855 -380 1889 -346
rect 2047 -380 2081 -346
rect 2239 -380 2273 -346
rect 2431 -380 2465 -346
rect 2623 -380 2657 -346
rect 2815 -380 2849 -346
rect 3007 -380 3041 -346
rect 3199 -380 3233 -346
rect 3391 -380 3425 -346
rect 3583 -380 3617 -346
rect 3775 -380 3809 -346
rect -3809 -890 -3775 -856
rect -3617 -890 -3583 -856
rect -3425 -890 -3391 -856
rect -3233 -890 -3199 -856
rect -3041 -890 -3007 -856
rect -2849 -890 -2815 -856
rect -2657 -890 -2623 -856
rect -2465 -890 -2431 -856
rect -2273 -890 -2239 -856
rect -2081 -890 -2047 -856
rect -1889 -890 -1855 -856
rect -1697 -890 -1663 -856
rect -1505 -890 -1471 -856
rect -1313 -890 -1279 -856
rect -1121 -890 -1087 -856
rect -929 -890 -895 -856
rect -737 -890 -703 -856
rect -545 -890 -511 -856
rect -353 -890 -319 -856
rect -161 -890 -127 -856
rect 31 -890 65 -856
rect 223 -890 257 -856
rect 415 -890 449 -856
rect 607 -890 641 -856
rect 799 -890 833 -856
rect 991 -890 1025 -856
rect 1183 -890 1217 -856
rect 1375 -890 1409 -856
rect 1567 -890 1601 -856
rect 1759 -890 1793 -856
rect 1951 -890 1985 -856
rect 2143 -890 2177 -856
rect 2335 -890 2369 -856
rect 2527 -890 2561 -856
rect 2719 -890 2753 -856
rect 2911 -890 2945 -856
rect 3103 -890 3137 -856
rect 3295 -890 3329 -856
rect 3487 -890 3521 -856
rect 3679 -890 3713 -856
<< locali >>
rect -3971 958 -3875 992
rect 3875 958 3971 992
rect -3971 896 -3937 958
rect 3937 896 3971 958
rect -3729 856 -3713 890
rect -3679 856 -3663 890
rect -3537 856 -3521 890
rect -3487 856 -3471 890
rect -3345 856 -3329 890
rect -3295 856 -3279 890
rect -3153 856 -3137 890
rect -3103 856 -3087 890
rect -2961 856 -2945 890
rect -2911 856 -2895 890
rect -2769 856 -2753 890
rect -2719 856 -2703 890
rect -2577 856 -2561 890
rect -2527 856 -2511 890
rect -2385 856 -2369 890
rect -2335 856 -2319 890
rect -2193 856 -2177 890
rect -2143 856 -2127 890
rect -2001 856 -1985 890
rect -1951 856 -1935 890
rect -1809 856 -1793 890
rect -1759 856 -1743 890
rect -1617 856 -1601 890
rect -1567 856 -1551 890
rect -1425 856 -1409 890
rect -1375 856 -1359 890
rect -1233 856 -1217 890
rect -1183 856 -1167 890
rect -1041 856 -1025 890
rect -991 856 -975 890
rect -849 856 -833 890
rect -799 856 -783 890
rect -657 856 -641 890
rect -607 856 -591 890
rect -465 856 -449 890
rect -415 856 -399 890
rect -273 856 -257 890
rect -223 856 -207 890
rect -81 856 -65 890
rect -31 856 -15 890
rect 111 856 127 890
rect 161 856 177 890
rect 303 856 319 890
rect 353 856 369 890
rect 495 856 511 890
rect 545 856 561 890
rect 687 856 703 890
rect 737 856 753 890
rect 879 856 895 890
rect 929 856 945 890
rect 1071 856 1087 890
rect 1121 856 1137 890
rect 1263 856 1279 890
rect 1313 856 1329 890
rect 1455 856 1471 890
rect 1505 856 1521 890
rect 1647 856 1663 890
rect 1697 856 1713 890
rect 1839 856 1855 890
rect 1889 856 1905 890
rect 2031 856 2047 890
rect 2081 856 2097 890
rect 2223 856 2239 890
rect 2273 856 2289 890
rect 2415 856 2431 890
rect 2465 856 2481 890
rect 2607 856 2623 890
rect 2657 856 2673 890
rect 2799 856 2815 890
rect 2849 856 2865 890
rect 2991 856 3007 890
rect 3041 856 3057 890
rect 3183 856 3199 890
rect 3233 856 3249 890
rect 3375 856 3391 890
rect 3425 856 3441 890
rect 3567 856 3583 890
rect 3617 856 3633 890
rect 3759 856 3775 890
rect 3809 856 3825 890
rect -3857 806 -3823 822
rect -3857 414 -3823 430
rect -3761 806 -3727 822
rect -3761 414 -3727 430
rect -3665 806 -3631 822
rect -3665 414 -3631 430
rect -3569 806 -3535 822
rect -3569 414 -3535 430
rect -3473 806 -3439 822
rect -3473 414 -3439 430
rect -3377 806 -3343 822
rect -3377 414 -3343 430
rect -3281 806 -3247 822
rect -3281 414 -3247 430
rect -3185 806 -3151 822
rect -3185 414 -3151 430
rect -3089 806 -3055 822
rect -3089 414 -3055 430
rect -2993 806 -2959 822
rect -2993 414 -2959 430
rect -2897 806 -2863 822
rect -2897 414 -2863 430
rect -2801 806 -2767 822
rect -2801 414 -2767 430
rect -2705 806 -2671 822
rect -2705 414 -2671 430
rect -2609 806 -2575 822
rect -2609 414 -2575 430
rect -2513 806 -2479 822
rect -2513 414 -2479 430
rect -2417 806 -2383 822
rect -2417 414 -2383 430
rect -2321 806 -2287 822
rect -2321 414 -2287 430
rect -2225 806 -2191 822
rect -2225 414 -2191 430
rect -2129 806 -2095 822
rect -2129 414 -2095 430
rect -2033 806 -1999 822
rect -2033 414 -1999 430
rect -1937 806 -1903 822
rect -1937 414 -1903 430
rect -1841 806 -1807 822
rect -1841 414 -1807 430
rect -1745 806 -1711 822
rect -1745 414 -1711 430
rect -1649 806 -1615 822
rect -1649 414 -1615 430
rect -1553 806 -1519 822
rect -1553 414 -1519 430
rect -1457 806 -1423 822
rect -1457 414 -1423 430
rect -1361 806 -1327 822
rect -1361 414 -1327 430
rect -1265 806 -1231 822
rect -1265 414 -1231 430
rect -1169 806 -1135 822
rect -1169 414 -1135 430
rect -1073 806 -1039 822
rect -1073 414 -1039 430
rect -977 806 -943 822
rect -977 414 -943 430
rect -881 806 -847 822
rect -881 414 -847 430
rect -785 806 -751 822
rect -785 414 -751 430
rect -689 806 -655 822
rect -689 414 -655 430
rect -593 806 -559 822
rect -593 414 -559 430
rect -497 806 -463 822
rect -497 414 -463 430
rect -401 806 -367 822
rect -401 414 -367 430
rect -305 806 -271 822
rect -305 414 -271 430
rect -209 806 -175 822
rect -209 414 -175 430
rect -113 806 -79 822
rect -113 414 -79 430
rect -17 806 17 822
rect -17 414 17 430
rect 79 806 113 822
rect 79 414 113 430
rect 175 806 209 822
rect 175 414 209 430
rect 271 806 305 822
rect 271 414 305 430
rect 367 806 401 822
rect 367 414 401 430
rect 463 806 497 822
rect 463 414 497 430
rect 559 806 593 822
rect 559 414 593 430
rect 655 806 689 822
rect 655 414 689 430
rect 751 806 785 822
rect 751 414 785 430
rect 847 806 881 822
rect 847 414 881 430
rect 943 806 977 822
rect 943 414 977 430
rect 1039 806 1073 822
rect 1039 414 1073 430
rect 1135 806 1169 822
rect 1135 414 1169 430
rect 1231 806 1265 822
rect 1231 414 1265 430
rect 1327 806 1361 822
rect 1327 414 1361 430
rect 1423 806 1457 822
rect 1423 414 1457 430
rect 1519 806 1553 822
rect 1519 414 1553 430
rect 1615 806 1649 822
rect 1615 414 1649 430
rect 1711 806 1745 822
rect 1711 414 1745 430
rect 1807 806 1841 822
rect 1807 414 1841 430
rect 1903 806 1937 822
rect 1903 414 1937 430
rect 1999 806 2033 822
rect 1999 414 2033 430
rect 2095 806 2129 822
rect 2095 414 2129 430
rect 2191 806 2225 822
rect 2191 414 2225 430
rect 2287 806 2321 822
rect 2287 414 2321 430
rect 2383 806 2417 822
rect 2383 414 2417 430
rect 2479 806 2513 822
rect 2479 414 2513 430
rect 2575 806 2609 822
rect 2575 414 2609 430
rect 2671 806 2705 822
rect 2671 414 2705 430
rect 2767 806 2801 822
rect 2767 414 2801 430
rect 2863 806 2897 822
rect 2863 414 2897 430
rect 2959 806 2993 822
rect 2959 414 2993 430
rect 3055 806 3089 822
rect 3055 414 3089 430
rect 3151 806 3185 822
rect 3151 414 3185 430
rect 3247 806 3281 822
rect 3247 414 3281 430
rect 3343 806 3377 822
rect 3343 414 3377 430
rect 3439 806 3473 822
rect 3439 414 3473 430
rect 3535 806 3569 822
rect 3535 414 3569 430
rect 3631 806 3665 822
rect 3631 414 3665 430
rect 3727 806 3761 822
rect 3727 414 3761 430
rect 3823 806 3857 822
rect 3823 414 3857 430
rect -3825 346 -3809 380
rect -3775 346 -3759 380
rect -3633 346 -3617 380
rect -3583 346 -3567 380
rect -3441 346 -3425 380
rect -3391 346 -3375 380
rect -3249 346 -3233 380
rect -3199 346 -3183 380
rect -3057 346 -3041 380
rect -3007 346 -2991 380
rect -2865 346 -2849 380
rect -2815 346 -2799 380
rect -2673 346 -2657 380
rect -2623 346 -2607 380
rect -2481 346 -2465 380
rect -2431 346 -2415 380
rect -2289 346 -2273 380
rect -2239 346 -2223 380
rect -2097 346 -2081 380
rect -2047 346 -2031 380
rect -1905 346 -1889 380
rect -1855 346 -1839 380
rect -1713 346 -1697 380
rect -1663 346 -1647 380
rect -1521 346 -1505 380
rect -1471 346 -1455 380
rect -1329 346 -1313 380
rect -1279 346 -1263 380
rect -1137 346 -1121 380
rect -1087 346 -1071 380
rect -945 346 -929 380
rect -895 346 -879 380
rect -753 346 -737 380
rect -703 346 -687 380
rect -561 346 -545 380
rect -511 346 -495 380
rect -369 346 -353 380
rect -319 346 -303 380
rect -177 346 -161 380
rect -127 346 -111 380
rect 15 346 31 380
rect 65 346 81 380
rect 207 346 223 380
rect 257 346 273 380
rect 399 346 415 380
rect 449 346 465 380
rect 591 346 607 380
rect 641 346 657 380
rect 783 346 799 380
rect 833 346 849 380
rect 975 346 991 380
rect 1025 346 1041 380
rect 1167 346 1183 380
rect 1217 346 1233 380
rect 1359 346 1375 380
rect 1409 346 1425 380
rect 1551 346 1567 380
rect 1601 346 1617 380
rect 1743 346 1759 380
rect 1793 346 1809 380
rect 1935 346 1951 380
rect 1985 346 2001 380
rect 2127 346 2143 380
rect 2177 346 2193 380
rect 2319 346 2335 380
rect 2369 346 2385 380
rect 2511 346 2527 380
rect 2561 346 2577 380
rect 2703 346 2719 380
rect 2753 346 2769 380
rect 2895 346 2911 380
rect 2945 346 2961 380
rect 3087 346 3103 380
rect 3137 346 3153 380
rect 3279 346 3295 380
rect 3329 346 3345 380
rect 3471 346 3487 380
rect 3521 346 3537 380
rect 3663 346 3679 380
rect 3713 346 3729 380
rect -3825 238 -3809 272
rect -3775 238 -3759 272
rect -3633 238 -3617 272
rect -3583 238 -3567 272
rect -3441 238 -3425 272
rect -3391 238 -3375 272
rect -3249 238 -3233 272
rect -3199 238 -3183 272
rect -3057 238 -3041 272
rect -3007 238 -2991 272
rect -2865 238 -2849 272
rect -2815 238 -2799 272
rect -2673 238 -2657 272
rect -2623 238 -2607 272
rect -2481 238 -2465 272
rect -2431 238 -2415 272
rect -2289 238 -2273 272
rect -2239 238 -2223 272
rect -2097 238 -2081 272
rect -2047 238 -2031 272
rect -1905 238 -1889 272
rect -1855 238 -1839 272
rect -1713 238 -1697 272
rect -1663 238 -1647 272
rect -1521 238 -1505 272
rect -1471 238 -1455 272
rect -1329 238 -1313 272
rect -1279 238 -1263 272
rect -1137 238 -1121 272
rect -1087 238 -1071 272
rect -945 238 -929 272
rect -895 238 -879 272
rect -753 238 -737 272
rect -703 238 -687 272
rect -561 238 -545 272
rect -511 238 -495 272
rect -369 238 -353 272
rect -319 238 -303 272
rect -177 238 -161 272
rect -127 238 -111 272
rect 15 238 31 272
rect 65 238 81 272
rect 207 238 223 272
rect 257 238 273 272
rect 399 238 415 272
rect 449 238 465 272
rect 591 238 607 272
rect 641 238 657 272
rect 783 238 799 272
rect 833 238 849 272
rect 975 238 991 272
rect 1025 238 1041 272
rect 1167 238 1183 272
rect 1217 238 1233 272
rect 1359 238 1375 272
rect 1409 238 1425 272
rect 1551 238 1567 272
rect 1601 238 1617 272
rect 1743 238 1759 272
rect 1793 238 1809 272
rect 1935 238 1951 272
rect 1985 238 2001 272
rect 2127 238 2143 272
rect 2177 238 2193 272
rect 2319 238 2335 272
rect 2369 238 2385 272
rect 2511 238 2527 272
rect 2561 238 2577 272
rect 2703 238 2719 272
rect 2753 238 2769 272
rect 2895 238 2911 272
rect 2945 238 2961 272
rect 3087 238 3103 272
rect 3137 238 3153 272
rect 3279 238 3295 272
rect 3329 238 3345 272
rect 3471 238 3487 272
rect 3521 238 3537 272
rect 3663 238 3679 272
rect 3713 238 3729 272
rect -3857 188 -3823 204
rect -3857 -204 -3823 -188
rect -3761 188 -3727 204
rect -3761 -204 -3727 -188
rect -3665 188 -3631 204
rect -3665 -204 -3631 -188
rect -3569 188 -3535 204
rect -3569 -204 -3535 -188
rect -3473 188 -3439 204
rect -3473 -204 -3439 -188
rect -3377 188 -3343 204
rect -3377 -204 -3343 -188
rect -3281 188 -3247 204
rect -3281 -204 -3247 -188
rect -3185 188 -3151 204
rect -3185 -204 -3151 -188
rect -3089 188 -3055 204
rect -3089 -204 -3055 -188
rect -2993 188 -2959 204
rect -2993 -204 -2959 -188
rect -2897 188 -2863 204
rect -2897 -204 -2863 -188
rect -2801 188 -2767 204
rect -2801 -204 -2767 -188
rect -2705 188 -2671 204
rect -2705 -204 -2671 -188
rect -2609 188 -2575 204
rect -2609 -204 -2575 -188
rect -2513 188 -2479 204
rect -2513 -204 -2479 -188
rect -2417 188 -2383 204
rect -2417 -204 -2383 -188
rect -2321 188 -2287 204
rect -2321 -204 -2287 -188
rect -2225 188 -2191 204
rect -2225 -204 -2191 -188
rect -2129 188 -2095 204
rect -2129 -204 -2095 -188
rect -2033 188 -1999 204
rect -2033 -204 -1999 -188
rect -1937 188 -1903 204
rect -1937 -204 -1903 -188
rect -1841 188 -1807 204
rect -1841 -204 -1807 -188
rect -1745 188 -1711 204
rect -1745 -204 -1711 -188
rect -1649 188 -1615 204
rect -1649 -204 -1615 -188
rect -1553 188 -1519 204
rect -1553 -204 -1519 -188
rect -1457 188 -1423 204
rect -1457 -204 -1423 -188
rect -1361 188 -1327 204
rect -1361 -204 -1327 -188
rect -1265 188 -1231 204
rect -1265 -204 -1231 -188
rect -1169 188 -1135 204
rect -1169 -204 -1135 -188
rect -1073 188 -1039 204
rect -1073 -204 -1039 -188
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect 1039 188 1073 204
rect 1039 -204 1073 -188
rect 1135 188 1169 204
rect 1135 -204 1169 -188
rect 1231 188 1265 204
rect 1231 -204 1265 -188
rect 1327 188 1361 204
rect 1327 -204 1361 -188
rect 1423 188 1457 204
rect 1423 -204 1457 -188
rect 1519 188 1553 204
rect 1519 -204 1553 -188
rect 1615 188 1649 204
rect 1615 -204 1649 -188
rect 1711 188 1745 204
rect 1711 -204 1745 -188
rect 1807 188 1841 204
rect 1807 -204 1841 -188
rect 1903 188 1937 204
rect 1903 -204 1937 -188
rect 1999 188 2033 204
rect 1999 -204 2033 -188
rect 2095 188 2129 204
rect 2095 -204 2129 -188
rect 2191 188 2225 204
rect 2191 -204 2225 -188
rect 2287 188 2321 204
rect 2287 -204 2321 -188
rect 2383 188 2417 204
rect 2383 -204 2417 -188
rect 2479 188 2513 204
rect 2479 -204 2513 -188
rect 2575 188 2609 204
rect 2575 -204 2609 -188
rect 2671 188 2705 204
rect 2671 -204 2705 -188
rect 2767 188 2801 204
rect 2767 -204 2801 -188
rect 2863 188 2897 204
rect 2863 -204 2897 -188
rect 2959 188 2993 204
rect 2959 -204 2993 -188
rect 3055 188 3089 204
rect 3055 -204 3089 -188
rect 3151 188 3185 204
rect 3151 -204 3185 -188
rect 3247 188 3281 204
rect 3247 -204 3281 -188
rect 3343 188 3377 204
rect 3343 -204 3377 -188
rect 3439 188 3473 204
rect 3439 -204 3473 -188
rect 3535 188 3569 204
rect 3535 -204 3569 -188
rect 3631 188 3665 204
rect 3631 -204 3665 -188
rect 3727 188 3761 204
rect 3727 -204 3761 -188
rect 3823 188 3857 204
rect 3823 -204 3857 -188
rect -3729 -272 -3713 -238
rect -3679 -272 -3663 -238
rect -3537 -272 -3521 -238
rect -3487 -272 -3471 -238
rect -3345 -272 -3329 -238
rect -3295 -272 -3279 -238
rect -3153 -272 -3137 -238
rect -3103 -272 -3087 -238
rect -2961 -272 -2945 -238
rect -2911 -272 -2895 -238
rect -2769 -272 -2753 -238
rect -2719 -272 -2703 -238
rect -2577 -272 -2561 -238
rect -2527 -272 -2511 -238
rect -2385 -272 -2369 -238
rect -2335 -272 -2319 -238
rect -2193 -272 -2177 -238
rect -2143 -272 -2127 -238
rect -2001 -272 -1985 -238
rect -1951 -272 -1935 -238
rect -1809 -272 -1793 -238
rect -1759 -272 -1743 -238
rect -1617 -272 -1601 -238
rect -1567 -272 -1551 -238
rect -1425 -272 -1409 -238
rect -1375 -272 -1359 -238
rect -1233 -272 -1217 -238
rect -1183 -272 -1167 -238
rect -1041 -272 -1025 -238
rect -991 -272 -975 -238
rect -849 -272 -833 -238
rect -799 -272 -783 -238
rect -657 -272 -641 -238
rect -607 -272 -591 -238
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 495 -272 511 -238
rect 545 -272 561 -238
rect 687 -272 703 -238
rect 737 -272 753 -238
rect 879 -272 895 -238
rect 929 -272 945 -238
rect 1071 -272 1087 -238
rect 1121 -272 1137 -238
rect 1263 -272 1279 -238
rect 1313 -272 1329 -238
rect 1455 -272 1471 -238
rect 1505 -272 1521 -238
rect 1647 -272 1663 -238
rect 1697 -272 1713 -238
rect 1839 -272 1855 -238
rect 1889 -272 1905 -238
rect 2031 -272 2047 -238
rect 2081 -272 2097 -238
rect 2223 -272 2239 -238
rect 2273 -272 2289 -238
rect 2415 -272 2431 -238
rect 2465 -272 2481 -238
rect 2607 -272 2623 -238
rect 2657 -272 2673 -238
rect 2799 -272 2815 -238
rect 2849 -272 2865 -238
rect 2991 -272 3007 -238
rect 3041 -272 3057 -238
rect 3183 -272 3199 -238
rect 3233 -272 3249 -238
rect 3375 -272 3391 -238
rect 3425 -272 3441 -238
rect 3567 -272 3583 -238
rect 3617 -272 3633 -238
rect 3759 -272 3775 -238
rect 3809 -272 3825 -238
rect -3729 -380 -3713 -346
rect -3679 -380 -3663 -346
rect -3537 -380 -3521 -346
rect -3487 -380 -3471 -346
rect -3345 -380 -3329 -346
rect -3295 -380 -3279 -346
rect -3153 -380 -3137 -346
rect -3103 -380 -3087 -346
rect -2961 -380 -2945 -346
rect -2911 -380 -2895 -346
rect -2769 -380 -2753 -346
rect -2719 -380 -2703 -346
rect -2577 -380 -2561 -346
rect -2527 -380 -2511 -346
rect -2385 -380 -2369 -346
rect -2335 -380 -2319 -346
rect -2193 -380 -2177 -346
rect -2143 -380 -2127 -346
rect -2001 -380 -1985 -346
rect -1951 -380 -1935 -346
rect -1809 -380 -1793 -346
rect -1759 -380 -1743 -346
rect -1617 -380 -1601 -346
rect -1567 -380 -1551 -346
rect -1425 -380 -1409 -346
rect -1375 -380 -1359 -346
rect -1233 -380 -1217 -346
rect -1183 -380 -1167 -346
rect -1041 -380 -1025 -346
rect -991 -380 -975 -346
rect -849 -380 -833 -346
rect -799 -380 -783 -346
rect -657 -380 -641 -346
rect -607 -380 -591 -346
rect -465 -380 -449 -346
rect -415 -380 -399 -346
rect -273 -380 -257 -346
rect -223 -380 -207 -346
rect -81 -380 -65 -346
rect -31 -380 -15 -346
rect 111 -380 127 -346
rect 161 -380 177 -346
rect 303 -380 319 -346
rect 353 -380 369 -346
rect 495 -380 511 -346
rect 545 -380 561 -346
rect 687 -380 703 -346
rect 737 -380 753 -346
rect 879 -380 895 -346
rect 929 -380 945 -346
rect 1071 -380 1087 -346
rect 1121 -380 1137 -346
rect 1263 -380 1279 -346
rect 1313 -380 1329 -346
rect 1455 -380 1471 -346
rect 1505 -380 1521 -346
rect 1647 -380 1663 -346
rect 1697 -380 1713 -346
rect 1839 -380 1855 -346
rect 1889 -380 1905 -346
rect 2031 -380 2047 -346
rect 2081 -380 2097 -346
rect 2223 -380 2239 -346
rect 2273 -380 2289 -346
rect 2415 -380 2431 -346
rect 2465 -380 2481 -346
rect 2607 -380 2623 -346
rect 2657 -380 2673 -346
rect 2799 -380 2815 -346
rect 2849 -380 2865 -346
rect 2991 -380 3007 -346
rect 3041 -380 3057 -346
rect 3183 -380 3199 -346
rect 3233 -380 3249 -346
rect 3375 -380 3391 -346
rect 3425 -380 3441 -346
rect 3567 -380 3583 -346
rect 3617 -380 3633 -346
rect 3759 -380 3775 -346
rect 3809 -380 3825 -346
rect -3857 -430 -3823 -414
rect -3857 -822 -3823 -806
rect -3761 -430 -3727 -414
rect -3761 -822 -3727 -806
rect -3665 -430 -3631 -414
rect -3665 -822 -3631 -806
rect -3569 -430 -3535 -414
rect -3569 -822 -3535 -806
rect -3473 -430 -3439 -414
rect -3473 -822 -3439 -806
rect -3377 -430 -3343 -414
rect -3377 -822 -3343 -806
rect -3281 -430 -3247 -414
rect -3281 -822 -3247 -806
rect -3185 -430 -3151 -414
rect -3185 -822 -3151 -806
rect -3089 -430 -3055 -414
rect -3089 -822 -3055 -806
rect -2993 -430 -2959 -414
rect -2993 -822 -2959 -806
rect -2897 -430 -2863 -414
rect -2897 -822 -2863 -806
rect -2801 -430 -2767 -414
rect -2801 -822 -2767 -806
rect -2705 -430 -2671 -414
rect -2705 -822 -2671 -806
rect -2609 -430 -2575 -414
rect -2609 -822 -2575 -806
rect -2513 -430 -2479 -414
rect -2513 -822 -2479 -806
rect -2417 -430 -2383 -414
rect -2417 -822 -2383 -806
rect -2321 -430 -2287 -414
rect -2321 -822 -2287 -806
rect -2225 -430 -2191 -414
rect -2225 -822 -2191 -806
rect -2129 -430 -2095 -414
rect -2129 -822 -2095 -806
rect -2033 -430 -1999 -414
rect -2033 -822 -1999 -806
rect -1937 -430 -1903 -414
rect -1937 -822 -1903 -806
rect -1841 -430 -1807 -414
rect -1841 -822 -1807 -806
rect -1745 -430 -1711 -414
rect -1745 -822 -1711 -806
rect -1649 -430 -1615 -414
rect -1649 -822 -1615 -806
rect -1553 -430 -1519 -414
rect -1553 -822 -1519 -806
rect -1457 -430 -1423 -414
rect -1457 -822 -1423 -806
rect -1361 -430 -1327 -414
rect -1361 -822 -1327 -806
rect -1265 -430 -1231 -414
rect -1265 -822 -1231 -806
rect -1169 -430 -1135 -414
rect -1169 -822 -1135 -806
rect -1073 -430 -1039 -414
rect -1073 -822 -1039 -806
rect -977 -430 -943 -414
rect -977 -822 -943 -806
rect -881 -430 -847 -414
rect -881 -822 -847 -806
rect -785 -430 -751 -414
rect -785 -822 -751 -806
rect -689 -430 -655 -414
rect -689 -822 -655 -806
rect -593 -430 -559 -414
rect -593 -822 -559 -806
rect -497 -430 -463 -414
rect -497 -822 -463 -806
rect -401 -430 -367 -414
rect -401 -822 -367 -806
rect -305 -430 -271 -414
rect -305 -822 -271 -806
rect -209 -430 -175 -414
rect -209 -822 -175 -806
rect -113 -430 -79 -414
rect -113 -822 -79 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 79 -430 113 -414
rect 79 -822 113 -806
rect 175 -430 209 -414
rect 175 -822 209 -806
rect 271 -430 305 -414
rect 271 -822 305 -806
rect 367 -430 401 -414
rect 367 -822 401 -806
rect 463 -430 497 -414
rect 463 -822 497 -806
rect 559 -430 593 -414
rect 559 -822 593 -806
rect 655 -430 689 -414
rect 655 -822 689 -806
rect 751 -430 785 -414
rect 751 -822 785 -806
rect 847 -430 881 -414
rect 847 -822 881 -806
rect 943 -430 977 -414
rect 943 -822 977 -806
rect 1039 -430 1073 -414
rect 1039 -822 1073 -806
rect 1135 -430 1169 -414
rect 1135 -822 1169 -806
rect 1231 -430 1265 -414
rect 1231 -822 1265 -806
rect 1327 -430 1361 -414
rect 1327 -822 1361 -806
rect 1423 -430 1457 -414
rect 1423 -822 1457 -806
rect 1519 -430 1553 -414
rect 1519 -822 1553 -806
rect 1615 -430 1649 -414
rect 1615 -822 1649 -806
rect 1711 -430 1745 -414
rect 1711 -822 1745 -806
rect 1807 -430 1841 -414
rect 1807 -822 1841 -806
rect 1903 -430 1937 -414
rect 1903 -822 1937 -806
rect 1999 -430 2033 -414
rect 1999 -822 2033 -806
rect 2095 -430 2129 -414
rect 2095 -822 2129 -806
rect 2191 -430 2225 -414
rect 2191 -822 2225 -806
rect 2287 -430 2321 -414
rect 2287 -822 2321 -806
rect 2383 -430 2417 -414
rect 2383 -822 2417 -806
rect 2479 -430 2513 -414
rect 2479 -822 2513 -806
rect 2575 -430 2609 -414
rect 2575 -822 2609 -806
rect 2671 -430 2705 -414
rect 2671 -822 2705 -806
rect 2767 -430 2801 -414
rect 2767 -822 2801 -806
rect 2863 -430 2897 -414
rect 2863 -822 2897 -806
rect 2959 -430 2993 -414
rect 2959 -822 2993 -806
rect 3055 -430 3089 -414
rect 3055 -822 3089 -806
rect 3151 -430 3185 -414
rect 3151 -822 3185 -806
rect 3247 -430 3281 -414
rect 3247 -822 3281 -806
rect 3343 -430 3377 -414
rect 3343 -822 3377 -806
rect 3439 -430 3473 -414
rect 3439 -822 3473 -806
rect 3535 -430 3569 -414
rect 3535 -822 3569 -806
rect 3631 -430 3665 -414
rect 3631 -822 3665 -806
rect 3727 -430 3761 -414
rect 3727 -822 3761 -806
rect 3823 -430 3857 -414
rect 3823 -822 3857 -806
rect -3825 -890 -3809 -856
rect -3775 -890 -3759 -856
rect -3633 -890 -3617 -856
rect -3583 -890 -3567 -856
rect -3441 -890 -3425 -856
rect -3391 -890 -3375 -856
rect -3249 -890 -3233 -856
rect -3199 -890 -3183 -856
rect -3057 -890 -3041 -856
rect -3007 -890 -2991 -856
rect -2865 -890 -2849 -856
rect -2815 -890 -2799 -856
rect -2673 -890 -2657 -856
rect -2623 -890 -2607 -856
rect -2481 -890 -2465 -856
rect -2431 -890 -2415 -856
rect -2289 -890 -2273 -856
rect -2239 -890 -2223 -856
rect -2097 -890 -2081 -856
rect -2047 -890 -2031 -856
rect -1905 -890 -1889 -856
rect -1855 -890 -1839 -856
rect -1713 -890 -1697 -856
rect -1663 -890 -1647 -856
rect -1521 -890 -1505 -856
rect -1471 -890 -1455 -856
rect -1329 -890 -1313 -856
rect -1279 -890 -1263 -856
rect -1137 -890 -1121 -856
rect -1087 -890 -1071 -856
rect -945 -890 -929 -856
rect -895 -890 -879 -856
rect -753 -890 -737 -856
rect -703 -890 -687 -856
rect -561 -890 -545 -856
rect -511 -890 -495 -856
rect -369 -890 -353 -856
rect -319 -890 -303 -856
rect -177 -890 -161 -856
rect -127 -890 -111 -856
rect 15 -890 31 -856
rect 65 -890 81 -856
rect 207 -890 223 -856
rect 257 -890 273 -856
rect 399 -890 415 -856
rect 449 -890 465 -856
rect 591 -890 607 -856
rect 641 -890 657 -856
rect 783 -890 799 -856
rect 833 -890 849 -856
rect 975 -890 991 -856
rect 1025 -890 1041 -856
rect 1167 -890 1183 -856
rect 1217 -890 1233 -856
rect 1359 -890 1375 -856
rect 1409 -890 1425 -856
rect 1551 -890 1567 -856
rect 1601 -890 1617 -856
rect 1743 -890 1759 -856
rect 1793 -890 1809 -856
rect 1935 -890 1951 -856
rect 1985 -890 2001 -856
rect 2127 -890 2143 -856
rect 2177 -890 2193 -856
rect 2319 -890 2335 -856
rect 2369 -890 2385 -856
rect 2511 -890 2527 -856
rect 2561 -890 2577 -856
rect 2703 -890 2719 -856
rect 2753 -890 2769 -856
rect 2895 -890 2911 -856
rect 2945 -890 2961 -856
rect 3087 -890 3103 -856
rect 3137 -890 3153 -856
rect 3279 -890 3295 -856
rect 3329 -890 3345 -856
rect 3471 -890 3487 -856
rect 3521 -890 3537 -856
rect 3663 -890 3679 -856
rect 3713 -890 3729 -856
rect -3971 -958 -3937 -896
rect 3937 -958 3971 -896
rect -3971 -992 -3875 -958
rect 3875 -992 3971 -958
<< viali >>
rect -3713 856 -3679 890
rect -3521 856 -3487 890
rect -3329 856 -3295 890
rect -3137 856 -3103 890
rect -2945 856 -2911 890
rect -2753 856 -2719 890
rect -2561 856 -2527 890
rect -2369 856 -2335 890
rect -2177 856 -2143 890
rect -1985 856 -1951 890
rect -1793 856 -1759 890
rect -1601 856 -1567 890
rect -1409 856 -1375 890
rect -1217 856 -1183 890
rect -1025 856 -991 890
rect -833 856 -799 890
rect -641 856 -607 890
rect -449 856 -415 890
rect -257 856 -223 890
rect -65 856 -31 890
rect 127 856 161 890
rect 319 856 353 890
rect 511 856 545 890
rect 703 856 737 890
rect 895 856 929 890
rect 1087 856 1121 890
rect 1279 856 1313 890
rect 1471 856 1505 890
rect 1663 856 1697 890
rect 1855 856 1889 890
rect 2047 856 2081 890
rect 2239 856 2273 890
rect 2431 856 2465 890
rect 2623 856 2657 890
rect 2815 856 2849 890
rect 3007 856 3041 890
rect 3199 856 3233 890
rect 3391 856 3425 890
rect 3583 856 3617 890
rect 3775 856 3809 890
rect -3857 430 -3823 806
rect -3761 430 -3727 806
rect -3665 430 -3631 806
rect -3569 430 -3535 806
rect -3473 430 -3439 806
rect -3377 430 -3343 806
rect -3281 430 -3247 806
rect -3185 430 -3151 806
rect -3089 430 -3055 806
rect -2993 430 -2959 806
rect -2897 430 -2863 806
rect -2801 430 -2767 806
rect -2705 430 -2671 806
rect -2609 430 -2575 806
rect -2513 430 -2479 806
rect -2417 430 -2383 806
rect -2321 430 -2287 806
rect -2225 430 -2191 806
rect -2129 430 -2095 806
rect -2033 430 -1999 806
rect -1937 430 -1903 806
rect -1841 430 -1807 806
rect -1745 430 -1711 806
rect -1649 430 -1615 806
rect -1553 430 -1519 806
rect -1457 430 -1423 806
rect -1361 430 -1327 806
rect -1265 430 -1231 806
rect -1169 430 -1135 806
rect -1073 430 -1039 806
rect -977 430 -943 806
rect -881 430 -847 806
rect -785 430 -751 806
rect -689 430 -655 806
rect -593 430 -559 806
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect 559 430 593 806
rect 655 430 689 806
rect 751 430 785 806
rect 847 430 881 806
rect 943 430 977 806
rect 1039 430 1073 806
rect 1135 430 1169 806
rect 1231 430 1265 806
rect 1327 430 1361 806
rect 1423 430 1457 806
rect 1519 430 1553 806
rect 1615 430 1649 806
rect 1711 430 1745 806
rect 1807 430 1841 806
rect 1903 430 1937 806
rect 1999 430 2033 806
rect 2095 430 2129 806
rect 2191 430 2225 806
rect 2287 430 2321 806
rect 2383 430 2417 806
rect 2479 430 2513 806
rect 2575 430 2609 806
rect 2671 430 2705 806
rect 2767 430 2801 806
rect 2863 430 2897 806
rect 2959 430 2993 806
rect 3055 430 3089 806
rect 3151 430 3185 806
rect 3247 430 3281 806
rect 3343 430 3377 806
rect 3439 430 3473 806
rect 3535 430 3569 806
rect 3631 430 3665 806
rect 3727 430 3761 806
rect 3823 430 3857 806
rect -3809 346 -3775 380
rect -3617 346 -3583 380
rect -3425 346 -3391 380
rect -3233 346 -3199 380
rect -3041 346 -3007 380
rect -2849 346 -2815 380
rect -2657 346 -2623 380
rect -2465 346 -2431 380
rect -2273 346 -2239 380
rect -2081 346 -2047 380
rect -1889 346 -1855 380
rect -1697 346 -1663 380
rect -1505 346 -1471 380
rect -1313 346 -1279 380
rect -1121 346 -1087 380
rect -929 346 -895 380
rect -737 346 -703 380
rect -545 346 -511 380
rect -353 346 -319 380
rect -161 346 -127 380
rect 31 346 65 380
rect 223 346 257 380
rect 415 346 449 380
rect 607 346 641 380
rect 799 346 833 380
rect 991 346 1025 380
rect 1183 346 1217 380
rect 1375 346 1409 380
rect 1567 346 1601 380
rect 1759 346 1793 380
rect 1951 346 1985 380
rect 2143 346 2177 380
rect 2335 346 2369 380
rect 2527 346 2561 380
rect 2719 346 2753 380
rect 2911 346 2945 380
rect 3103 346 3137 380
rect 3295 346 3329 380
rect 3487 346 3521 380
rect 3679 346 3713 380
rect -3809 238 -3775 272
rect -3617 238 -3583 272
rect -3425 238 -3391 272
rect -3233 238 -3199 272
rect -3041 238 -3007 272
rect -2849 238 -2815 272
rect -2657 238 -2623 272
rect -2465 238 -2431 272
rect -2273 238 -2239 272
rect -2081 238 -2047 272
rect -1889 238 -1855 272
rect -1697 238 -1663 272
rect -1505 238 -1471 272
rect -1313 238 -1279 272
rect -1121 238 -1087 272
rect -929 238 -895 272
rect -737 238 -703 272
rect -545 238 -511 272
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect 607 238 641 272
rect 799 238 833 272
rect 991 238 1025 272
rect 1183 238 1217 272
rect 1375 238 1409 272
rect 1567 238 1601 272
rect 1759 238 1793 272
rect 1951 238 1985 272
rect 2143 238 2177 272
rect 2335 238 2369 272
rect 2527 238 2561 272
rect 2719 238 2753 272
rect 2911 238 2945 272
rect 3103 238 3137 272
rect 3295 238 3329 272
rect 3487 238 3521 272
rect 3679 238 3713 272
rect -3857 -188 -3823 188
rect -3761 -188 -3727 188
rect -3665 -188 -3631 188
rect -3569 -188 -3535 188
rect -3473 -188 -3439 188
rect -3377 -188 -3343 188
rect -3281 -188 -3247 188
rect -3185 -188 -3151 188
rect -3089 -188 -3055 188
rect -2993 -188 -2959 188
rect -2897 -188 -2863 188
rect -2801 -188 -2767 188
rect -2705 -188 -2671 188
rect -2609 -188 -2575 188
rect -2513 -188 -2479 188
rect -2417 -188 -2383 188
rect -2321 -188 -2287 188
rect -2225 -188 -2191 188
rect -2129 -188 -2095 188
rect -2033 -188 -1999 188
rect -1937 -188 -1903 188
rect -1841 -188 -1807 188
rect -1745 -188 -1711 188
rect -1649 -188 -1615 188
rect -1553 -188 -1519 188
rect -1457 -188 -1423 188
rect -1361 -188 -1327 188
rect -1265 -188 -1231 188
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect 1231 -188 1265 188
rect 1327 -188 1361 188
rect 1423 -188 1457 188
rect 1519 -188 1553 188
rect 1615 -188 1649 188
rect 1711 -188 1745 188
rect 1807 -188 1841 188
rect 1903 -188 1937 188
rect 1999 -188 2033 188
rect 2095 -188 2129 188
rect 2191 -188 2225 188
rect 2287 -188 2321 188
rect 2383 -188 2417 188
rect 2479 -188 2513 188
rect 2575 -188 2609 188
rect 2671 -188 2705 188
rect 2767 -188 2801 188
rect 2863 -188 2897 188
rect 2959 -188 2993 188
rect 3055 -188 3089 188
rect 3151 -188 3185 188
rect 3247 -188 3281 188
rect 3343 -188 3377 188
rect 3439 -188 3473 188
rect 3535 -188 3569 188
rect 3631 -188 3665 188
rect 3727 -188 3761 188
rect 3823 -188 3857 188
rect -3713 -272 -3679 -238
rect -3521 -272 -3487 -238
rect -3329 -272 -3295 -238
rect -3137 -272 -3103 -238
rect -2945 -272 -2911 -238
rect -2753 -272 -2719 -238
rect -2561 -272 -2527 -238
rect -2369 -272 -2335 -238
rect -2177 -272 -2143 -238
rect -1985 -272 -1951 -238
rect -1793 -272 -1759 -238
rect -1601 -272 -1567 -238
rect -1409 -272 -1375 -238
rect -1217 -272 -1183 -238
rect -1025 -272 -991 -238
rect -833 -272 -799 -238
rect -641 -272 -607 -238
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect 511 -272 545 -238
rect 703 -272 737 -238
rect 895 -272 929 -238
rect 1087 -272 1121 -238
rect 1279 -272 1313 -238
rect 1471 -272 1505 -238
rect 1663 -272 1697 -238
rect 1855 -272 1889 -238
rect 2047 -272 2081 -238
rect 2239 -272 2273 -238
rect 2431 -272 2465 -238
rect 2623 -272 2657 -238
rect 2815 -272 2849 -238
rect 3007 -272 3041 -238
rect 3199 -272 3233 -238
rect 3391 -272 3425 -238
rect 3583 -272 3617 -238
rect 3775 -272 3809 -238
rect -3713 -380 -3679 -346
rect -3521 -380 -3487 -346
rect -3329 -380 -3295 -346
rect -3137 -380 -3103 -346
rect -2945 -380 -2911 -346
rect -2753 -380 -2719 -346
rect -2561 -380 -2527 -346
rect -2369 -380 -2335 -346
rect -2177 -380 -2143 -346
rect -1985 -380 -1951 -346
rect -1793 -380 -1759 -346
rect -1601 -380 -1567 -346
rect -1409 -380 -1375 -346
rect -1217 -380 -1183 -346
rect -1025 -380 -991 -346
rect -833 -380 -799 -346
rect -641 -380 -607 -346
rect -449 -380 -415 -346
rect -257 -380 -223 -346
rect -65 -380 -31 -346
rect 127 -380 161 -346
rect 319 -380 353 -346
rect 511 -380 545 -346
rect 703 -380 737 -346
rect 895 -380 929 -346
rect 1087 -380 1121 -346
rect 1279 -380 1313 -346
rect 1471 -380 1505 -346
rect 1663 -380 1697 -346
rect 1855 -380 1889 -346
rect 2047 -380 2081 -346
rect 2239 -380 2273 -346
rect 2431 -380 2465 -346
rect 2623 -380 2657 -346
rect 2815 -380 2849 -346
rect 3007 -380 3041 -346
rect 3199 -380 3233 -346
rect 3391 -380 3425 -346
rect 3583 -380 3617 -346
rect 3775 -380 3809 -346
rect -3857 -806 -3823 -430
rect -3761 -806 -3727 -430
rect -3665 -806 -3631 -430
rect -3569 -806 -3535 -430
rect -3473 -806 -3439 -430
rect -3377 -806 -3343 -430
rect -3281 -806 -3247 -430
rect -3185 -806 -3151 -430
rect -3089 -806 -3055 -430
rect -2993 -806 -2959 -430
rect -2897 -806 -2863 -430
rect -2801 -806 -2767 -430
rect -2705 -806 -2671 -430
rect -2609 -806 -2575 -430
rect -2513 -806 -2479 -430
rect -2417 -806 -2383 -430
rect -2321 -806 -2287 -430
rect -2225 -806 -2191 -430
rect -2129 -806 -2095 -430
rect -2033 -806 -1999 -430
rect -1937 -806 -1903 -430
rect -1841 -806 -1807 -430
rect -1745 -806 -1711 -430
rect -1649 -806 -1615 -430
rect -1553 -806 -1519 -430
rect -1457 -806 -1423 -430
rect -1361 -806 -1327 -430
rect -1265 -806 -1231 -430
rect -1169 -806 -1135 -430
rect -1073 -806 -1039 -430
rect -977 -806 -943 -430
rect -881 -806 -847 -430
rect -785 -806 -751 -430
rect -689 -806 -655 -430
rect -593 -806 -559 -430
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect 559 -806 593 -430
rect 655 -806 689 -430
rect 751 -806 785 -430
rect 847 -806 881 -430
rect 943 -806 977 -430
rect 1039 -806 1073 -430
rect 1135 -806 1169 -430
rect 1231 -806 1265 -430
rect 1327 -806 1361 -430
rect 1423 -806 1457 -430
rect 1519 -806 1553 -430
rect 1615 -806 1649 -430
rect 1711 -806 1745 -430
rect 1807 -806 1841 -430
rect 1903 -806 1937 -430
rect 1999 -806 2033 -430
rect 2095 -806 2129 -430
rect 2191 -806 2225 -430
rect 2287 -806 2321 -430
rect 2383 -806 2417 -430
rect 2479 -806 2513 -430
rect 2575 -806 2609 -430
rect 2671 -806 2705 -430
rect 2767 -806 2801 -430
rect 2863 -806 2897 -430
rect 2959 -806 2993 -430
rect 3055 -806 3089 -430
rect 3151 -806 3185 -430
rect 3247 -806 3281 -430
rect 3343 -806 3377 -430
rect 3439 -806 3473 -430
rect 3535 -806 3569 -430
rect 3631 -806 3665 -430
rect 3727 -806 3761 -430
rect 3823 -806 3857 -430
rect -3809 -890 -3775 -856
rect -3617 -890 -3583 -856
rect -3425 -890 -3391 -856
rect -3233 -890 -3199 -856
rect -3041 -890 -3007 -856
rect -2849 -890 -2815 -856
rect -2657 -890 -2623 -856
rect -2465 -890 -2431 -856
rect -2273 -890 -2239 -856
rect -2081 -890 -2047 -856
rect -1889 -890 -1855 -856
rect -1697 -890 -1663 -856
rect -1505 -890 -1471 -856
rect -1313 -890 -1279 -856
rect -1121 -890 -1087 -856
rect -929 -890 -895 -856
rect -737 -890 -703 -856
rect -545 -890 -511 -856
rect -353 -890 -319 -856
rect -161 -890 -127 -856
rect 31 -890 65 -856
rect 223 -890 257 -856
rect 415 -890 449 -856
rect 607 -890 641 -856
rect 799 -890 833 -856
rect 991 -890 1025 -856
rect 1183 -890 1217 -856
rect 1375 -890 1409 -856
rect 1567 -890 1601 -856
rect 1759 -890 1793 -856
rect 1951 -890 1985 -856
rect 2143 -890 2177 -856
rect 2335 -890 2369 -856
rect 2527 -890 2561 -856
rect 2719 -890 2753 -856
rect 2911 -890 2945 -856
rect 3103 -890 3137 -856
rect 3295 -890 3329 -856
rect 3487 -890 3521 -856
rect 3679 -890 3713 -856
<< metal1 >>
rect -3725 890 -3667 896
rect -3725 856 -3713 890
rect -3679 856 -3667 890
rect -3725 850 -3667 856
rect -3533 890 -3475 896
rect -3533 856 -3521 890
rect -3487 856 -3475 890
rect -3533 850 -3475 856
rect -3341 890 -3283 896
rect -3341 856 -3329 890
rect -3295 856 -3283 890
rect -3341 850 -3283 856
rect -3149 890 -3091 896
rect -3149 856 -3137 890
rect -3103 856 -3091 890
rect -3149 850 -3091 856
rect -2957 890 -2899 896
rect -2957 856 -2945 890
rect -2911 856 -2899 890
rect -2957 850 -2899 856
rect -2765 890 -2707 896
rect -2765 856 -2753 890
rect -2719 856 -2707 890
rect -2765 850 -2707 856
rect -2573 890 -2515 896
rect -2573 856 -2561 890
rect -2527 856 -2515 890
rect -2573 850 -2515 856
rect -2381 890 -2323 896
rect -2381 856 -2369 890
rect -2335 856 -2323 890
rect -2381 850 -2323 856
rect -2189 890 -2131 896
rect -2189 856 -2177 890
rect -2143 856 -2131 890
rect -2189 850 -2131 856
rect -1997 890 -1939 896
rect -1997 856 -1985 890
rect -1951 856 -1939 890
rect -1997 850 -1939 856
rect -1805 890 -1747 896
rect -1805 856 -1793 890
rect -1759 856 -1747 890
rect -1805 850 -1747 856
rect -1613 890 -1555 896
rect -1613 856 -1601 890
rect -1567 856 -1555 890
rect -1613 850 -1555 856
rect -1421 890 -1363 896
rect -1421 856 -1409 890
rect -1375 856 -1363 890
rect -1421 850 -1363 856
rect -1229 890 -1171 896
rect -1229 856 -1217 890
rect -1183 856 -1171 890
rect -1229 850 -1171 856
rect -1037 890 -979 896
rect -1037 856 -1025 890
rect -991 856 -979 890
rect -1037 850 -979 856
rect -845 890 -787 896
rect -845 856 -833 890
rect -799 856 -787 890
rect -845 850 -787 856
rect -653 890 -595 896
rect -653 856 -641 890
rect -607 856 -595 890
rect -653 850 -595 856
rect -461 890 -403 896
rect -461 856 -449 890
rect -415 856 -403 890
rect -461 850 -403 856
rect -269 890 -211 896
rect -269 856 -257 890
rect -223 856 -211 890
rect -269 850 -211 856
rect -77 890 -19 896
rect -77 856 -65 890
rect -31 856 -19 890
rect -77 850 -19 856
rect 115 890 173 896
rect 115 856 127 890
rect 161 856 173 890
rect 115 850 173 856
rect 307 890 365 896
rect 307 856 319 890
rect 353 856 365 890
rect 307 850 365 856
rect 499 890 557 896
rect 499 856 511 890
rect 545 856 557 890
rect 499 850 557 856
rect 691 890 749 896
rect 691 856 703 890
rect 737 856 749 890
rect 691 850 749 856
rect 883 890 941 896
rect 883 856 895 890
rect 929 856 941 890
rect 883 850 941 856
rect 1075 890 1133 896
rect 1075 856 1087 890
rect 1121 856 1133 890
rect 1075 850 1133 856
rect 1267 890 1325 896
rect 1267 856 1279 890
rect 1313 856 1325 890
rect 1267 850 1325 856
rect 1459 890 1517 896
rect 1459 856 1471 890
rect 1505 856 1517 890
rect 1459 850 1517 856
rect 1651 890 1709 896
rect 1651 856 1663 890
rect 1697 856 1709 890
rect 1651 850 1709 856
rect 1843 890 1901 896
rect 1843 856 1855 890
rect 1889 856 1901 890
rect 1843 850 1901 856
rect 2035 890 2093 896
rect 2035 856 2047 890
rect 2081 856 2093 890
rect 2035 850 2093 856
rect 2227 890 2285 896
rect 2227 856 2239 890
rect 2273 856 2285 890
rect 2227 850 2285 856
rect 2419 890 2477 896
rect 2419 856 2431 890
rect 2465 856 2477 890
rect 2419 850 2477 856
rect 2611 890 2669 896
rect 2611 856 2623 890
rect 2657 856 2669 890
rect 2611 850 2669 856
rect 2803 890 2861 896
rect 2803 856 2815 890
rect 2849 856 2861 890
rect 2803 850 2861 856
rect 2995 890 3053 896
rect 2995 856 3007 890
rect 3041 856 3053 890
rect 2995 850 3053 856
rect 3187 890 3245 896
rect 3187 856 3199 890
rect 3233 856 3245 890
rect 3187 850 3245 856
rect 3379 890 3437 896
rect 3379 856 3391 890
rect 3425 856 3437 890
rect 3379 850 3437 856
rect 3571 890 3629 896
rect 3571 856 3583 890
rect 3617 856 3629 890
rect 3571 850 3629 856
rect 3763 890 3821 896
rect 3763 856 3775 890
rect 3809 856 3821 890
rect 3763 850 3821 856
rect -3863 806 -3817 818
rect -3863 430 -3857 806
rect -3823 430 -3817 806
rect -3863 418 -3817 430
rect -3767 806 -3721 818
rect -3767 430 -3761 806
rect -3727 430 -3721 806
rect -3767 418 -3721 430
rect -3671 806 -3625 818
rect -3671 430 -3665 806
rect -3631 430 -3625 806
rect -3671 418 -3625 430
rect -3575 806 -3529 818
rect -3575 430 -3569 806
rect -3535 430 -3529 806
rect -3575 418 -3529 430
rect -3479 806 -3433 818
rect -3479 430 -3473 806
rect -3439 430 -3433 806
rect -3479 418 -3433 430
rect -3383 806 -3337 818
rect -3383 430 -3377 806
rect -3343 430 -3337 806
rect -3383 418 -3337 430
rect -3287 806 -3241 818
rect -3287 430 -3281 806
rect -3247 430 -3241 806
rect -3287 418 -3241 430
rect -3191 806 -3145 818
rect -3191 430 -3185 806
rect -3151 430 -3145 806
rect -3191 418 -3145 430
rect -3095 806 -3049 818
rect -3095 430 -3089 806
rect -3055 430 -3049 806
rect -3095 418 -3049 430
rect -2999 806 -2953 818
rect -2999 430 -2993 806
rect -2959 430 -2953 806
rect -2999 418 -2953 430
rect -2903 806 -2857 818
rect -2903 430 -2897 806
rect -2863 430 -2857 806
rect -2903 418 -2857 430
rect -2807 806 -2761 818
rect -2807 430 -2801 806
rect -2767 430 -2761 806
rect -2807 418 -2761 430
rect -2711 806 -2665 818
rect -2711 430 -2705 806
rect -2671 430 -2665 806
rect -2711 418 -2665 430
rect -2615 806 -2569 818
rect -2615 430 -2609 806
rect -2575 430 -2569 806
rect -2615 418 -2569 430
rect -2519 806 -2473 818
rect -2519 430 -2513 806
rect -2479 430 -2473 806
rect -2519 418 -2473 430
rect -2423 806 -2377 818
rect -2423 430 -2417 806
rect -2383 430 -2377 806
rect -2423 418 -2377 430
rect -2327 806 -2281 818
rect -2327 430 -2321 806
rect -2287 430 -2281 806
rect -2327 418 -2281 430
rect -2231 806 -2185 818
rect -2231 430 -2225 806
rect -2191 430 -2185 806
rect -2231 418 -2185 430
rect -2135 806 -2089 818
rect -2135 430 -2129 806
rect -2095 430 -2089 806
rect -2135 418 -2089 430
rect -2039 806 -1993 818
rect -2039 430 -2033 806
rect -1999 430 -1993 806
rect -2039 418 -1993 430
rect -1943 806 -1897 818
rect -1943 430 -1937 806
rect -1903 430 -1897 806
rect -1943 418 -1897 430
rect -1847 806 -1801 818
rect -1847 430 -1841 806
rect -1807 430 -1801 806
rect -1847 418 -1801 430
rect -1751 806 -1705 818
rect -1751 430 -1745 806
rect -1711 430 -1705 806
rect -1751 418 -1705 430
rect -1655 806 -1609 818
rect -1655 430 -1649 806
rect -1615 430 -1609 806
rect -1655 418 -1609 430
rect -1559 806 -1513 818
rect -1559 430 -1553 806
rect -1519 430 -1513 806
rect -1559 418 -1513 430
rect -1463 806 -1417 818
rect -1463 430 -1457 806
rect -1423 430 -1417 806
rect -1463 418 -1417 430
rect -1367 806 -1321 818
rect -1367 430 -1361 806
rect -1327 430 -1321 806
rect -1367 418 -1321 430
rect -1271 806 -1225 818
rect -1271 430 -1265 806
rect -1231 430 -1225 806
rect -1271 418 -1225 430
rect -1175 806 -1129 818
rect -1175 430 -1169 806
rect -1135 430 -1129 806
rect -1175 418 -1129 430
rect -1079 806 -1033 818
rect -1079 430 -1073 806
rect -1039 430 -1033 806
rect -1079 418 -1033 430
rect -983 806 -937 818
rect -983 430 -977 806
rect -943 430 -937 806
rect -983 418 -937 430
rect -887 806 -841 818
rect -887 430 -881 806
rect -847 430 -841 806
rect -887 418 -841 430
rect -791 806 -745 818
rect -791 430 -785 806
rect -751 430 -745 806
rect -791 418 -745 430
rect -695 806 -649 818
rect -695 430 -689 806
rect -655 430 -649 806
rect -695 418 -649 430
rect -599 806 -553 818
rect -599 430 -593 806
rect -559 430 -553 806
rect -599 418 -553 430
rect -503 806 -457 818
rect -503 430 -497 806
rect -463 430 -457 806
rect -503 418 -457 430
rect -407 806 -361 818
rect -407 430 -401 806
rect -367 430 -361 806
rect -407 418 -361 430
rect -311 806 -265 818
rect -311 430 -305 806
rect -271 430 -265 806
rect -311 418 -265 430
rect -215 806 -169 818
rect -215 430 -209 806
rect -175 430 -169 806
rect -215 418 -169 430
rect -119 806 -73 818
rect -119 430 -113 806
rect -79 430 -73 806
rect -119 418 -73 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 73 806 119 818
rect 73 430 79 806
rect 113 430 119 806
rect 73 418 119 430
rect 169 806 215 818
rect 169 430 175 806
rect 209 430 215 806
rect 169 418 215 430
rect 265 806 311 818
rect 265 430 271 806
rect 305 430 311 806
rect 265 418 311 430
rect 361 806 407 818
rect 361 430 367 806
rect 401 430 407 806
rect 361 418 407 430
rect 457 806 503 818
rect 457 430 463 806
rect 497 430 503 806
rect 457 418 503 430
rect 553 806 599 818
rect 553 430 559 806
rect 593 430 599 806
rect 553 418 599 430
rect 649 806 695 818
rect 649 430 655 806
rect 689 430 695 806
rect 649 418 695 430
rect 745 806 791 818
rect 745 430 751 806
rect 785 430 791 806
rect 745 418 791 430
rect 841 806 887 818
rect 841 430 847 806
rect 881 430 887 806
rect 841 418 887 430
rect 937 806 983 818
rect 937 430 943 806
rect 977 430 983 806
rect 937 418 983 430
rect 1033 806 1079 818
rect 1033 430 1039 806
rect 1073 430 1079 806
rect 1033 418 1079 430
rect 1129 806 1175 818
rect 1129 430 1135 806
rect 1169 430 1175 806
rect 1129 418 1175 430
rect 1225 806 1271 818
rect 1225 430 1231 806
rect 1265 430 1271 806
rect 1225 418 1271 430
rect 1321 806 1367 818
rect 1321 430 1327 806
rect 1361 430 1367 806
rect 1321 418 1367 430
rect 1417 806 1463 818
rect 1417 430 1423 806
rect 1457 430 1463 806
rect 1417 418 1463 430
rect 1513 806 1559 818
rect 1513 430 1519 806
rect 1553 430 1559 806
rect 1513 418 1559 430
rect 1609 806 1655 818
rect 1609 430 1615 806
rect 1649 430 1655 806
rect 1609 418 1655 430
rect 1705 806 1751 818
rect 1705 430 1711 806
rect 1745 430 1751 806
rect 1705 418 1751 430
rect 1801 806 1847 818
rect 1801 430 1807 806
rect 1841 430 1847 806
rect 1801 418 1847 430
rect 1897 806 1943 818
rect 1897 430 1903 806
rect 1937 430 1943 806
rect 1897 418 1943 430
rect 1993 806 2039 818
rect 1993 430 1999 806
rect 2033 430 2039 806
rect 1993 418 2039 430
rect 2089 806 2135 818
rect 2089 430 2095 806
rect 2129 430 2135 806
rect 2089 418 2135 430
rect 2185 806 2231 818
rect 2185 430 2191 806
rect 2225 430 2231 806
rect 2185 418 2231 430
rect 2281 806 2327 818
rect 2281 430 2287 806
rect 2321 430 2327 806
rect 2281 418 2327 430
rect 2377 806 2423 818
rect 2377 430 2383 806
rect 2417 430 2423 806
rect 2377 418 2423 430
rect 2473 806 2519 818
rect 2473 430 2479 806
rect 2513 430 2519 806
rect 2473 418 2519 430
rect 2569 806 2615 818
rect 2569 430 2575 806
rect 2609 430 2615 806
rect 2569 418 2615 430
rect 2665 806 2711 818
rect 2665 430 2671 806
rect 2705 430 2711 806
rect 2665 418 2711 430
rect 2761 806 2807 818
rect 2761 430 2767 806
rect 2801 430 2807 806
rect 2761 418 2807 430
rect 2857 806 2903 818
rect 2857 430 2863 806
rect 2897 430 2903 806
rect 2857 418 2903 430
rect 2953 806 2999 818
rect 2953 430 2959 806
rect 2993 430 2999 806
rect 2953 418 2999 430
rect 3049 806 3095 818
rect 3049 430 3055 806
rect 3089 430 3095 806
rect 3049 418 3095 430
rect 3145 806 3191 818
rect 3145 430 3151 806
rect 3185 430 3191 806
rect 3145 418 3191 430
rect 3241 806 3287 818
rect 3241 430 3247 806
rect 3281 430 3287 806
rect 3241 418 3287 430
rect 3337 806 3383 818
rect 3337 430 3343 806
rect 3377 430 3383 806
rect 3337 418 3383 430
rect 3433 806 3479 818
rect 3433 430 3439 806
rect 3473 430 3479 806
rect 3433 418 3479 430
rect 3529 806 3575 818
rect 3529 430 3535 806
rect 3569 430 3575 806
rect 3529 418 3575 430
rect 3625 806 3671 818
rect 3625 430 3631 806
rect 3665 430 3671 806
rect 3625 418 3671 430
rect 3721 806 3767 818
rect 3721 430 3727 806
rect 3761 430 3767 806
rect 3721 418 3767 430
rect 3817 806 3863 818
rect 3817 430 3823 806
rect 3857 430 3863 806
rect 3817 418 3863 430
rect -3821 380 -3763 386
rect -3821 346 -3809 380
rect -3775 346 -3763 380
rect -3821 340 -3763 346
rect -3629 380 -3571 386
rect -3629 346 -3617 380
rect -3583 346 -3571 380
rect -3629 340 -3571 346
rect -3437 380 -3379 386
rect -3437 346 -3425 380
rect -3391 346 -3379 380
rect -3437 340 -3379 346
rect -3245 380 -3187 386
rect -3245 346 -3233 380
rect -3199 346 -3187 380
rect -3245 340 -3187 346
rect -3053 380 -2995 386
rect -3053 346 -3041 380
rect -3007 346 -2995 380
rect -3053 340 -2995 346
rect -2861 380 -2803 386
rect -2861 346 -2849 380
rect -2815 346 -2803 380
rect -2861 340 -2803 346
rect -2669 380 -2611 386
rect -2669 346 -2657 380
rect -2623 346 -2611 380
rect -2669 340 -2611 346
rect -2477 380 -2419 386
rect -2477 346 -2465 380
rect -2431 346 -2419 380
rect -2477 340 -2419 346
rect -2285 380 -2227 386
rect -2285 346 -2273 380
rect -2239 346 -2227 380
rect -2285 340 -2227 346
rect -2093 380 -2035 386
rect -2093 346 -2081 380
rect -2047 346 -2035 380
rect -2093 340 -2035 346
rect -1901 380 -1843 386
rect -1901 346 -1889 380
rect -1855 346 -1843 380
rect -1901 340 -1843 346
rect -1709 380 -1651 386
rect -1709 346 -1697 380
rect -1663 346 -1651 380
rect -1709 340 -1651 346
rect -1517 380 -1459 386
rect -1517 346 -1505 380
rect -1471 346 -1459 380
rect -1517 340 -1459 346
rect -1325 380 -1267 386
rect -1325 346 -1313 380
rect -1279 346 -1267 380
rect -1325 340 -1267 346
rect -1133 380 -1075 386
rect -1133 346 -1121 380
rect -1087 346 -1075 380
rect -1133 340 -1075 346
rect -941 380 -883 386
rect -941 346 -929 380
rect -895 346 -883 380
rect -941 340 -883 346
rect -749 380 -691 386
rect -749 346 -737 380
rect -703 346 -691 380
rect -749 340 -691 346
rect -557 380 -499 386
rect -557 346 -545 380
rect -511 346 -499 380
rect -557 340 -499 346
rect -365 380 -307 386
rect -365 346 -353 380
rect -319 346 -307 380
rect -365 340 -307 346
rect -173 380 -115 386
rect -173 346 -161 380
rect -127 346 -115 380
rect -173 340 -115 346
rect 19 380 77 386
rect 19 346 31 380
rect 65 346 77 380
rect 19 340 77 346
rect 211 380 269 386
rect 211 346 223 380
rect 257 346 269 380
rect 211 340 269 346
rect 403 380 461 386
rect 403 346 415 380
rect 449 346 461 380
rect 403 340 461 346
rect 595 380 653 386
rect 595 346 607 380
rect 641 346 653 380
rect 595 340 653 346
rect 787 380 845 386
rect 787 346 799 380
rect 833 346 845 380
rect 787 340 845 346
rect 979 380 1037 386
rect 979 346 991 380
rect 1025 346 1037 380
rect 979 340 1037 346
rect 1171 380 1229 386
rect 1171 346 1183 380
rect 1217 346 1229 380
rect 1171 340 1229 346
rect 1363 380 1421 386
rect 1363 346 1375 380
rect 1409 346 1421 380
rect 1363 340 1421 346
rect 1555 380 1613 386
rect 1555 346 1567 380
rect 1601 346 1613 380
rect 1555 340 1613 346
rect 1747 380 1805 386
rect 1747 346 1759 380
rect 1793 346 1805 380
rect 1747 340 1805 346
rect 1939 380 1997 386
rect 1939 346 1951 380
rect 1985 346 1997 380
rect 1939 340 1997 346
rect 2131 380 2189 386
rect 2131 346 2143 380
rect 2177 346 2189 380
rect 2131 340 2189 346
rect 2323 380 2381 386
rect 2323 346 2335 380
rect 2369 346 2381 380
rect 2323 340 2381 346
rect 2515 380 2573 386
rect 2515 346 2527 380
rect 2561 346 2573 380
rect 2515 340 2573 346
rect 2707 380 2765 386
rect 2707 346 2719 380
rect 2753 346 2765 380
rect 2707 340 2765 346
rect 2899 380 2957 386
rect 2899 346 2911 380
rect 2945 346 2957 380
rect 2899 340 2957 346
rect 3091 380 3149 386
rect 3091 346 3103 380
rect 3137 346 3149 380
rect 3091 340 3149 346
rect 3283 380 3341 386
rect 3283 346 3295 380
rect 3329 346 3341 380
rect 3283 340 3341 346
rect 3475 380 3533 386
rect 3475 346 3487 380
rect 3521 346 3533 380
rect 3475 340 3533 346
rect 3667 380 3725 386
rect 3667 346 3679 380
rect 3713 346 3725 380
rect 3667 340 3725 346
rect -3821 272 -3763 278
rect -3821 238 -3809 272
rect -3775 238 -3763 272
rect -3821 232 -3763 238
rect -3629 272 -3571 278
rect -3629 238 -3617 272
rect -3583 238 -3571 272
rect -3629 232 -3571 238
rect -3437 272 -3379 278
rect -3437 238 -3425 272
rect -3391 238 -3379 272
rect -3437 232 -3379 238
rect -3245 272 -3187 278
rect -3245 238 -3233 272
rect -3199 238 -3187 272
rect -3245 232 -3187 238
rect -3053 272 -2995 278
rect -3053 238 -3041 272
rect -3007 238 -2995 272
rect -3053 232 -2995 238
rect -2861 272 -2803 278
rect -2861 238 -2849 272
rect -2815 238 -2803 272
rect -2861 232 -2803 238
rect -2669 272 -2611 278
rect -2669 238 -2657 272
rect -2623 238 -2611 272
rect -2669 232 -2611 238
rect -2477 272 -2419 278
rect -2477 238 -2465 272
rect -2431 238 -2419 272
rect -2477 232 -2419 238
rect -2285 272 -2227 278
rect -2285 238 -2273 272
rect -2239 238 -2227 272
rect -2285 232 -2227 238
rect -2093 272 -2035 278
rect -2093 238 -2081 272
rect -2047 238 -2035 272
rect -2093 232 -2035 238
rect -1901 272 -1843 278
rect -1901 238 -1889 272
rect -1855 238 -1843 272
rect -1901 232 -1843 238
rect -1709 272 -1651 278
rect -1709 238 -1697 272
rect -1663 238 -1651 272
rect -1709 232 -1651 238
rect -1517 272 -1459 278
rect -1517 238 -1505 272
rect -1471 238 -1459 272
rect -1517 232 -1459 238
rect -1325 272 -1267 278
rect -1325 238 -1313 272
rect -1279 238 -1267 272
rect -1325 232 -1267 238
rect -1133 272 -1075 278
rect -1133 238 -1121 272
rect -1087 238 -1075 272
rect -1133 232 -1075 238
rect -941 272 -883 278
rect -941 238 -929 272
rect -895 238 -883 272
rect -941 232 -883 238
rect -749 272 -691 278
rect -749 238 -737 272
rect -703 238 -691 272
rect -749 232 -691 238
rect -557 272 -499 278
rect -557 238 -545 272
rect -511 238 -499 272
rect -557 232 -499 238
rect -365 272 -307 278
rect -365 238 -353 272
rect -319 238 -307 272
rect -365 232 -307 238
rect -173 272 -115 278
rect -173 238 -161 272
rect -127 238 -115 272
rect -173 232 -115 238
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect 211 272 269 278
rect 211 238 223 272
rect 257 238 269 272
rect 211 232 269 238
rect 403 272 461 278
rect 403 238 415 272
rect 449 238 461 272
rect 403 232 461 238
rect 595 272 653 278
rect 595 238 607 272
rect 641 238 653 272
rect 595 232 653 238
rect 787 272 845 278
rect 787 238 799 272
rect 833 238 845 272
rect 787 232 845 238
rect 979 272 1037 278
rect 979 238 991 272
rect 1025 238 1037 272
rect 979 232 1037 238
rect 1171 272 1229 278
rect 1171 238 1183 272
rect 1217 238 1229 272
rect 1171 232 1229 238
rect 1363 272 1421 278
rect 1363 238 1375 272
rect 1409 238 1421 272
rect 1363 232 1421 238
rect 1555 272 1613 278
rect 1555 238 1567 272
rect 1601 238 1613 272
rect 1555 232 1613 238
rect 1747 272 1805 278
rect 1747 238 1759 272
rect 1793 238 1805 272
rect 1747 232 1805 238
rect 1939 272 1997 278
rect 1939 238 1951 272
rect 1985 238 1997 272
rect 1939 232 1997 238
rect 2131 272 2189 278
rect 2131 238 2143 272
rect 2177 238 2189 272
rect 2131 232 2189 238
rect 2323 272 2381 278
rect 2323 238 2335 272
rect 2369 238 2381 272
rect 2323 232 2381 238
rect 2515 272 2573 278
rect 2515 238 2527 272
rect 2561 238 2573 272
rect 2515 232 2573 238
rect 2707 272 2765 278
rect 2707 238 2719 272
rect 2753 238 2765 272
rect 2707 232 2765 238
rect 2899 272 2957 278
rect 2899 238 2911 272
rect 2945 238 2957 272
rect 2899 232 2957 238
rect 3091 272 3149 278
rect 3091 238 3103 272
rect 3137 238 3149 272
rect 3091 232 3149 238
rect 3283 272 3341 278
rect 3283 238 3295 272
rect 3329 238 3341 272
rect 3283 232 3341 238
rect 3475 272 3533 278
rect 3475 238 3487 272
rect 3521 238 3533 272
rect 3475 232 3533 238
rect 3667 272 3725 278
rect 3667 238 3679 272
rect 3713 238 3725 272
rect 3667 232 3725 238
rect -3863 188 -3817 200
rect -3863 -188 -3857 188
rect -3823 -188 -3817 188
rect -3863 -200 -3817 -188
rect -3767 188 -3721 200
rect -3767 -188 -3761 188
rect -3727 -188 -3721 188
rect -3767 -200 -3721 -188
rect -3671 188 -3625 200
rect -3671 -188 -3665 188
rect -3631 -188 -3625 188
rect -3671 -200 -3625 -188
rect -3575 188 -3529 200
rect -3575 -188 -3569 188
rect -3535 -188 -3529 188
rect -3575 -200 -3529 -188
rect -3479 188 -3433 200
rect -3479 -188 -3473 188
rect -3439 -188 -3433 188
rect -3479 -200 -3433 -188
rect -3383 188 -3337 200
rect -3383 -188 -3377 188
rect -3343 -188 -3337 188
rect -3383 -200 -3337 -188
rect -3287 188 -3241 200
rect -3287 -188 -3281 188
rect -3247 -188 -3241 188
rect -3287 -200 -3241 -188
rect -3191 188 -3145 200
rect -3191 -188 -3185 188
rect -3151 -188 -3145 188
rect -3191 -200 -3145 -188
rect -3095 188 -3049 200
rect -3095 -188 -3089 188
rect -3055 -188 -3049 188
rect -3095 -200 -3049 -188
rect -2999 188 -2953 200
rect -2999 -188 -2993 188
rect -2959 -188 -2953 188
rect -2999 -200 -2953 -188
rect -2903 188 -2857 200
rect -2903 -188 -2897 188
rect -2863 -188 -2857 188
rect -2903 -200 -2857 -188
rect -2807 188 -2761 200
rect -2807 -188 -2801 188
rect -2767 -188 -2761 188
rect -2807 -200 -2761 -188
rect -2711 188 -2665 200
rect -2711 -188 -2705 188
rect -2671 -188 -2665 188
rect -2711 -200 -2665 -188
rect -2615 188 -2569 200
rect -2615 -188 -2609 188
rect -2575 -188 -2569 188
rect -2615 -200 -2569 -188
rect -2519 188 -2473 200
rect -2519 -188 -2513 188
rect -2479 -188 -2473 188
rect -2519 -200 -2473 -188
rect -2423 188 -2377 200
rect -2423 -188 -2417 188
rect -2383 -188 -2377 188
rect -2423 -200 -2377 -188
rect -2327 188 -2281 200
rect -2327 -188 -2321 188
rect -2287 -188 -2281 188
rect -2327 -200 -2281 -188
rect -2231 188 -2185 200
rect -2231 -188 -2225 188
rect -2191 -188 -2185 188
rect -2231 -200 -2185 -188
rect -2135 188 -2089 200
rect -2135 -188 -2129 188
rect -2095 -188 -2089 188
rect -2135 -200 -2089 -188
rect -2039 188 -1993 200
rect -2039 -188 -2033 188
rect -1999 -188 -1993 188
rect -2039 -200 -1993 -188
rect -1943 188 -1897 200
rect -1943 -188 -1937 188
rect -1903 -188 -1897 188
rect -1943 -200 -1897 -188
rect -1847 188 -1801 200
rect -1847 -188 -1841 188
rect -1807 -188 -1801 188
rect -1847 -200 -1801 -188
rect -1751 188 -1705 200
rect -1751 -188 -1745 188
rect -1711 -188 -1705 188
rect -1751 -200 -1705 -188
rect -1655 188 -1609 200
rect -1655 -188 -1649 188
rect -1615 -188 -1609 188
rect -1655 -200 -1609 -188
rect -1559 188 -1513 200
rect -1559 -188 -1553 188
rect -1519 -188 -1513 188
rect -1559 -200 -1513 -188
rect -1463 188 -1417 200
rect -1463 -188 -1457 188
rect -1423 -188 -1417 188
rect -1463 -200 -1417 -188
rect -1367 188 -1321 200
rect -1367 -188 -1361 188
rect -1327 -188 -1321 188
rect -1367 -200 -1321 -188
rect -1271 188 -1225 200
rect -1271 -188 -1265 188
rect -1231 -188 -1225 188
rect -1271 -200 -1225 -188
rect -1175 188 -1129 200
rect -1175 -188 -1169 188
rect -1135 -188 -1129 188
rect -1175 -200 -1129 -188
rect -1079 188 -1033 200
rect -1079 -188 -1073 188
rect -1039 -188 -1033 188
rect -1079 -200 -1033 -188
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect 1033 188 1079 200
rect 1033 -188 1039 188
rect 1073 -188 1079 188
rect 1033 -200 1079 -188
rect 1129 188 1175 200
rect 1129 -188 1135 188
rect 1169 -188 1175 188
rect 1129 -200 1175 -188
rect 1225 188 1271 200
rect 1225 -188 1231 188
rect 1265 -188 1271 188
rect 1225 -200 1271 -188
rect 1321 188 1367 200
rect 1321 -188 1327 188
rect 1361 -188 1367 188
rect 1321 -200 1367 -188
rect 1417 188 1463 200
rect 1417 -188 1423 188
rect 1457 -188 1463 188
rect 1417 -200 1463 -188
rect 1513 188 1559 200
rect 1513 -188 1519 188
rect 1553 -188 1559 188
rect 1513 -200 1559 -188
rect 1609 188 1655 200
rect 1609 -188 1615 188
rect 1649 -188 1655 188
rect 1609 -200 1655 -188
rect 1705 188 1751 200
rect 1705 -188 1711 188
rect 1745 -188 1751 188
rect 1705 -200 1751 -188
rect 1801 188 1847 200
rect 1801 -188 1807 188
rect 1841 -188 1847 188
rect 1801 -200 1847 -188
rect 1897 188 1943 200
rect 1897 -188 1903 188
rect 1937 -188 1943 188
rect 1897 -200 1943 -188
rect 1993 188 2039 200
rect 1993 -188 1999 188
rect 2033 -188 2039 188
rect 1993 -200 2039 -188
rect 2089 188 2135 200
rect 2089 -188 2095 188
rect 2129 -188 2135 188
rect 2089 -200 2135 -188
rect 2185 188 2231 200
rect 2185 -188 2191 188
rect 2225 -188 2231 188
rect 2185 -200 2231 -188
rect 2281 188 2327 200
rect 2281 -188 2287 188
rect 2321 -188 2327 188
rect 2281 -200 2327 -188
rect 2377 188 2423 200
rect 2377 -188 2383 188
rect 2417 -188 2423 188
rect 2377 -200 2423 -188
rect 2473 188 2519 200
rect 2473 -188 2479 188
rect 2513 -188 2519 188
rect 2473 -200 2519 -188
rect 2569 188 2615 200
rect 2569 -188 2575 188
rect 2609 -188 2615 188
rect 2569 -200 2615 -188
rect 2665 188 2711 200
rect 2665 -188 2671 188
rect 2705 -188 2711 188
rect 2665 -200 2711 -188
rect 2761 188 2807 200
rect 2761 -188 2767 188
rect 2801 -188 2807 188
rect 2761 -200 2807 -188
rect 2857 188 2903 200
rect 2857 -188 2863 188
rect 2897 -188 2903 188
rect 2857 -200 2903 -188
rect 2953 188 2999 200
rect 2953 -188 2959 188
rect 2993 -188 2999 188
rect 2953 -200 2999 -188
rect 3049 188 3095 200
rect 3049 -188 3055 188
rect 3089 -188 3095 188
rect 3049 -200 3095 -188
rect 3145 188 3191 200
rect 3145 -188 3151 188
rect 3185 -188 3191 188
rect 3145 -200 3191 -188
rect 3241 188 3287 200
rect 3241 -188 3247 188
rect 3281 -188 3287 188
rect 3241 -200 3287 -188
rect 3337 188 3383 200
rect 3337 -188 3343 188
rect 3377 -188 3383 188
rect 3337 -200 3383 -188
rect 3433 188 3479 200
rect 3433 -188 3439 188
rect 3473 -188 3479 188
rect 3433 -200 3479 -188
rect 3529 188 3575 200
rect 3529 -188 3535 188
rect 3569 -188 3575 188
rect 3529 -200 3575 -188
rect 3625 188 3671 200
rect 3625 -188 3631 188
rect 3665 -188 3671 188
rect 3625 -200 3671 -188
rect 3721 188 3767 200
rect 3721 -188 3727 188
rect 3761 -188 3767 188
rect 3721 -200 3767 -188
rect 3817 188 3863 200
rect 3817 -188 3823 188
rect 3857 -188 3863 188
rect 3817 -200 3863 -188
rect -3725 -238 -3667 -232
rect -3725 -272 -3713 -238
rect -3679 -272 -3667 -238
rect -3725 -278 -3667 -272
rect -3533 -238 -3475 -232
rect -3533 -272 -3521 -238
rect -3487 -272 -3475 -238
rect -3533 -278 -3475 -272
rect -3341 -238 -3283 -232
rect -3341 -272 -3329 -238
rect -3295 -272 -3283 -238
rect -3341 -278 -3283 -272
rect -3149 -238 -3091 -232
rect -3149 -272 -3137 -238
rect -3103 -272 -3091 -238
rect -3149 -278 -3091 -272
rect -2957 -238 -2899 -232
rect -2957 -272 -2945 -238
rect -2911 -272 -2899 -238
rect -2957 -278 -2899 -272
rect -2765 -238 -2707 -232
rect -2765 -272 -2753 -238
rect -2719 -272 -2707 -238
rect -2765 -278 -2707 -272
rect -2573 -238 -2515 -232
rect -2573 -272 -2561 -238
rect -2527 -272 -2515 -238
rect -2573 -278 -2515 -272
rect -2381 -238 -2323 -232
rect -2381 -272 -2369 -238
rect -2335 -272 -2323 -238
rect -2381 -278 -2323 -272
rect -2189 -238 -2131 -232
rect -2189 -272 -2177 -238
rect -2143 -272 -2131 -238
rect -2189 -278 -2131 -272
rect -1997 -238 -1939 -232
rect -1997 -272 -1985 -238
rect -1951 -272 -1939 -238
rect -1997 -278 -1939 -272
rect -1805 -238 -1747 -232
rect -1805 -272 -1793 -238
rect -1759 -272 -1747 -238
rect -1805 -278 -1747 -272
rect -1613 -238 -1555 -232
rect -1613 -272 -1601 -238
rect -1567 -272 -1555 -238
rect -1613 -278 -1555 -272
rect -1421 -238 -1363 -232
rect -1421 -272 -1409 -238
rect -1375 -272 -1363 -238
rect -1421 -278 -1363 -272
rect -1229 -238 -1171 -232
rect -1229 -272 -1217 -238
rect -1183 -272 -1171 -238
rect -1229 -278 -1171 -272
rect -1037 -238 -979 -232
rect -1037 -272 -1025 -238
rect -991 -272 -979 -238
rect -1037 -278 -979 -272
rect -845 -238 -787 -232
rect -845 -272 -833 -238
rect -799 -272 -787 -238
rect -845 -278 -787 -272
rect -653 -238 -595 -232
rect -653 -272 -641 -238
rect -607 -272 -595 -238
rect -653 -278 -595 -272
rect -461 -238 -403 -232
rect -461 -272 -449 -238
rect -415 -272 -403 -238
rect -461 -278 -403 -272
rect -269 -238 -211 -232
rect -269 -272 -257 -238
rect -223 -272 -211 -238
rect -269 -278 -211 -272
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
rect 115 -238 173 -232
rect 115 -272 127 -238
rect 161 -272 173 -238
rect 115 -278 173 -272
rect 307 -238 365 -232
rect 307 -272 319 -238
rect 353 -272 365 -238
rect 307 -278 365 -272
rect 499 -238 557 -232
rect 499 -272 511 -238
rect 545 -272 557 -238
rect 499 -278 557 -272
rect 691 -238 749 -232
rect 691 -272 703 -238
rect 737 -272 749 -238
rect 691 -278 749 -272
rect 883 -238 941 -232
rect 883 -272 895 -238
rect 929 -272 941 -238
rect 883 -278 941 -272
rect 1075 -238 1133 -232
rect 1075 -272 1087 -238
rect 1121 -272 1133 -238
rect 1075 -278 1133 -272
rect 1267 -238 1325 -232
rect 1267 -272 1279 -238
rect 1313 -272 1325 -238
rect 1267 -278 1325 -272
rect 1459 -238 1517 -232
rect 1459 -272 1471 -238
rect 1505 -272 1517 -238
rect 1459 -278 1517 -272
rect 1651 -238 1709 -232
rect 1651 -272 1663 -238
rect 1697 -272 1709 -238
rect 1651 -278 1709 -272
rect 1843 -238 1901 -232
rect 1843 -272 1855 -238
rect 1889 -272 1901 -238
rect 1843 -278 1901 -272
rect 2035 -238 2093 -232
rect 2035 -272 2047 -238
rect 2081 -272 2093 -238
rect 2035 -278 2093 -272
rect 2227 -238 2285 -232
rect 2227 -272 2239 -238
rect 2273 -272 2285 -238
rect 2227 -278 2285 -272
rect 2419 -238 2477 -232
rect 2419 -272 2431 -238
rect 2465 -272 2477 -238
rect 2419 -278 2477 -272
rect 2611 -238 2669 -232
rect 2611 -272 2623 -238
rect 2657 -272 2669 -238
rect 2611 -278 2669 -272
rect 2803 -238 2861 -232
rect 2803 -272 2815 -238
rect 2849 -272 2861 -238
rect 2803 -278 2861 -272
rect 2995 -238 3053 -232
rect 2995 -272 3007 -238
rect 3041 -272 3053 -238
rect 2995 -278 3053 -272
rect 3187 -238 3245 -232
rect 3187 -272 3199 -238
rect 3233 -272 3245 -238
rect 3187 -278 3245 -272
rect 3379 -238 3437 -232
rect 3379 -272 3391 -238
rect 3425 -272 3437 -238
rect 3379 -278 3437 -272
rect 3571 -238 3629 -232
rect 3571 -272 3583 -238
rect 3617 -272 3629 -238
rect 3571 -278 3629 -272
rect 3763 -238 3821 -232
rect 3763 -272 3775 -238
rect 3809 -272 3821 -238
rect 3763 -278 3821 -272
rect -3725 -346 -3667 -340
rect -3725 -380 -3713 -346
rect -3679 -380 -3667 -346
rect -3725 -386 -3667 -380
rect -3533 -346 -3475 -340
rect -3533 -380 -3521 -346
rect -3487 -380 -3475 -346
rect -3533 -386 -3475 -380
rect -3341 -346 -3283 -340
rect -3341 -380 -3329 -346
rect -3295 -380 -3283 -346
rect -3341 -386 -3283 -380
rect -3149 -346 -3091 -340
rect -3149 -380 -3137 -346
rect -3103 -380 -3091 -346
rect -3149 -386 -3091 -380
rect -2957 -346 -2899 -340
rect -2957 -380 -2945 -346
rect -2911 -380 -2899 -346
rect -2957 -386 -2899 -380
rect -2765 -346 -2707 -340
rect -2765 -380 -2753 -346
rect -2719 -380 -2707 -346
rect -2765 -386 -2707 -380
rect -2573 -346 -2515 -340
rect -2573 -380 -2561 -346
rect -2527 -380 -2515 -346
rect -2573 -386 -2515 -380
rect -2381 -346 -2323 -340
rect -2381 -380 -2369 -346
rect -2335 -380 -2323 -346
rect -2381 -386 -2323 -380
rect -2189 -346 -2131 -340
rect -2189 -380 -2177 -346
rect -2143 -380 -2131 -346
rect -2189 -386 -2131 -380
rect -1997 -346 -1939 -340
rect -1997 -380 -1985 -346
rect -1951 -380 -1939 -346
rect -1997 -386 -1939 -380
rect -1805 -346 -1747 -340
rect -1805 -380 -1793 -346
rect -1759 -380 -1747 -346
rect -1805 -386 -1747 -380
rect -1613 -346 -1555 -340
rect -1613 -380 -1601 -346
rect -1567 -380 -1555 -346
rect -1613 -386 -1555 -380
rect -1421 -346 -1363 -340
rect -1421 -380 -1409 -346
rect -1375 -380 -1363 -346
rect -1421 -386 -1363 -380
rect -1229 -346 -1171 -340
rect -1229 -380 -1217 -346
rect -1183 -380 -1171 -346
rect -1229 -386 -1171 -380
rect -1037 -346 -979 -340
rect -1037 -380 -1025 -346
rect -991 -380 -979 -346
rect -1037 -386 -979 -380
rect -845 -346 -787 -340
rect -845 -380 -833 -346
rect -799 -380 -787 -346
rect -845 -386 -787 -380
rect -653 -346 -595 -340
rect -653 -380 -641 -346
rect -607 -380 -595 -346
rect -653 -386 -595 -380
rect -461 -346 -403 -340
rect -461 -380 -449 -346
rect -415 -380 -403 -346
rect -461 -386 -403 -380
rect -269 -346 -211 -340
rect -269 -380 -257 -346
rect -223 -380 -211 -346
rect -269 -386 -211 -380
rect -77 -346 -19 -340
rect -77 -380 -65 -346
rect -31 -380 -19 -346
rect -77 -386 -19 -380
rect 115 -346 173 -340
rect 115 -380 127 -346
rect 161 -380 173 -346
rect 115 -386 173 -380
rect 307 -346 365 -340
rect 307 -380 319 -346
rect 353 -380 365 -346
rect 307 -386 365 -380
rect 499 -346 557 -340
rect 499 -380 511 -346
rect 545 -380 557 -346
rect 499 -386 557 -380
rect 691 -346 749 -340
rect 691 -380 703 -346
rect 737 -380 749 -346
rect 691 -386 749 -380
rect 883 -346 941 -340
rect 883 -380 895 -346
rect 929 -380 941 -346
rect 883 -386 941 -380
rect 1075 -346 1133 -340
rect 1075 -380 1087 -346
rect 1121 -380 1133 -346
rect 1075 -386 1133 -380
rect 1267 -346 1325 -340
rect 1267 -380 1279 -346
rect 1313 -380 1325 -346
rect 1267 -386 1325 -380
rect 1459 -346 1517 -340
rect 1459 -380 1471 -346
rect 1505 -380 1517 -346
rect 1459 -386 1517 -380
rect 1651 -346 1709 -340
rect 1651 -380 1663 -346
rect 1697 -380 1709 -346
rect 1651 -386 1709 -380
rect 1843 -346 1901 -340
rect 1843 -380 1855 -346
rect 1889 -380 1901 -346
rect 1843 -386 1901 -380
rect 2035 -346 2093 -340
rect 2035 -380 2047 -346
rect 2081 -380 2093 -346
rect 2035 -386 2093 -380
rect 2227 -346 2285 -340
rect 2227 -380 2239 -346
rect 2273 -380 2285 -346
rect 2227 -386 2285 -380
rect 2419 -346 2477 -340
rect 2419 -380 2431 -346
rect 2465 -380 2477 -346
rect 2419 -386 2477 -380
rect 2611 -346 2669 -340
rect 2611 -380 2623 -346
rect 2657 -380 2669 -346
rect 2611 -386 2669 -380
rect 2803 -346 2861 -340
rect 2803 -380 2815 -346
rect 2849 -380 2861 -346
rect 2803 -386 2861 -380
rect 2995 -346 3053 -340
rect 2995 -380 3007 -346
rect 3041 -380 3053 -346
rect 2995 -386 3053 -380
rect 3187 -346 3245 -340
rect 3187 -380 3199 -346
rect 3233 -380 3245 -346
rect 3187 -386 3245 -380
rect 3379 -346 3437 -340
rect 3379 -380 3391 -346
rect 3425 -380 3437 -346
rect 3379 -386 3437 -380
rect 3571 -346 3629 -340
rect 3571 -380 3583 -346
rect 3617 -380 3629 -346
rect 3571 -386 3629 -380
rect 3763 -346 3821 -340
rect 3763 -380 3775 -346
rect 3809 -380 3821 -346
rect 3763 -386 3821 -380
rect -3863 -430 -3817 -418
rect -3863 -806 -3857 -430
rect -3823 -806 -3817 -430
rect -3863 -818 -3817 -806
rect -3767 -430 -3721 -418
rect -3767 -806 -3761 -430
rect -3727 -806 -3721 -430
rect -3767 -818 -3721 -806
rect -3671 -430 -3625 -418
rect -3671 -806 -3665 -430
rect -3631 -806 -3625 -430
rect -3671 -818 -3625 -806
rect -3575 -430 -3529 -418
rect -3575 -806 -3569 -430
rect -3535 -806 -3529 -430
rect -3575 -818 -3529 -806
rect -3479 -430 -3433 -418
rect -3479 -806 -3473 -430
rect -3439 -806 -3433 -430
rect -3479 -818 -3433 -806
rect -3383 -430 -3337 -418
rect -3383 -806 -3377 -430
rect -3343 -806 -3337 -430
rect -3383 -818 -3337 -806
rect -3287 -430 -3241 -418
rect -3287 -806 -3281 -430
rect -3247 -806 -3241 -430
rect -3287 -818 -3241 -806
rect -3191 -430 -3145 -418
rect -3191 -806 -3185 -430
rect -3151 -806 -3145 -430
rect -3191 -818 -3145 -806
rect -3095 -430 -3049 -418
rect -3095 -806 -3089 -430
rect -3055 -806 -3049 -430
rect -3095 -818 -3049 -806
rect -2999 -430 -2953 -418
rect -2999 -806 -2993 -430
rect -2959 -806 -2953 -430
rect -2999 -818 -2953 -806
rect -2903 -430 -2857 -418
rect -2903 -806 -2897 -430
rect -2863 -806 -2857 -430
rect -2903 -818 -2857 -806
rect -2807 -430 -2761 -418
rect -2807 -806 -2801 -430
rect -2767 -806 -2761 -430
rect -2807 -818 -2761 -806
rect -2711 -430 -2665 -418
rect -2711 -806 -2705 -430
rect -2671 -806 -2665 -430
rect -2711 -818 -2665 -806
rect -2615 -430 -2569 -418
rect -2615 -806 -2609 -430
rect -2575 -806 -2569 -430
rect -2615 -818 -2569 -806
rect -2519 -430 -2473 -418
rect -2519 -806 -2513 -430
rect -2479 -806 -2473 -430
rect -2519 -818 -2473 -806
rect -2423 -430 -2377 -418
rect -2423 -806 -2417 -430
rect -2383 -806 -2377 -430
rect -2423 -818 -2377 -806
rect -2327 -430 -2281 -418
rect -2327 -806 -2321 -430
rect -2287 -806 -2281 -430
rect -2327 -818 -2281 -806
rect -2231 -430 -2185 -418
rect -2231 -806 -2225 -430
rect -2191 -806 -2185 -430
rect -2231 -818 -2185 -806
rect -2135 -430 -2089 -418
rect -2135 -806 -2129 -430
rect -2095 -806 -2089 -430
rect -2135 -818 -2089 -806
rect -2039 -430 -1993 -418
rect -2039 -806 -2033 -430
rect -1999 -806 -1993 -430
rect -2039 -818 -1993 -806
rect -1943 -430 -1897 -418
rect -1943 -806 -1937 -430
rect -1903 -806 -1897 -430
rect -1943 -818 -1897 -806
rect -1847 -430 -1801 -418
rect -1847 -806 -1841 -430
rect -1807 -806 -1801 -430
rect -1847 -818 -1801 -806
rect -1751 -430 -1705 -418
rect -1751 -806 -1745 -430
rect -1711 -806 -1705 -430
rect -1751 -818 -1705 -806
rect -1655 -430 -1609 -418
rect -1655 -806 -1649 -430
rect -1615 -806 -1609 -430
rect -1655 -818 -1609 -806
rect -1559 -430 -1513 -418
rect -1559 -806 -1553 -430
rect -1519 -806 -1513 -430
rect -1559 -818 -1513 -806
rect -1463 -430 -1417 -418
rect -1463 -806 -1457 -430
rect -1423 -806 -1417 -430
rect -1463 -818 -1417 -806
rect -1367 -430 -1321 -418
rect -1367 -806 -1361 -430
rect -1327 -806 -1321 -430
rect -1367 -818 -1321 -806
rect -1271 -430 -1225 -418
rect -1271 -806 -1265 -430
rect -1231 -806 -1225 -430
rect -1271 -818 -1225 -806
rect -1175 -430 -1129 -418
rect -1175 -806 -1169 -430
rect -1135 -806 -1129 -430
rect -1175 -818 -1129 -806
rect -1079 -430 -1033 -418
rect -1079 -806 -1073 -430
rect -1039 -806 -1033 -430
rect -1079 -818 -1033 -806
rect -983 -430 -937 -418
rect -983 -806 -977 -430
rect -943 -806 -937 -430
rect -983 -818 -937 -806
rect -887 -430 -841 -418
rect -887 -806 -881 -430
rect -847 -806 -841 -430
rect -887 -818 -841 -806
rect -791 -430 -745 -418
rect -791 -806 -785 -430
rect -751 -806 -745 -430
rect -791 -818 -745 -806
rect -695 -430 -649 -418
rect -695 -806 -689 -430
rect -655 -806 -649 -430
rect -695 -818 -649 -806
rect -599 -430 -553 -418
rect -599 -806 -593 -430
rect -559 -806 -553 -430
rect -599 -818 -553 -806
rect -503 -430 -457 -418
rect -503 -806 -497 -430
rect -463 -806 -457 -430
rect -503 -818 -457 -806
rect -407 -430 -361 -418
rect -407 -806 -401 -430
rect -367 -806 -361 -430
rect -407 -818 -361 -806
rect -311 -430 -265 -418
rect -311 -806 -305 -430
rect -271 -806 -265 -430
rect -311 -818 -265 -806
rect -215 -430 -169 -418
rect -215 -806 -209 -430
rect -175 -806 -169 -430
rect -215 -818 -169 -806
rect -119 -430 -73 -418
rect -119 -806 -113 -430
rect -79 -806 -73 -430
rect -119 -818 -73 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 73 -430 119 -418
rect 73 -806 79 -430
rect 113 -806 119 -430
rect 73 -818 119 -806
rect 169 -430 215 -418
rect 169 -806 175 -430
rect 209 -806 215 -430
rect 169 -818 215 -806
rect 265 -430 311 -418
rect 265 -806 271 -430
rect 305 -806 311 -430
rect 265 -818 311 -806
rect 361 -430 407 -418
rect 361 -806 367 -430
rect 401 -806 407 -430
rect 361 -818 407 -806
rect 457 -430 503 -418
rect 457 -806 463 -430
rect 497 -806 503 -430
rect 457 -818 503 -806
rect 553 -430 599 -418
rect 553 -806 559 -430
rect 593 -806 599 -430
rect 553 -818 599 -806
rect 649 -430 695 -418
rect 649 -806 655 -430
rect 689 -806 695 -430
rect 649 -818 695 -806
rect 745 -430 791 -418
rect 745 -806 751 -430
rect 785 -806 791 -430
rect 745 -818 791 -806
rect 841 -430 887 -418
rect 841 -806 847 -430
rect 881 -806 887 -430
rect 841 -818 887 -806
rect 937 -430 983 -418
rect 937 -806 943 -430
rect 977 -806 983 -430
rect 937 -818 983 -806
rect 1033 -430 1079 -418
rect 1033 -806 1039 -430
rect 1073 -806 1079 -430
rect 1033 -818 1079 -806
rect 1129 -430 1175 -418
rect 1129 -806 1135 -430
rect 1169 -806 1175 -430
rect 1129 -818 1175 -806
rect 1225 -430 1271 -418
rect 1225 -806 1231 -430
rect 1265 -806 1271 -430
rect 1225 -818 1271 -806
rect 1321 -430 1367 -418
rect 1321 -806 1327 -430
rect 1361 -806 1367 -430
rect 1321 -818 1367 -806
rect 1417 -430 1463 -418
rect 1417 -806 1423 -430
rect 1457 -806 1463 -430
rect 1417 -818 1463 -806
rect 1513 -430 1559 -418
rect 1513 -806 1519 -430
rect 1553 -806 1559 -430
rect 1513 -818 1559 -806
rect 1609 -430 1655 -418
rect 1609 -806 1615 -430
rect 1649 -806 1655 -430
rect 1609 -818 1655 -806
rect 1705 -430 1751 -418
rect 1705 -806 1711 -430
rect 1745 -806 1751 -430
rect 1705 -818 1751 -806
rect 1801 -430 1847 -418
rect 1801 -806 1807 -430
rect 1841 -806 1847 -430
rect 1801 -818 1847 -806
rect 1897 -430 1943 -418
rect 1897 -806 1903 -430
rect 1937 -806 1943 -430
rect 1897 -818 1943 -806
rect 1993 -430 2039 -418
rect 1993 -806 1999 -430
rect 2033 -806 2039 -430
rect 1993 -818 2039 -806
rect 2089 -430 2135 -418
rect 2089 -806 2095 -430
rect 2129 -806 2135 -430
rect 2089 -818 2135 -806
rect 2185 -430 2231 -418
rect 2185 -806 2191 -430
rect 2225 -806 2231 -430
rect 2185 -818 2231 -806
rect 2281 -430 2327 -418
rect 2281 -806 2287 -430
rect 2321 -806 2327 -430
rect 2281 -818 2327 -806
rect 2377 -430 2423 -418
rect 2377 -806 2383 -430
rect 2417 -806 2423 -430
rect 2377 -818 2423 -806
rect 2473 -430 2519 -418
rect 2473 -806 2479 -430
rect 2513 -806 2519 -430
rect 2473 -818 2519 -806
rect 2569 -430 2615 -418
rect 2569 -806 2575 -430
rect 2609 -806 2615 -430
rect 2569 -818 2615 -806
rect 2665 -430 2711 -418
rect 2665 -806 2671 -430
rect 2705 -806 2711 -430
rect 2665 -818 2711 -806
rect 2761 -430 2807 -418
rect 2761 -806 2767 -430
rect 2801 -806 2807 -430
rect 2761 -818 2807 -806
rect 2857 -430 2903 -418
rect 2857 -806 2863 -430
rect 2897 -806 2903 -430
rect 2857 -818 2903 -806
rect 2953 -430 2999 -418
rect 2953 -806 2959 -430
rect 2993 -806 2999 -430
rect 2953 -818 2999 -806
rect 3049 -430 3095 -418
rect 3049 -806 3055 -430
rect 3089 -806 3095 -430
rect 3049 -818 3095 -806
rect 3145 -430 3191 -418
rect 3145 -806 3151 -430
rect 3185 -806 3191 -430
rect 3145 -818 3191 -806
rect 3241 -430 3287 -418
rect 3241 -806 3247 -430
rect 3281 -806 3287 -430
rect 3241 -818 3287 -806
rect 3337 -430 3383 -418
rect 3337 -806 3343 -430
rect 3377 -806 3383 -430
rect 3337 -818 3383 -806
rect 3433 -430 3479 -418
rect 3433 -806 3439 -430
rect 3473 -806 3479 -430
rect 3433 -818 3479 -806
rect 3529 -430 3575 -418
rect 3529 -806 3535 -430
rect 3569 -806 3575 -430
rect 3529 -818 3575 -806
rect 3625 -430 3671 -418
rect 3625 -806 3631 -430
rect 3665 -806 3671 -430
rect 3625 -818 3671 -806
rect 3721 -430 3767 -418
rect 3721 -806 3727 -430
rect 3761 -806 3767 -430
rect 3721 -818 3767 -806
rect 3817 -430 3863 -418
rect 3817 -806 3823 -430
rect 3857 -806 3863 -430
rect 3817 -818 3863 -806
rect -3821 -856 -3763 -850
rect -3821 -890 -3809 -856
rect -3775 -890 -3763 -856
rect -3821 -896 -3763 -890
rect -3629 -856 -3571 -850
rect -3629 -890 -3617 -856
rect -3583 -890 -3571 -856
rect -3629 -896 -3571 -890
rect -3437 -856 -3379 -850
rect -3437 -890 -3425 -856
rect -3391 -890 -3379 -856
rect -3437 -896 -3379 -890
rect -3245 -856 -3187 -850
rect -3245 -890 -3233 -856
rect -3199 -890 -3187 -856
rect -3245 -896 -3187 -890
rect -3053 -856 -2995 -850
rect -3053 -890 -3041 -856
rect -3007 -890 -2995 -856
rect -3053 -896 -2995 -890
rect -2861 -856 -2803 -850
rect -2861 -890 -2849 -856
rect -2815 -890 -2803 -856
rect -2861 -896 -2803 -890
rect -2669 -856 -2611 -850
rect -2669 -890 -2657 -856
rect -2623 -890 -2611 -856
rect -2669 -896 -2611 -890
rect -2477 -856 -2419 -850
rect -2477 -890 -2465 -856
rect -2431 -890 -2419 -856
rect -2477 -896 -2419 -890
rect -2285 -856 -2227 -850
rect -2285 -890 -2273 -856
rect -2239 -890 -2227 -856
rect -2285 -896 -2227 -890
rect -2093 -856 -2035 -850
rect -2093 -890 -2081 -856
rect -2047 -890 -2035 -856
rect -2093 -896 -2035 -890
rect -1901 -856 -1843 -850
rect -1901 -890 -1889 -856
rect -1855 -890 -1843 -856
rect -1901 -896 -1843 -890
rect -1709 -856 -1651 -850
rect -1709 -890 -1697 -856
rect -1663 -890 -1651 -856
rect -1709 -896 -1651 -890
rect -1517 -856 -1459 -850
rect -1517 -890 -1505 -856
rect -1471 -890 -1459 -856
rect -1517 -896 -1459 -890
rect -1325 -856 -1267 -850
rect -1325 -890 -1313 -856
rect -1279 -890 -1267 -856
rect -1325 -896 -1267 -890
rect -1133 -856 -1075 -850
rect -1133 -890 -1121 -856
rect -1087 -890 -1075 -856
rect -1133 -896 -1075 -890
rect -941 -856 -883 -850
rect -941 -890 -929 -856
rect -895 -890 -883 -856
rect -941 -896 -883 -890
rect -749 -856 -691 -850
rect -749 -890 -737 -856
rect -703 -890 -691 -856
rect -749 -896 -691 -890
rect -557 -856 -499 -850
rect -557 -890 -545 -856
rect -511 -890 -499 -856
rect -557 -896 -499 -890
rect -365 -856 -307 -850
rect -365 -890 -353 -856
rect -319 -890 -307 -856
rect -365 -896 -307 -890
rect -173 -856 -115 -850
rect -173 -890 -161 -856
rect -127 -890 -115 -856
rect -173 -896 -115 -890
rect 19 -856 77 -850
rect 19 -890 31 -856
rect 65 -890 77 -856
rect 19 -896 77 -890
rect 211 -856 269 -850
rect 211 -890 223 -856
rect 257 -890 269 -856
rect 211 -896 269 -890
rect 403 -856 461 -850
rect 403 -890 415 -856
rect 449 -890 461 -856
rect 403 -896 461 -890
rect 595 -856 653 -850
rect 595 -890 607 -856
rect 641 -890 653 -856
rect 595 -896 653 -890
rect 787 -856 845 -850
rect 787 -890 799 -856
rect 833 -890 845 -856
rect 787 -896 845 -890
rect 979 -856 1037 -850
rect 979 -890 991 -856
rect 1025 -890 1037 -856
rect 979 -896 1037 -890
rect 1171 -856 1229 -850
rect 1171 -890 1183 -856
rect 1217 -890 1229 -856
rect 1171 -896 1229 -890
rect 1363 -856 1421 -850
rect 1363 -890 1375 -856
rect 1409 -890 1421 -856
rect 1363 -896 1421 -890
rect 1555 -856 1613 -850
rect 1555 -890 1567 -856
rect 1601 -890 1613 -856
rect 1555 -896 1613 -890
rect 1747 -856 1805 -850
rect 1747 -890 1759 -856
rect 1793 -890 1805 -856
rect 1747 -896 1805 -890
rect 1939 -856 1997 -850
rect 1939 -890 1951 -856
rect 1985 -890 1997 -856
rect 1939 -896 1997 -890
rect 2131 -856 2189 -850
rect 2131 -890 2143 -856
rect 2177 -890 2189 -856
rect 2131 -896 2189 -890
rect 2323 -856 2381 -850
rect 2323 -890 2335 -856
rect 2369 -890 2381 -856
rect 2323 -896 2381 -890
rect 2515 -856 2573 -850
rect 2515 -890 2527 -856
rect 2561 -890 2573 -856
rect 2515 -896 2573 -890
rect 2707 -856 2765 -850
rect 2707 -890 2719 -856
rect 2753 -890 2765 -856
rect 2707 -896 2765 -890
rect 2899 -856 2957 -850
rect 2899 -890 2911 -856
rect 2945 -890 2957 -856
rect 2899 -896 2957 -890
rect 3091 -856 3149 -850
rect 3091 -890 3103 -856
rect 3137 -890 3149 -856
rect 3091 -896 3149 -890
rect 3283 -856 3341 -850
rect 3283 -890 3295 -856
rect 3329 -890 3341 -856
rect 3283 -896 3341 -890
rect 3475 -856 3533 -850
rect 3475 -890 3487 -856
rect 3521 -890 3533 -856
rect 3475 -896 3533 -890
rect 3667 -856 3725 -850
rect 3667 -890 3679 -856
rect 3713 -890 3725 -856
rect 3667 -896 3725 -890
<< properties >>
string FIXED_BBOX -3954 -975 3954 975
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 3 nf 80 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
