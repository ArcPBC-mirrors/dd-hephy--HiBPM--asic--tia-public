magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< locali >>
rect -1352 -2420 -752 -2180
rect 442 -2210 1042 -2180
rect 1654 -2192 2864 -2178
rect 2242 -2200 2864 -2192
rect 442 -2420 1048 -2210
rect 2242 -2380 2858 -2200
rect -1036 -4140 -752 -2420
rect 764 -4140 1048 -2420
rect 2572 -4140 2856 -2380
rect -2560 -4340 -2260 -4140
rect -1036 -4340 -460 -4140
rect 764 -4340 1340 -4140
rect 2572 -4340 3140 -4140
rect -1036 -7960 -752 -4340
rect 764 -7952 1048 -4340
rect 764 -7960 836 -7952
rect -1040 -8160 -980 -7960
rect -800 -8160 -740 -7960
rect 760 -8160 836 -7960
rect 780 -8164 836 -8160
rect 1016 -7960 1048 -7952
rect 2572 -7952 2856 -4340
rect 2572 -7960 2612 -7952
rect 1016 -8164 1060 -7960
rect 2560 -8160 2612 -7960
rect 780 -8180 1060 -8164
rect 2576 -8164 2612 -8160
rect 2792 -7960 2856 -7952
rect 2792 -8160 2860 -7960
rect 2792 -8164 2852 -8160
rect 2576 -8188 2852 -8164
<< viali >>
rect -980 -8160 -800 -7960
rect 836 -8164 1016 -7952
rect 2612 -8164 2792 -7952
<< metal1 >>
rect -2646 -2320 3988 -2176
rect -2646 -2792 -2592 -2320
rect -1408 -2792 -1176 -2320
rect 396 -2792 628 -2320
rect 2196 -2792 2428 -2320
rect -2646 -2936 3988 -2792
rect -2646 -3408 -2592 -2936
rect -1408 -3408 -1176 -2936
rect 396 -3408 628 -2936
rect 2196 -3408 2428 -2936
rect -2646 -3552 3988 -3408
rect -2646 -4032 -2592 -3552
rect -1408 -4032 -1176 -3552
rect 396 -4032 628 -3552
rect 2196 -4032 2428 -3552
rect 3996 -4032 4228 -2244
rect -2646 -4440 4232 -4032
rect -986 -7960 -794 -7948
rect 830 -7952 1022 -7940
rect 2606 -7952 2798 -7940
rect -990 -8160 -980 -7960
rect -800 -8160 -790 -7960
rect -986 -8172 -794 -8160
rect 826 -8164 836 -7952
rect 1016 -8164 1026 -7952
rect 2602 -8164 2612 -7952
rect 2792 -8164 2802 -7952
rect 830 -8176 1022 -8164
rect 2606 -8176 2798 -8164
<< via1 >>
rect -980 -8160 -800 -7960
rect 836 -8164 1016 -7952
rect 2612 -8164 2792 -7952
<< metal2 >>
rect -2374 -2510 4296 -2174
rect -1440 -4680 4036 -4464
rect -980 -7960 -800 -7950
rect -980 -8170 -800 -8160
rect 836 -7952 1016 -7942
rect 836 -8174 1016 -8164
rect 2612 -7952 2792 -7942
rect 2612 -8174 2792 -8164
<< via2 >>
rect -980 -8160 -800 -7960
rect 2612 -8164 2792 -7952
<< metal3 >>
rect -1710 -7988 -1700 -7548
rect -1128 -7988 -1118 -7548
rect -990 -7960 -790 -7955
rect -990 -8160 -980 -7960
rect -800 -8160 -790 -7960
rect 90 -7988 100 -7548
rect 672 -7988 682 -7548
rect -990 -8165 -790 -8160
rect 826 -8164 836 -7952
rect 1016 -8164 1026 -7952
rect 1886 -7992 1896 -7552
rect 2468 -7992 2478 -7552
rect 2602 -7952 2802 -7947
rect 2602 -8164 2612 -7952
rect 2792 -8164 2802 -7952
rect 3686 -7992 3696 -7552
rect 4268 -7992 4278 -7552
rect 2602 -8169 2802 -8164
<< via3 >>
rect -1700 -7988 -1128 -7548
rect -980 -8160 -800 -7960
rect 100 -7988 672 -7548
rect 836 -8164 1016 -7952
rect 1896 -7992 2468 -7552
rect 2612 -8164 2792 -7952
rect 3696 -7992 4268 -7552
<< metal4 >>
rect -1716 -7548 -1116 -7540
rect -1716 -7988 -1700 -7548
rect -1128 -7900 -1116 -7548
rect 84 -7548 684 -7540
rect -1128 -7960 -740 -7900
rect -1128 -7988 -980 -7960
rect -1716 -8160 -980 -7988
rect -800 -8160 -740 -7960
rect -1716 -8320 -740 -8160
rect 84 -7988 100 -7548
rect 672 -7904 684 -7548
rect 1884 -7552 2484 -7540
rect 672 -7952 1036 -7904
rect 672 -7988 836 -7952
rect 84 -8164 836 -7988
rect 1016 -8164 1036 -7952
rect 84 -8320 1036 -8164
rect 1884 -7992 1896 -7552
rect 2468 -7876 2484 -7552
rect 3684 -7552 4284 -7544
rect 2468 -7952 2820 -7876
rect 2468 -7992 2612 -7952
rect 1884 -8164 2612 -7992
rect 2792 -8164 2820 -7952
rect 1884 -8320 2820 -8164
rect 3684 -7992 3696 -7552
rect 4268 -7992 4284 -7552
rect 3684 -8320 4284 -7992
use curr_m  curr_m_0
timestamp 1686659968
transform 1 0 -800 0 1 -3800
box 0 -4400 1624 1656
use curr_m  curr_m_1
timestamp 1686659968
transform 1 0 -2600 0 1 -3800
box 0 -4400 1624 1656
use curr_m  curr_m_2
timestamp 1686659968
transform 1 0 1000 0 1 -3800
box 0 -4400 1624 1656
use curr_m  curr_m_3
timestamp 1686659968
transform 1 0 2800 0 1 -3800
box 0 -4400 1624 1656
<< end >>
