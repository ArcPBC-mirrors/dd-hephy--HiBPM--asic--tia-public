magic
tech sky130A
magscale 1 2
timestamp 1685096196
<< metal3 >>
rect -1186 2512 1186 2540
rect -1186 -2512 1102 2512
rect 1166 -2512 1186 2512
rect -1186 -2540 1186 -2512
<< via3 >>
rect 1102 -2512 1166 2512
<< mimcap >>
rect -1146 2460 854 2500
rect -1146 -2460 -1106 2460
rect 814 -2460 854 2460
rect -1146 -2500 854 -2460
<< mimcapcontact >>
rect -1106 -2460 814 2460
<< metal4 >>
rect 1086 2512 1182 2528
rect -1107 2460 815 2461
rect -1107 -2460 -1106 2460
rect 814 -2460 815 2460
rect -1107 -2461 815 -2460
rect 1086 -2512 1102 2512
rect 1166 -2512 1182 2512
rect 1086 -2528 1182 -2512
<< properties >>
string FIXED_BBOX -1186 -2540 894 2540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 25 val 513.299 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
