magic
tech sky130A
magscale 1 2
timestamp 1683553987
<< error_p >>
rect -365 917 -307 923
rect -173 917 -115 923
rect 19 917 77 923
rect 211 917 269 923
rect 403 917 461 923
rect -365 883 -353 917
rect -173 883 -161 917
rect 19 883 31 917
rect 211 883 223 917
rect 403 883 415 917
rect -365 877 -307 883
rect -173 877 -115 883
rect 19 877 77 883
rect 211 877 269 883
rect 403 877 461 883
rect -461 389 -403 395
rect -269 389 -211 395
rect -77 389 -19 395
rect 115 389 173 395
rect 307 389 365 395
rect -461 355 -449 389
rect -269 355 -257 389
rect -77 355 -65 389
rect 115 355 127 389
rect 307 355 319 389
rect -461 349 -403 355
rect -269 349 -211 355
rect -77 349 -19 355
rect 115 349 173 355
rect 307 349 365 355
rect -461 281 -403 287
rect -269 281 -211 287
rect -77 281 -19 287
rect 115 281 173 287
rect 307 281 365 287
rect -461 247 -449 281
rect -269 247 -257 281
rect -77 247 -65 281
rect 115 247 127 281
rect 307 247 319 281
rect -461 241 -403 247
rect -269 241 -211 247
rect -77 241 -19 247
rect 115 241 173 247
rect 307 241 365 247
rect -365 -247 -307 -241
rect -173 -247 -115 -241
rect 19 -247 77 -241
rect 211 -247 269 -241
rect 403 -247 461 -241
rect -365 -281 -353 -247
rect -173 -281 -161 -247
rect 19 -281 31 -247
rect 211 -281 223 -247
rect 403 -281 415 -247
rect -365 -287 -307 -281
rect -173 -287 -115 -281
rect 19 -287 77 -281
rect 211 -287 269 -281
rect 403 -287 461 -281
rect -365 -355 -307 -349
rect -173 -355 -115 -349
rect 19 -355 77 -349
rect 211 -355 269 -349
rect 403 -355 461 -349
rect -365 -389 -353 -355
rect -173 -389 -161 -355
rect 19 -389 31 -355
rect 211 -389 223 -355
rect 403 -389 415 -355
rect -365 -395 -307 -389
rect -173 -395 -115 -389
rect 19 -395 77 -389
rect 211 -395 269 -389
rect 403 -395 461 -389
rect -461 -883 -403 -877
rect -269 -883 -211 -877
rect -77 -883 -19 -877
rect 115 -883 173 -877
rect 307 -883 365 -877
rect -461 -917 -449 -883
rect -269 -917 -257 -883
rect -77 -917 -65 -883
rect 115 -917 127 -883
rect 307 -917 319 -883
rect -461 -923 -403 -917
rect -269 -923 -211 -917
rect -77 -923 -19 -917
rect 115 -923 173 -917
rect 307 -923 365 -917
<< nwell >>
rect -647 -1055 647 1055
<< pmos >>
rect -447 436 -417 836
rect -351 436 -321 836
rect -255 436 -225 836
rect -159 436 -129 836
rect -63 436 -33 836
rect 33 436 63 836
rect 129 436 159 836
rect 225 436 255 836
rect 321 436 351 836
rect 417 436 447 836
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect -447 -836 -417 -436
rect -351 -836 -321 -436
rect -255 -836 -225 -436
rect -159 -836 -129 -436
rect -63 -836 -33 -436
rect 33 -836 63 -436
rect 129 -836 159 -436
rect 225 -836 255 -436
rect 321 -836 351 -436
rect 417 -836 447 -436
<< pdiff >>
rect -509 824 -447 836
rect -509 448 -497 824
rect -463 448 -447 824
rect -509 436 -447 448
rect -417 824 -351 836
rect -417 448 -401 824
rect -367 448 -351 824
rect -417 436 -351 448
rect -321 824 -255 836
rect -321 448 -305 824
rect -271 448 -255 824
rect -321 436 -255 448
rect -225 824 -159 836
rect -225 448 -209 824
rect -175 448 -159 824
rect -225 436 -159 448
rect -129 824 -63 836
rect -129 448 -113 824
rect -79 448 -63 824
rect -129 436 -63 448
rect -33 824 33 836
rect -33 448 -17 824
rect 17 448 33 824
rect -33 436 33 448
rect 63 824 129 836
rect 63 448 79 824
rect 113 448 129 824
rect 63 436 129 448
rect 159 824 225 836
rect 159 448 175 824
rect 209 448 225 824
rect 159 436 225 448
rect 255 824 321 836
rect 255 448 271 824
rect 305 448 321 824
rect 255 436 321 448
rect 351 824 417 836
rect 351 448 367 824
rect 401 448 417 824
rect 351 436 417 448
rect 447 824 509 836
rect 447 448 463 824
rect 497 448 509 824
rect 447 436 509 448
rect -509 188 -447 200
rect -509 -188 -497 188
rect -463 -188 -447 188
rect -509 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 509 200
rect 447 -188 463 188
rect 497 -188 509 188
rect 447 -200 509 -188
rect -509 -448 -447 -436
rect -509 -824 -497 -448
rect -463 -824 -447 -448
rect -509 -836 -447 -824
rect -417 -448 -351 -436
rect -417 -824 -401 -448
rect -367 -824 -351 -448
rect -417 -836 -351 -824
rect -321 -448 -255 -436
rect -321 -824 -305 -448
rect -271 -824 -255 -448
rect -321 -836 -255 -824
rect -225 -448 -159 -436
rect -225 -824 -209 -448
rect -175 -824 -159 -448
rect -225 -836 -159 -824
rect -129 -448 -63 -436
rect -129 -824 -113 -448
rect -79 -824 -63 -448
rect -129 -836 -63 -824
rect -33 -448 33 -436
rect -33 -824 -17 -448
rect 17 -824 33 -448
rect -33 -836 33 -824
rect 63 -448 129 -436
rect 63 -824 79 -448
rect 113 -824 129 -448
rect 63 -836 129 -824
rect 159 -448 225 -436
rect 159 -824 175 -448
rect 209 -824 225 -448
rect 159 -836 225 -824
rect 255 -448 321 -436
rect 255 -824 271 -448
rect 305 -824 321 -448
rect 255 -836 321 -824
rect 351 -448 417 -436
rect 351 -824 367 -448
rect 401 -824 417 -448
rect 351 -836 417 -824
rect 447 -448 509 -436
rect 447 -824 463 -448
rect 497 -824 509 -448
rect 447 -836 509 -824
<< pdiffc >>
rect -497 448 -463 824
rect -401 448 -367 824
rect -305 448 -271 824
rect -209 448 -175 824
rect -113 448 -79 824
rect -17 448 17 824
rect 79 448 113 824
rect 175 448 209 824
rect 271 448 305 824
rect 367 448 401 824
rect 463 448 497 824
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -497 -824 -463 -448
rect -401 -824 -367 -448
rect -305 -824 -271 -448
rect -209 -824 -175 -448
rect -113 -824 -79 -448
rect -17 -824 17 -448
rect 79 -824 113 -448
rect 175 -824 209 -448
rect 271 -824 305 -448
rect 367 -824 401 -448
rect 463 -824 497 -448
<< nsubdiff >>
rect -611 985 -515 1019
rect 515 985 611 1019
rect -611 923 -577 985
rect 577 923 611 985
rect -611 -985 -577 -923
rect 577 -985 611 -923
rect -611 -1019 -515 -985
rect 515 -1019 611 -985
<< nsubdiffcont >>
rect -515 985 515 1019
rect -611 -923 -577 923
rect 577 -923 611 923
rect -515 -1019 515 -985
<< poly >>
rect -369 917 -303 933
rect -369 883 -353 917
rect -319 883 -303 917
rect -369 867 -303 883
rect -177 917 -111 933
rect -177 883 -161 917
rect -127 883 -111 917
rect -177 867 -111 883
rect 15 917 81 933
rect 15 883 31 917
rect 65 883 81 917
rect 15 867 81 883
rect 207 917 273 933
rect 207 883 223 917
rect 257 883 273 917
rect 207 867 273 883
rect 399 917 465 933
rect 399 883 415 917
rect 449 883 465 917
rect 399 867 465 883
rect -447 836 -417 862
rect -351 836 -321 867
rect -255 836 -225 862
rect -159 836 -129 867
rect -63 836 -33 862
rect 33 836 63 867
rect 129 836 159 862
rect 225 836 255 867
rect 321 836 351 862
rect 417 836 447 867
rect -447 405 -417 436
rect -351 410 -321 436
rect -255 405 -225 436
rect -159 410 -129 436
rect -63 405 -33 436
rect 33 410 63 436
rect 129 405 159 436
rect 225 410 255 436
rect 321 405 351 436
rect 417 410 447 436
rect -465 389 -399 405
rect -465 355 -449 389
rect -415 355 -399 389
rect -465 339 -399 355
rect -273 389 -207 405
rect -273 355 -257 389
rect -223 355 -207 389
rect -273 339 -207 355
rect -81 389 -15 405
rect -81 355 -65 389
rect -31 355 -15 389
rect -81 339 -15 355
rect 111 389 177 405
rect 111 355 127 389
rect 161 355 177 389
rect 111 339 177 355
rect 303 389 369 405
rect 303 355 319 389
rect 353 355 369 389
rect 303 339 369 355
rect -465 281 -399 297
rect -465 247 -449 281
rect -415 247 -399 281
rect -465 231 -399 247
rect -273 281 -207 297
rect -273 247 -257 281
rect -223 247 -207 281
rect -273 231 -207 247
rect -81 281 -15 297
rect -81 247 -65 281
rect -31 247 -15 281
rect -81 231 -15 247
rect 111 281 177 297
rect 111 247 127 281
rect 161 247 177 281
rect 111 231 177 247
rect 303 281 369 297
rect 303 247 319 281
rect 353 247 369 281
rect 303 231 369 247
rect -447 200 -417 231
rect -351 200 -321 226
rect -255 200 -225 231
rect -159 200 -129 226
rect -63 200 -33 231
rect 33 200 63 226
rect 129 200 159 231
rect 225 200 255 226
rect 321 200 351 231
rect 417 200 447 226
rect -447 -226 -417 -200
rect -351 -231 -321 -200
rect -255 -226 -225 -200
rect -159 -231 -129 -200
rect -63 -226 -33 -200
rect 33 -231 63 -200
rect 129 -226 159 -200
rect 225 -231 255 -200
rect 321 -226 351 -200
rect 417 -231 447 -200
rect -369 -247 -303 -231
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -369 -297 -303 -281
rect -177 -247 -111 -231
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect -177 -297 -111 -281
rect 15 -247 81 -231
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 15 -297 81 -281
rect 207 -247 273 -231
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 207 -297 273 -281
rect 399 -247 465 -231
rect 399 -281 415 -247
rect 449 -281 465 -247
rect 399 -297 465 -281
rect -369 -355 -303 -339
rect -369 -389 -353 -355
rect -319 -389 -303 -355
rect -369 -405 -303 -389
rect -177 -355 -111 -339
rect -177 -389 -161 -355
rect -127 -389 -111 -355
rect -177 -405 -111 -389
rect 15 -355 81 -339
rect 15 -389 31 -355
rect 65 -389 81 -355
rect 15 -405 81 -389
rect 207 -355 273 -339
rect 207 -389 223 -355
rect 257 -389 273 -355
rect 207 -405 273 -389
rect 399 -355 465 -339
rect 399 -389 415 -355
rect 449 -389 465 -355
rect 399 -405 465 -389
rect -447 -436 -417 -410
rect -351 -436 -321 -405
rect -255 -436 -225 -410
rect -159 -436 -129 -405
rect -63 -436 -33 -410
rect 33 -436 63 -405
rect 129 -436 159 -410
rect 225 -436 255 -405
rect 321 -436 351 -410
rect 417 -436 447 -405
rect -447 -867 -417 -836
rect -351 -862 -321 -836
rect -255 -867 -225 -836
rect -159 -862 -129 -836
rect -63 -867 -33 -836
rect 33 -862 63 -836
rect 129 -867 159 -836
rect 225 -862 255 -836
rect 321 -867 351 -836
rect 417 -862 447 -836
rect -465 -883 -399 -867
rect -465 -917 -449 -883
rect -415 -917 -399 -883
rect -465 -933 -399 -917
rect -273 -883 -207 -867
rect -273 -917 -257 -883
rect -223 -917 -207 -883
rect -273 -933 -207 -917
rect -81 -883 -15 -867
rect -81 -917 -65 -883
rect -31 -917 -15 -883
rect -81 -933 -15 -917
rect 111 -883 177 -867
rect 111 -917 127 -883
rect 161 -917 177 -883
rect 111 -933 177 -917
rect 303 -883 369 -867
rect 303 -917 319 -883
rect 353 -917 369 -883
rect 303 -933 369 -917
<< polycont >>
rect -353 883 -319 917
rect -161 883 -127 917
rect 31 883 65 917
rect 223 883 257 917
rect 415 883 449 917
rect -449 355 -415 389
rect -257 355 -223 389
rect -65 355 -31 389
rect 127 355 161 389
rect 319 355 353 389
rect -449 247 -415 281
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
rect 415 -281 449 -247
rect -353 -389 -319 -355
rect -161 -389 -127 -355
rect 31 -389 65 -355
rect 223 -389 257 -355
rect 415 -389 449 -355
rect -449 -917 -415 -883
rect -257 -917 -223 -883
rect -65 -917 -31 -883
rect 127 -917 161 -883
rect 319 -917 353 -883
<< locali >>
rect -611 985 -515 1019
rect 515 985 611 1019
rect -611 923 -577 985
rect 577 923 611 985
rect -369 883 -353 917
rect -319 883 -303 917
rect -177 883 -161 917
rect -127 883 -111 917
rect 15 883 31 917
rect 65 883 81 917
rect 207 883 223 917
rect 257 883 273 917
rect 399 883 415 917
rect 449 883 465 917
rect -497 824 -463 840
rect -497 432 -463 448
rect -401 824 -367 840
rect -401 432 -367 448
rect -305 824 -271 840
rect -305 432 -271 448
rect -209 824 -175 840
rect -209 432 -175 448
rect -113 824 -79 840
rect -113 432 -79 448
rect -17 824 17 840
rect -17 432 17 448
rect 79 824 113 840
rect 79 432 113 448
rect 175 824 209 840
rect 175 432 209 448
rect 271 824 305 840
rect 271 432 305 448
rect 367 824 401 840
rect 367 432 401 448
rect 463 824 497 840
rect 463 432 497 448
rect -465 355 -449 389
rect -415 355 -399 389
rect -273 355 -257 389
rect -223 355 -207 389
rect -81 355 -65 389
rect -31 355 -15 389
rect 111 355 127 389
rect 161 355 177 389
rect 303 355 319 389
rect 353 355 369 389
rect -465 247 -449 281
rect -415 247 -399 281
rect -273 247 -257 281
rect -223 247 -207 281
rect -81 247 -65 281
rect -31 247 -15 281
rect 111 247 127 281
rect 161 247 177 281
rect 303 247 319 281
rect 353 247 369 281
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 399 -281 415 -247
rect 449 -281 465 -247
rect -369 -389 -353 -355
rect -319 -389 -303 -355
rect -177 -389 -161 -355
rect -127 -389 -111 -355
rect 15 -389 31 -355
rect 65 -389 81 -355
rect 207 -389 223 -355
rect 257 -389 273 -355
rect 399 -389 415 -355
rect 449 -389 465 -355
rect -497 -448 -463 -432
rect -497 -840 -463 -824
rect -401 -448 -367 -432
rect -401 -840 -367 -824
rect -305 -448 -271 -432
rect -305 -840 -271 -824
rect -209 -448 -175 -432
rect -209 -840 -175 -824
rect -113 -448 -79 -432
rect -113 -840 -79 -824
rect -17 -448 17 -432
rect -17 -840 17 -824
rect 79 -448 113 -432
rect 79 -840 113 -824
rect 175 -448 209 -432
rect 175 -840 209 -824
rect 271 -448 305 -432
rect 271 -840 305 -824
rect 367 -448 401 -432
rect 367 -840 401 -824
rect 463 -448 497 -432
rect 463 -840 497 -824
rect -465 -917 -449 -883
rect -415 -917 -399 -883
rect -273 -917 -257 -883
rect -223 -917 -207 -883
rect -81 -917 -65 -883
rect -31 -917 -15 -883
rect 111 -917 127 -883
rect 161 -917 177 -883
rect 303 -917 319 -883
rect 353 -917 369 -883
rect -611 -985 -577 -923
rect 577 -985 611 -923
rect -611 -1019 -515 -985
rect 515 -1019 611 -985
<< viali >>
rect -353 883 -319 917
rect -161 883 -127 917
rect 31 883 65 917
rect 223 883 257 917
rect 415 883 449 917
rect -497 448 -463 824
rect -401 448 -367 824
rect -305 448 -271 824
rect -209 448 -175 824
rect -113 448 -79 824
rect -17 448 17 824
rect 79 448 113 824
rect 175 448 209 824
rect 271 448 305 824
rect 367 448 401 824
rect 463 448 497 824
rect -449 355 -415 389
rect -257 355 -223 389
rect -65 355 -31 389
rect 127 355 161 389
rect 319 355 353 389
rect -449 247 -415 281
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
rect 415 -281 449 -247
rect -353 -389 -319 -355
rect -161 -389 -127 -355
rect 31 -389 65 -355
rect 223 -389 257 -355
rect 415 -389 449 -355
rect -497 -824 -463 -448
rect -401 -824 -367 -448
rect -305 -824 -271 -448
rect -209 -824 -175 -448
rect -113 -824 -79 -448
rect -17 -824 17 -448
rect 79 -824 113 -448
rect 175 -824 209 -448
rect 271 -824 305 -448
rect 367 -824 401 -448
rect 463 -824 497 -448
rect -449 -917 -415 -883
rect -257 -917 -223 -883
rect -65 -917 -31 -883
rect 127 -917 161 -883
rect 319 -917 353 -883
<< metal1 >>
rect -365 917 -307 923
rect -365 883 -353 917
rect -319 883 -307 917
rect -365 877 -307 883
rect -173 917 -115 923
rect -173 883 -161 917
rect -127 883 -115 917
rect -173 877 -115 883
rect 19 917 77 923
rect 19 883 31 917
rect 65 883 77 917
rect 19 877 77 883
rect 211 917 269 923
rect 211 883 223 917
rect 257 883 269 917
rect 211 877 269 883
rect 403 917 461 923
rect 403 883 415 917
rect 449 883 461 917
rect 403 877 461 883
rect -503 824 -457 836
rect -503 448 -497 824
rect -463 448 -457 824
rect -503 436 -457 448
rect -407 824 -361 836
rect -407 448 -401 824
rect -367 448 -361 824
rect -407 436 -361 448
rect -311 824 -265 836
rect -311 448 -305 824
rect -271 448 -265 824
rect -311 436 -265 448
rect -215 824 -169 836
rect -215 448 -209 824
rect -175 448 -169 824
rect -215 436 -169 448
rect -119 824 -73 836
rect -119 448 -113 824
rect -79 448 -73 824
rect -119 436 -73 448
rect -23 824 23 836
rect -23 448 -17 824
rect 17 448 23 824
rect -23 436 23 448
rect 73 824 119 836
rect 73 448 79 824
rect 113 448 119 824
rect 73 436 119 448
rect 169 824 215 836
rect 169 448 175 824
rect 209 448 215 824
rect 169 436 215 448
rect 265 824 311 836
rect 265 448 271 824
rect 305 448 311 824
rect 265 436 311 448
rect 361 824 407 836
rect 361 448 367 824
rect 401 448 407 824
rect 361 436 407 448
rect 457 824 503 836
rect 457 448 463 824
rect 497 448 503 824
rect 457 436 503 448
rect -461 389 -403 395
rect -461 355 -449 389
rect -415 355 -403 389
rect -461 349 -403 355
rect -269 389 -211 395
rect -269 355 -257 389
rect -223 355 -211 389
rect -269 349 -211 355
rect -77 389 -19 395
rect -77 355 -65 389
rect -31 355 -19 389
rect -77 349 -19 355
rect 115 389 173 395
rect 115 355 127 389
rect 161 355 173 389
rect 115 349 173 355
rect 307 389 365 395
rect 307 355 319 389
rect 353 355 365 389
rect 307 349 365 355
rect -461 281 -403 287
rect -461 247 -449 281
rect -415 247 -403 281
rect -461 241 -403 247
rect -269 281 -211 287
rect -269 247 -257 281
rect -223 247 -211 281
rect -269 241 -211 247
rect -77 281 -19 287
rect -77 247 -65 281
rect -31 247 -19 281
rect -77 241 -19 247
rect 115 281 173 287
rect 115 247 127 281
rect 161 247 173 281
rect 115 241 173 247
rect 307 281 365 287
rect 307 247 319 281
rect 353 247 365 281
rect 307 241 365 247
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect -365 -247 -307 -241
rect -365 -281 -353 -247
rect -319 -281 -307 -247
rect -365 -287 -307 -281
rect -173 -247 -115 -241
rect -173 -281 -161 -247
rect -127 -281 -115 -247
rect -173 -287 -115 -281
rect 19 -247 77 -241
rect 19 -281 31 -247
rect 65 -281 77 -247
rect 19 -287 77 -281
rect 211 -247 269 -241
rect 211 -281 223 -247
rect 257 -281 269 -247
rect 211 -287 269 -281
rect 403 -247 461 -241
rect 403 -281 415 -247
rect 449 -281 461 -247
rect 403 -287 461 -281
rect -365 -355 -307 -349
rect -365 -389 -353 -355
rect -319 -389 -307 -355
rect -365 -395 -307 -389
rect -173 -355 -115 -349
rect -173 -389 -161 -355
rect -127 -389 -115 -355
rect -173 -395 -115 -389
rect 19 -355 77 -349
rect 19 -389 31 -355
rect 65 -389 77 -355
rect 19 -395 77 -389
rect 211 -355 269 -349
rect 211 -389 223 -355
rect 257 -389 269 -355
rect 211 -395 269 -389
rect 403 -355 461 -349
rect 403 -389 415 -355
rect 449 -389 461 -355
rect 403 -395 461 -389
rect -503 -448 -457 -436
rect -503 -824 -497 -448
rect -463 -824 -457 -448
rect -503 -836 -457 -824
rect -407 -448 -361 -436
rect -407 -824 -401 -448
rect -367 -824 -361 -448
rect -407 -836 -361 -824
rect -311 -448 -265 -436
rect -311 -824 -305 -448
rect -271 -824 -265 -448
rect -311 -836 -265 -824
rect -215 -448 -169 -436
rect -215 -824 -209 -448
rect -175 -824 -169 -448
rect -215 -836 -169 -824
rect -119 -448 -73 -436
rect -119 -824 -113 -448
rect -79 -824 -73 -448
rect -119 -836 -73 -824
rect -23 -448 23 -436
rect -23 -824 -17 -448
rect 17 -824 23 -448
rect -23 -836 23 -824
rect 73 -448 119 -436
rect 73 -824 79 -448
rect 113 -824 119 -448
rect 73 -836 119 -824
rect 169 -448 215 -436
rect 169 -824 175 -448
rect 209 -824 215 -448
rect 169 -836 215 -824
rect 265 -448 311 -436
rect 265 -824 271 -448
rect 305 -824 311 -448
rect 265 -836 311 -824
rect 361 -448 407 -436
rect 361 -824 367 -448
rect 401 -824 407 -448
rect 361 -836 407 -824
rect 457 -448 503 -436
rect 457 -824 463 -448
rect 497 -824 503 -448
rect 457 -836 503 -824
rect -461 -883 -403 -877
rect -461 -917 -449 -883
rect -415 -917 -403 -883
rect -461 -923 -403 -917
rect -269 -883 -211 -877
rect -269 -917 -257 -883
rect -223 -917 -211 -883
rect -269 -923 -211 -917
rect -77 -883 -19 -877
rect -77 -917 -65 -883
rect -31 -917 -19 -883
rect -77 -923 -19 -917
rect 115 -883 173 -877
rect 115 -917 127 -883
rect 161 -917 173 -883
rect 115 -923 173 -917
rect 307 -883 365 -877
rect 307 -917 319 -883
rect 353 -917 365 -883
rect 307 -923 365 -917
<< properties >>
string FIXED_BBOX -594 -1002 594 1002
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 3 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
