magic
tech sky130A
magscale 1 2
timestamp 1689773955
<< psubdiff >>
rect -8900 -4720 -8160 -4696
rect -8900 -5604 -8160 -5580
<< psubdiffcont >>
rect -8900 -5580 -8160 -4720
<< locali >>
rect -10240 4380 -7200 4500
rect -10280 3560 -7240 3680
rect -10380 1320 -7340 1440
rect -9560 -100 -9420 1320
rect -6900 1220 -6840 6760
rect -5100 4420 1500 4520
rect -5140 3540 1580 3700
rect -3580 680 -3440 3540
rect -1840 680 -1700 3540
rect -100 680 40 3540
rect 2760 1820 3800 1920
rect -5100 560 1640 680
rect 3400 440 3800 1820
rect 3400 400 3840 440
rect -5080 -320 2580 -140
rect -5080 -420 2600 -320
rect -9560 -2320 -9420 -800
rect -8900 -4720 -8160 -4704
rect -4820 -4820 -4700 -420
rect -3760 -4820 -3640 -420
rect -2740 -4820 -2620 -420
rect -1680 -4820 -1560 -420
rect -640 -4820 -520 -420
rect 400 -4820 520 -420
rect 1440 -4820 1560 -420
rect 2480 -4820 2600 -420
rect 3520 -4820 3840 400
rect -5760 -4860 3840 -4820
rect -5760 -4960 -5040 -4860
rect -4620 -4960 -860 -4860
rect -440 -4960 3300 -4860
rect 3780 -4960 3840 -4860
rect -8900 -5596 -8160 -5580
<< viali >>
rect -6900 6760 -6840 6860
rect -10140 -3340 -9860 -3060
rect -8900 -5580 -8160 -4720
rect -5040 -4980 -4620 -4860
rect -860 -4980 -440 -4860
rect 3300 -4980 3780 -4860
<< metal1 >>
rect -10520 8320 16620 8440
rect -10520 8220 6640 8320
rect -10520 7500 3280 8220
rect -10520 6860 -6700 7500
rect -10520 6760 -6900 6860
rect -6840 6760 -6700 6860
rect -6906 6748 -6700 6760
rect -6880 5860 -6700 6748
rect -5400 6960 3280 7500
rect 4100 6960 6640 8220
rect -5400 6760 6640 6960
rect -5400 5880 -5390 6760
rect 1660 5880 2720 6760
rect -5400 5860 2720 5880
rect -6880 5220 2720 5860
rect 6500 6560 6640 6760
rect 16540 6560 16620 8320
rect 6500 5580 16620 6560
rect -10340 4260 -9896 4376
rect -7336 4360 -7052 4376
rect -7336 4260 -7100 4360
rect -10340 3800 -10180 4260
rect -7152 3800 -7100 4260
rect -10340 3684 -10024 3800
rect -7360 3684 -7100 3800
rect -7110 3680 -7100 3684
rect -6980 3680 -6970 4360
rect -6880 3520 -5400 5220
rect 1660 4680 2720 5220
rect 1660 4160 1720 4680
rect 3320 4160 3330 4680
rect 1660 3520 2720 4160
rect -6880 2700 2720 3520
rect -6880 2040 -5400 2700
rect 1700 2040 2720 2700
rect -6880 1900 2720 2040
rect -10228 1418 -7336 1558
rect -6880 1420 2540 1900
rect 3000 1740 3300 2020
rect 7130 1700 7140 2480
rect 7300 2320 11320 2480
rect 12400 2320 16520 2480
rect 7300 1820 7380 2320
rect 12400 2240 12600 2320
rect 12010 2040 12020 2240
rect 12540 2040 12600 2240
rect 12400 1820 12600 2040
rect 7300 1700 11220 1820
rect 12400 1700 16420 1820
rect -9480 -716 -9264 1418
rect -7520 1100 -7360 1418
rect -6660 1320 2540 1420
rect -7520 920 -6060 1100
rect -7450 740 -7440 820
rect -7260 740 -7250 820
rect -9480 -2990 -9262 -716
rect -6220 -800 -6060 920
rect -6230 -940 -6220 -800
rect -6060 -940 -6050 -800
rect -6220 -1040 -6060 -940
rect -6220 -1160 -5540 -1040
rect -10152 -3060 -9848 -3054
rect -10152 -3340 -10140 -3060
rect -9860 -3340 -9848 -3060
rect -10152 -3346 -9848 -3340
rect -4860 -4120 -4680 -1920
rect -3820 -4120 -3640 -1920
rect -2760 -2440 -2600 -1920
rect -1720 -2440 -1560 -1920
rect -700 -1940 -520 -1920
rect 340 -1940 520 -1920
rect 1380 -1940 1560 -1920
rect 2420 -1940 2600 -1920
rect -2780 -4120 -2600 -2440
rect -1740 -4120 -1560 -2440
rect -680 -2460 -520 -1940
rect 360 -2460 520 -1940
rect 1400 -2460 1560 -1940
rect 2440 -2460 2600 -1940
rect -700 -4120 -520 -2460
rect 340 -4120 520 -2460
rect 1380 -4120 1560 -2460
rect 2420 -4120 2600 -2460
rect 3480 -4040 3660 320
rect 7220 -4040 7340 -2680
rect 3480 -4120 7340 -4040
rect -5620 -4220 7340 -4120
rect -8906 -4720 -8154 -4708
rect -8910 -5580 -8900 -4720
rect -8160 -5580 -8150 -4720
rect -5052 -4860 -4608 -4854
rect -5052 -4980 -5040 -4860
rect -4620 -4980 -4608 -4860
rect -5052 -4986 -4608 -4980
rect -872 -4860 -428 -4854
rect -872 -4980 -860 -4860
rect -440 -4980 -428 -4860
rect -872 -4986 -428 -4980
rect 3288 -4860 3792 -4854
rect 3288 -4980 3300 -4860
rect 3780 -4980 3792 -4860
rect 3288 -4986 3792 -4980
rect 7220 -5140 7340 -4220
rect -8906 -5592 -8154 -5580
<< via1 >>
rect -6700 5860 -5400 7500
rect 3280 6960 4100 8220
rect 6640 6560 16540 8320
rect -7100 3680 -6980 4360
rect 1720 4160 3320 4680
rect 7140 1700 7300 2480
rect 12020 2040 12540 2240
rect -7440 740 -7260 820
rect -6220 -940 -6060 -800
rect -10140 -3340 -9860 -3060
rect -8900 -5580 -8160 -4720
rect -5040 -4980 -4620 -4860
rect -860 -4980 -440 -4860
rect 3300 -4980 3780 -4860
<< metal2 >>
rect -10520 8320 16620 8440
rect -10520 8220 6640 8320
rect -10520 7500 3280 8220
rect -10520 6760 -6700 7500
rect -6880 5860 -6700 6760
rect -5400 6960 3280 7500
rect 4100 6960 6640 8220
rect -5400 6760 6640 6960
rect 1660 5880 2720 6760
rect -5400 5860 2720 5880
rect -6880 5220 2720 5860
rect -7100 4360 -6980 4370
rect -10130 3926 -8950 3936
rect -10130 3660 -8950 3670
rect -8944 3928 -7208 3938
rect -8944 3672 -8388 3928
rect -8944 3662 -8080 3672
rect -8944 3660 -8342 3662
rect -7610 3662 -7208 3672
rect -7100 3670 -6980 3680
rect -8080 3650 -7610 3660
rect -6880 3520 -5400 5220
rect 1660 4690 2720 5220
rect 4440 6560 6640 6760
rect 16540 6560 16620 8320
rect 4440 5580 16620 6560
rect 1660 4680 3320 4690
rect 1660 4160 1720 4680
rect 1660 4150 3320 4160
rect 1660 3520 2720 4150
rect -10156 3172 -9754 3182
rect -10156 2640 -9754 2650
rect -9116 3172 -8714 3182
rect -9116 2640 -8714 2650
rect -8084 3168 -7682 3178
rect -8084 2636 -7682 2646
rect -6880 2700 2720 3520
rect 3040 3660 3440 3670
rect 3040 3130 3440 3140
rect -10418 1078 -10330 2402
rect -9552 2288 -8202 2364
rect -6880 2040 -5400 2700
rect 1700 2040 2720 2700
rect -6880 1900 2720 2040
rect -10280 1704 -7440 1742
rect -10280 1452 -9520 1704
rect -9134 1452 -8012 1704
rect -9520 1322 -9134 1374
rect -7636 1452 -7440 1704
rect -7636 1336 -7446 1452
rect -8012 1326 -7446 1336
rect -10168 928 -9766 938
rect -10168 396 -9766 406
rect -10420 -1078 -10330 116
rect -9484 0 -9134 1322
rect -7880 1324 -7446 1326
rect -7880 1270 -7520 1324
rect -6880 1320 2460 1900
rect 2780 1700 2860 2780
rect 4440 2580 6800 5580
rect 3300 2080 3800 2090
rect 4440 2040 4520 2580
rect 6700 2040 6800 2580
rect 4440 1980 6800 2040
rect 7140 2480 7300 2490
rect 3300 1870 3800 1880
rect 12000 2240 12560 2260
rect 12000 2220 12020 2240
rect 12540 2040 12560 2240
rect 12000 2020 12560 2040
rect 7140 1690 7300 1700
rect 2800 1420 3200 1430
rect 2800 890 3200 900
rect -7440 820 -7260 830
rect -7440 738 -7438 740
rect -7262 738 -7260 740
rect -7440 730 -7260 738
rect -7438 728 -7262 730
rect -9520 -488 -9134 0
rect -9660 -498 -9130 -488
rect -9660 -892 -9130 -882
rect -6220 -800 -6060 -790
rect -9520 -972 -9134 -892
rect -6220 -950 -6060 -940
rect -10174 -1320 -9772 -1310
rect -10174 -1852 -9772 -1842
rect -9476 -2252 -9134 -972
rect -9520 -2694 -9134 -2252
rect -9526 -2724 -9134 -2694
rect -9554 -2740 -9134 -2724
rect -9672 -2750 -9134 -2740
rect -10140 -3060 -9860 -3050
rect -9142 -3132 -9134 -2750
rect -9672 -3142 -9134 -3132
rect -10140 -3350 -9860 -3340
rect -9520 -4316 -9134 -3142
rect -5900 -1600 -5760 -540
rect 2520 -620 2600 600
rect 3300 -20 3800 -10
rect 3720 -280 3800 -20
rect 3300 -290 3800 -280
rect -5540 -840 -5140 -830
rect -5540 -1370 -5140 -1360
rect -4500 -840 -4100 -830
rect -4500 -1370 -4100 -1360
rect -3460 -840 -3060 -830
rect -3460 -1370 -3060 -1360
rect -2420 -840 -2020 -830
rect -2420 -1370 -2020 -1360
rect -1380 -840 -980 -830
rect -1380 -1370 -980 -1360
rect -320 -840 80 -830
rect -320 -1370 80 -1360
rect 720 -840 1120 -830
rect 720 -1370 1120 -1360
rect 1760 -840 2160 -830
rect 1760 -1370 2160 -1360
rect 2800 -840 3200 -830
rect 2800 -1370 3200 -1360
rect -5900 -1720 3200 -1600
rect -8860 -3420 -8120 -3410
rect -8320 -3690 -8120 -3420
rect -8860 -3710 -8320 -3700
rect -5900 -3840 -5760 -1720
rect 3300 -2260 3800 -2250
rect -4664 -2270 -4600 -2260
rect -3608 -2270 -3544 -2264
rect -2564 -2270 -2500 -2264
rect -1524 -2270 -1460 -2260
rect -484 -2270 -420 -2264
rect 560 -2270 624 -2264
rect 1600 -2270 1664 -2260
rect 2644 -2270 2708 -2260
rect -5040 -2280 -4600 -2270
rect -4640 -2500 -4600 -2280
rect -5040 -2510 -4600 -2500
rect -3980 -2280 -3544 -2270
rect -3580 -2500 -3544 -2280
rect -3980 -2510 -3544 -2500
rect -2940 -2280 -2500 -2270
rect -2540 -2500 -2500 -2280
rect -2940 -2510 -2500 -2500
rect -1900 -2280 -1460 -2270
rect -1500 -2500 -1460 -2280
rect -1900 -2510 -1460 -2500
rect -860 -2280 -420 -2270
rect -460 -2500 -420 -2280
rect -860 -2510 -420 -2500
rect 180 -2280 624 -2270
rect 580 -2500 624 -2280
rect 180 -2510 624 -2500
rect 1220 -2280 1664 -2270
rect 1620 -2500 1664 -2280
rect 1220 -2510 1664 -2500
rect 2260 -2280 2708 -2270
rect 2660 -2500 2708 -2280
rect 2260 -2510 2708 -2500
rect -4664 -2516 -4600 -2510
rect -3608 -2520 -3544 -2510
rect -2564 -2520 -2500 -2510
rect -1524 -2516 -1460 -2510
rect -484 -2520 -420 -2510
rect 560 -2520 624 -2510
rect 1600 -2516 1664 -2510
rect 2644 -2516 2708 -2510
rect 3720 -2520 3800 -2260
rect 3300 -2530 3800 -2520
rect -5540 -3080 -5140 -3070
rect -5540 -3610 -5140 -3600
rect -4500 -3080 -4100 -3070
rect -4500 -3610 -4100 -3600
rect -3460 -3080 -3060 -3070
rect -3460 -3610 -3060 -3600
rect -2420 -3080 -2020 -3070
rect -2420 -3610 -2020 -3600
rect -1380 -3080 -980 -3070
rect -1380 -3610 -980 -3600
rect -320 -3080 80 -3070
rect -320 -3610 80 -3600
rect 720 -3080 1120 -3070
rect 720 -3610 1120 -3600
rect 1740 -3080 2140 -3070
rect 1740 -3610 2140 -3600
rect 2800 -3080 3200 -3070
rect 2800 -3610 3200 -3600
rect -5900 -3960 3420 -3840
rect -9684 -4326 -9124 -4316
rect -10160 -5420 -9684 -5180
rect -10180 -5512 -9684 -5420
rect -4656 -4510 -4604 -4484
rect -5040 -4520 -4604 -4510
rect -8900 -4720 -8160 -4710
rect -9124 -5512 -8900 -5180
rect -10180 -5580 -8900 -5512
rect -4640 -4792 -4604 -4520
rect -3604 -4530 -3552 -4496
rect -2560 -4530 -2508 -4488
rect -1520 -4530 -1468 -4484
rect -480 -4530 -428 -4496
rect 560 -4530 612 -4488
rect 1600 -4530 1684 -4484
rect 2620 -4530 2704 -4480
rect -3980 -4540 -3552 -4530
rect -4640 -4860 -4620 -4850
rect -3580 -4788 -3552 -4540
rect -2940 -4540 -2508 -4530
rect -3980 -4970 -3580 -4960
rect -2540 -4780 -2508 -4540
rect -1900 -4540 -1468 -4530
rect -2940 -4970 -2540 -4960
rect -1500 -4776 -1468 -4540
rect -860 -4540 -428 -4530
rect -1900 -4970 -1500 -4960
rect -460 -4788 -428 -4540
rect 180 -4540 612 -4530
rect -460 -4860 -440 -4850
rect -5040 -4990 -4620 -4980
rect 580 -4780 612 -4540
rect 1220 -4540 1684 -4530
rect 180 -4970 580 -4960
rect 1620 -4776 1684 -4540
rect 2260 -4540 2704 -4530
rect 1220 -4970 1620 -4960
rect 2660 -4772 2704 -4540
rect 3300 -4540 3800 -4530
rect 2260 -4970 2660 -4960
rect 3720 -4820 3800 -4540
rect 3300 -4860 3780 -4820
rect -860 -4990 -440 -4980
rect 3300 -4990 3780 -4980
rect -8160 -5460 7200 -5180
rect 7260 -5460 7860 -5450
rect -8160 -5580 7260 -5460
rect -10180 -5900 7260 -5580
rect -10180 -7600 -8980 -5900
rect -6180 -7600 7260 -5900
rect -10180 -7820 7260 -7600
rect 7260 -7830 7860 -7820
<< via2 >>
rect -6700 5860 -5400 7500
rect 3280 6960 4100 8220
rect -10130 3670 -8950 3926
rect -8388 3672 -7208 3928
rect -8080 3660 -7610 3672
rect -7100 3860 -6980 4360
rect 6640 6560 16540 8320
rect 1720 4160 3320 4680
rect -10156 2650 -9754 3172
rect -9116 2650 -8714 3172
rect -8084 2646 -7682 3168
rect 3040 3140 3440 3660
rect -9520 1374 -9134 1704
rect -8012 1336 -7636 1704
rect -10168 406 -9766 928
rect 3300 1880 3800 2080
rect 4520 2040 6700 2580
rect 7140 1700 7300 2480
rect 12000 2040 12020 2220
rect 12020 2040 12380 2220
rect 2800 900 3200 1420
rect -7438 740 -7262 810
rect -7438 738 -7262 740
rect -9660 -882 -9130 -498
rect -6220 -940 -6060 -800
rect -10174 -1842 -9772 -1320
rect -10140 -3340 -9860 -3060
rect -9672 -3132 -9142 -2750
rect 3300 -280 3720 -20
rect -5540 -1360 -5140 -840
rect -4500 -1360 -4100 -840
rect -3460 -1360 -3060 -840
rect -2420 -1360 -2020 -840
rect -1380 -1360 -980 -840
rect -320 -1360 80 -840
rect 720 -1360 1120 -840
rect 1760 -1360 2160 -840
rect 2800 -1360 3200 -840
rect -8860 -3700 -8320 -3420
rect -5040 -2500 -4640 -2280
rect -3980 -2500 -3580 -2280
rect -2940 -2500 -2540 -2280
rect -1900 -2500 -1500 -2280
rect -860 -2500 -460 -2280
rect 180 -2500 580 -2280
rect 1220 -2500 1620 -2280
rect 2260 -2500 2660 -2280
rect 3300 -2520 3720 -2260
rect -5540 -3600 -5140 -3080
rect -4500 -3600 -4100 -3080
rect -3460 -3600 -3060 -3080
rect -2420 -3600 -2020 -3080
rect -1380 -3600 -980 -3080
rect -320 -3600 80 -3080
rect 720 -3600 1120 -3080
rect 1740 -3600 2140 -3080
rect 2800 -3600 3200 -3080
rect -9684 -5512 -9124 -4326
rect -8900 -5580 -8160 -4720
rect -5040 -4860 -4640 -4520
rect -5040 -4980 -4620 -4860
rect -3980 -4960 -3580 -4540
rect -2940 -4960 -2540 -4540
rect -1900 -4960 -1500 -4540
rect -860 -4860 -460 -4540
rect -860 -4980 -440 -4860
rect 180 -4960 580 -4540
rect 1220 -4960 1620 -4540
rect 2260 -4960 2660 -4540
rect 3300 -4820 3720 -4540
rect -8980 -7600 -6180 -5900
rect 7260 -7820 7860 -5460
<< metal3 >>
rect 6620 8440 16620 8520
rect -10520 8320 16620 8440
rect -10520 8220 6640 8320
rect -10520 7500 3280 8220
rect -10520 7496 -6700 7500
rect -10522 6762 -6700 7496
rect -10520 6760 -6700 6762
rect -6710 5860 -6700 6760
rect -5400 6960 3280 7500
rect 4100 6960 6640 8220
rect -5400 6760 6640 6960
rect -5400 5860 -5390 6760
rect -6710 5855 -5390 5860
rect -9130 4600 -9120 5060
rect -8820 4600 -8810 5060
rect -7390 4580 -7380 5040
rect -7080 4580 -7070 5040
rect -5130 4620 -5120 5060
rect 1520 4620 1530 5060
rect 1960 4685 3380 6760
rect 1710 4680 3380 4685
rect -7110 4360 -6970 4365
rect -10172 3931 -9748 3980
rect -8080 3933 -7680 3978
rect -10172 3930 -8940 3931
rect -8398 3930 -7198 3933
rect -10172 3928 -7198 3930
rect -10172 3926 -8388 3928
rect -10172 3670 -10130 3926
rect -8950 3672 -8388 3926
rect -7208 3672 -7198 3928
rect -7110 3860 -7100 4360
rect -6980 3860 -6760 4360
rect 1710 4160 1720 4680
rect 3320 4160 3380 4680
rect 1710 4155 3380 4160
rect 1960 4120 3380 4155
rect 4420 6560 6640 6760
rect 16540 6560 16620 8320
rect 4420 6340 16620 6560
rect -7110 3855 -6760 3860
rect -8950 3670 -8080 3672
rect -10172 3667 -8080 3670
rect -10172 3665 -8356 3667
rect -10172 3177 -9748 3665
rect -8972 3664 -8356 3665
rect -8090 3660 -8080 3667
rect -7610 3667 -7198 3672
rect -7610 3660 -7600 3667
rect -8090 3655 -7600 3660
rect -10172 3172 -9744 3177
rect -10174 2650 -10156 3172
rect -9754 3170 -9744 3172
rect -9126 3172 -8704 3177
rect -8080 3173 -7680 3655
rect -7100 3460 -6760 3855
rect -5880 3998 -3696 4000
rect 1380 3998 1460 4000
rect -5880 3540 -5010 3998
rect 2640 3660 2660 4000
rect 3030 3660 3450 3665
rect -5880 3520 1680 3540
rect -9126 3170 -9116 3172
rect -9754 2650 -9116 3170
rect -8714 3170 -8704 3172
rect -8094 3170 -7672 3173
rect -8714 3168 -7672 3170
rect -8714 2650 -8084 3168
rect -10174 2645 -9744 2650
rect -9126 2645 -8704 2650
rect -8094 2646 -8084 2650
rect -7682 2646 -7672 3168
rect -10174 933 -9750 2645
rect -8094 2641 -7672 2646
rect -9682 1709 -7636 1728
rect -9682 1708 -7626 1709
rect -9684 1704 -7626 1708
rect -9684 1700 -9520 1704
rect -9690 1320 -9680 1700
rect -9134 1374 -8012 1704
rect -9140 1336 -8012 1374
rect -7636 1336 -7626 1704
rect -9140 1332 -7626 1336
rect -9140 1320 -9124 1332
rect -8022 1331 -7626 1332
rect -10178 928 -9750 933
rect -10178 406 -10168 928
rect -9766 406 -9750 928
rect -10178 401 -9750 406
rect -10174 -1315 -9750 401
rect -10184 -1320 -9750 -1315
rect -10184 -1842 -10174 -1320
rect -9772 -1842 -9750 -1320
rect -9684 -493 -9124 1320
rect -7448 810 -6728 882
rect -7448 738 -7438 810
rect -7262 802 -6728 810
rect -7262 738 -7252 802
rect -7448 733 -7252 738
rect -8492 384 -8124 510
rect -9684 -498 -9120 -493
rect -9684 -882 -9660 -498
rect -9130 -500 -9120 -498
rect -9120 -880 -9110 -500
rect -9130 -882 -9120 -880
rect -9684 -887 -9120 -882
rect -10184 -1847 -9762 -1842
rect -9684 -2750 -9124 -887
rect -6862 -1220 -6730 802
rect -5880 156 -5240 3520
rect -5100 2774 1540 3422
rect 1680 2780 1720 3520
rect 2640 3140 3040 3660
rect 3440 3140 3450 3660
rect 2640 2780 2660 3140
rect 3030 3135 3450 3140
rect -4718 2160 -4708 2578
rect -4060 2160 -4050 2578
rect -2978 2162 -2968 2580
rect -2320 2162 -2310 2580
rect -1238 2162 -1228 2580
rect -580 2162 -570 2580
rect 502 2162 512 2580
rect 1160 2162 1170 2580
rect 1680 2020 2660 2780
rect 4420 2580 6780 6340
rect 13150 3860 13160 4820
rect 13420 3860 13430 4820
rect 13890 3860 13900 4820
rect 14160 3860 14170 4820
rect 14650 3860 14660 4820
rect 14920 3860 14930 4820
rect 15410 3860 15420 4820
rect 15680 3860 15690 4820
rect 16170 3860 16180 4820
rect 16440 3860 16450 4820
rect 6950 2780 6960 3360
rect 7280 2780 7290 3360
rect 1680 158 1700 2020
rect 2620 1424 2660 2020
rect 3290 2080 3810 2085
rect 3290 1880 3300 2080
rect 3800 1880 3810 2080
rect 3290 1875 3810 1880
rect 4420 2040 4520 2580
rect 6700 2040 6780 2580
rect 2790 1424 3210 1425
rect 2620 1420 3210 1424
rect 2620 900 2800 1420
rect 3200 900 3210 1420
rect -4988 156 -4978 158
rect -5880 120 -4978 156
rect -6230 -800 -6050 -795
rect -6230 -940 -6220 -800
rect -6060 -940 -6050 -800
rect -5880 -800 -5860 120
rect 2620 -200 2660 900
rect 2790 895 3210 900
rect 3300 1320 3800 1875
rect 3300 -15 3720 1320
rect 3290 -20 3730 -15
rect 2620 -300 3200 -200
rect 3290 -280 3300 -20
rect 3720 -280 3730 -20
rect 3290 -285 3730 -280
rect 2600 -800 3200 -300
rect -5880 -820 3200 -800
rect -5860 -835 3200 -820
rect -5860 -840 3210 -835
rect -5860 -900 -5540 -840
rect -6230 -945 -6050 -940
rect -6220 -1220 -6060 -945
rect -6862 -1340 -6060 -1220
rect -8840 -1440 -8700 -1380
rect -6862 -1400 -6140 -1340
rect -5550 -1360 -5540 -900
rect -5140 -900 -4500 -840
rect -5140 -1360 -5130 -900
rect -5550 -1365 -5130 -1360
rect -4510 -1360 -4500 -900
rect -4100 -900 -3460 -840
rect -4100 -1360 -4090 -900
rect -4510 -1365 -4090 -1360
rect -3470 -1360 -3460 -900
rect -3060 -900 -2420 -840
rect -3060 -1360 -3050 -900
rect -3470 -1365 -3050 -1360
rect -2430 -1360 -2420 -900
rect -2020 -900 -1380 -840
rect -2020 -1360 -2010 -900
rect -2430 -1365 -2010 -1360
rect -1390 -1360 -1380 -900
rect -980 -900 -320 -840
rect -980 -1360 -970 -900
rect -1390 -1365 -970 -1360
rect -330 -1360 -320 -900
rect 80 -900 720 -840
rect 80 -1360 90 -900
rect -330 -1365 90 -1360
rect 710 -1360 720 -900
rect 1120 -900 1760 -840
rect 1120 -1360 1130 -900
rect 710 -1365 1130 -1360
rect 1740 -1360 1760 -900
rect 2160 -900 2800 -840
rect 2160 -1360 2170 -900
rect 1740 -1365 2170 -1360
rect 2790 -1360 2800 -900
rect 3200 -1360 3210 -840
rect 2790 -1365 3210 -1360
rect -6862 -1926 -6730 -1400
rect -10150 -3060 -9850 -3055
rect -10150 -3340 -10140 -3060
rect -9860 -3340 -9850 -3060
rect -10150 -3345 -9850 -3340
rect -9684 -3132 -9672 -2750
rect -9142 -3132 -9124 -2750
rect -5540 -3075 -5140 -1365
rect -5040 -2275 -4640 -2240
rect -5050 -2280 -4630 -2275
rect -5050 -2500 -5040 -2280
rect -4640 -2500 -4630 -2280
rect -5050 -2505 -4630 -2500
rect -9684 -4321 -9124 -3132
rect -5550 -3080 -5130 -3075
rect -8870 -3420 -8310 -3415
rect -8870 -4040 -8860 -3420
rect -8320 -4040 -8310 -3420
rect -5550 -3600 -5540 -3080
rect -5140 -3600 -5130 -3080
rect -5550 -3605 -5130 -3600
rect -9694 -4326 -9114 -4321
rect -9694 -5512 -9684 -4326
rect -9124 -5512 -9114 -4326
rect -5040 -4515 -4640 -2505
rect -4500 -3075 -4100 -1365
rect -3980 -2275 -3580 -2240
rect -3990 -2280 -3570 -2275
rect -3990 -2500 -3980 -2280
rect -3580 -2500 -3570 -2280
rect -3990 -2505 -3570 -2500
rect -4510 -3080 -4090 -3075
rect -4510 -3600 -4500 -3080
rect -4100 -3600 -4090 -3080
rect -4510 -3605 -4090 -3600
rect -5050 -4520 -4630 -4515
rect -9694 -5517 -9114 -5512
rect -8910 -4720 -8150 -4715
rect -8910 -5580 -8900 -4720
rect -8160 -5580 -8150 -4720
rect -5050 -4980 -5040 -4520
rect -4640 -4855 -4630 -4520
rect -3980 -4535 -3580 -2505
rect -3460 -3075 -3060 -1365
rect -2940 -2275 -2540 -2240
rect -2950 -2280 -2530 -2275
rect -2950 -2500 -2940 -2280
rect -2540 -2500 -2530 -2280
rect -2950 -2505 -2530 -2500
rect -3470 -3080 -3050 -3075
rect -3470 -3600 -3460 -3080
rect -3060 -3600 -3050 -3080
rect -3470 -3605 -3050 -3600
rect -2940 -4535 -2540 -2505
rect -2420 -3075 -2020 -1365
rect -1900 -2275 -1500 -2240
rect -1910 -2280 -1490 -2275
rect -1910 -2500 -1900 -2280
rect -1500 -2500 -1490 -2280
rect -1910 -2505 -1490 -2500
rect -2430 -3080 -2010 -3075
rect -2430 -3600 -2420 -3080
rect -2020 -3600 -2010 -3080
rect -2430 -3605 -2010 -3600
rect -1900 -4535 -1500 -2505
rect -1380 -3075 -980 -1365
rect -860 -2275 -460 -2240
rect -870 -2280 -450 -2275
rect -870 -2500 -860 -2280
rect -460 -2500 -450 -2280
rect -870 -2505 -450 -2500
rect -1390 -3080 -970 -3075
rect -1390 -3600 -1380 -3080
rect -980 -3600 -970 -3080
rect -1390 -3605 -970 -3600
rect -860 -4535 -460 -2505
rect -320 -3075 80 -1365
rect 180 -2275 580 -2240
rect 170 -2280 590 -2275
rect 170 -2500 180 -2280
rect 580 -2500 590 -2280
rect 170 -2505 590 -2500
rect -330 -3080 90 -3075
rect -330 -3600 -320 -3080
rect 80 -3600 90 -3080
rect -330 -3605 90 -3600
rect 180 -4535 580 -2505
rect 720 -3075 1120 -1365
rect 1220 -2275 1620 -2240
rect 1210 -2280 1630 -2275
rect 1210 -2500 1220 -2280
rect 1620 -2500 1630 -2280
rect 1210 -2505 1630 -2500
rect 710 -3080 1130 -3075
rect 710 -3600 720 -3080
rect 1120 -3600 1130 -3080
rect 710 -3605 1130 -3600
rect 1220 -4535 1620 -2505
rect 1740 -3075 2140 -1365
rect 2260 -2275 2660 -2240
rect 2250 -2280 2670 -2275
rect 2250 -2500 2260 -2280
rect 2660 -2500 2670 -2280
rect 2250 -2505 2670 -2500
rect 1730 -3080 2150 -3075
rect 1730 -3600 1740 -3080
rect 2140 -3600 2150 -3080
rect 1730 -3605 2150 -3600
rect 2260 -4535 2660 -2505
rect 2800 -3075 3200 -1365
rect 3300 -2255 3720 -285
rect 4420 -1420 6780 2040
rect 6960 2485 7280 2780
rect 6960 2480 7310 2485
rect 6960 1700 7140 2480
rect 7300 1700 7310 2480
rect 7950 2340 7960 3300
rect 8220 2340 8230 3300
rect 8690 2340 8700 3300
rect 8960 2340 8970 3300
rect 9450 2340 9460 3300
rect 9720 2340 9730 3300
rect 10210 2340 10220 3300
rect 10480 2340 10490 3300
rect 10970 2340 10980 3300
rect 11240 2340 11250 3300
rect 11990 2220 12390 2225
rect 11990 2040 12000 2220
rect 12380 2040 12390 2220
rect 11990 2035 12390 2040
rect 7130 1695 7310 1700
rect 3290 -2260 3730 -2255
rect 3290 -2520 3300 -2260
rect 3720 -2520 3730 -2260
rect 3290 -2525 3730 -2520
rect 2790 -3080 3210 -3075
rect 2790 -3600 2800 -3080
rect 3200 -3600 3210 -3080
rect 2790 -3605 3210 -3600
rect 3300 -4535 3720 -2525
rect -3990 -4540 -3570 -4535
rect -4640 -4860 -4610 -4855
rect -4620 -4980 -4610 -4860
rect -3990 -4960 -3980 -4540
rect -3580 -4960 -3570 -4540
rect -3990 -4965 -3570 -4960
rect -2950 -4540 -2530 -4535
rect -2950 -4960 -2940 -4540
rect -2540 -4960 -2530 -4540
rect -2950 -4965 -2530 -4960
rect -1910 -4540 -1490 -4535
rect -1910 -4960 -1900 -4540
rect -1500 -4960 -1490 -4540
rect -1910 -4965 -1490 -4960
rect -870 -4540 -450 -4535
rect -5050 -4985 -4610 -4980
rect -870 -4980 -860 -4540
rect -460 -4855 -450 -4540
rect 170 -4540 590 -4535
rect -460 -4860 -430 -4855
rect -440 -4980 -430 -4860
rect 170 -4960 180 -4540
rect 580 -4960 590 -4540
rect 170 -4965 590 -4960
rect 1210 -4540 1630 -4535
rect 1210 -4960 1220 -4540
rect 1620 -4960 1630 -4540
rect 1210 -4965 1630 -4960
rect 2250 -4540 2670 -4535
rect 2250 -4960 2260 -4540
rect 2660 -4960 2670 -4540
rect 3290 -4540 3730 -4535
rect 3290 -4820 3300 -4540
rect 3720 -4820 3730 -4540
rect 3290 -4825 3730 -4820
rect 2250 -4965 2670 -4960
rect -870 -4985 -430 -4980
rect -8910 -5585 -8150 -5580
rect 4240 -5780 5980 -3680
rect 7250 -5460 7870 -5455
rect -8990 -5900 -6170 -5895
rect -8990 -7600 -8980 -5900
rect -6180 -7600 -6170 -5900
rect -80 -7220 1620 -5920
rect -8990 -7605 -6170 -7600
rect 7250 -7820 7260 -5460
rect 7860 -6200 7870 -5460
rect 7860 -7380 16180 -6200
rect 7860 -7740 8080 -7380
rect 16060 -7740 16180 -7380
rect 7860 -7820 16180 -7740
rect 7250 -7825 7870 -7820
<< via3 >>
rect -6700 5860 -5400 7500
rect -9120 4600 -8820 5060
rect -7380 4580 -7080 5040
rect -5120 4620 1520 5060
rect 1460 3998 2640 4000
rect -5010 3540 2640 3998
rect 1680 3520 2640 3540
rect -9680 1374 -9520 1700
rect -9520 1374 -9140 1700
rect -9680 1320 -9140 1374
rect -8012 1336 -7636 1704
rect -9660 -880 -9130 -500
rect -9130 -880 -9120 -500
rect 1720 2780 2640 3520
rect -4708 2160 -4060 2578
rect -2968 2162 -2320 2580
rect -1228 2162 -580 2580
rect 512 2162 1160 2580
rect 13160 3860 13420 4820
rect 13900 3860 14160 4820
rect 14660 3860 14920 4820
rect 15420 3860 15680 4820
rect 16180 3860 16440 4820
rect 6960 2780 7280 3360
rect 1700 158 2620 2020
rect -4978 120 2620 158
rect -5860 -300 2620 120
rect -5860 -800 2600 -300
rect -10140 -3340 -9860 -3060
rect -9660 -3120 -9160 -2760
rect -8860 -3700 -8320 -3420
rect -8860 -4040 -8320 -3700
rect -9684 -5512 -9124 -4326
rect -8900 -5580 -8160 -4720
rect -5040 -4960 -4640 -4600
rect 7960 2340 8220 3300
rect 8700 2340 8960 3300
rect 9460 2340 9720 3300
rect 10220 2340 10480 3300
rect 10980 2340 11240 3300
rect 12000 2040 12380 2220
rect -3980 -4960 -3580 -4600
rect -2940 -4960 -2540 -4600
rect -1900 -4960 -1500 -4600
rect -860 -4960 -460 -4600
rect 180 -4960 580 -4600
rect 1220 -4960 1620 -4600
rect 2260 -4960 2660 -4600
rect 3300 -4820 3720 -4600
rect -8980 -7600 -6180 -5900
rect 7260 -7820 7860 -5460
rect 8080 -7740 16060 -7380
<< metal4 >>
rect -6701 7500 -5399 7501
rect -6701 5860 -6700 7500
rect -5400 5860 -5399 7500
rect -6701 5859 -5399 5860
rect -9120 5736 -5300 5740
rect -9120 5320 -5286 5736
rect -9120 5061 -8760 5320
rect -9121 5060 -8760 5061
rect -9121 4600 -9120 5060
rect -8820 4600 -8760 5060
rect -7381 5040 -7079 5041
rect -9121 4599 -8819 4600
rect -7381 4580 -7380 5040
rect -7080 5018 -5620 5040
rect -7080 4580 -5618 5018
rect -7381 4579 -7079 4580
rect -10200 1701 -9140 1720
rect -8013 1704 -7635 1705
rect -10200 1700 -9139 1701
rect -10200 1320 -9680 1700
rect -9140 1320 -8994 1700
rect -8013 1336 -8012 1704
rect -7636 1700 -7635 1704
rect -7636 1336 -6100 1700
rect -8013 1335 -6100 1336
rect -10200 840 -8994 1320
rect -8012 840 -6100 1335
rect -10200 -499 -9140 840
rect -10200 -500 -9119 -499
rect -10200 -880 -9660 -500
rect -9120 -880 -9119 -500
rect -10200 -881 -9119 -880
rect -10200 -2760 -9140 -881
rect -6760 -1960 -6100 840
rect -5942 556 -5618 4580
rect -5546 4402 -5286 5320
rect -5121 5060 1521 5061
rect -5121 4620 -5120 5060
rect 1520 4620 3960 5060
rect -5121 4619 1521 4620
rect -5546 4128 -4930 4402
rect 1834 4001 2318 4004
rect 1459 4000 2641 4001
rect 1459 3999 1460 4000
rect -5011 3998 1460 3999
rect -5011 3540 -5010 3998
rect -5011 3520 1680 3540
rect -5011 3514 1720 3520
rect 1680 2780 1720 3514
rect 2640 2780 2660 4000
rect 3580 3360 3960 4620
rect 13140 4820 17040 4840
rect 13140 3860 13160 4820
rect 13420 3860 13900 4820
rect 14160 3860 14660 4820
rect 14920 3860 15420 4820
rect 15680 3860 16180 4820
rect 16440 3860 17040 4820
rect 13140 3840 17040 3860
rect 6959 3360 7281 3361
rect 3580 2900 6960 3360
rect 1680 2740 2660 2780
rect 6959 2780 6960 2900
rect 7280 2780 7281 3360
rect 6959 2779 7281 2780
rect 7940 3300 17040 3320
rect -4720 2580 7200 2600
rect -4720 2578 -2968 2580
rect -4720 2160 -4708 2578
rect -4060 2162 -2968 2578
rect -2320 2162 -1228 2580
rect -580 2162 512 2580
rect 1160 2162 7200 2580
rect 7940 2340 7960 3300
rect 8220 2340 8700 3300
rect 8960 2340 9460 3300
rect 9720 2340 10220 3300
rect 10480 2340 10980 3300
rect 11240 2340 17040 3300
rect 7940 2320 17040 2340
rect -4060 2160 7200 2162
rect -4720 2140 7200 2160
rect 1699 2020 2621 2021
rect -5946 282 -3652 556
rect 1699 159 1700 2020
rect -4979 158 1700 159
rect -4979 121 -4978 158
rect -5861 120 -4978 121
rect -5861 -260 -5860 120
rect -5880 -800 -5860 -260
rect 2620 -300 2621 2020
rect 6820 1680 7200 2140
rect 11999 2220 12381 2221
rect 11999 2040 12000 2220
rect 12380 2040 12381 2220
rect 11999 2039 12381 2040
rect 12000 1680 12380 2039
rect 6820 1320 12380 1680
rect 2600 -301 2621 -300
rect 2600 -800 2620 -301
rect -5880 -820 2620 -800
rect -10200 -3060 -9660 -2760
rect -10200 -3340 -10140 -3060
rect -9860 -3120 -9660 -3060
rect -9160 -3120 -9140 -2760
rect -9860 -3340 -9140 -3120
rect -10200 -3380 -9140 -3340
rect -10200 -3419 -8320 -3380
rect -10200 -3420 -8319 -3419
rect -10200 -4040 -8860 -3420
rect -8320 -4040 -8319 -3420
rect -10200 -4041 -8319 -4040
rect -10200 -4100 -8320 -4041
rect -10200 -4325 -9140 -4100
rect -10200 -4326 -9123 -4325
rect -10200 -5512 -9684 -4326
rect -9124 -4598 -9123 -4326
rect -7100 -4598 -6380 -4280
rect -9124 -4600 -6020 -4598
rect -5500 -4600 3872 -4598
rect -9124 -4720 -5040 -4600
rect -9124 -5512 -8900 -4720
rect -10200 -5580 -8900 -5512
rect -8160 -4960 -5040 -4720
rect -4640 -4960 -3980 -4600
rect -3580 -4960 -2940 -4600
rect -2540 -4960 -1900 -4600
rect -1500 -4960 -860 -4600
rect -460 -4960 180 -4600
rect 580 -4960 1220 -4600
rect 1620 -4960 2260 -4600
rect 2660 -4820 3300 -4600
rect 3720 -4820 3920 -4600
rect 2660 -4960 3920 -4820
rect -8160 -5200 3920 -4960
rect 4280 -5200 6100 -2640
rect -8160 -5460 16180 -5200
rect -8160 -5580 7260 -5460
rect -10200 -5900 7260 -5580
rect -10200 -7600 -8980 -5900
rect -6180 -7600 7260 -5900
rect -10200 -7800 7260 -7600
rect -10180 -7820 7260 -7800
rect 7860 -7380 16180 -5460
rect 7860 -7740 8080 -7380
rect 16060 -7740 16180 -7380
rect 7860 -7820 16180 -7740
rect 7259 -7821 7861 -7820
use outd_curm  outd_curm_0
timestamp 1683888831
transform 1 0 2816 0 1 952
box -40 916 1002 3158
use outd_curm  outd_curm_1
timestamp 1683888831
transform 1 0 -9340 0 1 464
box -40 916 1002 3158
use outd_curm  outd_curm_2
timestamp 1683888831
transform 1 0 -8300 0 1 464
box -40 916 1002 3158
use outd_curm  outd_curm_3
timestamp 1683888831
transform 1 0 -10380 0 1 -1776
box -40 916 1002 3158
use outd_curm  outd_curm_4
timestamp 1683888831
transform 1 0 -10382 0 1 -4020
box -40 916 1002 3158
use outd_curm  outd_curm_5
timestamp 1683888831
transform 1 0 492 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_6
timestamp 1683888831
transform 1 0 -1592 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_7
timestamp 1683888831
transform 1 0 -2634 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_8
timestamp 1683888831
transform 1 0 -4718 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_9
timestamp 1683888831
transform 1 0 -10380 0 1 464
box -40 916 1002 3158
use outd_curm  outd_curm_10
timestamp 1683888831
transform 1 0 -5760 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_11
timestamp 1683888831
transform 1 0 -3676 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_12
timestamp 1683888831
transform 1 0 -2634 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_13
timestamp 1683888831
transform 1 0 -1592 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_14
timestamp 1683888831
transform 1 0 2576 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_15
timestamp 1683888831
transform 1 0 -550 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_16
timestamp 1683888831
transform 1 0 2576 0 1 -1292
box -40 916 1002 3158
use outd_curm  outd_curm_17
timestamp 1683888831
transform 1 0 1534 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_18
timestamp 1683888831
transform 1 0 -550 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_19
timestamp 1683888831
transform 1 0 492 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_20
timestamp 1683888831
transform 1 0 1534 0 1 -5776
box -40 916 1002 3158
use outd_curm  outd_curm_21
timestamp 1683888831
transform 1 0 -5760 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_22
timestamp 1683888831
transform 1 0 -3676 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_23
timestamp 1683888831
transform 1 0 -4718 0 1 -3534
box -40 916 1002 3158
use outd_curm  outd_curm_24
timestamp 1683888831
transform 1 0 2576 0 1 -5776
box -40 916 1002 3158
use outd_diffamp_12  outd_diffamp_12_0
timestamp 1689773955
transform 1 0 -10340 0 1 3600
box -80 20 1668 3804
use outd_diffamp_12  outd_diffamp_12_1
timestamp 1689773955
transform 1 0 -8600 0 1 3600
box -80 20 1668 3804
use outd_diffamp_50ohm_top  outd_diffamp_50ohm_top_0
timestamp 1687207134
transform 1 0 518 0 1 -202
box 6740 -7100 16178 6720
use outd_diffamp_quad  outd_diffamp_quad_0
timestamp 1689773955
transform 1 0 -498 0 1 -3820
box -4760 3612 2208 7404
use outd_diffamp_quad  outd_diffamp_quad_2
timestamp 1689773955
transform 1 0 -530 0 1 24
box -4760 3612 2208 7404
use outd_filter  outd_filter_0
timestamp 1684930430
transform 1 0 -12000 0 1 -4650
box 2696 870 5300 5940
use sky130_fd_pr__cap_mim_m3_1_2YC3NK  sky130_fd_pr__cap_mim_m3_1_2YC3NK_0
timestamp 1685108691
transform 1 0 5626 0 1 -1920
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_2YC3NK  sky130_fd_pr__cap_mim_m3_1_2YC3NK_1
timestamp 1685108691
transform 0 1 -2380 -1 0 -6894
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_2YC3NK  sky130_fd_pr__cap_mim_m3_1_2YC3NK_2
timestamp 1685108691
transform 0 1 3940 -1 0 -6894
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_0
timestamp 1684833579
transform 0 -1 -6652 1 0 2380
box -1186 -640 1186 640
use sky130_fd_pr__cap_mim_m3_1_5KPPX9  sky130_fd_pr__cap_mim_m3_1_5KPPX9_0
timestamp 1684929745
transform 1 0 -6834 0 1 -2880
box -1186 -1640 1186 1640
<< labels >>
rlabel metal4 -9960 -6980 -9240 -4660 1 VN
port 4 n
rlabel metal1 -10318 3778 -10268 4194 1 InputSignal
port 5 n
rlabel metal3 -7068 3922 -6994 4080 1 InputRef
port 6 n
rlabel metal3 -10306 7624 -9980 7986 1 VP
port 7 n
rlabel metal3 -8412 406 -8214 500 1 I_Bias
port 8 n
rlabel metal4 -5340 4200 -5220 4300 1 V_da2_P
rlabel metal4 -5200 340 -5140 460 1 V_da2_N
rlabel metal4 3980 2280 4120 2440 1 V_da3_N
rlabel metal3 -8840 -1440 -8700 -1380 1 VM18D
rlabel metal1 -6040 -1140 -5920 -1060 1 VM6D
rlabel metal4 3776 3042 3904 3208 1 V_da3_P
rlabel metal4 16720 2580 16920 3060 1 OutP
port 9 n
rlabel metal4 16700 4040 16900 4520 1 OutN
port 10 n
<< end >>
