magic
tech sky130A
magscale 1 2
timestamp 1685110944
<< pwell >>
rect -1063 -2082 1063 2082
<< psubdiff >>
rect -1027 2012 -931 2046
rect 931 2012 1027 2046
rect -1027 1950 -993 2012
rect 993 1950 1027 2012
rect -1027 -2012 -993 -1950
rect 993 -2012 1027 -1950
rect -1027 -2046 -931 -2012
rect 931 -2046 1027 -2012
<< psubdiffcont >>
rect -931 2012 931 2046
rect -1027 -1950 -993 1950
rect 993 -1950 1027 1950
rect -931 -2046 931 -2012
<< xpolycontact >>
rect -897 1484 -615 1916
rect -897 52 -615 484
rect -519 1484 -237 1916
rect -519 52 -237 484
rect -141 1484 141 1916
rect -141 52 141 484
rect 237 1484 519 1916
rect 237 52 519 484
rect 615 1484 897 1916
rect 615 52 897 484
rect -897 -484 -615 -52
rect -897 -1916 -615 -1484
rect -519 -484 -237 -52
rect -519 -1916 -237 -1484
rect -141 -484 141 -52
rect -141 -1916 141 -1484
rect 237 -484 519 -52
rect 237 -1916 519 -1484
rect 615 -484 897 -52
rect 615 -1916 897 -1484
<< ppolyres >>
rect -897 484 -615 1484
rect -519 484 -237 1484
rect -141 484 141 1484
rect 237 484 519 1484
rect 615 484 897 1484
rect -897 -1484 -615 -484
rect -519 -1484 -237 -484
rect -141 -1484 141 -484
rect 237 -1484 519 -484
rect 615 -1484 897 -484
<< locali >>
rect -1027 2012 -931 2046
rect 931 2012 1027 2046
rect -1027 1950 -993 2012
rect 993 1950 1027 2012
rect -1027 -2012 -993 -1950
rect 993 -2012 1027 -1950
rect -1027 -2046 -931 -2012
rect 931 -2046 1027 -2012
<< viali >>
rect -881 1501 -631 1898
rect -503 1501 -253 1898
rect -125 1501 125 1898
rect 253 1501 503 1898
rect 631 1501 881 1898
rect -881 70 -631 467
rect -503 70 -253 467
rect -125 70 125 467
rect 253 70 503 467
rect 631 70 881 467
rect -881 -467 -631 -70
rect -503 -467 -253 -70
rect -125 -467 125 -70
rect 253 -467 503 -70
rect 631 -467 881 -70
rect -881 -1898 -631 -1501
rect -503 -1898 -253 -1501
rect -125 -1898 125 -1501
rect 253 -1898 503 -1501
rect 631 -1898 881 -1501
<< metal1 >>
rect -887 1898 -625 1910
rect -887 1501 -881 1898
rect -631 1501 -625 1898
rect -887 1489 -625 1501
rect -509 1898 -247 1910
rect -509 1501 -503 1898
rect -253 1501 -247 1898
rect -509 1489 -247 1501
rect -131 1898 131 1910
rect -131 1501 -125 1898
rect 125 1501 131 1898
rect -131 1489 131 1501
rect 247 1898 509 1910
rect 247 1501 253 1898
rect 503 1501 509 1898
rect 247 1489 509 1501
rect 625 1898 887 1910
rect 625 1501 631 1898
rect 881 1501 887 1898
rect 625 1489 887 1501
rect -887 467 -625 479
rect -887 70 -881 467
rect -631 70 -625 467
rect -887 58 -625 70
rect -509 467 -247 479
rect -509 70 -503 467
rect -253 70 -247 467
rect -509 58 -247 70
rect -131 467 131 479
rect -131 70 -125 467
rect 125 70 131 467
rect -131 58 131 70
rect 247 467 509 479
rect 247 70 253 467
rect 503 70 509 467
rect 247 58 509 70
rect 625 467 887 479
rect 625 70 631 467
rect 881 70 887 467
rect 625 58 887 70
rect -887 -70 -625 -58
rect -887 -467 -881 -70
rect -631 -467 -625 -70
rect -887 -479 -625 -467
rect -509 -70 -247 -58
rect -509 -467 -503 -70
rect -253 -467 -247 -70
rect -509 -479 -247 -467
rect -131 -70 131 -58
rect -131 -467 -125 -70
rect 125 -467 131 -70
rect -131 -479 131 -467
rect 247 -70 509 -58
rect 247 -467 253 -70
rect 503 -467 509 -70
rect 247 -479 509 -467
rect 625 -70 887 -58
rect 625 -467 631 -70
rect 881 -467 887 -70
rect 625 -479 887 -467
rect -887 -1501 -625 -1489
rect -887 -1898 -881 -1501
rect -631 -1898 -625 -1501
rect -887 -1910 -625 -1898
rect -509 -1501 -247 -1489
rect -509 -1898 -503 -1501
rect -253 -1898 -247 -1501
rect -509 -1910 -247 -1898
rect -131 -1501 131 -1489
rect -131 -1898 -125 -1501
rect 125 -1898 131 -1501
rect -131 -1910 131 -1898
rect 247 -1501 509 -1489
rect 247 -1898 253 -1501
rect 503 -1898 509 -1501
rect 247 -1910 509 -1898
rect 625 -1501 887 -1489
rect 625 -1898 631 -1501
rect 881 -1898 887 -1501
rect 625 -1910 887 -1898
<< res1p41 >>
rect -899 482 -613 1486
rect -521 482 -235 1486
rect -143 482 143 1486
rect 235 482 521 1486
rect 613 482 899 1486
rect -899 -1486 -613 -482
rect -521 -1486 -235 -482
rect -143 -1486 143 -482
rect 235 -1486 521 -482
rect 613 -1486 899 -482
<< properties >>
string FIXED_BBOX -1010 -2029 1010 2029
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.41 l 5.0 m 2 nx 5 wmin 1.410 lmin 0.50 rho 319.8 val 1.41k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
