magic
tech sky130A
magscale 1 2
timestamp 1683537326
<< error_p >>
rect -845 890 -787 896
rect -653 890 -595 896
rect -461 890 -403 896
rect -269 890 -211 896
rect -77 890 -19 896
rect 115 890 173 896
rect 307 890 365 896
rect 499 890 557 896
rect 691 890 749 896
rect 883 890 941 896
rect -845 856 -833 890
rect -653 856 -641 890
rect -461 856 -449 890
rect -269 856 -257 890
rect -77 856 -65 890
rect 115 856 127 890
rect 307 856 319 890
rect 499 856 511 890
rect 691 856 703 890
rect 883 856 895 890
rect -845 850 -787 856
rect -653 850 -595 856
rect -461 850 -403 856
rect -269 850 -211 856
rect -77 850 -19 856
rect 115 850 173 856
rect 307 850 365 856
rect 499 850 557 856
rect 691 850 749 856
rect 883 850 941 856
rect -941 380 -883 386
rect -749 380 -691 386
rect -557 380 -499 386
rect -365 380 -307 386
rect -173 380 -115 386
rect 19 380 77 386
rect 211 380 269 386
rect 403 380 461 386
rect 595 380 653 386
rect 787 380 845 386
rect -941 346 -929 380
rect -749 346 -737 380
rect -557 346 -545 380
rect -365 346 -353 380
rect -173 346 -161 380
rect 19 346 31 380
rect 211 346 223 380
rect 403 346 415 380
rect 595 346 607 380
rect 787 346 799 380
rect -941 340 -883 346
rect -749 340 -691 346
rect -557 340 -499 346
rect -365 340 -307 346
rect -173 340 -115 346
rect 19 340 77 346
rect 211 340 269 346
rect 403 340 461 346
rect 595 340 653 346
rect 787 340 845 346
rect -941 272 -883 278
rect -749 272 -691 278
rect -557 272 -499 278
rect -365 272 -307 278
rect -173 272 -115 278
rect 19 272 77 278
rect 211 272 269 278
rect 403 272 461 278
rect 595 272 653 278
rect 787 272 845 278
rect -941 238 -929 272
rect -749 238 -737 272
rect -557 238 -545 272
rect -365 238 -353 272
rect -173 238 -161 272
rect 19 238 31 272
rect 211 238 223 272
rect 403 238 415 272
rect 595 238 607 272
rect 787 238 799 272
rect -941 232 -883 238
rect -749 232 -691 238
rect -557 232 -499 238
rect -365 232 -307 238
rect -173 232 -115 238
rect 19 232 77 238
rect 211 232 269 238
rect 403 232 461 238
rect 595 232 653 238
rect 787 232 845 238
rect -845 -238 -787 -232
rect -653 -238 -595 -232
rect -461 -238 -403 -232
rect -269 -238 -211 -232
rect -77 -238 -19 -232
rect 115 -238 173 -232
rect 307 -238 365 -232
rect 499 -238 557 -232
rect 691 -238 749 -232
rect 883 -238 941 -232
rect -845 -272 -833 -238
rect -653 -272 -641 -238
rect -461 -272 -449 -238
rect -269 -272 -257 -238
rect -77 -272 -65 -238
rect 115 -272 127 -238
rect 307 -272 319 -238
rect 499 -272 511 -238
rect 691 -272 703 -238
rect 883 -272 895 -238
rect -845 -278 -787 -272
rect -653 -278 -595 -272
rect -461 -278 -403 -272
rect -269 -278 -211 -272
rect -77 -278 -19 -272
rect 115 -278 173 -272
rect 307 -278 365 -272
rect 499 -278 557 -272
rect 691 -278 749 -272
rect 883 -278 941 -272
rect -845 -346 -787 -340
rect -653 -346 -595 -340
rect -461 -346 -403 -340
rect -269 -346 -211 -340
rect -77 -346 -19 -340
rect 115 -346 173 -340
rect 307 -346 365 -340
rect 499 -346 557 -340
rect 691 -346 749 -340
rect 883 -346 941 -340
rect -845 -380 -833 -346
rect -653 -380 -641 -346
rect -461 -380 -449 -346
rect -269 -380 -257 -346
rect -77 -380 -65 -346
rect 115 -380 127 -346
rect 307 -380 319 -346
rect 499 -380 511 -346
rect 691 -380 703 -346
rect 883 -380 895 -346
rect -845 -386 -787 -380
rect -653 -386 -595 -380
rect -461 -386 -403 -380
rect -269 -386 -211 -380
rect -77 -386 -19 -380
rect 115 -386 173 -380
rect 307 -386 365 -380
rect 499 -386 557 -380
rect 691 -386 749 -380
rect 883 -386 941 -380
rect -941 -856 -883 -850
rect -749 -856 -691 -850
rect -557 -856 -499 -850
rect -365 -856 -307 -850
rect -173 -856 -115 -850
rect 19 -856 77 -850
rect 211 -856 269 -850
rect 403 -856 461 -850
rect 595 -856 653 -850
rect 787 -856 845 -850
rect -941 -890 -929 -856
rect -749 -890 -737 -856
rect -557 -890 -545 -856
rect -365 -890 -353 -856
rect -173 -890 -161 -856
rect 19 -890 31 -856
rect 211 -890 223 -856
rect 403 -890 415 -856
rect 595 -890 607 -856
rect 787 -890 799 -856
rect -941 -896 -883 -890
rect -749 -896 -691 -890
rect -557 -896 -499 -890
rect -365 -896 -307 -890
rect -173 -896 -115 -890
rect 19 -896 77 -890
rect 211 -896 269 -890
rect 403 -896 461 -890
rect 595 -896 653 -890
rect 787 -896 845 -890
<< pwell >>
rect -1127 -1028 1127 1028
<< nmoslvt >>
rect -927 418 -897 818
rect -831 418 -801 818
rect -735 418 -705 818
rect -639 418 -609 818
rect -543 418 -513 818
rect -447 418 -417 818
rect -351 418 -321 818
rect -255 418 -225 818
rect -159 418 -129 818
rect -63 418 -33 818
rect 33 418 63 818
rect 129 418 159 818
rect 225 418 255 818
rect 321 418 351 818
rect 417 418 447 818
rect 513 418 543 818
rect 609 418 639 818
rect 705 418 735 818
rect 801 418 831 818
rect 897 418 927 818
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
rect -927 -818 -897 -418
rect -831 -818 -801 -418
rect -735 -818 -705 -418
rect -639 -818 -609 -418
rect -543 -818 -513 -418
rect -447 -818 -417 -418
rect -351 -818 -321 -418
rect -255 -818 -225 -418
rect -159 -818 -129 -418
rect -63 -818 -33 -418
rect 33 -818 63 -418
rect 129 -818 159 -418
rect 225 -818 255 -418
rect 321 -818 351 -418
rect 417 -818 447 -418
rect 513 -818 543 -418
rect 609 -818 639 -418
rect 705 -818 735 -418
rect 801 -818 831 -418
rect 897 -818 927 -418
<< ndiff >>
rect -989 806 -927 818
rect -989 430 -977 806
rect -943 430 -927 806
rect -989 418 -927 430
rect -897 806 -831 818
rect -897 430 -881 806
rect -847 430 -831 806
rect -897 418 -831 430
rect -801 806 -735 818
rect -801 430 -785 806
rect -751 430 -735 806
rect -801 418 -735 430
rect -705 806 -639 818
rect -705 430 -689 806
rect -655 430 -639 806
rect -705 418 -639 430
rect -609 806 -543 818
rect -609 430 -593 806
rect -559 430 -543 806
rect -609 418 -543 430
rect -513 806 -447 818
rect -513 430 -497 806
rect -463 430 -447 806
rect -513 418 -447 430
rect -417 806 -351 818
rect -417 430 -401 806
rect -367 430 -351 806
rect -417 418 -351 430
rect -321 806 -255 818
rect -321 430 -305 806
rect -271 430 -255 806
rect -321 418 -255 430
rect -225 806 -159 818
rect -225 430 -209 806
rect -175 430 -159 806
rect -225 418 -159 430
rect -129 806 -63 818
rect -129 430 -113 806
rect -79 430 -63 806
rect -129 418 -63 430
rect -33 806 33 818
rect -33 430 -17 806
rect 17 430 33 806
rect -33 418 33 430
rect 63 806 129 818
rect 63 430 79 806
rect 113 430 129 806
rect 63 418 129 430
rect 159 806 225 818
rect 159 430 175 806
rect 209 430 225 806
rect 159 418 225 430
rect 255 806 321 818
rect 255 430 271 806
rect 305 430 321 806
rect 255 418 321 430
rect 351 806 417 818
rect 351 430 367 806
rect 401 430 417 806
rect 351 418 417 430
rect 447 806 513 818
rect 447 430 463 806
rect 497 430 513 806
rect 447 418 513 430
rect 543 806 609 818
rect 543 430 559 806
rect 593 430 609 806
rect 543 418 609 430
rect 639 806 705 818
rect 639 430 655 806
rect 689 430 705 806
rect 639 418 705 430
rect 735 806 801 818
rect 735 430 751 806
rect 785 430 801 806
rect 735 418 801 430
rect 831 806 897 818
rect 831 430 847 806
rect 881 430 897 806
rect 831 418 897 430
rect 927 806 989 818
rect 927 430 943 806
rect 977 430 989 806
rect 927 418 989 430
rect -989 188 -927 200
rect -989 -188 -977 188
rect -943 -188 -927 188
rect -989 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 989 200
rect 927 -188 943 188
rect 977 -188 989 188
rect 927 -200 989 -188
rect -989 -430 -927 -418
rect -989 -806 -977 -430
rect -943 -806 -927 -430
rect -989 -818 -927 -806
rect -897 -430 -831 -418
rect -897 -806 -881 -430
rect -847 -806 -831 -430
rect -897 -818 -831 -806
rect -801 -430 -735 -418
rect -801 -806 -785 -430
rect -751 -806 -735 -430
rect -801 -818 -735 -806
rect -705 -430 -639 -418
rect -705 -806 -689 -430
rect -655 -806 -639 -430
rect -705 -818 -639 -806
rect -609 -430 -543 -418
rect -609 -806 -593 -430
rect -559 -806 -543 -430
rect -609 -818 -543 -806
rect -513 -430 -447 -418
rect -513 -806 -497 -430
rect -463 -806 -447 -430
rect -513 -818 -447 -806
rect -417 -430 -351 -418
rect -417 -806 -401 -430
rect -367 -806 -351 -430
rect -417 -818 -351 -806
rect -321 -430 -255 -418
rect -321 -806 -305 -430
rect -271 -806 -255 -430
rect -321 -818 -255 -806
rect -225 -430 -159 -418
rect -225 -806 -209 -430
rect -175 -806 -159 -430
rect -225 -818 -159 -806
rect -129 -430 -63 -418
rect -129 -806 -113 -430
rect -79 -806 -63 -430
rect -129 -818 -63 -806
rect -33 -430 33 -418
rect -33 -806 -17 -430
rect 17 -806 33 -430
rect -33 -818 33 -806
rect 63 -430 129 -418
rect 63 -806 79 -430
rect 113 -806 129 -430
rect 63 -818 129 -806
rect 159 -430 225 -418
rect 159 -806 175 -430
rect 209 -806 225 -430
rect 159 -818 225 -806
rect 255 -430 321 -418
rect 255 -806 271 -430
rect 305 -806 321 -430
rect 255 -818 321 -806
rect 351 -430 417 -418
rect 351 -806 367 -430
rect 401 -806 417 -430
rect 351 -818 417 -806
rect 447 -430 513 -418
rect 447 -806 463 -430
rect 497 -806 513 -430
rect 447 -818 513 -806
rect 543 -430 609 -418
rect 543 -806 559 -430
rect 593 -806 609 -430
rect 543 -818 609 -806
rect 639 -430 705 -418
rect 639 -806 655 -430
rect 689 -806 705 -430
rect 639 -818 705 -806
rect 735 -430 801 -418
rect 735 -806 751 -430
rect 785 -806 801 -430
rect 735 -818 801 -806
rect 831 -430 897 -418
rect 831 -806 847 -430
rect 881 -806 897 -430
rect 831 -818 897 -806
rect 927 -430 989 -418
rect 927 -806 943 -430
rect 977 -806 989 -430
rect 927 -818 989 -806
<< ndiffc >>
rect -977 430 -943 806
rect -881 430 -847 806
rect -785 430 -751 806
rect -689 430 -655 806
rect -593 430 -559 806
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect 559 430 593 806
rect 655 430 689 806
rect 751 430 785 806
rect 847 430 881 806
rect 943 430 977 806
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect -977 -806 -943 -430
rect -881 -806 -847 -430
rect -785 -806 -751 -430
rect -689 -806 -655 -430
rect -593 -806 -559 -430
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect 559 -806 593 -430
rect 655 -806 689 -430
rect 751 -806 785 -430
rect 847 -806 881 -430
rect 943 -806 977 -430
<< psubdiff >>
rect -1091 958 -995 992
rect 995 958 1091 992
rect -1091 896 -1057 958
rect 1057 896 1091 958
rect -1091 -958 -1057 -896
rect 1057 -958 1091 -896
rect -1091 -992 -995 -958
rect 995 -992 1091 -958
<< psubdiffcont >>
rect -995 958 995 992
rect -1091 -896 -1057 896
rect 1057 -896 1091 896
rect -995 -992 995 -958
<< poly >>
rect -849 890 -783 906
rect -849 856 -833 890
rect -799 856 -783 890
rect -927 818 -897 844
rect -849 840 -783 856
rect -657 890 -591 906
rect -657 856 -641 890
rect -607 856 -591 890
rect -831 818 -801 840
rect -735 818 -705 844
rect -657 840 -591 856
rect -465 890 -399 906
rect -465 856 -449 890
rect -415 856 -399 890
rect -639 818 -609 840
rect -543 818 -513 844
rect -465 840 -399 856
rect -273 890 -207 906
rect -273 856 -257 890
rect -223 856 -207 890
rect -447 818 -417 840
rect -351 818 -321 844
rect -273 840 -207 856
rect -81 890 -15 906
rect -81 856 -65 890
rect -31 856 -15 890
rect -255 818 -225 840
rect -159 818 -129 844
rect -81 840 -15 856
rect 111 890 177 906
rect 111 856 127 890
rect 161 856 177 890
rect -63 818 -33 840
rect 33 818 63 844
rect 111 840 177 856
rect 303 890 369 906
rect 303 856 319 890
rect 353 856 369 890
rect 129 818 159 840
rect 225 818 255 844
rect 303 840 369 856
rect 495 890 561 906
rect 495 856 511 890
rect 545 856 561 890
rect 321 818 351 840
rect 417 818 447 844
rect 495 840 561 856
rect 687 890 753 906
rect 687 856 703 890
rect 737 856 753 890
rect 513 818 543 840
rect 609 818 639 844
rect 687 840 753 856
rect 879 890 945 906
rect 879 856 895 890
rect 929 856 945 890
rect 705 818 735 840
rect 801 818 831 844
rect 879 840 945 856
rect 897 818 927 840
rect -927 396 -897 418
rect -945 380 -879 396
rect -831 392 -801 418
rect -735 396 -705 418
rect -945 346 -929 380
rect -895 346 -879 380
rect -945 330 -879 346
rect -753 380 -687 396
rect -639 392 -609 418
rect -543 396 -513 418
rect -753 346 -737 380
rect -703 346 -687 380
rect -753 330 -687 346
rect -561 380 -495 396
rect -447 392 -417 418
rect -351 396 -321 418
rect -561 346 -545 380
rect -511 346 -495 380
rect -561 330 -495 346
rect -369 380 -303 396
rect -255 392 -225 418
rect -159 396 -129 418
rect -369 346 -353 380
rect -319 346 -303 380
rect -369 330 -303 346
rect -177 380 -111 396
rect -63 392 -33 418
rect 33 396 63 418
rect -177 346 -161 380
rect -127 346 -111 380
rect -177 330 -111 346
rect 15 380 81 396
rect 129 392 159 418
rect 225 396 255 418
rect 15 346 31 380
rect 65 346 81 380
rect 15 330 81 346
rect 207 380 273 396
rect 321 392 351 418
rect 417 396 447 418
rect 207 346 223 380
rect 257 346 273 380
rect 207 330 273 346
rect 399 380 465 396
rect 513 392 543 418
rect 609 396 639 418
rect 399 346 415 380
rect 449 346 465 380
rect 399 330 465 346
rect 591 380 657 396
rect 705 392 735 418
rect 801 396 831 418
rect 591 346 607 380
rect 641 346 657 380
rect 591 330 657 346
rect 783 380 849 396
rect 897 392 927 418
rect 783 346 799 380
rect 833 346 849 380
rect 783 330 849 346
rect -945 272 -879 288
rect -945 238 -929 272
rect -895 238 -879 272
rect -945 222 -879 238
rect -753 272 -687 288
rect -753 238 -737 272
rect -703 238 -687 272
rect -927 200 -897 222
rect -831 200 -801 226
rect -753 222 -687 238
rect -561 272 -495 288
rect -561 238 -545 272
rect -511 238 -495 272
rect -735 200 -705 222
rect -639 200 -609 226
rect -561 222 -495 238
rect -369 272 -303 288
rect -369 238 -353 272
rect -319 238 -303 272
rect -543 200 -513 222
rect -447 200 -417 226
rect -369 222 -303 238
rect -177 272 -111 288
rect -177 238 -161 272
rect -127 238 -111 272
rect -351 200 -321 222
rect -255 200 -225 226
rect -177 222 -111 238
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -159 200 -129 222
rect -63 200 -33 226
rect 15 222 81 238
rect 207 272 273 288
rect 207 238 223 272
rect 257 238 273 272
rect 33 200 63 222
rect 129 200 159 226
rect 207 222 273 238
rect 399 272 465 288
rect 399 238 415 272
rect 449 238 465 272
rect 225 200 255 222
rect 321 200 351 226
rect 399 222 465 238
rect 591 272 657 288
rect 591 238 607 272
rect 641 238 657 272
rect 417 200 447 222
rect 513 200 543 226
rect 591 222 657 238
rect 783 272 849 288
rect 783 238 799 272
rect 833 238 849 272
rect 609 200 639 222
rect 705 200 735 226
rect 783 222 849 238
rect 801 200 831 222
rect 897 200 927 226
rect -927 -226 -897 -200
rect -831 -222 -801 -200
rect -849 -238 -783 -222
rect -735 -226 -705 -200
rect -639 -222 -609 -200
rect -849 -272 -833 -238
rect -799 -272 -783 -238
rect -849 -288 -783 -272
rect -657 -238 -591 -222
rect -543 -226 -513 -200
rect -447 -222 -417 -200
rect -657 -272 -641 -238
rect -607 -272 -591 -238
rect -657 -288 -591 -272
rect -465 -238 -399 -222
rect -351 -226 -321 -200
rect -255 -222 -225 -200
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -465 -288 -399 -272
rect -273 -238 -207 -222
rect -159 -226 -129 -200
rect -63 -222 -33 -200
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -273 -288 -207 -272
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect 129 -222 159 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
rect 111 -238 177 -222
rect 225 -226 255 -200
rect 321 -222 351 -200
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 111 -288 177 -272
rect 303 -238 369 -222
rect 417 -226 447 -200
rect 513 -222 543 -200
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 303 -288 369 -272
rect 495 -238 561 -222
rect 609 -226 639 -200
rect 705 -222 735 -200
rect 495 -272 511 -238
rect 545 -272 561 -238
rect 495 -288 561 -272
rect 687 -238 753 -222
rect 801 -226 831 -200
rect 897 -222 927 -200
rect 687 -272 703 -238
rect 737 -272 753 -238
rect 687 -288 753 -272
rect 879 -238 945 -222
rect 879 -272 895 -238
rect 929 -272 945 -238
rect 879 -288 945 -272
rect -849 -346 -783 -330
rect -849 -380 -833 -346
rect -799 -380 -783 -346
rect -927 -418 -897 -392
rect -849 -396 -783 -380
rect -657 -346 -591 -330
rect -657 -380 -641 -346
rect -607 -380 -591 -346
rect -831 -418 -801 -396
rect -735 -418 -705 -392
rect -657 -396 -591 -380
rect -465 -346 -399 -330
rect -465 -380 -449 -346
rect -415 -380 -399 -346
rect -639 -418 -609 -396
rect -543 -418 -513 -392
rect -465 -396 -399 -380
rect -273 -346 -207 -330
rect -273 -380 -257 -346
rect -223 -380 -207 -346
rect -447 -418 -417 -396
rect -351 -418 -321 -392
rect -273 -396 -207 -380
rect -81 -346 -15 -330
rect -81 -380 -65 -346
rect -31 -380 -15 -346
rect -255 -418 -225 -396
rect -159 -418 -129 -392
rect -81 -396 -15 -380
rect 111 -346 177 -330
rect 111 -380 127 -346
rect 161 -380 177 -346
rect -63 -418 -33 -396
rect 33 -418 63 -392
rect 111 -396 177 -380
rect 303 -346 369 -330
rect 303 -380 319 -346
rect 353 -380 369 -346
rect 129 -418 159 -396
rect 225 -418 255 -392
rect 303 -396 369 -380
rect 495 -346 561 -330
rect 495 -380 511 -346
rect 545 -380 561 -346
rect 321 -418 351 -396
rect 417 -418 447 -392
rect 495 -396 561 -380
rect 687 -346 753 -330
rect 687 -380 703 -346
rect 737 -380 753 -346
rect 513 -418 543 -396
rect 609 -418 639 -392
rect 687 -396 753 -380
rect 879 -346 945 -330
rect 879 -380 895 -346
rect 929 -380 945 -346
rect 705 -418 735 -396
rect 801 -418 831 -392
rect 879 -396 945 -380
rect 897 -418 927 -396
rect -927 -840 -897 -818
rect -945 -856 -879 -840
rect -831 -844 -801 -818
rect -735 -840 -705 -818
rect -945 -890 -929 -856
rect -895 -890 -879 -856
rect -945 -906 -879 -890
rect -753 -856 -687 -840
rect -639 -844 -609 -818
rect -543 -840 -513 -818
rect -753 -890 -737 -856
rect -703 -890 -687 -856
rect -753 -906 -687 -890
rect -561 -856 -495 -840
rect -447 -844 -417 -818
rect -351 -840 -321 -818
rect -561 -890 -545 -856
rect -511 -890 -495 -856
rect -561 -906 -495 -890
rect -369 -856 -303 -840
rect -255 -844 -225 -818
rect -159 -840 -129 -818
rect -369 -890 -353 -856
rect -319 -890 -303 -856
rect -369 -906 -303 -890
rect -177 -856 -111 -840
rect -63 -844 -33 -818
rect 33 -840 63 -818
rect -177 -890 -161 -856
rect -127 -890 -111 -856
rect -177 -906 -111 -890
rect 15 -856 81 -840
rect 129 -844 159 -818
rect 225 -840 255 -818
rect 15 -890 31 -856
rect 65 -890 81 -856
rect 15 -906 81 -890
rect 207 -856 273 -840
rect 321 -844 351 -818
rect 417 -840 447 -818
rect 207 -890 223 -856
rect 257 -890 273 -856
rect 207 -906 273 -890
rect 399 -856 465 -840
rect 513 -844 543 -818
rect 609 -840 639 -818
rect 399 -890 415 -856
rect 449 -890 465 -856
rect 399 -906 465 -890
rect 591 -856 657 -840
rect 705 -844 735 -818
rect 801 -840 831 -818
rect 591 -890 607 -856
rect 641 -890 657 -856
rect 591 -906 657 -890
rect 783 -856 849 -840
rect 897 -844 927 -818
rect 783 -890 799 -856
rect 833 -890 849 -856
rect 783 -906 849 -890
<< polycont >>
rect -833 856 -799 890
rect -641 856 -607 890
rect -449 856 -415 890
rect -257 856 -223 890
rect -65 856 -31 890
rect 127 856 161 890
rect 319 856 353 890
rect 511 856 545 890
rect 703 856 737 890
rect 895 856 929 890
rect -929 346 -895 380
rect -737 346 -703 380
rect -545 346 -511 380
rect -353 346 -319 380
rect -161 346 -127 380
rect 31 346 65 380
rect 223 346 257 380
rect 415 346 449 380
rect 607 346 641 380
rect 799 346 833 380
rect -929 238 -895 272
rect -737 238 -703 272
rect -545 238 -511 272
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect 607 238 641 272
rect 799 238 833 272
rect -833 -272 -799 -238
rect -641 -272 -607 -238
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect 511 -272 545 -238
rect 703 -272 737 -238
rect 895 -272 929 -238
rect -833 -380 -799 -346
rect -641 -380 -607 -346
rect -449 -380 -415 -346
rect -257 -380 -223 -346
rect -65 -380 -31 -346
rect 127 -380 161 -346
rect 319 -380 353 -346
rect 511 -380 545 -346
rect 703 -380 737 -346
rect 895 -380 929 -346
rect -929 -890 -895 -856
rect -737 -890 -703 -856
rect -545 -890 -511 -856
rect -353 -890 -319 -856
rect -161 -890 -127 -856
rect 31 -890 65 -856
rect 223 -890 257 -856
rect 415 -890 449 -856
rect 607 -890 641 -856
rect 799 -890 833 -856
<< locali >>
rect -1091 958 -995 992
rect 995 958 1091 992
rect -1091 896 -1057 958
rect 1057 896 1091 958
rect -849 856 -833 890
rect -799 856 -783 890
rect -657 856 -641 890
rect -607 856 -591 890
rect -465 856 -449 890
rect -415 856 -399 890
rect -273 856 -257 890
rect -223 856 -207 890
rect -81 856 -65 890
rect -31 856 -15 890
rect 111 856 127 890
rect 161 856 177 890
rect 303 856 319 890
rect 353 856 369 890
rect 495 856 511 890
rect 545 856 561 890
rect 687 856 703 890
rect 737 856 753 890
rect 879 856 895 890
rect 929 856 945 890
rect -977 806 -943 822
rect -977 414 -943 430
rect -881 806 -847 822
rect -881 414 -847 430
rect -785 806 -751 822
rect -785 414 -751 430
rect -689 806 -655 822
rect -689 414 -655 430
rect -593 806 -559 822
rect -593 414 -559 430
rect -497 806 -463 822
rect -497 414 -463 430
rect -401 806 -367 822
rect -401 414 -367 430
rect -305 806 -271 822
rect -305 414 -271 430
rect -209 806 -175 822
rect -209 414 -175 430
rect -113 806 -79 822
rect -113 414 -79 430
rect -17 806 17 822
rect -17 414 17 430
rect 79 806 113 822
rect 79 414 113 430
rect 175 806 209 822
rect 175 414 209 430
rect 271 806 305 822
rect 271 414 305 430
rect 367 806 401 822
rect 367 414 401 430
rect 463 806 497 822
rect 463 414 497 430
rect 559 806 593 822
rect 559 414 593 430
rect 655 806 689 822
rect 655 414 689 430
rect 751 806 785 822
rect 751 414 785 430
rect 847 806 881 822
rect 847 414 881 430
rect 943 806 977 822
rect 943 414 977 430
rect -945 346 -929 380
rect -895 346 -879 380
rect -753 346 -737 380
rect -703 346 -687 380
rect -561 346 -545 380
rect -511 346 -495 380
rect -369 346 -353 380
rect -319 346 -303 380
rect -177 346 -161 380
rect -127 346 -111 380
rect 15 346 31 380
rect 65 346 81 380
rect 207 346 223 380
rect 257 346 273 380
rect 399 346 415 380
rect 449 346 465 380
rect 591 346 607 380
rect 641 346 657 380
rect 783 346 799 380
rect 833 346 849 380
rect -945 238 -929 272
rect -895 238 -879 272
rect -753 238 -737 272
rect -703 238 -687 272
rect -561 238 -545 272
rect -511 238 -495 272
rect -369 238 -353 272
rect -319 238 -303 272
rect -177 238 -161 272
rect -127 238 -111 272
rect 15 238 31 272
rect 65 238 81 272
rect 207 238 223 272
rect 257 238 273 272
rect 399 238 415 272
rect 449 238 465 272
rect 591 238 607 272
rect 641 238 657 272
rect 783 238 799 272
rect 833 238 849 272
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect -849 -272 -833 -238
rect -799 -272 -783 -238
rect -657 -272 -641 -238
rect -607 -272 -591 -238
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 495 -272 511 -238
rect 545 -272 561 -238
rect 687 -272 703 -238
rect 737 -272 753 -238
rect 879 -272 895 -238
rect 929 -272 945 -238
rect -849 -380 -833 -346
rect -799 -380 -783 -346
rect -657 -380 -641 -346
rect -607 -380 -591 -346
rect -465 -380 -449 -346
rect -415 -380 -399 -346
rect -273 -380 -257 -346
rect -223 -380 -207 -346
rect -81 -380 -65 -346
rect -31 -380 -15 -346
rect 111 -380 127 -346
rect 161 -380 177 -346
rect 303 -380 319 -346
rect 353 -380 369 -346
rect 495 -380 511 -346
rect 545 -380 561 -346
rect 687 -380 703 -346
rect 737 -380 753 -346
rect 879 -380 895 -346
rect 929 -380 945 -346
rect -977 -430 -943 -414
rect -977 -822 -943 -806
rect -881 -430 -847 -414
rect -881 -822 -847 -806
rect -785 -430 -751 -414
rect -785 -822 -751 -806
rect -689 -430 -655 -414
rect -689 -822 -655 -806
rect -593 -430 -559 -414
rect -593 -822 -559 -806
rect -497 -430 -463 -414
rect -497 -822 -463 -806
rect -401 -430 -367 -414
rect -401 -822 -367 -806
rect -305 -430 -271 -414
rect -305 -822 -271 -806
rect -209 -430 -175 -414
rect -209 -822 -175 -806
rect -113 -430 -79 -414
rect -113 -822 -79 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 79 -430 113 -414
rect 79 -822 113 -806
rect 175 -430 209 -414
rect 175 -822 209 -806
rect 271 -430 305 -414
rect 271 -822 305 -806
rect 367 -430 401 -414
rect 367 -822 401 -806
rect 463 -430 497 -414
rect 463 -822 497 -806
rect 559 -430 593 -414
rect 559 -822 593 -806
rect 655 -430 689 -414
rect 655 -822 689 -806
rect 751 -430 785 -414
rect 751 -822 785 -806
rect 847 -430 881 -414
rect 847 -822 881 -806
rect 943 -430 977 -414
rect 943 -822 977 -806
rect -945 -890 -929 -856
rect -895 -890 -879 -856
rect -753 -890 -737 -856
rect -703 -890 -687 -856
rect -561 -890 -545 -856
rect -511 -890 -495 -856
rect -369 -890 -353 -856
rect -319 -890 -303 -856
rect -177 -890 -161 -856
rect -127 -890 -111 -856
rect 15 -890 31 -856
rect 65 -890 81 -856
rect 207 -890 223 -856
rect 257 -890 273 -856
rect 399 -890 415 -856
rect 449 -890 465 -856
rect 591 -890 607 -856
rect 641 -890 657 -856
rect 783 -890 799 -856
rect 833 -890 849 -856
rect -1091 -958 -1057 -896
rect 1057 -958 1091 -896
rect -1091 -992 -995 -958
rect 995 -992 1091 -958
<< viali >>
rect -833 856 -799 890
rect -641 856 -607 890
rect -449 856 -415 890
rect -257 856 -223 890
rect -65 856 -31 890
rect 127 856 161 890
rect 319 856 353 890
rect 511 856 545 890
rect 703 856 737 890
rect 895 856 929 890
rect -977 430 -943 806
rect -881 430 -847 806
rect -785 430 -751 806
rect -689 430 -655 806
rect -593 430 -559 806
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect 559 430 593 806
rect 655 430 689 806
rect 751 430 785 806
rect 847 430 881 806
rect 943 430 977 806
rect -929 346 -895 380
rect -737 346 -703 380
rect -545 346 -511 380
rect -353 346 -319 380
rect -161 346 -127 380
rect 31 346 65 380
rect 223 346 257 380
rect 415 346 449 380
rect 607 346 641 380
rect 799 346 833 380
rect -929 238 -895 272
rect -737 238 -703 272
rect -545 238 -511 272
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect 607 238 641 272
rect 799 238 833 272
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect -833 -272 -799 -238
rect -641 -272 -607 -238
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect 511 -272 545 -238
rect 703 -272 737 -238
rect 895 -272 929 -238
rect -833 -380 -799 -346
rect -641 -380 -607 -346
rect -449 -380 -415 -346
rect -257 -380 -223 -346
rect -65 -380 -31 -346
rect 127 -380 161 -346
rect 319 -380 353 -346
rect 511 -380 545 -346
rect 703 -380 737 -346
rect 895 -380 929 -346
rect -977 -806 -943 -430
rect -881 -806 -847 -430
rect -785 -806 -751 -430
rect -689 -806 -655 -430
rect -593 -806 -559 -430
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect 559 -806 593 -430
rect 655 -806 689 -430
rect 751 -806 785 -430
rect 847 -806 881 -430
rect 943 -806 977 -430
rect -929 -890 -895 -856
rect -737 -890 -703 -856
rect -545 -890 -511 -856
rect -353 -890 -319 -856
rect -161 -890 -127 -856
rect 31 -890 65 -856
rect 223 -890 257 -856
rect 415 -890 449 -856
rect 607 -890 641 -856
rect 799 -890 833 -856
<< metal1 >>
rect -845 890 -787 896
rect -845 856 -833 890
rect -799 856 -787 890
rect -845 850 -787 856
rect -653 890 -595 896
rect -653 856 -641 890
rect -607 856 -595 890
rect -653 850 -595 856
rect -461 890 -403 896
rect -461 856 -449 890
rect -415 856 -403 890
rect -461 850 -403 856
rect -269 890 -211 896
rect -269 856 -257 890
rect -223 856 -211 890
rect -269 850 -211 856
rect -77 890 -19 896
rect -77 856 -65 890
rect -31 856 -19 890
rect -77 850 -19 856
rect 115 890 173 896
rect 115 856 127 890
rect 161 856 173 890
rect 115 850 173 856
rect 307 890 365 896
rect 307 856 319 890
rect 353 856 365 890
rect 307 850 365 856
rect 499 890 557 896
rect 499 856 511 890
rect 545 856 557 890
rect 499 850 557 856
rect 691 890 749 896
rect 691 856 703 890
rect 737 856 749 890
rect 691 850 749 856
rect 883 890 941 896
rect 883 856 895 890
rect 929 856 941 890
rect 883 850 941 856
rect -983 806 -937 818
rect -983 430 -977 806
rect -943 430 -937 806
rect -983 418 -937 430
rect -887 806 -841 818
rect -887 430 -881 806
rect -847 430 -841 806
rect -887 418 -841 430
rect -791 806 -745 818
rect -791 430 -785 806
rect -751 430 -745 806
rect -791 418 -745 430
rect -695 806 -649 818
rect -695 430 -689 806
rect -655 430 -649 806
rect -695 418 -649 430
rect -599 806 -553 818
rect -599 430 -593 806
rect -559 430 -553 806
rect -599 418 -553 430
rect -503 806 -457 818
rect -503 430 -497 806
rect -463 430 -457 806
rect -503 418 -457 430
rect -407 806 -361 818
rect -407 430 -401 806
rect -367 430 -361 806
rect -407 418 -361 430
rect -311 806 -265 818
rect -311 430 -305 806
rect -271 430 -265 806
rect -311 418 -265 430
rect -215 806 -169 818
rect -215 430 -209 806
rect -175 430 -169 806
rect -215 418 -169 430
rect -119 806 -73 818
rect -119 430 -113 806
rect -79 430 -73 806
rect -119 418 -73 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 73 806 119 818
rect 73 430 79 806
rect 113 430 119 806
rect 73 418 119 430
rect 169 806 215 818
rect 169 430 175 806
rect 209 430 215 806
rect 169 418 215 430
rect 265 806 311 818
rect 265 430 271 806
rect 305 430 311 806
rect 265 418 311 430
rect 361 806 407 818
rect 361 430 367 806
rect 401 430 407 806
rect 361 418 407 430
rect 457 806 503 818
rect 457 430 463 806
rect 497 430 503 806
rect 457 418 503 430
rect 553 806 599 818
rect 553 430 559 806
rect 593 430 599 806
rect 553 418 599 430
rect 649 806 695 818
rect 649 430 655 806
rect 689 430 695 806
rect 649 418 695 430
rect 745 806 791 818
rect 745 430 751 806
rect 785 430 791 806
rect 745 418 791 430
rect 841 806 887 818
rect 841 430 847 806
rect 881 430 887 806
rect 841 418 887 430
rect 937 806 983 818
rect 937 430 943 806
rect 977 430 983 806
rect 937 418 983 430
rect -941 380 -883 386
rect -941 346 -929 380
rect -895 346 -883 380
rect -941 340 -883 346
rect -749 380 -691 386
rect -749 346 -737 380
rect -703 346 -691 380
rect -749 340 -691 346
rect -557 380 -499 386
rect -557 346 -545 380
rect -511 346 -499 380
rect -557 340 -499 346
rect -365 380 -307 386
rect -365 346 -353 380
rect -319 346 -307 380
rect -365 340 -307 346
rect -173 380 -115 386
rect -173 346 -161 380
rect -127 346 -115 380
rect -173 340 -115 346
rect 19 380 77 386
rect 19 346 31 380
rect 65 346 77 380
rect 19 340 77 346
rect 211 380 269 386
rect 211 346 223 380
rect 257 346 269 380
rect 211 340 269 346
rect 403 380 461 386
rect 403 346 415 380
rect 449 346 461 380
rect 403 340 461 346
rect 595 380 653 386
rect 595 346 607 380
rect 641 346 653 380
rect 595 340 653 346
rect 787 380 845 386
rect 787 346 799 380
rect 833 346 845 380
rect 787 340 845 346
rect -941 272 -883 278
rect -941 238 -929 272
rect -895 238 -883 272
rect -941 232 -883 238
rect -749 272 -691 278
rect -749 238 -737 272
rect -703 238 -691 272
rect -749 232 -691 238
rect -557 272 -499 278
rect -557 238 -545 272
rect -511 238 -499 272
rect -557 232 -499 238
rect -365 272 -307 278
rect -365 238 -353 272
rect -319 238 -307 272
rect -365 232 -307 238
rect -173 272 -115 278
rect -173 238 -161 272
rect -127 238 -115 272
rect -173 232 -115 238
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect 211 272 269 278
rect 211 238 223 272
rect 257 238 269 272
rect 211 232 269 238
rect 403 272 461 278
rect 403 238 415 272
rect 449 238 461 272
rect 403 232 461 238
rect 595 272 653 278
rect 595 238 607 272
rect 641 238 653 272
rect 595 232 653 238
rect 787 272 845 278
rect 787 238 799 272
rect 833 238 845 272
rect 787 232 845 238
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect -845 -238 -787 -232
rect -845 -272 -833 -238
rect -799 -272 -787 -238
rect -845 -278 -787 -272
rect -653 -238 -595 -232
rect -653 -272 -641 -238
rect -607 -272 -595 -238
rect -653 -278 -595 -272
rect -461 -238 -403 -232
rect -461 -272 -449 -238
rect -415 -272 -403 -238
rect -461 -278 -403 -272
rect -269 -238 -211 -232
rect -269 -272 -257 -238
rect -223 -272 -211 -238
rect -269 -278 -211 -272
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
rect 115 -238 173 -232
rect 115 -272 127 -238
rect 161 -272 173 -238
rect 115 -278 173 -272
rect 307 -238 365 -232
rect 307 -272 319 -238
rect 353 -272 365 -238
rect 307 -278 365 -272
rect 499 -238 557 -232
rect 499 -272 511 -238
rect 545 -272 557 -238
rect 499 -278 557 -272
rect 691 -238 749 -232
rect 691 -272 703 -238
rect 737 -272 749 -238
rect 691 -278 749 -272
rect 883 -238 941 -232
rect 883 -272 895 -238
rect 929 -272 941 -238
rect 883 -278 941 -272
rect -845 -346 -787 -340
rect -845 -380 -833 -346
rect -799 -380 -787 -346
rect -845 -386 -787 -380
rect -653 -346 -595 -340
rect -653 -380 -641 -346
rect -607 -380 -595 -346
rect -653 -386 -595 -380
rect -461 -346 -403 -340
rect -461 -380 -449 -346
rect -415 -380 -403 -346
rect -461 -386 -403 -380
rect -269 -346 -211 -340
rect -269 -380 -257 -346
rect -223 -380 -211 -346
rect -269 -386 -211 -380
rect -77 -346 -19 -340
rect -77 -380 -65 -346
rect -31 -380 -19 -346
rect -77 -386 -19 -380
rect 115 -346 173 -340
rect 115 -380 127 -346
rect 161 -380 173 -346
rect 115 -386 173 -380
rect 307 -346 365 -340
rect 307 -380 319 -346
rect 353 -380 365 -346
rect 307 -386 365 -380
rect 499 -346 557 -340
rect 499 -380 511 -346
rect 545 -380 557 -346
rect 499 -386 557 -380
rect 691 -346 749 -340
rect 691 -380 703 -346
rect 737 -380 749 -346
rect 691 -386 749 -380
rect 883 -346 941 -340
rect 883 -380 895 -346
rect 929 -380 941 -346
rect 883 -386 941 -380
rect -983 -430 -937 -418
rect -983 -806 -977 -430
rect -943 -806 -937 -430
rect -983 -818 -937 -806
rect -887 -430 -841 -418
rect -887 -806 -881 -430
rect -847 -806 -841 -430
rect -887 -818 -841 -806
rect -791 -430 -745 -418
rect -791 -806 -785 -430
rect -751 -806 -745 -430
rect -791 -818 -745 -806
rect -695 -430 -649 -418
rect -695 -806 -689 -430
rect -655 -806 -649 -430
rect -695 -818 -649 -806
rect -599 -430 -553 -418
rect -599 -806 -593 -430
rect -559 -806 -553 -430
rect -599 -818 -553 -806
rect -503 -430 -457 -418
rect -503 -806 -497 -430
rect -463 -806 -457 -430
rect -503 -818 -457 -806
rect -407 -430 -361 -418
rect -407 -806 -401 -430
rect -367 -806 -361 -430
rect -407 -818 -361 -806
rect -311 -430 -265 -418
rect -311 -806 -305 -430
rect -271 -806 -265 -430
rect -311 -818 -265 -806
rect -215 -430 -169 -418
rect -215 -806 -209 -430
rect -175 -806 -169 -430
rect -215 -818 -169 -806
rect -119 -430 -73 -418
rect -119 -806 -113 -430
rect -79 -806 -73 -430
rect -119 -818 -73 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 73 -430 119 -418
rect 73 -806 79 -430
rect 113 -806 119 -430
rect 73 -818 119 -806
rect 169 -430 215 -418
rect 169 -806 175 -430
rect 209 -806 215 -430
rect 169 -818 215 -806
rect 265 -430 311 -418
rect 265 -806 271 -430
rect 305 -806 311 -430
rect 265 -818 311 -806
rect 361 -430 407 -418
rect 361 -806 367 -430
rect 401 -806 407 -430
rect 361 -818 407 -806
rect 457 -430 503 -418
rect 457 -806 463 -430
rect 497 -806 503 -430
rect 457 -818 503 -806
rect 553 -430 599 -418
rect 553 -806 559 -430
rect 593 -806 599 -430
rect 553 -818 599 -806
rect 649 -430 695 -418
rect 649 -806 655 -430
rect 689 -806 695 -430
rect 649 -818 695 -806
rect 745 -430 791 -418
rect 745 -806 751 -430
rect 785 -806 791 -430
rect 745 -818 791 -806
rect 841 -430 887 -418
rect 841 -806 847 -430
rect 881 -806 887 -430
rect 841 -818 887 -806
rect 937 -430 983 -418
rect 937 -806 943 -430
rect 977 -806 983 -430
rect 937 -818 983 -806
rect -941 -856 -883 -850
rect -941 -890 -929 -856
rect -895 -890 -883 -856
rect -941 -896 -883 -890
rect -749 -856 -691 -850
rect -749 -890 -737 -856
rect -703 -890 -691 -856
rect -749 -896 -691 -890
rect -557 -856 -499 -850
rect -557 -890 -545 -856
rect -511 -890 -499 -856
rect -557 -896 -499 -890
rect -365 -856 -307 -850
rect -365 -890 -353 -856
rect -319 -890 -307 -856
rect -365 -896 -307 -890
rect -173 -856 -115 -850
rect -173 -890 -161 -856
rect -127 -890 -115 -856
rect -173 -896 -115 -890
rect 19 -856 77 -850
rect 19 -890 31 -856
rect 65 -890 77 -856
rect 19 -896 77 -890
rect 211 -856 269 -850
rect 211 -890 223 -856
rect 257 -890 269 -856
rect 211 -896 269 -890
rect 403 -856 461 -850
rect 403 -890 415 -856
rect 449 -890 461 -856
rect 403 -896 461 -890
rect 595 -856 653 -850
rect 595 -890 607 -856
rect 641 -890 653 -856
rect 595 -896 653 -890
rect 787 -856 845 -850
rect 787 -890 799 -856
rect 833 -890 845 -856
rect 787 -896 845 -890
<< properties >>
string FIXED_BBOX -1074 -975 1074 975
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 3 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
