magic
tech sky130A
magscale 1 2
timestamp 1684500887
<< locali >>
rect 1688 376 3976 452
rect 1688 -336 1764 376
rect 3888 -336 3976 376
rect 1688 -444 3976 -336
rect 1688 -1148 1764 -444
rect 3888 -1148 3976 -444
rect 1688 -1248 3976 -1148
rect 1688 -1952 1764 -1248
rect 3888 -1952 3976 -1248
rect 1688 -2028 3976 -1952
<< metal1 >>
rect 1976 260 4224 368
rect 1926 52 1936 232
rect 1988 52 1998 232
rect 2118 52 2128 232
rect 2180 52 2190 232
rect 2310 52 2320 232
rect 2372 52 2382 232
rect 2502 52 2512 232
rect 2564 52 2574 232
rect 2694 52 2704 232
rect 2756 52 2766 232
rect 2886 52 2896 232
rect 2948 52 2958 232
rect 3078 52 3088 232
rect 3140 52 3150 232
rect 3270 52 3280 232
rect 3332 52 3342 232
rect 3462 52 3472 232
rect 3524 52 3534 232
rect 3654 52 3664 232
rect 3716 52 3726 232
rect 1830 -172 1840 8
rect 1892 -172 1902 8
rect 2022 -172 2032 8
rect 2084 -172 2094 8
rect 2214 -172 2224 8
rect 2276 -172 2286 8
rect 2406 -172 2416 8
rect 2468 -172 2478 8
rect 2598 -172 2608 8
rect 2660 -172 2670 8
rect 2790 -172 2800 8
rect 2852 -172 2862 8
rect 2982 -172 2992 8
rect 3044 -172 3054 8
rect 3174 -172 3184 8
rect 3236 -172 3246 8
rect 3366 -172 3376 8
rect 3428 -172 3438 8
rect 3558 -172 3568 8
rect 3620 -172 3630 8
rect 3750 -172 3760 8
rect 3812 -172 3822 8
rect 4088 -200 4224 260
rect 1884 -308 4224 -200
rect 4088 -456 4224 -308
rect 1980 -560 4224 -456
rect 1926 -768 1936 -588
rect 1988 -768 1998 -588
rect 2118 -768 2128 -588
rect 2180 -768 2190 -588
rect 2310 -768 2320 -588
rect 2372 -768 2382 -588
rect 2502 -768 2512 -588
rect 2564 -768 2574 -588
rect 2694 -768 2704 -588
rect 2756 -768 2766 -588
rect 2886 -768 2896 -588
rect 2948 -768 2958 -588
rect 3078 -768 3088 -588
rect 3140 -768 3150 -588
rect 3270 -768 3280 -588
rect 3332 -768 3342 -588
rect 3462 -768 3472 -588
rect 3524 -768 3534 -588
rect 3654 -768 3664 -588
rect 3716 -768 3726 -588
rect 1830 -992 1840 -812
rect 1892 -992 1902 -812
rect 2022 -992 2032 -812
rect 2084 -992 2094 -812
rect 2214 -992 2224 -812
rect 2276 -992 2286 -812
rect 2406 -992 2416 -812
rect 2468 -992 2478 -812
rect 2598 -992 2608 -812
rect 2660 -992 2670 -812
rect 2790 -992 2800 -812
rect 2852 -992 2862 -812
rect 2982 -992 2992 -812
rect 3044 -992 3054 -812
rect 3174 -992 3184 -812
rect 3236 -992 3246 -812
rect 3366 -992 3376 -812
rect 3428 -992 3438 -812
rect 3558 -992 3568 -812
rect 3620 -992 3630 -812
rect 3750 -992 3760 -812
rect 3812 -992 3822 -812
rect 4088 -1020 4224 -560
rect 1880 -1128 4224 -1020
rect 4088 -1272 4224 -1128
rect 1976 -1380 4224 -1272
rect 1926 -1588 1936 -1408
rect 1988 -1588 1998 -1408
rect 2118 -1588 2128 -1408
rect 2180 -1588 2190 -1408
rect 2310 -1588 2320 -1408
rect 2372 -1588 2382 -1408
rect 2502 -1588 2512 -1408
rect 2564 -1588 2574 -1408
rect 2694 -1588 2704 -1408
rect 2756 -1588 2766 -1408
rect 2886 -1588 2896 -1408
rect 2948 -1588 2958 -1408
rect 3078 -1588 3088 -1408
rect 3140 -1588 3150 -1408
rect 3270 -1588 3280 -1408
rect 3332 -1588 3342 -1408
rect 3462 -1588 3472 -1408
rect 3524 -1588 3534 -1408
rect 3654 -1588 3664 -1408
rect 3716 -1588 3726 -1408
rect 1830 -1812 1840 -1632
rect 1892 -1812 1902 -1632
rect 2022 -1812 2032 -1632
rect 2084 -1812 2094 -1632
rect 2214 -1812 2224 -1632
rect 2276 -1812 2286 -1632
rect 2406 -1812 2416 -1632
rect 2468 -1812 2478 -1632
rect 2598 -1812 2608 -1632
rect 2660 -1812 2670 -1632
rect 2790 -1812 2800 -1632
rect 2852 -1812 2862 -1632
rect 2982 -1812 2992 -1632
rect 3044 -1812 3054 -1632
rect 3174 -1812 3184 -1632
rect 3236 -1812 3246 -1632
rect 3366 -1812 3376 -1632
rect 3428 -1812 3438 -1632
rect 3558 -1812 3568 -1632
rect 3620 -1812 3630 -1632
rect 3750 -1812 3760 -1632
rect 3812 -1812 3822 -1632
rect 4088 -1840 4224 -1380
rect 1884 -1948 4224 -1840
<< via1 >>
rect 1936 52 1988 232
rect 2128 52 2180 232
rect 2320 52 2372 232
rect 2512 52 2564 232
rect 2704 52 2756 232
rect 2896 52 2948 232
rect 3088 52 3140 232
rect 3280 52 3332 232
rect 3472 52 3524 232
rect 3664 52 3716 232
rect 1840 -172 1892 8
rect 2032 -172 2084 8
rect 2224 -172 2276 8
rect 2416 -172 2468 8
rect 2608 -172 2660 8
rect 2800 -172 2852 8
rect 2992 -172 3044 8
rect 3184 -172 3236 8
rect 3376 -172 3428 8
rect 3568 -172 3620 8
rect 3760 -172 3812 8
rect 1936 -768 1988 -588
rect 2128 -768 2180 -588
rect 2320 -768 2372 -588
rect 2512 -768 2564 -588
rect 2704 -768 2756 -588
rect 2896 -768 2948 -588
rect 3088 -768 3140 -588
rect 3280 -768 3332 -588
rect 3472 -768 3524 -588
rect 3664 -768 3716 -588
rect 1840 -992 1892 -812
rect 2032 -992 2084 -812
rect 2224 -992 2276 -812
rect 2416 -992 2468 -812
rect 2608 -992 2660 -812
rect 2800 -992 2852 -812
rect 2992 -992 3044 -812
rect 3184 -992 3236 -812
rect 3376 -992 3428 -812
rect 3568 -992 3620 -812
rect 3760 -992 3812 -812
rect 1936 -1588 1988 -1408
rect 2128 -1588 2180 -1408
rect 2320 -1588 2372 -1408
rect 2512 -1588 2564 -1408
rect 2704 -1588 2756 -1408
rect 2896 -1588 2948 -1408
rect 3088 -1588 3140 -1408
rect 3280 -1588 3332 -1408
rect 3472 -1588 3524 -1408
rect 3664 -1588 3716 -1408
rect 1840 -1812 1892 -1632
rect 2032 -1812 2084 -1632
rect 2224 -1812 2276 -1632
rect 2416 -1812 2468 -1632
rect 2608 -1812 2660 -1632
rect 2800 -1812 2852 -1632
rect 2992 -1812 3044 -1632
rect 3184 -1812 3236 -1632
rect 3376 -1812 3428 -1632
rect 3568 -1812 3620 -1632
rect 3760 -1812 3812 -1632
<< metal2 >>
rect 1936 232 1988 242
rect 1936 42 1988 52
rect 2128 232 2180 242
rect 2128 42 2180 52
rect 2320 232 2372 242
rect 2320 42 2372 52
rect 2512 232 2564 242
rect 2512 42 2564 52
rect 2704 232 2756 242
rect 2704 42 2756 52
rect 2896 232 2948 242
rect 2896 42 2948 52
rect 3088 232 3140 242
rect 3088 42 3140 52
rect 3280 232 3332 242
rect 3280 42 3332 52
rect 3472 232 3524 242
rect 3472 42 3524 52
rect 3664 232 3716 242
rect 3664 42 3716 52
rect 1840 8 1892 18
rect 1840 -182 1892 -172
rect 2032 8 2084 18
rect 2032 -182 2084 -172
rect 2224 8 2276 18
rect 2224 -182 2276 -172
rect 2416 8 2468 18
rect 2416 -182 2468 -172
rect 2608 8 2660 18
rect 2608 -182 2660 -172
rect 2800 8 2852 18
rect 2800 -182 2852 -172
rect 2992 8 3044 18
rect 2992 -182 3044 -172
rect 3184 8 3236 18
rect 3184 -182 3236 -172
rect 3376 8 3428 18
rect 3376 -182 3428 -172
rect 3568 8 3620 18
rect 3568 -182 3620 -172
rect 3760 8 3812 18
rect 3760 -182 3812 -172
rect 1936 -588 1988 -578
rect 1936 -778 1988 -768
rect 2128 -588 2180 -578
rect 2128 -778 2180 -768
rect 2320 -588 2372 -578
rect 2320 -778 2372 -768
rect 2512 -588 2564 -578
rect 2512 -778 2564 -768
rect 2704 -588 2756 -578
rect 2704 -778 2756 -768
rect 2896 -588 2948 -578
rect 2896 -778 2948 -768
rect 3088 -588 3140 -578
rect 3088 -778 3140 -768
rect 3280 -588 3332 -578
rect 3280 -778 3332 -768
rect 3472 -588 3524 -578
rect 3472 -778 3524 -768
rect 3664 -588 3716 -578
rect 3664 -778 3716 -768
rect 1840 -812 1892 -802
rect 1840 -1002 1892 -992
rect 2032 -812 2084 -802
rect 2032 -1002 2084 -992
rect 2224 -812 2276 -802
rect 2224 -1002 2276 -992
rect 2416 -812 2468 -802
rect 2416 -1002 2468 -992
rect 2608 -812 2660 -802
rect 2608 -1002 2660 -992
rect 2800 -812 2852 -802
rect 2800 -1002 2852 -992
rect 2992 -812 3044 -802
rect 2992 -1002 3044 -992
rect 3184 -812 3236 -802
rect 3184 -1002 3236 -992
rect 3376 -812 3428 -802
rect 3376 -1002 3428 -992
rect 3568 -812 3620 -802
rect 3568 -1002 3620 -992
rect 3760 -812 3812 -802
rect 3760 -1002 3812 -992
rect 1936 -1408 1988 -1398
rect 1936 -1598 1988 -1588
rect 2128 -1408 2180 -1398
rect 2128 -1598 2180 -1588
rect 2320 -1408 2372 -1398
rect 2320 -1598 2372 -1588
rect 2512 -1408 2564 -1398
rect 2512 -1598 2564 -1588
rect 2704 -1408 2756 -1398
rect 2704 -1598 2756 -1588
rect 2896 -1408 2948 -1398
rect 2896 -1598 2948 -1588
rect 3088 -1408 3140 -1398
rect 3088 -1598 3140 -1588
rect 3280 -1408 3332 -1398
rect 3280 -1598 3332 -1588
rect 3472 -1408 3524 -1398
rect 3472 -1598 3524 -1588
rect 3664 -1408 3716 -1398
rect 3664 -1598 3716 -1588
rect 1840 -1632 1892 -1622
rect 1840 -1822 1892 -1812
rect 2032 -1632 2084 -1622
rect 2032 -1822 2084 -1812
rect 2224 -1632 2276 -1622
rect 2224 -1822 2276 -1812
rect 2416 -1632 2468 -1622
rect 2416 -1822 2468 -1812
rect 2608 -1632 2660 -1622
rect 2608 -1822 2660 -1812
rect 2800 -1632 2852 -1622
rect 2800 -1822 2852 -1812
rect 2992 -1632 3044 -1622
rect 2992 -1822 3044 -1812
rect 3184 -1632 3236 -1622
rect 3184 -1822 3236 -1812
rect 3376 -1632 3428 -1622
rect 3376 -1822 3428 -1812
rect 3568 -1632 3620 -1622
rect 3568 -1822 3620 -1812
rect 3760 -1632 3812 -1622
rect 3760 -1822 3812 -1812
use sky130_fd_pr__nfet_01v8_lvt_SDPJLJ  sky130_fd_pr__nfet_01v8_lvt_SDPJLJ_0
timestamp 1684252655
transform 1 0 2827 0 1 -790
box -1127 -410 1127 410
use sky130_fd_pr__nfet_01v8_lvt_SDPJLJ  sky130_fd_pr__nfet_01v8_lvt_SDPJLJ_1
timestamp 1684252655
transform 1 0 2827 0 1 -1610
box -1127 -410 1127 410
use sky130_fd_pr__nfet_01v8_lvt_SDPJLJ  sky130_fd_pr__nfet_01v8_lvt_SDPJLJ_2
timestamp 1684252655
transform 1 0 2827 0 1 30
box -1127 -410 1127 410
<< end >>
