magic
tech sky130A
magscale 1 2
timestamp 1685007810
<< metal4 >>
tri 1934 33739 2266 34071 se
rect 2266 34047 12734 34071
tri 12734 34047 12758 34071 sw
rect 2266 34027 2589 34047
rect 2266 33791 2269 34027
rect 2505 33811 2589 34027
rect 2825 33811 2909 34047
rect 3145 33811 3229 34047
rect 3465 33811 3549 34047
rect 3785 33811 3869 34047
rect 4105 33811 4189 34047
rect 4425 33811 4509 34047
rect 4745 33811 4829 34047
rect 5065 33811 5149 34047
rect 5385 33811 5469 34047
rect 5705 33811 5789 34047
rect 6025 33811 6109 34047
rect 6345 33811 6429 34047
rect 6665 33811 6749 34047
rect 6985 33811 7069 34047
rect 7305 33811 7389 34047
rect 7625 33811 7709 34047
rect 7945 33811 8029 34047
rect 8265 33811 8349 34047
rect 8585 33811 8669 34047
rect 8905 33811 8989 34047
rect 9225 33811 9309 34047
rect 9545 33811 9629 34047
rect 9865 33811 9949 34047
rect 10185 33811 10269 34047
rect 10505 33811 10589 34047
rect 10825 33811 10909 34047
rect 11145 33811 11229 34047
rect 11465 33811 11549 34047
rect 11785 33811 11869 34047
rect 12105 33811 12189 34047
rect 12425 34015 12758 34047
rect 12425 33811 12509 34015
rect 2505 33791 12509 33811
rect 2266 33779 12509 33791
rect 12745 33779 12758 34015
rect 2266 33739 12758 33779
tri 1726 33531 1934 33739 se
rect 1934 33723 12758 33739
rect 1934 33531 1950 33723
tri 1614 33419 1726 33531 se
rect 1726 33487 1950 33531
rect 2186 33685 12758 33723
tri 12758 33685 13120 34047 sw
rect 2186 33669 13120 33685
rect 2186 33531 12868 33669
rect 2186 33487 2378 33531
rect 1726 33419 2378 33487
tri 2378 33419 2490 33531 nw
tri 1500 33305 1614 33419 se
rect 1614 33403 2142 33419
rect 1614 33305 1630 33403
tri 1294 33099 1500 33305 se
rect 1500 33167 1630 33305
rect 1866 33183 2142 33403
tri 2142 33183 2378 33419 nw
tri 12510 33183 12858 33531 ne
rect 12858 33433 12868 33531
rect 13104 33433 13120 33669
rect 12858 33365 13120 33433
tri 13120 33365 13440 33685 sw
rect 12858 33349 13440 33365
rect 12858 33183 13188 33349
rect 1866 33180 2139 33183
tri 2139 33180 2142 33183 nw
rect 1866 33167 2126 33180
tri 2126 33167 2139 33180 nw
rect 1500 33099 1726 33167
tri 971 32776 1294 33099 se
rect 1294 33083 1726 33099
rect 1294 32847 1333 33083
rect 1569 32847 1726 33083
rect 1294 32776 1726 32847
tri 960 32765 971 32776 se
rect 971 32765 1048 32776
rect 960 32540 1048 32765
rect 1284 32767 1726 32776
tri 1726 32767 2126 33167 nw
tri 12858 33129 12912 33183 ne
rect 12912 33129 13188 33183
tri 12912 33124 12917 33129 ne
rect 12917 33124 13188 33129
tri 12917 33113 12928 33124 ne
rect 12928 33113 13188 33124
rect 13424 33113 13440 33349
tri 12928 32767 13274 33113 ne
rect 13274 33045 13440 33113
tri 13440 33045 13760 33365 sw
rect 13274 33029 13760 33045
rect 13274 32793 13508 33029
rect 13744 32793 13760 33029
rect 13274 32767 13760 32793
rect 1284 32540 1500 32767
tri 1500 32541 1726 32767 nw
tri 13274 32541 13500 32767 ne
rect 13500 32765 13760 32767
tri 13760 32765 14040 33045 sw
rect 13500 32682 14040 32765
rect 960 32456 1500 32540
rect 960 32220 984 32456
rect 1220 32220 1500 32456
rect 960 32136 1500 32220
rect 960 31900 984 32136
rect 1220 31900 1500 32136
rect 960 31816 1500 31900
rect 960 31580 984 31816
rect 1220 31580 1500 31816
rect 960 31496 1500 31580
rect 960 31260 984 31496
rect 1220 31260 1500 31496
rect 960 31176 1500 31260
rect 960 30940 984 31176
rect 1220 30940 1500 31176
rect 960 30856 1500 30940
rect 960 30620 984 30856
rect 1220 30620 1500 30856
rect 960 30536 1500 30620
rect 960 30300 984 30536
rect 1220 30300 1500 30536
rect 960 30216 1500 30300
rect 960 29980 984 30216
rect 1220 29980 1500 30216
rect 960 29896 1500 29980
rect 960 29660 984 29896
rect 1220 29660 1500 29896
rect 960 29576 1500 29660
rect 960 29340 984 29576
rect 1220 29340 1500 29576
rect 960 29256 1500 29340
rect 960 29020 984 29256
rect 1220 29020 1500 29256
rect 960 28936 1500 29020
rect 960 28700 984 28936
rect 1220 28700 1500 28936
rect 960 28616 1500 28700
rect 960 28380 984 28616
rect 1220 28380 1500 28616
rect 960 28296 1500 28380
rect 960 28060 984 28296
rect 1220 28060 1500 28296
rect 960 27976 1500 28060
rect 960 27740 984 27976
rect 1220 27740 1500 27976
rect 960 27656 1500 27740
rect 960 27420 984 27656
rect 1220 27420 1500 27656
rect 960 27336 1500 27420
rect 960 27100 984 27336
rect 1220 27100 1500 27336
rect 960 27016 1500 27100
rect 960 26780 984 27016
rect 1220 26780 1500 27016
rect 960 26696 1500 26780
rect 960 26460 984 26696
rect 1220 26460 1500 26696
rect 960 26376 1500 26460
rect 960 26140 984 26376
rect 1220 26140 1500 26376
rect 960 26056 1500 26140
rect 960 25820 984 26056
rect 1220 25820 1500 26056
rect 960 25736 1500 25820
rect 960 25500 984 25736
rect 1220 25500 1500 25736
rect 960 25416 1500 25500
rect 960 25180 984 25416
rect 1220 25180 1500 25416
rect 960 25096 1500 25180
rect 960 24860 984 25096
rect 1220 24860 1500 25096
rect 960 24776 1500 24860
rect 960 24540 984 24776
rect 1220 24540 1500 24776
rect 960 24456 1500 24540
rect 960 24220 984 24456
rect 1220 24220 1500 24456
rect 960 24136 1500 24220
rect 960 23900 984 24136
rect 1220 23900 1500 24136
rect 960 23816 1500 23900
rect 960 23580 984 23816
rect 1220 23580 1500 23816
rect 960 23496 1500 23580
rect 960 23260 984 23496
rect 1220 23260 1500 23496
rect 960 23176 1500 23260
rect 960 22940 984 23176
rect 1220 22940 1500 23176
rect 960 22856 1500 22940
rect 960 22620 984 22856
rect 1220 22620 1500 22856
rect 960 22536 1500 22620
rect 960 22300 984 22536
rect 1220 22300 1500 22536
rect 960 22216 1500 22300
rect 960 21980 984 22216
rect 1220 21980 1500 22216
rect 960 21896 1500 21980
rect 960 21660 984 21896
rect 1220 21660 1500 21896
rect 960 21576 1500 21660
rect 960 21340 984 21576
rect 1220 21340 1500 21576
rect 960 21256 1500 21340
rect 960 21020 984 21256
rect 1220 21020 1500 21256
rect 960 20936 1500 21020
rect 960 20700 984 20936
rect 1220 20700 1500 20936
rect 960 20616 1500 20700
rect 960 20380 984 20616
rect 1220 20380 1500 20616
rect 13500 32446 13780 32682
rect 14016 32446 14040 32682
rect 13500 32362 14040 32446
rect 13500 32126 13780 32362
rect 14016 32126 14040 32362
rect 13500 32042 14040 32126
rect 13500 31806 13780 32042
rect 14016 31806 14040 32042
rect 13500 31722 14040 31806
rect 13500 31486 13780 31722
rect 14016 31486 14040 31722
rect 13500 31402 14040 31486
rect 13500 31166 13780 31402
rect 14016 31166 14040 31402
rect 13500 31082 14040 31166
rect 13500 30846 13780 31082
rect 14016 30846 14040 31082
rect 13500 30762 14040 30846
rect 13500 30526 13780 30762
rect 14016 30526 14040 30762
rect 13500 30442 14040 30526
rect 13500 30206 13780 30442
rect 14016 30206 14040 30442
rect 13500 30122 14040 30206
rect 13500 29886 13780 30122
rect 14016 29886 14040 30122
rect 13500 29802 14040 29886
rect 13500 29566 13780 29802
rect 14016 29566 14040 29802
rect 13500 29482 14040 29566
rect 13500 29246 13780 29482
rect 14016 29246 14040 29482
rect 13500 29162 14040 29246
rect 13500 28926 13780 29162
rect 14016 28926 14040 29162
rect 13500 28842 14040 28926
rect 13500 28606 13780 28842
rect 14016 28606 14040 28842
rect 13500 28522 14040 28606
rect 13500 28286 13780 28522
rect 14016 28286 14040 28522
rect 13500 28202 14040 28286
rect 13500 27966 13780 28202
rect 14016 27966 14040 28202
rect 13500 27882 14040 27966
rect 13500 27646 13780 27882
rect 14016 27646 14040 27882
rect 13500 27562 14040 27646
rect 13500 27326 13780 27562
rect 14016 27326 14040 27562
rect 13500 27242 14040 27326
rect 13500 27006 13780 27242
rect 14016 27006 14040 27242
rect 13500 26922 14040 27006
rect 13500 26686 13780 26922
rect 14016 26686 14040 26922
rect 13500 26602 14040 26686
rect 13500 26366 13780 26602
rect 14016 26366 14040 26602
rect 13500 26282 14040 26366
rect 13500 26046 13780 26282
rect 14016 26046 14040 26282
rect 13500 25962 14040 26046
rect 13500 25726 13780 25962
rect 14016 25726 14040 25962
rect 13500 25642 14040 25726
rect 13500 25406 13780 25642
rect 14016 25406 14040 25642
rect 13500 25322 14040 25406
rect 13500 25086 13780 25322
rect 14016 25086 14040 25322
rect 13500 25002 14040 25086
rect 13500 24766 13780 25002
rect 14016 24766 14040 25002
rect 13500 24682 14040 24766
rect 13500 24446 13780 24682
rect 14016 24446 14040 24682
rect 13500 24362 14040 24446
rect 13500 24126 13780 24362
rect 14016 24126 14040 24362
rect 13500 24042 14040 24126
rect 13500 23806 13780 24042
rect 14016 23806 14040 24042
rect 13500 23722 14040 23806
rect 13500 23486 13780 23722
rect 14016 23486 14040 23722
rect 13500 23402 14040 23486
rect 13500 23166 13780 23402
rect 14016 23166 14040 23402
rect 13500 23082 14040 23166
rect 13500 22846 13780 23082
rect 14016 22846 14040 23082
rect 13500 22762 14040 22846
rect 13500 22526 13780 22762
rect 14016 22526 14040 22762
rect 13500 22442 14040 22526
rect 13500 22206 13780 22442
rect 14016 22206 14040 22442
rect 13500 22122 14040 22206
rect 13500 21886 13780 22122
rect 14016 21886 14040 22122
rect 13500 21802 14040 21886
rect 13500 21566 13780 21802
rect 14016 21566 14040 21802
rect 13500 21482 14040 21566
rect 13500 21246 13780 21482
rect 14016 21246 14040 21482
rect 13500 21162 14040 21246
rect 13500 20926 13780 21162
rect 14016 20926 14040 21162
rect 13500 20842 14040 20926
rect 13500 20606 13780 20842
rect 14016 20606 14040 20842
rect 13500 20522 14040 20606
rect 960 20297 1500 20380
tri 960 20017 1240 20297 ne
rect 1240 20269 1500 20297
rect 1240 20033 1256 20269
rect 1492 20033 1500 20269
rect 1240 20017 1500 20033
tri 1240 20015 1242 20017 ne
rect 1242 20015 1500 20017
tri 1242 19757 1500 20015 ne
tri 1500 19943 2078 20521 sw
tri 13274 20295 13500 20521 se
rect 13500 20295 13761 20522
rect 1500 19757 1582 19943
tri 1500 19697 1560 19757 ne
rect 1560 19707 1582 19757
rect 1818 19933 2078 19943
tri 2078 19933 2088 19943 sw
rect 1818 19757 2088 19933
tri 2088 19757 2264 19933 sw
tri 12864 19885 13274 20295 se
rect 13274 20286 13761 20295
rect 13997 20297 14040 20522
rect 13997 20286 14029 20297
tri 14029 20286 14040 20297 nw
rect 13274 20280 14023 20286
tri 14023 20280 14029 20286 nw
rect 13274 20215 13700 20280
rect 13274 19979 13454 20215
rect 13690 19979 13700 20215
rect 13274 19957 13700 19979
tri 13700 19957 14023 20280 nw
rect 13274 19885 13386 19957
tri 12858 19879 12864 19885 se
rect 12864 19879 13124 19885
tri 12736 19757 12858 19879 se
rect 12858 19757 13124 19879
rect 1818 19707 2264 19757
rect 1560 19697 2264 19707
tri 1560 19377 1880 19697 ne
rect 1880 19629 2264 19697
rect 1880 19393 1896 19629
rect 2132 19531 2264 19629
tri 2264 19531 2490 19757 sw
tri 12510 19531 12736 19757 se
rect 12736 19649 13124 19757
rect 13360 19649 13386 19885
rect 12736 19643 13386 19649
tri 13386 19643 13700 19957 nw
rect 12736 19640 13383 19643
tri 13383 19640 13386 19643 nw
rect 12736 19575 13066 19640
rect 12736 19531 12814 19575
rect 2132 19393 12814 19531
rect 1880 19377 12814 19393
tri 1880 19375 1882 19377 ne
rect 1882 19375 12814 19377
tri 1882 19015 2242 19375 ne
rect 2242 19339 12814 19375
rect 13050 19339 13066 19575
rect 2242 19323 13066 19339
tri 13066 19323 13383 19640 nw
rect 2242 19274 12734 19323
rect 2242 19038 2255 19274
rect 2491 19268 12734 19274
rect 2491 19251 12495 19268
rect 2491 19038 2575 19251
rect 2242 19015 2575 19038
rect 2811 19015 2895 19251
rect 3131 19015 3215 19251
rect 3451 19015 3535 19251
rect 3771 19015 3855 19251
rect 4091 19015 4175 19251
rect 4411 19015 4495 19251
rect 4731 19015 4815 19251
rect 5051 19015 5135 19251
rect 5371 19015 5455 19251
rect 5691 19015 5775 19251
rect 6011 19015 6095 19251
rect 6331 19015 6415 19251
rect 6651 19015 6735 19251
rect 6971 19015 7055 19251
rect 7291 19015 7375 19251
rect 7611 19015 7695 19251
rect 7931 19015 8015 19251
rect 8251 19015 8335 19251
rect 8571 19015 8655 19251
rect 8891 19015 8975 19251
rect 9211 19015 9295 19251
rect 9531 19015 9615 19251
rect 9851 19015 9935 19251
rect 10171 19015 10255 19251
rect 10491 19015 10575 19251
rect 10811 19015 10895 19251
rect 11131 19015 11215 19251
rect 11451 19015 11535 19251
rect 11771 19015 11855 19251
rect 12091 19015 12175 19251
rect 12411 19032 12495 19251
rect 12731 19032 12734 19268
rect 12411 19015 12734 19032
tri 2242 18991 2266 19015 ne
rect 2266 18991 12734 19015
tri 12734 18991 13066 19323 nw
<< via4 >>
rect 2269 33791 2505 34027
rect 2589 33811 2825 34047
rect 2909 33811 3145 34047
rect 3229 33811 3465 34047
rect 3549 33811 3785 34047
rect 3869 33811 4105 34047
rect 4189 33811 4425 34047
rect 4509 33811 4745 34047
rect 4829 33811 5065 34047
rect 5149 33811 5385 34047
rect 5469 33811 5705 34047
rect 5789 33811 6025 34047
rect 6109 33811 6345 34047
rect 6429 33811 6665 34047
rect 6749 33811 6985 34047
rect 7069 33811 7305 34047
rect 7389 33811 7625 34047
rect 7709 33811 7945 34047
rect 8029 33811 8265 34047
rect 8349 33811 8585 34047
rect 8669 33811 8905 34047
rect 8989 33811 9225 34047
rect 9309 33811 9545 34047
rect 9629 33811 9865 34047
rect 9949 33811 10185 34047
rect 10269 33811 10505 34047
rect 10589 33811 10825 34047
rect 10909 33811 11145 34047
rect 11229 33811 11465 34047
rect 11549 33811 11785 34047
rect 11869 33811 12105 34047
rect 12189 33811 12425 34047
rect 12509 33779 12745 34015
rect 1950 33487 2186 33723
rect 1630 33167 1866 33403
rect 12868 33433 13104 33669
rect 1333 32847 1569 33083
rect 1048 32540 1284 32776
rect 13188 33113 13424 33349
rect 13508 32793 13744 33029
rect 984 32220 1220 32456
rect 984 31900 1220 32136
rect 984 31580 1220 31816
rect 984 31260 1220 31496
rect 984 30940 1220 31176
rect 984 30620 1220 30856
rect 984 30300 1220 30536
rect 984 29980 1220 30216
rect 984 29660 1220 29896
rect 984 29340 1220 29576
rect 984 29020 1220 29256
rect 984 28700 1220 28936
rect 984 28380 1220 28616
rect 984 28060 1220 28296
rect 984 27740 1220 27976
rect 984 27420 1220 27656
rect 984 27100 1220 27336
rect 984 26780 1220 27016
rect 984 26460 1220 26696
rect 984 26140 1220 26376
rect 984 25820 1220 26056
rect 984 25500 1220 25736
rect 984 25180 1220 25416
rect 984 24860 1220 25096
rect 984 24540 1220 24776
rect 984 24220 1220 24456
rect 984 23900 1220 24136
rect 984 23580 1220 23816
rect 984 23260 1220 23496
rect 984 22940 1220 23176
rect 984 22620 1220 22856
rect 984 22300 1220 22536
rect 984 21980 1220 22216
rect 984 21660 1220 21896
rect 984 21340 1220 21576
rect 984 21020 1220 21256
rect 984 20700 1220 20936
rect 984 20380 1220 20616
rect 13780 32446 14016 32682
rect 13780 32126 14016 32362
rect 13780 31806 14016 32042
rect 13780 31486 14016 31722
rect 13780 31166 14016 31402
rect 13780 30846 14016 31082
rect 13780 30526 14016 30762
rect 13780 30206 14016 30442
rect 13780 29886 14016 30122
rect 13780 29566 14016 29802
rect 13780 29246 14016 29482
rect 13780 28926 14016 29162
rect 13780 28606 14016 28842
rect 13780 28286 14016 28522
rect 13780 27966 14016 28202
rect 13780 27646 14016 27882
rect 13780 27326 14016 27562
rect 13780 27006 14016 27242
rect 13780 26686 14016 26922
rect 13780 26366 14016 26602
rect 13780 26046 14016 26282
rect 13780 25726 14016 25962
rect 13780 25406 14016 25642
rect 13780 25086 14016 25322
rect 13780 24766 14016 25002
rect 13780 24446 14016 24682
rect 13780 24126 14016 24362
rect 13780 23806 14016 24042
rect 13780 23486 14016 23722
rect 13780 23166 14016 23402
rect 13780 22846 14016 23082
rect 13780 22526 14016 22762
rect 13780 22206 14016 22442
rect 13780 21886 14016 22122
rect 13780 21566 14016 21802
rect 13780 21246 14016 21482
rect 13780 20926 14016 21162
rect 13780 20606 14016 20842
rect 1256 20033 1492 20269
rect 1582 19707 1818 19943
rect 13761 20286 13997 20522
rect 13454 19979 13690 20215
rect 1896 19393 2132 19629
rect 13124 19649 13360 19885
rect 12814 19339 13050 19575
rect 2255 19038 2491 19274
rect 2575 19015 2811 19251
rect 2895 19015 3131 19251
rect 3215 19015 3451 19251
rect 3535 19015 3771 19251
rect 3855 19015 4091 19251
rect 4175 19015 4411 19251
rect 4495 19015 4731 19251
rect 4815 19015 5051 19251
rect 5135 19015 5371 19251
rect 5455 19015 5691 19251
rect 5775 19015 6011 19251
rect 6095 19015 6331 19251
rect 6415 19015 6651 19251
rect 6735 19015 6971 19251
rect 7055 19015 7291 19251
rect 7375 19015 7611 19251
rect 7695 19015 7931 19251
rect 8015 19015 8251 19251
rect 8335 19015 8571 19251
rect 8655 19015 8891 19251
rect 8975 19015 9211 19251
rect 9295 19015 9531 19251
rect 9615 19015 9851 19251
rect 9935 19015 10171 19251
rect 10255 19015 10491 19251
rect 10575 19015 10811 19251
rect 10895 19015 11131 19251
rect 11215 19015 11451 19251
rect 11535 19015 11771 19251
rect 11855 19015 12091 19251
rect 12175 19015 12411 19251
rect 12495 19032 12731 19268
<< metal5 >>
tri 1934 33739 2266 34071 se
rect 2266 34047 12734 34071
tri 12734 34047 12758 34071 sw
rect 2266 34027 2589 34047
rect 2266 33791 2269 34027
rect 2505 33811 2589 34027
rect 2825 33811 2909 34047
rect 3145 33811 3229 34047
rect 3465 33811 3549 34047
rect 3785 33811 3869 34047
rect 4105 33811 4189 34047
rect 4425 33811 4509 34047
rect 4745 33811 4829 34047
rect 5065 33811 5149 34047
rect 5385 33811 5469 34047
rect 5705 33811 5789 34047
rect 6025 33811 6109 34047
rect 6345 33811 6429 34047
rect 6665 33811 6749 34047
rect 6985 33811 7069 34047
rect 7305 33811 7389 34047
rect 7625 33811 7709 34047
rect 7945 33811 8029 34047
rect 8265 33811 8349 34047
rect 8585 33811 8669 34047
rect 8905 33811 8989 34047
rect 9225 33811 9309 34047
rect 9545 33811 9629 34047
rect 9865 33811 9949 34047
rect 10185 33811 10269 34047
rect 10505 33811 10589 34047
rect 10825 33811 10909 34047
rect 11145 33811 11229 34047
rect 11465 33811 11549 34047
rect 11785 33811 11869 34047
rect 12105 33811 12189 34047
rect 12425 34015 12758 34047
rect 12425 33811 12509 34015
rect 2505 33791 12509 33811
rect 2266 33779 12509 33791
rect 12745 33779 12758 34015
rect 2266 33739 12758 33779
tri 1731 33536 1934 33739 se
rect 1934 33723 12758 33739
rect 1934 33536 1950 33723
tri 1614 33419 1731 33536 se
rect 1731 33487 1950 33536
rect 2186 33685 12758 33723
tri 12758 33685 13120 34047 sw
rect 2186 33683 13120 33685
rect 2186 33663 2405 33683
tri 2405 33663 2425 33683 nw
tri 12578 33663 12598 33683 ne
rect 12598 33669 13120 33683
rect 12598 33663 12868 33669
rect 2186 33648 2390 33663
tri 2390 33648 2405 33663 nw
rect 2186 33620 2362 33648
tri 2362 33620 2390 33648 nw
tri 2405 33635 2433 33663 se
rect 2433 33635 12570 33663
tri 12570 33635 12598 33663 sw
tri 12598 33635 12626 33663 ne
rect 12626 33635 12868 33663
tri 2390 33620 2405 33635 se
rect 2405 33620 12598 33635
rect 2186 33592 2334 33620
tri 2334 33592 2362 33620 nw
tri 2362 33592 2390 33620 se
rect 2390 33607 12598 33620
tri 12598 33607 12626 33635 sw
tri 12626 33607 12654 33635 ne
rect 12654 33607 12868 33635
rect 2390 33592 12626 33607
rect 2186 33564 2306 33592
tri 2306 33564 2334 33592 nw
tri 2334 33564 2362 33592 se
rect 2362 33579 12626 33592
tri 12626 33579 12654 33607 sw
tri 12654 33579 12682 33607 ne
rect 12682 33579 12868 33607
rect 2362 33564 12654 33579
rect 2186 33536 2278 33564
tri 2278 33536 2306 33564 nw
tri 2306 33536 2334 33564 se
rect 2334 33551 12654 33564
tri 12654 33551 12682 33579 sw
tri 12682 33551 12710 33579 ne
rect 12710 33551 12868 33579
rect 2334 33536 12682 33551
rect 2186 33508 2250 33536
tri 2250 33508 2278 33536 nw
tri 2278 33508 2306 33536 se
rect 2306 33523 12682 33536
tri 12682 33523 12710 33551 sw
tri 12710 33523 12738 33551 ne
rect 12738 33523 12868 33551
rect 2306 33508 12710 33523
rect 2186 33487 2222 33508
rect 1731 33480 2222 33487
tri 2222 33480 2250 33508 nw
tri 2250 33480 2278 33508 se
rect 2278 33495 12710 33508
tri 12710 33495 12738 33523 sw
tri 12738 33495 12766 33523 ne
rect 12766 33495 12868 33523
rect 2278 33480 12738 33495
rect 1731 33452 2194 33480
tri 2194 33452 2222 33480 nw
tri 2222 33452 2250 33480 se
rect 2250 33467 12738 33480
tri 12738 33467 12766 33495 sw
tri 12766 33467 12794 33495 ne
rect 12794 33467 12868 33495
rect 2250 33452 12766 33467
rect 1731 33424 2166 33452
tri 2166 33424 2194 33452 nw
tri 2194 33424 2222 33452 se
rect 2222 33439 12766 33452
tri 12766 33439 12794 33467 sw
tri 12794 33439 12822 33467 ne
rect 12822 33439 12868 33467
rect 2222 33424 12794 33439
rect 1731 33419 2138 33424
tri 1294 33099 1614 33419 se
rect 1614 33403 2138 33419
rect 1614 33167 1630 33403
rect 1866 33396 2138 33403
tri 2138 33396 2166 33424 nw
tri 2166 33396 2194 33424 se
rect 2194 33411 12794 33424
tri 12794 33411 12822 33439 sw
tri 12822 33411 12850 33439 ne
rect 12850 33433 12868 33439
rect 13104 33433 13120 33669
rect 12850 33411 13120 33433
rect 2194 33396 12822 33411
rect 1866 33368 2110 33396
tri 2110 33368 2138 33396 nw
tri 2138 33368 2166 33396 se
rect 2166 33383 12822 33396
tri 12822 33383 12850 33411 sw
tri 12850 33383 12878 33411 ne
rect 12878 33383 13120 33411
rect 2166 33368 12850 33383
rect 1866 33340 2082 33368
tri 2082 33340 2110 33368 nw
tri 2110 33340 2138 33368 se
rect 2138 33355 12850 33368
tri 12850 33355 12878 33383 sw
tri 12878 33355 12906 33383 ne
rect 12906 33365 13120 33383
tri 13120 33365 13440 33685 sw
rect 12906 33355 13440 33365
rect 2138 33340 12878 33355
rect 1866 33312 2054 33340
tri 2054 33312 2082 33340 nw
tri 2082 33312 2110 33340 se
rect 2110 33327 12878 33340
tri 12878 33327 12906 33355 sw
tri 12906 33327 12934 33355 ne
rect 12934 33349 13440 33355
rect 12934 33327 13188 33349
rect 2110 33312 12906 33327
rect 1866 33284 2026 33312
tri 2026 33284 2054 33312 nw
tri 2054 33284 2082 33312 se
rect 2082 33299 12906 33312
tri 12906 33299 12934 33327 sw
tri 12934 33299 12962 33327 ne
rect 12962 33299 13188 33327
rect 2082 33284 12934 33299
rect 1866 33256 1998 33284
tri 1998 33256 2026 33284 nw
tri 2026 33256 2054 33284 se
rect 2054 33271 12934 33284
tri 12934 33271 12962 33299 sw
tri 12962 33271 12990 33299 ne
rect 12990 33271 13188 33299
rect 2054 33256 12962 33271
rect 1866 33228 1970 33256
tri 1970 33228 1998 33256 nw
tri 1998 33228 2026 33256 se
rect 2026 33243 12962 33256
tri 12962 33243 12990 33271 sw
tri 12990 33243 13018 33271 ne
rect 13018 33243 13188 33271
rect 2026 33228 12990 33243
rect 1866 33200 1942 33228
tri 1942 33200 1970 33228 nw
tri 1970 33200 1998 33228 se
rect 1998 33215 12990 33228
tri 12990 33215 13018 33243 sw
tri 13018 33215 13046 33243 ne
rect 13046 33215 13188 33243
rect 1998 33200 13018 33215
rect 1866 33172 1914 33200
tri 1914 33172 1942 33200 nw
tri 1942 33172 1970 33200 se
rect 1970 33187 13018 33200
tri 13018 33187 13046 33215 sw
tri 13046 33187 13074 33215 ne
rect 13074 33187 13188 33215
rect 1970 33172 13046 33187
rect 1866 33167 1886 33172
rect 1614 33144 1886 33167
tri 1886 33144 1914 33172 nw
tri 1914 33144 1942 33172 se
rect 1942 33159 13046 33172
tri 13046 33159 13074 33187 sw
tri 13074 33159 13102 33187 ne
rect 13102 33159 13188 33187
rect 1942 33144 13074 33159
rect 1614 33116 1858 33144
tri 1858 33116 1886 33144 nw
tri 1886 33116 1914 33144 se
rect 1914 33131 13074 33144
tri 13074 33131 13102 33159 sw
tri 13102 33131 13130 33159 ne
rect 13130 33131 13188 33159
rect 1914 33116 13102 33131
rect 1614 33099 1830 33116
tri 1199 33004 1294 33099 se
rect 1294 33088 1830 33099
tri 1830 33088 1858 33116 nw
tri 1858 33088 1886 33116 se
rect 1886 33103 13102 33116
tri 13102 33103 13130 33131 sw
tri 13130 33103 13158 33131 ne
rect 13158 33113 13188 33131
rect 13424 33113 13440 33349
rect 13158 33103 13440 33113
rect 1886 33088 13130 33103
rect 1294 33083 1802 33088
rect 1294 33004 1333 33083
tri 971 32776 1199 33004 se
rect 1199 32847 1333 33004
rect 1569 33060 1802 33083
tri 1802 33060 1830 33088 nw
tri 1830 33060 1858 33088 se
rect 1858 33075 13130 33088
tri 13130 33075 13158 33103 sw
tri 13158 33075 13186 33103 ne
rect 13186 33075 13440 33103
rect 1858 33060 13158 33075
rect 1569 33032 1774 33060
tri 1774 33032 1802 33060 nw
tri 1802 33032 1830 33060 se
rect 1830 33047 13158 33060
tri 13158 33047 13186 33075 sw
tri 13186 33047 13214 33075 ne
rect 13214 33047 13440 33075
rect 1830 33032 13186 33047
rect 1569 33004 1746 33032
tri 1746 33004 1774 33032 nw
tri 1774 33004 1802 33032 se
rect 1802 33019 13186 33032
tri 13186 33019 13214 33047 sw
tri 13214 33019 13242 33047 ne
rect 13242 33045 13440 33047
tri 13440 33045 13760 33365 sw
rect 13242 33029 13760 33045
rect 13242 33019 13508 33029
rect 1802 33004 13214 33019
rect 1569 32976 1718 33004
tri 1718 32976 1746 33004 nw
tri 1746 32976 1774 33004 se
rect 1774 32991 13214 33004
tri 13214 32991 13242 33019 sw
tri 13242 32991 13270 33019 ne
rect 13270 32991 13508 33019
rect 1774 32976 13242 32991
rect 1569 32948 1690 32976
tri 1690 32948 1718 32976 nw
tri 1718 32948 1746 32976 se
rect 1746 32963 13242 32976
tri 13242 32963 13270 32991 sw
tri 13270 32963 13298 32991 ne
rect 13298 32963 13508 32991
rect 1746 32948 13270 32963
rect 1569 32920 1662 32948
tri 1662 32920 1690 32948 nw
tri 1690 32920 1718 32948 se
rect 1718 32935 13270 32948
tri 13270 32935 13298 32963 sw
tri 13298 32935 13326 32963 ne
rect 13326 32935 13508 32963
rect 1718 32920 13298 32935
rect 1569 32892 1634 32920
tri 1634 32892 1662 32920 nw
tri 1662 32892 1690 32920 se
rect 1690 32907 13298 32920
tri 13298 32907 13326 32935 sw
tri 13326 32907 13354 32935 ne
rect 13354 32907 13508 32935
rect 1690 32892 13326 32907
rect 1569 32864 1606 32892
tri 1606 32864 1634 32892 nw
tri 1634 32864 1662 32892 se
rect 1662 32879 13326 32892
tri 13326 32879 13354 32907 sw
tri 13354 32879 13382 32907 ne
rect 13382 32879 13508 32907
rect 1662 32864 13354 32879
rect 1569 32847 1578 32864
rect 1199 32836 1578 32847
tri 1578 32836 1606 32864 nw
tri 1606 32836 1634 32864 se
rect 1634 32851 13354 32864
tri 13354 32851 13382 32879 sw
tri 13382 32851 13410 32879 ne
rect 13410 32851 13508 32879
rect 1634 32836 13382 32851
rect 1199 32808 1550 32836
tri 1550 32808 1578 32836 nw
tri 1578 32808 1606 32836 se
rect 1606 32823 13382 32836
tri 13382 32823 13410 32851 sw
tri 13410 32823 13438 32851 ne
rect 13438 32823 13508 32851
rect 1606 32808 13410 32823
rect 1199 32780 1522 32808
tri 1522 32780 1550 32808 nw
tri 1550 32780 1578 32808 se
rect 1578 32795 13410 32808
tri 13410 32795 13438 32823 sw
tri 13438 32795 13466 32823 ne
rect 13466 32795 13508 32823
rect 1578 32780 13438 32795
rect 1199 32776 1494 32780
tri 960 32765 971 32776 se
rect 971 32765 1048 32776
rect 960 32540 1048 32765
rect 1284 32752 1494 32776
tri 1494 32752 1522 32780 nw
tri 1522 32752 1550 32780 se
rect 1550 32767 13438 32780
tri 13438 32767 13466 32795 sw
tri 13466 32767 13494 32795 ne
rect 13494 32793 13508 32795
rect 13744 32793 13760 33029
rect 13494 32767 13760 32793
rect 1550 32752 13466 32767
rect 1284 32724 1466 32752
tri 1466 32724 1494 32752 nw
tri 1494 32724 1522 32752 se
rect 1522 32739 13466 32752
tri 13466 32739 13494 32767 sw
tri 13494 32739 13522 32767 ne
rect 13522 32765 13760 32767
tri 13760 32765 14040 33045 sw
rect 13522 32739 14040 32765
rect 1522 32724 13494 32739
rect 1284 32696 1438 32724
tri 1438 32696 1466 32724 nw
tri 1466 32696 1494 32724 se
rect 1494 32711 13494 32724
tri 13494 32711 13522 32739 sw
tri 13522 32711 13550 32739 ne
rect 13550 32711 14040 32739
rect 1494 32696 13522 32711
rect 1284 32668 1410 32696
tri 1410 32668 1438 32696 nw
tri 1438 32668 1466 32696 se
rect 1466 32683 13522 32696
tri 13522 32683 13550 32711 sw
tri 13550 32683 13578 32711 ne
rect 13578 32683 14040 32711
rect 1466 32668 13550 32683
rect 1284 32640 1382 32668
tri 1382 32640 1410 32668 nw
tri 1410 32640 1438 32668 se
rect 1438 32655 13550 32668
tri 13550 32655 13578 32683 sw
tri 13578 32655 13606 32683 ne
rect 13606 32682 14040 32683
rect 13606 32655 13780 32682
rect 1438 32640 13578 32655
rect 1284 32612 1354 32640
tri 1354 32612 1382 32640 nw
tri 1382 32612 1410 32640 se
rect 1410 32629 13578 32640
tri 13578 32629 13604 32655 sw
tri 13606 32637 13624 32655 ne
rect 1410 32612 13604 32629
rect 1284 32540 1334 32612
tri 1334 32592 1354 32612 nw
rect 960 32456 1334 32540
rect 960 32220 984 32456
rect 1220 32220 1334 32456
rect 960 32136 1334 32220
rect 960 31900 984 32136
rect 1220 31900 1334 32136
rect 960 31816 1334 31900
rect 960 31580 984 31816
rect 1220 31580 1334 31816
rect 960 31496 1334 31580
rect 960 31260 984 31496
rect 1220 31260 1334 31496
rect 960 31176 1334 31260
rect 960 30940 984 31176
rect 1220 30940 1334 31176
rect 960 30856 1334 30940
rect 960 30620 984 30856
rect 1220 30620 1334 30856
rect 960 30536 1334 30620
rect 960 30300 984 30536
rect 1220 30300 1334 30536
rect 960 30216 1334 30300
rect 960 29980 984 30216
rect 1220 29980 1334 30216
rect 960 29896 1334 29980
rect 960 29660 984 29896
rect 1220 29660 1334 29896
rect 960 29576 1334 29660
rect 960 29340 984 29576
rect 1220 29340 1334 29576
rect 960 29256 1334 29340
rect 960 29020 984 29256
rect 1220 29020 1334 29256
rect 960 28936 1334 29020
rect 960 28700 984 28936
rect 1220 28700 1334 28936
rect 960 28616 1334 28700
rect 960 28380 984 28616
rect 1220 28380 1334 28616
rect 960 28296 1334 28380
rect 960 28060 984 28296
rect 1220 28060 1334 28296
rect 960 27976 1334 28060
rect 960 27740 984 27976
rect 1220 27740 1334 27976
rect 960 27656 1334 27740
rect 960 27420 984 27656
rect 1220 27420 1334 27656
rect 960 27336 1334 27420
rect 960 27100 984 27336
rect 1220 27100 1334 27336
rect 960 27016 1334 27100
rect 960 26780 984 27016
rect 1220 26780 1334 27016
rect 960 26696 1334 26780
rect 960 26460 984 26696
rect 1220 26460 1334 26696
rect 960 26376 1334 26460
rect 960 26140 984 26376
rect 1220 26140 1334 26376
rect 960 26056 1334 26140
rect 960 25820 984 26056
rect 1220 25820 1334 26056
rect 960 25736 1334 25820
rect 960 25500 984 25736
rect 1220 25500 1334 25736
rect 960 25416 1334 25500
rect 960 25180 984 25416
rect 1220 25180 1334 25416
rect 960 25096 1334 25180
rect 960 24860 984 25096
rect 1220 24860 1334 25096
rect 960 24776 1334 24860
rect 960 24540 984 24776
rect 1220 24540 1334 24776
rect 960 24456 1334 24540
rect 960 24220 984 24456
rect 1220 24220 1334 24456
rect 960 24136 1334 24220
rect 960 23900 984 24136
rect 1220 23900 1334 24136
rect 960 23816 1334 23900
rect 960 23580 984 23816
rect 1220 23580 1334 23816
rect 960 23496 1334 23580
rect 960 23260 984 23496
rect 1220 23260 1334 23496
rect 960 23176 1334 23260
rect 960 22940 984 23176
rect 1220 22940 1334 23176
rect 960 22856 1334 22940
rect 960 22620 984 22856
rect 1220 22620 1334 22856
rect 960 22536 1334 22620
rect 960 22300 984 22536
rect 1220 22300 1334 22536
rect 960 22216 1334 22300
rect 960 21980 984 22216
rect 1220 21980 1334 22216
rect 960 21896 1334 21980
rect 960 21660 984 21896
rect 1220 21660 1334 21896
rect 960 21576 1334 21660
rect 960 21340 984 21576
rect 1220 21340 1334 21576
rect 960 21256 1334 21340
rect 960 21020 984 21256
rect 1220 21020 1334 21256
rect 960 20936 1334 21020
rect 960 20700 984 20936
rect 1220 20700 1334 20936
rect 960 20616 1334 20700
rect 960 20380 984 20616
rect 1220 20500 1334 20616
tri 1354 32584 1382 32612 se
rect 1382 32584 13604 32612
rect 1354 20528 13604 32584
tri 1334 20500 1354 20520 sw
tri 1354 20500 1382 20528 ne
rect 1382 20500 13604 20528
rect 1220 20475 1354 20500
tri 1354 20475 1379 20500 sw
tri 1382 20475 1407 20500 ne
rect 1407 20475 13604 20500
rect 1220 20447 1379 20475
tri 1379 20447 1407 20475 sw
tri 1407 20447 1435 20475 ne
rect 1435 20473 13604 20475
rect 1435 20447 13576 20473
rect 1220 20419 1407 20447
tri 1407 20419 1435 20447 sw
tri 1435 20419 1463 20447 ne
rect 1463 20445 13576 20447
tri 13576 20445 13604 20473 nw
rect 13624 32446 13780 32655
rect 14016 32446 14040 32682
rect 13624 32362 14040 32446
rect 13624 32126 13780 32362
rect 14016 32126 14040 32362
rect 13624 32042 14040 32126
rect 13624 31806 13780 32042
rect 14016 31806 14040 32042
rect 13624 31722 14040 31806
rect 13624 31486 13780 31722
rect 14016 31486 14040 31722
rect 13624 31402 14040 31486
rect 13624 31166 13780 31402
rect 14016 31166 14040 31402
rect 13624 31082 14040 31166
rect 13624 30846 13780 31082
rect 14016 30846 14040 31082
rect 13624 30762 14040 30846
rect 13624 30526 13780 30762
rect 14016 30526 14040 30762
rect 13624 30442 14040 30526
rect 13624 30206 13780 30442
rect 14016 30206 14040 30442
rect 13624 30122 14040 30206
rect 13624 29886 13780 30122
rect 14016 29886 14040 30122
rect 13624 29802 14040 29886
rect 13624 29566 13780 29802
rect 14016 29566 14040 29802
rect 13624 29482 14040 29566
rect 13624 29246 13780 29482
rect 14016 29246 14040 29482
rect 13624 29162 14040 29246
rect 13624 28926 13780 29162
rect 14016 28926 14040 29162
rect 13624 28842 14040 28926
rect 13624 28606 13780 28842
rect 14016 28606 14040 28842
rect 13624 28522 14040 28606
rect 13624 28286 13780 28522
rect 14016 28286 14040 28522
rect 13624 28202 14040 28286
rect 13624 27966 13780 28202
rect 14016 27966 14040 28202
rect 13624 27882 14040 27966
rect 13624 27646 13780 27882
rect 14016 27646 14040 27882
rect 13624 27562 14040 27646
rect 13624 27326 13780 27562
rect 14016 27326 14040 27562
rect 13624 27242 14040 27326
rect 13624 27006 13780 27242
rect 14016 27006 14040 27242
rect 13624 26922 14040 27006
rect 13624 26686 13780 26922
rect 14016 26686 14040 26922
rect 13624 26602 14040 26686
rect 13624 26366 13780 26602
rect 14016 26366 14040 26602
rect 13624 26282 14040 26366
rect 13624 26046 13780 26282
rect 14016 26046 14040 26282
rect 13624 25962 14040 26046
rect 13624 25726 13780 25962
rect 14016 25726 14040 25962
rect 13624 25642 14040 25726
rect 13624 25406 13780 25642
rect 14016 25406 14040 25642
rect 13624 25322 14040 25406
rect 13624 25086 13780 25322
rect 14016 25086 14040 25322
rect 13624 25002 14040 25086
rect 13624 24766 13780 25002
rect 14016 24766 14040 25002
rect 13624 24682 14040 24766
rect 13624 24446 13780 24682
rect 14016 24446 14040 24682
rect 13624 24362 14040 24446
rect 13624 24126 13780 24362
rect 14016 24126 14040 24362
rect 13624 24042 14040 24126
rect 13624 23806 13780 24042
rect 14016 23806 14040 24042
rect 13624 23722 14040 23806
rect 13624 23486 13780 23722
rect 14016 23486 14040 23722
rect 13624 23402 14040 23486
rect 13624 23166 13780 23402
rect 14016 23166 14040 23402
rect 13624 23082 14040 23166
rect 13624 22846 13780 23082
rect 14016 22846 14040 23082
rect 13624 22762 14040 22846
rect 13624 22526 13780 22762
rect 14016 22526 14040 22762
rect 13624 22442 14040 22526
rect 13624 22206 13780 22442
rect 14016 22206 14040 22442
rect 13624 22122 14040 22206
rect 13624 21886 13780 22122
rect 14016 21886 14040 22122
rect 13624 21802 14040 21886
rect 13624 21566 13780 21802
rect 14016 21566 14040 21802
rect 13624 21482 14040 21566
rect 13624 21246 13780 21482
rect 14016 21246 14040 21482
rect 13624 21162 14040 21246
rect 13624 20926 13780 21162
rect 14016 20926 14040 21162
rect 13624 20842 14040 20926
rect 13624 20606 13780 20842
rect 14016 20606 14040 20842
rect 13624 20522 14040 20606
tri 13604 20445 13624 20465 se
rect 13624 20445 13761 20522
rect 1463 20419 13548 20445
rect 1220 20391 1435 20419
tri 1435 20391 1463 20419 sw
tri 1463 20391 1491 20419 ne
rect 1491 20417 13548 20419
tri 13548 20417 13576 20445 nw
tri 13576 20417 13604 20445 se
rect 13604 20417 13761 20445
rect 1491 20391 13520 20417
rect 1220 20380 1463 20391
rect 960 20363 1463 20380
tri 1463 20363 1491 20391 sw
tri 1491 20363 1519 20391 ne
rect 1519 20389 13520 20391
tri 13520 20389 13548 20417 nw
tri 13548 20389 13576 20417 se
rect 13576 20389 13761 20417
rect 1519 20363 13492 20389
rect 960 20335 1491 20363
tri 1491 20335 1519 20363 sw
tri 1519 20335 1547 20363 ne
rect 1547 20361 13492 20363
tri 13492 20361 13520 20389 nw
tri 13520 20361 13548 20389 se
rect 13548 20361 13761 20389
rect 1547 20335 13464 20361
rect 960 20307 1519 20335
tri 1519 20307 1547 20335 sw
tri 1547 20307 1575 20335 ne
rect 1575 20333 13464 20335
tri 13464 20333 13492 20361 nw
tri 13492 20333 13520 20361 se
rect 13520 20333 13761 20361
rect 1575 20307 13436 20333
rect 960 20297 1547 20307
tri 960 20017 1240 20297 ne
rect 1240 20279 1547 20297
tri 1547 20279 1575 20307 sw
tri 1575 20279 1603 20307 ne
rect 1603 20305 13436 20307
tri 13436 20305 13464 20333 nw
tri 13464 20305 13492 20333 se
rect 13492 20305 13761 20333
rect 1603 20279 13408 20305
rect 1240 20269 1575 20279
rect 1240 20033 1256 20269
rect 1492 20251 1575 20269
tri 1575 20251 1603 20279 sw
tri 1603 20251 1631 20279 ne
rect 1631 20277 13408 20279
tri 13408 20277 13436 20305 nw
tri 13436 20277 13464 20305 se
rect 13464 20286 13761 20305
rect 13997 20297 14040 20522
rect 13997 20286 14020 20297
rect 13464 20277 14020 20286
tri 14020 20277 14040 20297 nw
rect 1631 20251 13380 20277
rect 1492 20223 1603 20251
tri 1603 20223 1631 20251 sw
tri 1631 20223 1659 20251 ne
rect 1659 20249 13380 20251
tri 13380 20249 13408 20277 nw
tri 13408 20249 13436 20277 se
rect 13436 20249 13706 20277
rect 1659 20223 13352 20249
rect 1492 20195 1631 20223
tri 1631 20195 1659 20223 sw
tri 1659 20195 1687 20223 ne
rect 1687 20221 13352 20223
tri 13352 20221 13380 20249 nw
tri 13380 20221 13408 20249 se
rect 13408 20221 13706 20249
rect 1687 20195 13324 20221
rect 1492 20167 1659 20195
tri 1659 20167 1687 20195 sw
tri 1687 20167 1715 20195 ne
rect 1715 20193 13324 20195
tri 13324 20193 13352 20221 nw
tri 13352 20193 13380 20221 se
rect 13380 20215 13706 20221
rect 13380 20193 13454 20215
rect 1715 20167 13296 20193
rect 1492 20139 1687 20167
tri 1687 20139 1715 20167 sw
tri 1715 20139 1743 20167 ne
rect 1743 20165 13296 20167
tri 13296 20165 13324 20193 nw
tri 13324 20165 13352 20193 se
rect 13352 20165 13454 20193
rect 1743 20139 13268 20165
rect 1492 20111 1715 20139
tri 1715 20111 1743 20139 sw
tri 1743 20111 1771 20139 ne
rect 1771 20137 13268 20139
tri 13268 20137 13296 20165 nw
tri 13296 20137 13324 20165 se
rect 13324 20137 13454 20165
rect 1771 20111 13240 20137
rect 1492 20083 1743 20111
tri 1743 20083 1771 20111 sw
tri 1771 20083 1799 20111 ne
rect 1799 20109 13240 20111
tri 13240 20109 13268 20137 nw
tri 13268 20109 13296 20137 se
rect 13296 20109 13454 20137
rect 1799 20083 13212 20109
rect 1492 20055 1771 20083
tri 1771 20055 1799 20083 sw
tri 1799 20055 1827 20083 ne
rect 1827 20081 13212 20083
tri 13212 20081 13240 20109 nw
tri 13240 20081 13268 20109 se
rect 13268 20081 13454 20109
rect 1827 20055 13184 20081
rect 1492 20033 1799 20055
rect 1240 20027 1799 20033
tri 1799 20027 1827 20055 sw
tri 1827 20027 1855 20055 ne
rect 1855 20053 13184 20055
tri 13184 20053 13212 20081 nw
tri 13212 20053 13240 20081 se
rect 13240 20053 13454 20081
rect 1855 20027 13156 20053
rect 1240 20017 1827 20027
tri 1240 19691 1566 20017 ne
rect 1566 19999 1827 20017
tri 1827 19999 1855 20027 sw
tri 1855 19999 1883 20027 ne
rect 1883 20025 13156 20027
tri 13156 20025 13184 20053 nw
tri 13184 20025 13212 20053 se
rect 13212 20025 13454 20053
rect 1883 19999 13128 20025
rect 1566 19971 1855 19999
tri 1855 19971 1883 19999 sw
tri 1883 19971 1911 19999 ne
rect 1911 19997 13128 19999
tri 13128 19997 13156 20025 nw
tri 13156 19997 13184 20025 se
rect 13184 19997 13454 20025
rect 1911 19971 13100 19997
rect 1566 19943 1883 19971
tri 1883 19943 1911 19971 sw
tri 1911 19943 1939 19971 ne
rect 1939 19969 13100 19971
tri 13100 19969 13128 19997 nw
tri 13128 19969 13156 19997 se
rect 13156 19979 13454 19997
rect 13690 19979 13706 20215
rect 13156 19969 13706 19979
rect 1939 19943 13072 19969
rect 1566 19707 1582 19943
rect 1818 19915 1911 19943
tri 1911 19915 1939 19943 sw
tri 1939 19915 1967 19943 ne
rect 1967 19941 13072 19943
tri 13072 19941 13100 19969 nw
tri 13100 19941 13128 19969 se
rect 13128 19963 13706 19969
tri 13706 19963 14020 20277 nw
rect 13128 19941 13383 19963
rect 1967 19915 13044 19941
rect 1818 19887 1939 19915
tri 1939 19887 1967 19915 sw
tri 1967 19887 1995 19915 ne
rect 1995 19913 13044 19915
tri 13044 19913 13072 19941 nw
tri 13072 19913 13100 19941 se
rect 13100 19913 13383 19941
rect 1995 19887 13016 19913
rect 1818 19859 1967 19887
tri 1967 19859 1995 19887 sw
tri 1995 19859 2023 19887 ne
rect 2023 19885 13016 19887
tri 13016 19885 13044 19913 nw
tri 13044 19885 13072 19913 se
rect 13072 19885 13383 19913
rect 2023 19859 12988 19885
rect 1818 19831 1995 19859
tri 1995 19831 2023 19859 sw
tri 2023 19831 2051 19859 ne
rect 2051 19857 12988 19859
tri 12988 19857 13016 19885 nw
tri 13016 19857 13044 19885 se
rect 13044 19857 13124 19885
rect 2051 19831 12960 19857
rect 1818 19803 2023 19831
tri 2023 19803 2051 19831 sw
tri 2051 19803 2079 19831 ne
rect 2079 19829 12960 19831
tri 12960 19829 12988 19857 nw
tri 12988 19829 13016 19857 se
rect 13016 19829 13124 19857
rect 2079 19803 12932 19829
rect 1818 19775 2051 19803
tri 2051 19775 2079 19803 sw
tri 2079 19775 2107 19803 ne
rect 2107 19801 12932 19803
tri 12932 19801 12960 19829 nw
tri 12960 19801 12988 19829 se
rect 12988 19801 13124 19829
rect 2107 19775 12904 19801
rect 1818 19747 2079 19775
tri 2079 19747 2107 19775 sw
tri 2107 19747 2135 19775 ne
rect 2135 19773 12904 19775
tri 12904 19773 12932 19801 nw
tri 12932 19773 12960 19801 se
rect 12960 19773 13124 19801
rect 2135 19747 12876 19773
rect 1818 19719 2107 19747
tri 2107 19719 2135 19747 sw
tri 2135 19719 2163 19747 ne
rect 2163 19745 12876 19747
tri 12876 19745 12904 19773 nw
tri 12904 19745 12932 19773 se
rect 12932 19745 13124 19773
rect 2163 19719 12848 19745
rect 1818 19707 2135 19719
rect 1566 19691 2135 19707
tri 2135 19691 2163 19719 sw
tri 2163 19691 2191 19719 ne
rect 2191 19717 12848 19719
tri 12848 19717 12876 19745 nw
tri 12876 19717 12904 19745 se
rect 12904 19717 13124 19745
rect 2191 19691 12820 19717
tri 1566 19377 1880 19691 ne
rect 1880 19663 2163 19691
tri 2163 19663 2191 19691 sw
tri 2191 19663 2219 19691 ne
rect 2219 19689 12820 19691
tri 12820 19689 12848 19717 nw
tri 12848 19689 12876 19717 se
rect 12876 19689 13124 19717
rect 2219 19663 12792 19689
rect 1880 19635 2191 19663
tri 2191 19635 2219 19663 sw
tri 2219 19635 2247 19663 ne
rect 2247 19661 12792 19663
tri 12792 19661 12820 19689 nw
tri 12820 19661 12848 19689 se
rect 12848 19661 13124 19689
rect 2247 19635 12764 19661
rect 1880 19629 2219 19635
rect 1880 19393 1896 19629
rect 2132 19607 2219 19629
tri 2219 19607 2247 19635 sw
tri 2247 19607 2275 19635 ne
rect 2275 19633 12764 19635
tri 12764 19633 12792 19661 nw
tri 12792 19633 12820 19661 se
rect 12820 19649 13124 19661
rect 13360 19649 13383 19885
rect 12820 19640 13383 19649
tri 13383 19640 13706 19963 nw
rect 12820 19633 13066 19640
rect 2275 19607 12736 19633
rect 2132 19579 2247 19607
tri 2247 19579 2275 19607 sw
tri 2275 19579 2303 19607 ne
rect 2303 19605 12736 19607
tri 12736 19605 12764 19633 nw
tri 12764 19605 12792 19633 se
rect 12792 19605 13066 19633
rect 2303 19579 12708 19605
rect 2132 19551 2275 19579
tri 2275 19551 2303 19579 sw
tri 2303 19551 2331 19579 ne
rect 2331 19577 12708 19579
tri 12708 19577 12736 19605 nw
tri 12736 19577 12764 19605 se
rect 12764 19577 13066 19605
rect 2331 19551 12680 19577
rect 2132 19523 2303 19551
tri 2303 19523 2331 19551 sw
tri 2331 19523 2359 19551 ne
rect 2359 19549 12680 19551
tri 12680 19549 12708 19577 nw
tri 12708 19549 12736 19577 se
rect 12736 19575 13066 19577
rect 12736 19549 12814 19575
rect 2359 19523 12652 19549
rect 2132 19495 2331 19523
tri 2331 19495 2359 19523 sw
tri 2359 19495 2387 19523 ne
rect 2387 19521 12652 19523
tri 12652 19521 12680 19549 nw
tri 12680 19521 12708 19549 se
rect 12708 19521 12814 19549
rect 2387 19495 12624 19521
rect 2132 19467 2359 19495
tri 2359 19467 2387 19495 sw
tri 2387 19467 2415 19495 ne
rect 2415 19493 12624 19495
tri 12624 19493 12652 19521 nw
tri 12652 19493 12680 19521 se
rect 12680 19493 12814 19521
rect 2415 19467 12596 19493
rect 2132 19439 2387 19467
tri 2387 19439 2415 19467 sw
tri 2415 19439 2443 19467 ne
rect 2443 19465 12596 19467
tri 12596 19465 12624 19493 nw
tri 12624 19465 12652 19493 se
rect 12652 19465 12814 19493
rect 2443 19439 12568 19465
rect 2132 19411 2415 19439
tri 2415 19411 2443 19439 sw
tri 2443 19411 2471 19439 ne
rect 2471 19437 12568 19439
tri 12568 19437 12596 19465 nw
tri 12596 19437 12624 19465 se
rect 12624 19437 12814 19465
rect 2471 19411 12540 19437
rect 2132 19393 2443 19411
rect 1880 19383 2443 19393
tri 2443 19383 2471 19411 sw
tri 2471 19383 2499 19411 ne
rect 2499 19409 12540 19411
tri 12540 19409 12568 19437 nw
tri 12568 19409 12596 19437 se
rect 12596 19409 12814 19437
rect 2499 19383 12512 19409
rect 1880 19377 2471 19383
tri 1880 19015 2242 19377 ne
rect 2242 19355 2471 19377
tri 2471 19355 2499 19383 sw
tri 2499 19355 2527 19383 ne
rect 2527 19381 12512 19383
tri 12512 19381 12540 19409 nw
tri 12540 19381 12568 19409 se
rect 12568 19381 12814 19409
rect 2527 19355 12486 19381
tri 12486 19355 12512 19381 nw
tri 12514 19355 12540 19381 se
rect 12540 19355 12814 19381
rect 2242 19335 2499 19355
tri 2499 19335 2519 19355 sw
tri 12494 19335 12514 19355 se
rect 12514 19339 12814 19355
rect 13050 19339 13066 19575
rect 12514 19335 13066 19339
rect 2242 19323 13066 19335
tri 13066 19323 13383 19640 nw
rect 2242 19274 12734 19323
rect 2242 19038 2255 19274
rect 2491 19268 12734 19274
rect 2491 19251 12495 19268
rect 2491 19038 2575 19251
rect 2242 19015 2575 19038
rect 2811 19015 2895 19251
rect 3131 19015 3215 19251
rect 3451 19015 3535 19251
rect 3771 19015 3855 19251
rect 4091 19015 4175 19251
rect 4411 19015 4495 19251
rect 4731 19015 4815 19251
rect 5051 19015 5135 19251
rect 5371 19015 5455 19251
rect 5691 19015 5775 19251
rect 6011 19015 6095 19251
rect 6331 19015 6415 19251
rect 6651 19015 6735 19251
rect 6971 19015 7055 19251
rect 7291 19015 7375 19251
rect 7611 19015 7695 19251
rect 7931 19015 8015 19251
rect 8251 19015 8335 19251
rect 8571 19015 8655 19251
rect 8891 19015 8975 19251
rect 9211 19015 9295 19251
rect 9531 19015 9615 19251
rect 9851 19015 9935 19251
rect 10171 19015 10255 19251
rect 10491 19015 10575 19251
rect 10811 19015 10895 19251
rect 11131 19015 11215 19251
rect 11451 19015 11535 19251
rect 11771 19015 11855 19251
rect 12091 19015 12175 19251
rect 12411 19032 12495 19251
rect 12731 19032 12734 19268
rect 12411 19015 12734 19032
tri 2242 18991 2266 19015 ne
rect 2266 18991 12734 19015
tri 12734 18991 13066 19323 nw
<< rm5 >>
tri 2405 33663 2425 33683 se
rect 2425 33663 12578 33683
tri 12578 33663 12598 33683 sw
tri 2390 33648 2405 33663 se
tri 2362 33620 2390 33648 se
rect 2390 33635 2405 33648
tri 2405 33635 2433 33663 nw
tri 12570 33635 12598 33663 ne
tri 12598 33635 12626 33663 sw
tri 2390 33620 2405 33635 nw
tri 2334 33592 2362 33620 se
tri 2362 33592 2390 33620 nw
tri 12598 33607 12626 33635 ne
tri 12626 33607 12654 33635 sw
tri 2306 33564 2334 33592 se
tri 2334 33564 2362 33592 nw
tri 12626 33579 12654 33607 ne
tri 12654 33579 12682 33607 sw
tri 2278 33536 2306 33564 se
tri 2306 33536 2334 33564 nw
tri 12654 33551 12682 33579 ne
tri 12682 33551 12710 33579 sw
tri 2250 33508 2278 33536 se
tri 2278 33508 2306 33536 nw
tri 12682 33523 12710 33551 ne
tri 12710 33523 12738 33551 sw
tri 2222 33480 2250 33508 se
tri 2250 33480 2278 33508 nw
tri 12710 33495 12738 33523 ne
tri 12738 33495 12766 33523 sw
tri 2194 33452 2222 33480 se
tri 2222 33452 2250 33480 nw
tri 12738 33467 12766 33495 ne
tri 12766 33467 12794 33495 sw
tri 2166 33424 2194 33452 se
tri 2194 33424 2222 33452 nw
tri 12766 33439 12794 33467 ne
tri 12794 33439 12822 33467 sw
tri 2138 33396 2166 33424 se
tri 2166 33396 2194 33424 nw
tri 12794 33411 12822 33439 ne
tri 12822 33411 12850 33439 sw
tri 2110 33368 2138 33396 se
tri 2138 33368 2166 33396 nw
tri 12822 33383 12850 33411 ne
tri 12850 33383 12878 33411 sw
tri 2082 33340 2110 33368 se
tri 2110 33340 2138 33368 nw
tri 12850 33355 12878 33383 ne
tri 12878 33355 12906 33383 sw
tri 2054 33312 2082 33340 se
tri 2082 33312 2110 33340 nw
tri 12878 33327 12906 33355 ne
tri 12906 33327 12934 33355 sw
tri 2026 33284 2054 33312 se
tri 2054 33284 2082 33312 nw
tri 12906 33299 12934 33327 ne
tri 12934 33299 12962 33327 sw
tri 1998 33256 2026 33284 se
tri 2026 33256 2054 33284 nw
tri 12934 33271 12962 33299 ne
tri 12962 33271 12990 33299 sw
tri 1970 33228 1998 33256 se
tri 1998 33228 2026 33256 nw
tri 12962 33243 12990 33271 ne
tri 12990 33243 13018 33271 sw
tri 1942 33200 1970 33228 se
tri 1970 33200 1998 33228 nw
tri 12990 33215 13018 33243 ne
tri 13018 33215 13046 33243 sw
tri 1914 33172 1942 33200 se
tri 1942 33172 1970 33200 nw
tri 13018 33187 13046 33215 ne
tri 13046 33187 13074 33215 sw
tri 1886 33144 1914 33172 se
tri 1914 33144 1942 33172 nw
tri 13046 33159 13074 33187 ne
tri 13074 33159 13102 33187 sw
tri 1858 33116 1886 33144 se
tri 1886 33116 1914 33144 nw
tri 13074 33131 13102 33159 ne
tri 13102 33131 13130 33159 sw
tri 1830 33088 1858 33116 se
tri 1858 33088 1886 33116 nw
tri 13102 33103 13130 33131 ne
tri 13130 33103 13158 33131 sw
tri 1802 33060 1830 33088 se
tri 1830 33060 1858 33088 nw
tri 13130 33075 13158 33103 ne
tri 13158 33075 13186 33103 sw
tri 1774 33032 1802 33060 se
tri 1802 33032 1830 33060 nw
tri 13158 33047 13186 33075 ne
tri 13186 33047 13214 33075 sw
tri 1746 33004 1774 33032 se
tri 1774 33004 1802 33032 nw
tri 13186 33019 13214 33047 ne
tri 13214 33019 13242 33047 sw
tri 1718 32976 1746 33004 se
tri 1746 32976 1774 33004 nw
tri 13214 32991 13242 33019 ne
tri 13242 32991 13270 33019 sw
tri 1690 32948 1718 32976 se
tri 1718 32948 1746 32976 nw
tri 13242 32963 13270 32991 ne
tri 13270 32963 13298 32991 sw
tri 1662 32920 1690 32948 se
tri 1690 32920 1718 32948 nw
tri 13270 32935 13298 32963 ne
tri 13298 32935 13326 32963 sw
tri 1634 32892 1662 32920 se
tri 1662 32892 1690 32920 nw
tri 13298 32907 13326 32935 ne
tri 13326 32907 13354 32935 sw
tri 1606 32864 1634 32892 se
tri 1634 32864 1662 32892 nw
tri 13326 32879 13354 32907 ne
tri 13354 32879 13382 32907 sw
tri 1578 32836 1606 32864 se
tri 1606 32836 1634 32864 nw
tri 13354 32851 13382 32879 ne
tri 13382 32851 13410 32879 sw
tri 1550 32808 1578 32836 se
tri 1578 32808 1606 32836 nw
tri 13382 32823 13410 32851 ne
tri 13410 32823 13438 32851 sw
tri 1522 32780 1550 32808 se
tri 1550 32780 1578 32808 nw
tri 13410 32795 13438 32823 ne
tri 13438 32795 13466 32823 sw
tri 1494 32752 1522 32780 se
tri 1522 32752 1550 32780 nw
tri 13438 32767 13466 32795 ne
tri 13466 32767 13494 32795 sw
tri 1466 32724 1494 32752 se
tri 1494 32724 1522 32752 nw
tri 13466 32739 13494 32767 ne
tri 13494 32739 13522 32767 sw
tri 1438 32696 1466 32724 se
tri 1466 32696 1494 32724 nw
tri 13494 32711 13522 32739 ne
tri 13522 32711 13550 32739 sw
tri 1410 32668 1438 32696 se
tri 1438 32668 1466 32696 nw
tri 13522 32683 13550 32711 ne
tri 13550 32683 13578 32711 sw
tri 1382 32640 1410 32668 se
tri 1410 32640 1438 32668 nw
tri 13550 32655 13578 32683 ne
tri 13578 32655 13606 32683 sw
tri 1354 32612 1382 32640 se
tri 1382 32612 1410 32640 nw
tri 13578 32629 13604 32655 ne
rect 13604 32637 13606 32655
tri 13606 32637 13624 32655 sw
tri 1334 32592 1354 32612 se
rect 1334 20520 1354 32592
tri 1354 32584 1382 32612 nw
tri 1334 20500 1354 20520 ne
tri 1354 20500 1382 20528 sw
tri 1354 20475 1379 20500 ne
rect 1379 20475 1382 20500
tri 1382 20475 1407 20500 sw
tri 1379 20447 1407 20475 ne
tri 1407 20447 1435 20475 sw
tri 1407 20419 1435 20447 ne
tri 1435 20419 1463 20447 sw
tri 13576 20445 13604 20473 se
rect 13604 20465 13624 32637
tri 13604 20445 13624 20465 nw
tri 1435 20391 1463 20419 ne
tri 1463 20391 1491 20419 sw
tri 13548 20417 13576 20445 se
tri 13576 20417 13604 20445 nw
tri 1463 20363 1491 20391 ne
tri 1491 20363 1519 20391 sw
tri 13520 20389 13548 20417 se
tri 13548 20389 13576 20417 nw
tri 1491 20335 1519 20363 ne
tri 1519 20335 1547 20363 sw
tri 13492 20361 13520 20389 se
tri 13520 20361 13548 20389 nw
tri 1519 20307 1547 20335 ne
tri 1547 20307 1575 20335 sw
tri 13464 20333 13492 20361 se
tri 13492 20333 13520 20361 nw
tri 1547 20279 1575 20307 ne
tri 1575 20279 1603 20307 sw
tri 13436 20305 13464 20333 se
tri 13464 20305 13492 20333 nw
tri 1575 20251 1603 20279 ne
tri 1603 20251 1631 20279 sw
tri 13408 20277 13436 20305 se
tri 13436 20277 13464 20305 nw
tri 1603 20223 1631 20251 ne
tri 1631 20223 1659 20251 sw
tri 13380 20249 13408 20277 se
tri 13408 20249 13436 20277 nw
tri 1631 20195 1659 20223 ne
tri 1659 20195 1687 20223 sw
tri 13352 20221 13380 20249 se
tri 13380 20221 13408 20249 nw
tri 1659 20167 1687 20195 ne
tri 1687 20167 1715 20195 sw
tri 13324 20193 13352 20221 se
tri 13352 20193 13380 20221 nw
tri 1687 20139 1715 20167 ne
tri 1715 20139 1743 20167 sw
tri 13296 20165 13324 20193 se
tri 13324 20165 13352 20193 nw
tri 1715 20111 1743 20139 ne
tri 1743 20111 1771 20139 sw
tri 13268 20137 13296 20165 se
tri 13296 20137 13324 20165 nw
tri 1743 20083 1771 20111 ne
tri 1771 20083 1799 20111 sw
tri 13240 20109 13268 20137 se
tri 13268 20109 13296 20137 nw
tri 1771 20055 1799 20083 ne
tri 1799 20055 1827 20083 sw
tri 13212 20081 13240 20109 se
tri 13240 20081 13268 20109 nw
tri 1799 20027 1827 20055 ne
tri 1827 20027 1855 20055 sw
tri 13184 20053 13212 20081 se
tri 13212 20053 13240 20081 nw
tri 1827 19999 1855 20027 ne
tri 1855 19999 1883 20027 sw
tri 13156 20025 13184 20053 se
tri 13184 20025 13212 20053 nw
tri 1855 19971 1883 19999 ne
tri 1883 19971 1911 19999 sw
tri 13128 19997 13156 20025 se
tri 13156 19997 13184 20025 nw
tri 1883 19943 1911 19971 ne
tri 1911 19943 1939 19971 sw
tri 13100 19969 13128 19997 se
tri 13128 19969 13156 19997 nw
tri 1911 19915 1939 19943 ne
tri 1939 19915 1967 19943 sw
tri 13072 19941 13100 19969 se
tri 13100 19941 13128 19969 nw
tri 1939 19887 1967 19915 ne
tri 1967 19887 1995 19915 sw
tri 13044 19913 13072 19941 se
tri 13072 19913 13100 19941 nw
tri 1967 19859 1995 19887 ne
tri 1995 19859 2023 19887 sw
tri 13016 19885 13044 19913 se
tri 13044 19885 13072 19913 nw
tri 1995 19831 2023 19859 ne
tri 2023 19831 2051 19859 sw
tri 12988 19857 13016 19885 se
tri 13016 19857 13044 19885 nw
tri 2023 19803 2051 19831 ne
tri 2051 19803 2079 19831 sw
tri 12960 19829 12988 19857 se
tri 12988 19829 13016 19857 nw
tri 2051 19775 2079 19803 ne
tri 2079 19775 2107 19803 sw
tri 12932 19801 12960 19829 se
tri 12960 19801 12988 19829 nw
tri 2079 19747 2107 19775 ne
tri 2107 19747 2135 19775 sw
tri 12904 19773 12932 19801 se
tri 12932 19773 12960 19801 nw
tri 2107 19719 2135 19747 ne
tri 2135 19719 2163 19747 sw
tri 12876 19745 12904 19773 se
tri 12904 19745 12932 19773 nw
tri 2135 19691 2163 19719 ne
tri 2163 19691 2191 19719 sw
tri 12848 19717 12876 19745 se
tri 12876 19717 12904 19745 nw
tri 2163 19663 2191 19691 ne
tri 2191 19663 2219 19691 sw
tri 12820 19689 12848 19717 se
tri 12848 19689 12876 19717 nw
tri 2191 19635 2219 19663 ne
tri 2219 19635 2247 19663 sw
tri 12792 19661 12820 19689 se
tri 12820 19661 12848 19689 nw
tri 2219 19607 2247 19635 ne
tri 2247 19607 2275 19635 sw
tri 12764 19633 12792 19661 se
tri 12792 19633 12820 19661 nw
tri 2247 19579 2275 19607 ne
tri 2275 19579 2303 19607 sw
tri 12736 19605 12764 19633 se
tri 12764 19605 12792 19633 nw
tri 2275 19551 2303 19579 ne
tri 2303 19551 2331 19579 sw
tri 12708 19577 12736 19605 se
tri 12736 19577 12764 19605 nw
tri 2303 19523 2331 19551 ne
tri 2331 19523 2359 19551 sw
tri 12680 19549 12708 19577 se
tri 12708 19549 12736 19577 nw
tri 2331 19495 2359 19523 ne
tri 2359 19495 2387 19523 sw
tri 12652 19521 12680 19549 se
tri 12680 19521 12708 19549 nw
tri 2359 19467 2387 19495 ne
tri 2387 19467 2415 19495 sw
tri 12624 19493 12652 19521 se
tri 12652 19493 12680 19521 nw
tri 2387 19439 2415 19467 ne
tri 2415 19439 2443 19467 sw
tri 12596 19465 12624 19493 se
tri 12624 19465 12652 19493 nw
tri 2415 19411 2443 19439 ne
tri 2443 19411 2471 19439 sw
tri 12568 19437 12596 19465 se
tri 12596 19437 12624 19465 nw
tri 2443 19383 2471 19411 ne
tri 2471 19383 2499 19411 sw
tri 12540 19409 12568 19437 se
tri 12568 19409 12596 19437 nw
tri 2471 19355 2499 19383 ne
tri 2499 19355 2527 19383 sw
tri 12512 19381 12540 19409 se
tri 12540 19381 12568 19409 nw
tri 12486 19355 12512 19381 se
rect 12512 19355 12514 19381
tri 12514 19355 12540 19381 nw
tri 2499 19335 2519 19355 ne
rect 2519 19335 12494 19355
tri 12494 19335 12514 19355 nw
<< glass >>
tri 1500 32541 2490 33531 se
rect 2490 32541 12510 33531
tri 12510 32541 13500 33531 sw
rect 1500 20521 13500 32541
tri 1500 19531 2490 20521 ne
rect 2490 19531 12510 20521
tri 12510 19531 13500 20521 nw
use sky130_fd_pr__padplhp__example_559591418080  sky130_fd_pr__padplhp__example_559591418080_0
timestamp 1685007810
transform 1 0 1500 0 1 19531
box -478 -478 1 1
<< properties >>
string GDS_END 11194754
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11194490
<< end >>
