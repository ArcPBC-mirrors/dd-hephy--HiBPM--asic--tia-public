magic
tech sky130A
magscale 1 2
timestamp 1683564698
<< error_p >>
rect -6070 2745 -4010 2772
rect -3550 2745 -1490 2772
rect -1030 2745 1030 2772
rect 1490 2745 3550 2772
rect 4010 2745 6070 2772
rect -6070 1536 -4010 1563
rect -3550 1536 -1490 1563
rect -1030 1536 1030 1563
rect 1490 1536 3550 1563
rect 4010 1536 6070 1563
rect -6070 1309 -4010 1336
rect -3550 1309 -1490 1336
rect -1030 1309 1030 1336
rect 1490 1309 3550 1336
rect 4010 1309 6070 1336
rect -6070 100 -4010 127
rect -3550 100 -1490 127
rect -1030 100 1030 127
rect 1490 100 3550 127
rect 4010 100 6070 127
rect -6070 -127 -4010 -100
rect -3550 -127 -1490 -100
rect -1030 -127 1030 -100
rect 1490 -127 3550 -100
rect 4010 -127 6070 -100
rect -6070 -1336 -4010 -1309
rect -3550 -1336 -1490 -1309
rect -1030 -1336 1030 -1309
rect 1490 -1336 3550 -1309
rect 4010 -1336 6070 -1309
rect -6070 -1563 -4010 -1536
rect -3550 -1563 -1490 -1536
rect -1030 -1563 1030 -1536
rect 1490 -1563 3550 -1536
rect 4010 -1563 6070 -1536
rect -6070 -2772 -4010 -2745
rect -3550 -2772 -1490 -2745
rect -1030 -2772 1030 -2745
rect 1490 -2772 3550 -2745
rect 4010 -2772 6070 -2745
<< nwell >>
rect -6173 1563 -3907 2745
rect -3653 1563 -1387 2745
rect -1133 1563 1133 2745
rect 1387 1563 3653 2745
rect 3907 1563 6173 2745
rect -6173 127 -3907 1309
rect -3653 127 -1387 1309
rect -1133 127 1133 1309
rect 1387 127 3653 1309
rect 3907 127 6173 1309
rect -6173 -1309 -3907 -127
rect -3653 -1309 -1387 -127
rect -1133 -1309 1133 -127
rect 1387 -1309 3653 -127
rect 3907 -1309 6173 -127
rect -6173 -2745 -3907 -1563
rect -3653 -2745 -1387 -1563
rect -1133 -2745 1133 -1563
rect 1387 -2745 3653 -1563
rect 3907 -2745 6173 -1563
<< pwell >>
rect -6283 2745 6283 2855
rect -6283 1563 -6173 2745
rect -3907 1563 -3653 2745
rect -1387 1563 -1133 2745
rect 1133 1563 1387 2745
rect 3653 1563 3907 2745
rect 6173 1563 6283 2745
rect -6283 1309 6283 1563
rect -6283 127 -6173 1309
rect -3907 127 -3653 1309
rect -1387 127 -1133 1309
rect 1133 127 1387 1309
rect 3653 127 3907 1309
rect 6173 127 6283 1309
rect -6283 -127 6283 127
rect -6283 -1309 -6173 -127
rect -3907 -1309 -3653 -127
rect -1387 -1309 -1133 -127
rect 1133 -1309 1387 -127
rect 3653 -1309 3907 -127
rect 6173 -1309 6283 -127
rect -6283 -1563 6283 -1309
rect -6283 -2745 -6173 -1563
rect -3907 -2745 -3653 -1563
rect -1387 -2745 -1133 -1563
rect 1133 -2745 1387 -1563
rect 3653 -2745 3907 -1563
rect 6173 -2745 6283 -1563
rect -6283 -2855 6283 -2745
<< varactor >>
rect -6040 1654 -4040 2654
rect -3520 1654 -1520 2654
rect -1000 1654 1000 2654
rect 1520 1654 3520 2654
rect 4040 1654 6040 2654
rect -6040 218 -4040 1218
rect -3520 218 -1520 1218
rect -1000 218 1000 1218
rect 1520 218 3520 1218
rect 4040 218 6040 1218
rect -6040 -1218 -4040 -218
rect -3520 -1218 -1520 -218
rect -1000 -1218 1000 -218
rect 1520 -1218 3520 -218
rect 4040 -1218 6040 -218
rect -6040 -2654 -4040 -1654
rect -3520 -2654 -1520 -1654
rect -1000 -2654 1000 -1654
rect 1520 -2654 3520 -1654
rect 4040 -2654 6040 -1654
<< psubdiff >>
rect -6247 2785 -6151 2819
rect 6151 2785 6247 2819
rect -6247 2723 -6213 2785
rect 6213 2723 6247 2785
rect -6247 -2785 -6213 -2723
rect 6213 -2785 6247 -2723
rect -6247 -2819 -6151 -2785
rect 6151 -2819 6247 -2785
<< nsubdiff >>
rect -6137 2630 -6040 2654
rect -6137 1678 -6125 2630
rect -6091 1678 -6040 2630
rect -6137 1654 -6040 1678
rect -4040 2630 -3943 2654
rect -4040 1678 -3989 2630
rect -3955 1678 -3943 2630
rect -4040 1654 -3943 1678
rect -3617 2630 -3520 2654
rect -3617 1678 -3605 2630
rect -3571 1678 -3520 2630
rect -3617 1654 -3520 1678
rect -1520 2630 -1423 2654
rect -1520 1678 -1469 2630
rect -1435 1678 -1423 2630
rect -1520 1654 -1423 1678
rect -1097 2630 -1000 2654
rect -1097 1678 -1085 2630
rect -1051 1678 -1000 2630
rect -1097 1654 -1000 1678
rect 1000 2630 1097 2654
rect 1000 1678 1051 2630
rect 1085 1678 1097 2630
rect 1000 1654 1097 1678
rect 1423 2630 1520 2654
rect 1423 1678 1435 2630
rect 1469 1678 1520 2630
rect 1423 1654 1520 1678
rect 3520 2630 3617 2654
rect 3520 1678 3571 2630
rect 3605 1678 3617 2630
rect 3520 1654 3617 1678
rect 3943 2630 4040 2654
rect 3943 1678 3955 2630
rect 3989 1678 4040 2630
rect 3943 1654 4040 1678
rect 6040 2630 6137 2654
rect 6040 1678 6091 2630
rect 6125 1678 6137 2630
rect 6040 1654 6137 1678
rect -6137 1194 -6040 1218
rect -6137 242 -6125 1194
rect -6091 242 -6040 1194
rect -6137 218 -6040 242
rect -4040 1194 -3943 1218
rect -4040 242 -3989 1194
rect -3955 242 -3943 1194
rect -4040 218 -3943 242
rect -3617 1194 -3520 1218
rect -3617 242 -3605 1194
rect -3571 242 -3520 1194
rect -3617 218 -3520 242
rect -1520 1194 -1423 1218
rect -1520 242 -1469 1194
rect -1435 242 -1423 1194
rect -1520 218 -1423 242
rect -1097 1194 -1000 1218
rect -1097 242 -1085 1194
rect -1051 242 -1000 1194
rect -1097 218 -1000 242
rect 1000 1194 1097 1218
rect 1000 242 1051 1194
rect 1085 242 1097 1194
rect 1000 218 1097 242
rect 1423 1194 1520 1218
rect 1423 242 1435 1194
rect 1469 242 1520 1194
rect 1423 218 1520 242
rect 3520 1194 3617 1218
rect 3520 242 3571 1194
rect 3605 242 3617 1194
rect 3520 218 3617 242
rect 3943 1194 4040 1218
rect 3943 242 3955 1194
rect 3989 242 4040 1194
rect 3943 218 4040 242
rect 6040 1194 6137 1218
rect 6040 242 6091 1194
rect 6125 242 6137 1194
rect 6040 218 6137 242
rect -6137 -242 -6040 -218
rect -6137 -1194 -6125 -242
rect -6091 -1194 -6040 -242
rect -6137 -1218 -6040 -1194
rect -4040 -242 -3943 -218
rect -4040 -1194 -3989 -242
rect -3955 -1194 -3943 -242
rect -4040 -1218 -3943 -1194
rect -3617 -242 -3520 -218
rect -3617 -1194 -3605 -242
rect -3571 -1194 -3520 -242
rect -3617 -1218 -3520 -1194
rect -1520 -242 -1423 -218
rect -1520 -1194 -1469 -242
rect -1435 -1194 -1423 -242
rect -1520 -1218 -1423 -1194
rect -1097 -242 -1000 -218
rect -1097 -1194 -1085 -242
rect -1051 -1194 -1000 -242
rect -1097 -1218 -1000 -1194
rect 1000 -242 1097 -218
rect 1000 -1194 1051 -242
rect 1085 -1194 1097 -242
rect 1000 -1218 1097 -1194
rect 1423 -242 1520 -218
rect 1423 -1194 1435 -242
rect 1469 -1194 1520 -242
rect 1423 -1218 1520 -1194
rect 3520 -242 3617 -218
rect 3520 -1194 3571 -242
rect 3605 -1194 3617 -242
rect 3520 -1218 3617 -1194
rect 3943 -242 4040 -218
rect 3943 -1194 3955 -242
rect 3989 -1194 4040 -242
rect 3943 -1218 4040 -1194
rect 6040 -242 6137 -218
rect 6040 -1194 6091 -242
rect 6125 -1194 6137 -242
rect 6040 -1218 6137 -1194
rect -6137 -1678 -6040 -1654
rect -6137 -2630 -6125 -1678
rect -6091 -2630 -6040 -1678
rect -6137 -2654 -6040 -2630
rect -4040 -1678 -3943 -1654
rect -4040 -2630 -3989 -1678
rect -3955 -2630 -3943 -1678
rect -4040 -2654 -3943 -2630
rect -3617 -1678 -3520 -1654
rect -3617 -2630 -3605 -1678
rect -3571 -2630 -3520 -1678
rect -3617 -2654 -3520 -2630
rect -1520 -1678 -1423 -1654
rect -1520 -2630 -1469 -1678
rect -1435 -2630 -1423 -1678
rect -1520 -2654 -1423 -2630
rect -1097 -1678 -1000 -1654
rect -1097 -2630 -1085 -1678
rect -1051 -2630 -1000 -1678
rect -1097 -2654 -1000 -2630
rect 1000 -1678 1097 -1654
rect 1000 -2630 1051 -1678
rect 1085 -2630 1097 -1678
rect 1000 -2654 1097 -2630
rect 1423 -1678 1520 -1654
rect 1423 -2630 1435 -1678
rect 1469 -2630 1520 -1678
rect 1423 -2654 1520 -2630
rect 3520 -1678 3617 -1654
rect 3520 -2630 3571 -1678
rect 3605 -2630 3617 -1678
rect 3520 -2654 3617 -2630
rect 3943 -1678 4040 -1654
rect 3943 -2630 3955 -1678
rect 3989 -2630 4040 -1678
rect 3943 -2654 4040 -2630
rect 6040 -1678 6137 -1654
rect 6040 -2630 6091 -1678
rect 6125 -2630 6137 -1678
rect 6040 -2654 6137 -2630
<< psubdiffcont >>
rect -6151 2785 6151 2819
rect -6247 -2723 -6213 2723
rect 6213 -2723 6247 2723
rect -6151 -2819 6151 -2785
<< nsubdiffcont >>
rect -6125 1678 -6091 2630
rect -3989 1678 -3955 2630
rect -3605 1678 -3571 2630
rect -1469 1678 -1435 2630
rect -1085 1678 -1051 2630
rect 1051 1678 1085 2630
rect 1435 1678 1469 2630
rect 3571 1678 3605 2630
rect 3955 1678 3989 2630
rect 6091 1678 6125 2630
rect -6125 242 -6091 1194
rect -3989 242 -3955 1194
rect -3605 242 -3571 1194
rect -1469 242 -1435 1194
rect -1085 242 -1051 1194
rect 1051 242 1085 1194
rect 1435 242 1469 1194
rect 3571 242 3605 1194
rect 3955 242 3989 1194
rect 6091 242 6125 1194
rect -6125 -1194 -6091 -242
rect -3989 -1194 -3955 -242
rect -3605 -1194 -3571 -242
rect -1469 -1194 -1435 -242
rect -1085 -1194 -1051 -242
rect 1051 -1194 1085 -242
rect 1435 -1194 1469 -242
rect 3571 -1194 3605 -242
rect 3955 -1194 3989 -242
rect 6091 -1194 6125 -242
rect -6125 -2630 -6091 -1678
rect -3989 -2630 -3955 -1678
rect -3605 -2630 -3571 -1678
rect -1469 -2630 -1435 -1678
rect -1085 -2630 -1051 -1678
rect 1051 -2630 1085 -1678
rect 1435 -2630 1469 -1678
rect 3571 -2630 3605 -1678
rect 3955 -2630 3989 -1678
rect 6091 -2630 6125 -1678
<< poly >>
rect -6040 2726 -4040 2742
rect -6040 2692 -6024 2726
rect -4056 2692 -4040 2726
rect -6040 2654 -4040 2692
rect -3520 2726 -1520 2742
rect -3520 2692 -3504 2726
rect -1536 2692 -1520 2726
rect -3520 2654 -1520 2692
rect -1000 2726 1000 2742
rect -1000 2692 -984 2726
rect 984 2692 1000 2726
rect -1000 2654 1000 2692
rect 1520 2726 3520 2742
rect 1520 2692 1536 2726
rect 3504 2692 3520 2726
rect 1520 2654 3520 2692
rect 4040 2726 6040 2742
rect 4040 2692 4056 2726
rect 6024 2692 6040 2726
rect 4040 2654 6040 2692
rect -6040 1616 -4040 1654
rect -6040 1582 -6024 1616
rect -4056 1582 -4040 1616
rect -6040 1566 -4040 1582
rect -3520 1616 -1520 1654
rect -3520 1582 -3504 1616
rect -1536 1582 -1520 1616
rect -3520 1566 -1520 1582
rect -1000 1616 1000 1654
rect -1000 1582 -984 1616
rect 984 1582 1000 1616
rect -1000 1566 1000 1582
rect 1520 1616 3520 1654
rect 1520 1582 1536 1616
rect 3504 1582 3520 1616
rect 1520 1566 3520 1582
rect 4040 1616 6040 1654
rect 4040 1582 4056 1616
rect 6024 1582 6040 1616
rect 4040 1566 6040 1582
rect -6040 1290 -4040 1306
rect -6040 1256 -6024 1290
rect -4056 1256 -4040 1290
rect -6040 1218 -4040 1256
rect -3520 1290 -1520 1306
rect -3520 1256 -3504 1290
rect -1536 1256 -1520 1290
rect -3520 1218 -1520 1256
rect -1000 1290 1000 1306
rect -1000 1256 -984 1290
rect 984 1256 1000 1290
rect -1000 1218 1000 1256
rect 1520 1290 3520 1306
rect 1520 1256 1536 1290
rect 3504 1256 3520 1290
rect 1520 1218 3520 1256
rect 4040 1290 6040 1306
rect 4040 1256 4056 1290
rect 6024 1256 6040 1290
rect 4040 1218 6040 1256
rect -6040 180 -4040 218
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -6040 130 -4040 146
rect -3520 180 -1520 218
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -3520 130 -1520 146
rect -1000 180 1000 218
rect -1000 146 -984 180
rect 984 146 1000 180
rect -1000 130 1000 146
rect 1520 180 3520 218
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 1520 130 3520 146
rect 4040 180 6040 218
rect 4040 146 4056 180
rect 6024 146 6040 180
rect 4040 130 6040 146
rect -6040 -146 -4040 -130
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -6040 -218 -4040 -180
rect -3520 -146 -1520 -130
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -3520 -218 -1520 -180
rect -1000 -146 1000 -130
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect -1000 -218 1000 -180
rect 1520 -146 3520 -130
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 1520 -218 3520 -180
rect 4040 -146 6040 -130
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect 4040 -218 6040 -180
rect -6040 -1256 -4040 -1218
rect -6040 -1290 -6024 -1256
rect -4056 -1290 -4040 -1256
rect -6040 -1306 -4040 -1290
rect -3520 -1256 -1520 -1218
rect -3520 -1290 -3504 -1256
rect -1536 -1290 -1520 -1256
rect -3520 -1306 -1520 -1290
rect -1000 -1256 1000 -1218
rect -1000 -1290 -984 -1256
rect 984 -1290 1000 -1256
rect -1000 -1306 1000 -1290
rect 1520 -1256 3520 -1218
rect 1520 -1290 1536 -1256
rect 3504 -1290 3520 -1256
rect 1520 -1306 3520 -1290
rect 4040 -1256 6040 -1218
rect 4040 -1290 4056 -1256
rect 6024 -1290 6040 -1256
rect 4040 -1306 6040 -1290
rect -6040 -1582 -4040 -1566
rect -6040 -1616 -6024 -1582
rect -4056 -1616 -4040 -1582
rect -6040 -1654 -4040 -1616
rect -3520 -1582 -1520 -1566
rect -3520 -1616 -3504 -1582
rect -1536 -1616 -1520 -1582
rect -3520 -1654 -1520 -1616
rect -1000 -1582 1000 -1566
rect -1000 -1616 -984 -1582
rect 984 -1616 1000 -1582
rect -1000 -1654 1000 -1616
rect 1520 -1582 3520 -1566
rect 1520 -1616 1536 -1582
rect 3504 -1616 3520 -1582
rect 1520 -1654 3520 -1616
rect 4040 -1582 6040 -1566
rect 4040 -1616 4056 -1582
rect 6024 -1616 6040 -1582
rect 4040 -1654 6040 -1616
rect -6040 -2692 -4040 -2654
rect -6040 -2726 -6024 -2692
rect -4056 -2726 -4040 -2692
rect -6040 -2742 -4040 -2726
rect -3520 -2692 -1520 -2654
rect -3520 -2726 -3504 -2692
rect -1536 -2726 -1520 -2692
rect -3520 -2742 -1520 -2726
rect -1000 -2692 1000 -2654
rect -1000 -2726 -984 -2692
rect 984 -2726 1000 -2692
rect -1000 -2742 1000 -2726
rect 1520 -2692 3520 -2654
rect 1520 -2726 1536 -2692
rect 3504 -2726 3520 -2692
rect 1520 -2742 3520 -2726
rect 4040 -2692 6040 -2654
rect 4040 -2726 4056 -2692
rect 6024 -2726 6040 -2692
rect 4040 -2742 6040 -2726
<< polycont >>
rect -6024 2692 -4056 2726
rect -3504 2692 -1536 2726
rect -984 2692 984 2726
rect 1536 2692 3504 2726
rect 4056 2692 6024 2726
rect -6024 1582 -4056 1616
rect -3504 1582 -1536 1616
rect -984 1582 984 1616
rect 1536 1582 3504 1616
rect 4056 1582 6024 1616
rect -6024 1256 -4056 1290
rect -3504 1256 -1536 1290
rect -984 1256 984 1290
rect 1536 1256 3504 1290
rect 4056 1256 6024 1290
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6024 -1290 -4056 -1256
rect -3504 -1290 -1536 -1256
rect -984 -1290 984 -1256
rect 1536 -1290 3504 -1256
rect 4056 -1290 6024 -1256
rect -6024 -1616 -4056 -1582
rect -3504 -1616 -1536 -1582
rect -984 -1616 984 -1582
rect 1536 -1616 3504 -1582
rect 4056 -1616 6024 -1582
rect -6024 -2726 -4056 -2692
rect -3504 -2726 -1536 -2692
rect -984 -2726 984 -2692
rect 1536 -2726 3504 -2692
rect 4056 -2726 6024 -2692
<< locali >>
rect -6247 2785 -6151 2819
rect 6151 2785 6247 2819
rect -6247 2723 -6213 2785
rect -6040 2692 -6024 2726
rect -4056 2692 -4040 2726
rect -3520 2692 -3504 2726
rect -1536 2692 -1520 2726
rect -1000 2692 -984 2726
rect 984 2692 1000 2726
rect 1520 2692 1536 2726
rect 3504 2692 3520 2726
rect 4040 2692 4056 2726
rect 6024 2692 6040 2726
rect 6213 2723 6247 2785
rect -6125 2630 -6091 2646
rect -6125 1662 -6091 1678
rect -3989 2630 -3955 2646
rect -3989 1662 -3955 1678
rect -3605 2630 -3571 2646
rect -3605 1662 -3571 1678
rect -1469 2630 -1435 2646
rect -1469 1662 -1435 1678
rect -1085 2630 -1051 2646
rect -1085 1662 -1051 1678
rect 1051 2630 1085 2646
rect 1051 1662 1085 1678
rect 1435 2630 1469 2646
rect 1435 1662 1469 1678
rect 3571 2630 3605 2646
rect 3571 1662 3605 1678
rect 3955 2630 3989 2646
rect 3955 1662 3989 1678
rect 6091 2630 6125 2646
rect 6091 1662 6125 1678
rect -6040 1582 -6024 1616
rect -4056 1582 -4040 1616
rect -3520 1582 -3504 1616
rect -1536 1582 -1520 1616
rect -1000 1582 -984 1616
rect 984 1582 1000 1616
rect 1520 1582 1536 1616
rect 3504 1582 3520 1616
rect 4040 1582 4056 1616
rect 6024 1582 6040 1616
rect -6040 1256 -6024 1290
rect -4056 1256 -4040 1290
rect -3520 1256 -3504 1290
rect -1536 1256 -1520 1290
rect -1000 1256 -984 1290
rect 984 1256 1000 1290
rect 1520 1256 1536 1290
rect 3504 1256 3520 1290
rect 4040 1256 4056 1290
rect 6024 1256 6040 1290
rect -6125 1194 -6091 1210
rect -6125 226 -6091 242
rect -3989 1194 -3955 1210
rect -3989 226 -3955 242
rect -3605 1194 -3571 1210
rect -3605 226 -3571 242
rect -1469 1194 -1435 1210
rect -1469 226 -1435 242
rect -1085 1194 -1051 1210
rect -1085 226 -1051 242
rect 1051 1194 1085 1210
rect 1051 226 1085 242
rect 1435 1194 1469 1210
rect 1435 226 1469 242
rect 3571 1194 3605 1210
rect 3571 226 3605 242
rect 3955 1194 3989 1210
rect 3955 226 3989 242
rect 6091 1194 6125 1210
rect 6091 226 6125 242
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -1000 146 -984 180
rect 984 146 1000 180
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 4040 146 4056 180
rect 6024 146 6040 180
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect -6125 -242 -6091 -226
rect -6125 -1210 -6091 -1194
rect -3989 -242 -3955 -226
rect -3989 -1210 -3955 -1194
rect -3605 -242 -3571 -226
rect -3605 -1210 -3571 -1194
rect -1469 -242 -1435 -226
rect -1469 -1210 -1435 -1194
rect -1085 -242 -1051 -226
rect -1085 -1210 -1051 -1194
rect 1051 -242 1085 -226
rect 1051 -1210 1085 -1194
rect 1435 -242 1469 -226
rect 1435 -1210 1469 -1194
rect 3571 -242 3605 -226
rect 3571 -1210 3605 -1194
rect 3955 -242 3989 -226
rect 3955 -1210 3989 -1194
rect 6091 -242 6125 -226
rect 6091 -1210 6125 -1194
rect -6040 -1290 -6024 -1256
rect -4056 -1290 -4040 -1256
rect -3520 -1290 -3504 -1256
rect -1536 -1290 -1520 -1256
rect -1000 -1290 -984 -1256
rect 984 -1290 1000 -1256
rect 1520 -1290 1536 -1256
rect 3504 -1290 3520 -1256
rect 4040 -1290 4056 -1256
rect 6024 -1290 6040 -1256
rect -6040 -1616 -6024 -1582
rect -4056 -1616 -4040 -1582
rect -3520 -1616 -3504 -1582
rect -1536 -1616 -1520 -1582
rect -1000 -1616 -984 -1582
rect 984 -1616 1000 -1582
rect 1520 -1616 1536 -1582
rect 3504 -1616 3520 -1582
rect 4040 -1616 4056 -1582
rect 6024 -1616 6040 -1582
rect -6125 -1678 -6091 -1662
rect -6125 -2646 -6091 -2630
rect -3989 -1678 -3955 -1662
rect -3989 -2646 -3955 -2630
rect -3605 -1678 -3571 -1662
rect -3605 -2646 -3571 -2630
rect -1469 -1678 -1435 -1662
rect -1469 -2646 -1435 -2630
rect -1085 -1678 -1051 -1662
rect -1085 -2646 -1051 -2630
rect 1051 -1678 1085 -1662
rect 1051 -2646 1085 -2630
rect 1435 -1678 1469 -1662
rect 1435 -2646 1469 -2630
rect 3571 -1678 3605 -1662
rect 3571 -2646 3605 -2630
rect 3955 -1678 3989 -1662
rect 3955 -2646 3989 -2630
rect 6091 -1678 6125 -1662
rect 6091 -2646 6125 -2630
rect -6247 -2785 -6213 -2723
rect -6040 -2726 -6024 -2692
rect -4056 -2726 -4040 -2692
rect -3520 -2726 -3504 -2692
rect -1536 -2726 -1520 -2692
rect -1000 -2726 -984 -2692
rect 984 -2726 1000 -2692
rect 1520 -2726 1536 -2692
rect 3504 -2726 3520 -2692
rect 4040 -2726 4056 -2692
rect 6024 -2726 6040 -2692
rect 6213 -2785 6247 -2723
rect -6247 -2819 -6151 -2785
rect 6151 -2819 6247 -2785
<< viali >>
rect -6024 2692 -4056 2726
rect -3504 2692 -1536 2726
rect -984 2692 984 2726
rect 1536 2692 3504 2726
rect 4056 2692 6024 2726
rect -6125 1678 -6091 2630
rect -3989 1678 -3955 2630
rect -3605 1678 -3571 2630
rect -1469 1678 -1435 2630
rect -1085 1678 -1051 2630
rect 1051 1678 1085 2630
rect 1435 1678 1469 2630
rect 3571 1678 3605 2630
rect 3955 1678 3989 2630
rect 6091 1678 6125 2630
rect -6024 1582 -4056 1616
rect -3504 1582 -1536 1616
rect -984 1582 984 1616
rect 1536 1582 3504 1616
rect 4056 1582 6024 1616
rect -6024 1256 -4056 1290
rect -3504 1256 -1536 1290
rect -984 1256 984 1290
rect 1536 1256 3504 1290
rect 4056 1256 6024 1290
rect -6125 242 -6091 1194
rect -3989 242 -3955 1194
rect -3605 242 -3571 1194
rect -1469 242 -1435 1194
rect -1085 242 -1051 1194
rect 1051 242 1085 1194
rect 1435 242 1469 1194
rect 3571 242 3605 1194
rect 3955 242 3989 1194
rect 6091 242 6125 1194
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6125 -1194 -6091 -242
rect -3989 -1194 -3955 -242
rect -3605 -1194 -3571 -242
rect -1469 -1194 -1435 -242
rect -1085 -1194 -1051 -242
rect 1051 -1194 1085 -242
rect 1435 -1194 1469 -242
rect 3571 -1194 3605 -242
rect 3955 -1194 3989 -242
rect 6091 -1194 6125 -242
rect -6024 -1290 -4056 -1256
rect -3504 -1290 -1536 -1256
rect -984 -1290 984 -1256
rect 1536 -1290 3504 -1256
rect 4056 -1290 6024 -1256
rect -6024 -1616 -4056 -1582
rect -3504 -1616 -1536 -1582
rect -984 -1616 984 -1582
rect 1536 -1616 3504 -1582
rect 4056 -1616 6024 -1582
rect -6125 -2630 -6091 -1678
rect -3989 -2630 -3955 -1678
rect -3605 -2630 -3571 -1678
rect -1469 -2630 -1435 -1678
rect -1085 -2630 -1051 -1678
rect 1051 -2630 1085 -1678
rect 1435 -2630 1469 -1678
rect 3571 -2630 3605 -1678
rect 3955 -2630 3989 -1678
rect 6091 -2630 6125 -1678
rect -6024 -2726 -4056 -2692
rect -3504 -2726 -1536 -2692
rect -984 -2726 984 -2692
rect 1536 -2726 3504 -2692
rect 4056 -2726 6024 -2692
<< metal1 >>
rect -6036 2726 -4044 2732
rect -6036 2692 -6024 2726
rect -4056 2692 -4044 2726
rect -6036 2686 -4044 2692
rect -3516 2726 -1524 2732
rect -3516 2692 -3504 2726
rect -1536 2692 -1524 2726
rect -3516 2686 -1524 2692
rect -996 2726 996 2732
rect -996 2692 -984 2726
rect 984 2692 996 2726
rect -996 2686 996 2692
rect 1524 2726 3516 2732
rect 1524 2692 1536 2726
rect 3504 2692 3516 2726
rect 1524 2686 3516 2692
rect 4044 2726 6036 2732
rect 4044 2692 4056 2726
rect 6024 2692 6036 2726
rect 4044 2686 6036 2692
rect -6131 2630 -6085 2642
rect -3995 2630 -3949 2642
rect -6131 1678 -6125 2630
rect -6091 1678 -3989 2630
rect -3955 1678 -3949 2630
rect -6131 1666 -6085 1678
rect -3995 1666 -3949 1678
rect -3611 2630 -3565 2642
rect -1475 2630 -1429 2642
rect -3611 1678 -3605 2630
rect -3571 1678 -1469 2630
rect -1435 1678 -1429 2630
rect -3611 1666 -3565 1678
rect -1475 1666 -1429 1678
rect -1091 2630 -1045 2642
rect 1045 2630 1091 2642
rect -1091 1678 -1085 2630
rect -1051 1678 1051 2630
rect 1085 1678 1091 2630
rect -1091 1666 -1045 1678
rect 1045 1666 1091 1678
rect 1429 2630 1475 2642
rect 3565 2630 3611 2642
rect 1429 1678 1435 2630
rect 1469 1678 3571 2630
rect 3605 1678 3611 2630
rect 1429 1666 1475 1678
rect 3565 1666 3611 1678
rect 3949 2630 3995 2642
rect 6085 2630 6131 2642
rect 3949 1678 3955 2630
rect 3989 1678 6091 2630
rect 6125 1678 6131 2630
rect 3949 1666 3995 1678
rect 6085 1666 6131 1678
rect -6036 1616 -4044 1622
rect -6036 1582 -6024 1616
rect -4056 1582 -4044 1616
rect -6036 1576 -4044 1582
rect -3516 1616 -1524 1622
rect -3516 1582 -3504 1616
rect -1536 1582 -1524 1616
rect -3516 1576 -1524 1582
rect -996 1616 996 1622
rect -996 1582 -984 1616
rect 984 1582 996 1616
rect -996 1576 996 1582
rect 1524 1616 3516 1622
rect 1524 1582 1536 1616
rect 3504 1582 3516 1616
rect 1524 1576 3516 1582
rect 4044 1616 6036 1622
rect 4044 1582 4056 1616
rect 6024 1582 6036 1616
rect 4044 1576 6036 1582
rect -6036 1290 -4044 1296
rect -6036 1256 -6024 1290
rect -4056 1256 -4044 1290
rect -6036 1250 -4044 1256
rect -3516 1290 -1524 1296
rect -3516 1256 -3504 1290
rect -1536 1256 -1524 1290
rect -3516 1250 -1524 1256
rect -996 1290 996 1296
rect -996 1256 -984 1290
rect 984 1256 996 1290
rect -996 1250 996 1256
rect 1524 1290 3516 1296
rect 1524 1256 1536 1290
rect 3504 1256 3516 1290
rect 1524 1250 3516 1256
rect 4044 1290 6036 1296
rect 4044 1256 4056 1290
rect 6024 1256 6036 1290
rect 4044 1250 6036 1256
rect -6131 1194 -6085 1206
rect -3995 1194 -3949 1206
rect -6131 242 -6125 1194
rect -6091 242 -3989 1194
rect -3955 242 -3949 1194
rect -6131 230 -6085 242
rect -3995 230 -3949 242
rect -3611 1194 -3565 1206
rect -1475 1194 -1429 1206
rect -3611 242 -3605 1194
rect -3571 242 -1469 1194
rect -1435 242 -1429 1194
rect -3611 230 -3565 242
rect -1475 230 -1429 242
rect -1091 1194 -1045 1206
rect 1045 1194 1091 1206
rect -1091 242 -1085 1194
rect -1051 242 1051 1194
rect 1085 242 1091 1194
rect -1091 230 -1045 242
rect 1045 230 1091 242
rect 1429 1194 1475 1206
rect 3565 1194 3611 1206
rect 1429 242 1435 1194
rect 1469 242 3571 1194
rect 3605 242 3611 1194
rect 1429 230 1475 242
rect 3565 230 3611 242
rect 3949 1194 3995 1206
rect 6085 1194 6131 1206
rect 3949 242 3955 1194
rect 3989 242 6091 1194
rect 6125 242 6131 1194
rect 3949 230 3995 242
rect 6085 230 6131 242
rect -6036 180 -4044 186
rect -6036 146 -6024 180
rect -4056 146 -4044 180
rect -6036 140 -4044 146
rect -3516 180 -1524 186
rect -3516 146 -3504 180
rect -1536 146 -1524 180
rect -3516 140 -1524 146
rect -996 180 996 186
rect -996 146 -984 180
rect 984 146 996 180
rect -996 140 996 146
rect 1524 180 3516 186
rect 1524 146 1536 180
rect 3504 146 3516 180
rect 1524 140 3516 146
rect 4044 180 6036 186
rect 4044 146 4056 180
rect 6024 146 6036 180
rect 4044 140 6036 146
rect -6036 -146 -4044 -140
rect -6036 -180 -6024 -146
rect -4056 -180 -4044 -146
rect -6036 -186 -4044 -180
rect -3516 -146 -1524 -140
rect -3516 -180 -3504 -146
rect -1536 -180 -1524 -146
rect -3516 -186 -1524 -180
rect -996 -146 996 -140
rect -996 -180 -984 -146
rect 984 -180 996 -146
rect -996 -186 996 -180
rect 1524 -146 3516 -140
rect 1524 -180 1536 -146
rect 3504 -180 3516 -146
rect 1524 -186 3516 -180
rect 4044 -146 6036 -140
rect 4044 -180 4056 -146
rect 6024 -180 6036 -146
rect 4044 -186 6036 -180
rect -6131 -242 -6085 -230
rect -3995 -242 -3949 -230
rect -6131 -1194 -6125 -242
rect -6091 -1194 -3989 -242
rect -3955 -1194 -3949 -242
rect -6131 -1206 -6085 -1194
rect -3995 -1206 -3949 -1194
rect -3611 -242 -3565 -230
rect -1475 -242 -1429 -230
rect -3611 -1194 -3605 -242
rect -3571 -1194 -1469 -242
rect -1435 -1194 -1429 -242
rect -3611 -1206 -3565 -1194
rect -1475 -1206 -1429 -1194
rect -1091 -242 -1045 -230
rect 1045 -242 1091 -230
rect -1091 -1194 -1085 -242
rect -1051 -1194 1051 -242
rect 1085 -1194 1091 -242
rect -1091 -1206 -1045 -1194
rect 1045 -1206 1091 -1194
rect 1429 -242 1475 -230
rect 3565 -242 3611 -230
rect 1429 -1194 1435 -242
rect 1469 -1194 3571 -242
rect 3605 -1194 3611 -242
rect 1429 -1206 1475 -1194
rect 3565 -1206 3611 -1194
rect 3949 -242 3995 -230
rect 6085 -242 6131 -230
rect 3949 -1194 3955 -242
rect 3989 -1194 6091 -242
rect 6125 -1194 6131 -242
rect 3949 -1206 3995 -1194
rect 6085 -1206 6131 -1194
rect -6036 -1256 -4044 -1250
rect -6036 -1290 -6024 -1256
rect -4056 -1290 -4044 -1256
rect -6036 -1296 -4044 -1290
rect -3516 -1256 -1524 -1250
rect -3516 -1290 -3504 -1256
rect -1536 -1290 -1524 -1256
rect -3516 -1296 -1524 -1290
rect -996 -1256 996 -1250
rect -996 -1290 -984 -1256
rect 984 -1290 996 -1256
rect -996 -1296 996 -1290
rect 1524 -1256 3516 -1250
rect 1524 -1290 1536 -1256
rect 3504 -1290 3516 -1256
rect 1524 -1296 3516 -1290
rect 4044 -1256 6036 -1250
rect 4044 -1290 4056 -1256
rect 6024 -1290 6036 -1256
rect 4044 -1296 6036 -1290
rect -6036 -1582 -4044 -1576
rect -6036 -1616 -6024 -1582
rect -4056 -1616 -4044 -1582
rect -6036 -1622 -4044 -1616
rect -3516 -1582 -1524 -1576
rect -3516 -1616 -3504 -1582
rect -1536 -1616 -1524 -1582
rect -3516 -1622 -1524 -1616
rect -996 -1582 996 -1576
rect -996 -1616 -984 -1582
rect 984 -1616 996 -1582
rect -996 -1622 996 -1616
rect 1524 -1582 3516 -1576
rect 1524 -1616 1536 -1582
rect 3504 -1616 3516 -1582
rect 1524 -1622 3516 -1616
rect 4044 -1582 6036 -1576
rect 4044 -1616 4056 -1582
rect 6024 -1616 6036 -1582
rect 4044 -1622 6036 -1616
rect -6131 -1678 -6085 -1666
rect -3995 -1678 -3949 -1666
rect -6131 -2630 -6125 -1678
rect -6091 -2630 -3989 -1678
rect -3955 -2630 -3949 -1678
rect -6131 -2642 -6085 -2630
rect -3995 -2642 -3949 -2630
rect -3611 -1678 -3565 -1666
rect -1475 -1678 -1429 -1666
rect -3611 -2630 -3605 -1678
rect -3571 -2630 -1469 -1678
rect -1435 -2630 -1429 -1678
rect -3611 -2642 -3565 -2630
rect -1475 -2642 -1429 -2630
rect -1091 -1678 -1045 -1666
rect 1045 -1678 1091 -1666
rect -1091 -2630 -1085 -1678
rect -1051 -2630 1051 -1678
rect 1085 -2630 1091 -1678
rect -1091 -2642 -1045 -2630
rect 1045 -2642 1091 -2630
rect 1429 -1678 1475 -1666
rect 3565 -1678 3611 -1666
rect 1429 -2630 1435 -1678
rect 1469 -2630 3571 -1678
rect 3605 -2630 3611 -1678
rect 1429 -2642 1475 -2630
rect 3565 -2642 3611 -2630
rect 3949 -1678 3995 -1666
rect 6085 -1678 6131 -1666
rect 3949 -2630 3955 -1678
rect 3989 -2630 6091 -1678
rect 6125 -2630 6131 -1678
rect 3949 -2642 3995 -2630
rect 6085 -2642 6131 -2630
rect -6036 -2692 -4044 -2686
rect -6036 -2726 -6024 -2692
rect -4056 -2726 -4044 -2692
rect -6036 -2732 -4044 -2726
rect -3516 -2692 -1524 -2686
rect -3516 -2726 -3504 -2692
rect -1536 -2726 -1524 -2692
rect -3516 -2732 -1524 -2726
rect -996 -2692 996 -2686
rect -996 -2726 -984 -2692
rect 984 -2726 996 -2692
rect -996 -2732 996 -2726
rect 1524 -2692 3516 -2686
rect 1524 -2726 1536 -2692
rect 3504 -2726 3516 -2692
rect 1524 -2732 3516 -2726
rect 4044 -2692 6036 -2686
rect 4044 -2726 4056 -2692
rect 6024 -2726 6036 -2692
rect 4044 -2732 6036 -2726
<< properties >>
string FIXED_BBOX -6230 -2802 6230 2802
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 10 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
