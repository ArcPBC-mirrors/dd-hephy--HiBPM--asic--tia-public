magic
tech sky130A
magscale 1 2
timestamp 1684252655
<< locali >>
rect 840 4100 1000 4220
rect -160 2220 0 2320
rect -160 1300 -80 2220
rect 860 2120 980 2220
rect -160 1100 -20 1300
rect 320 -240 460 -80
rect 260 -2920 460 -2800
<< viali >>
rect 840 4220 1000 4360
rect 260 -3020 460 -2920
<< metal1 >>
rect 828 4360 1012 4366
rect 120 4220 840 4360
rect 1000 4220 1012 4360
rect 120 3960 360 4220
rect 828 4214 1012 4220
rect 98 2344 108 2776
rect 468 2344 478 2776
rect 684 2080 780 3960
rect 814 2288 824 2372
rect 1012 2288 1022 2372
rect 672 2072 780 2080
rect 1060 2072 1156 3956
rect -32 1992 1192 2072
rect -32 1504 40 1992
rect 166 1768 176 1948
rect 228 1768 238 1948
rect 358 1768 368 1948
rect 420 1768 430 1948
rect 550 1768 560 1948
rect 612 1768 622 1948
rect 742 1768 752 1948
rect 804 1768 814 1948
rect 934 1768 944 1948
rect 996 1768 1006 1948
rect 70 1544 80 1724
rect 132 1544 142 1724
rect 262 1544 272 1724
rect 324 1544 334 1724
rect 454 1544 464 1724
rect 516 1544 526 1724
rect 646 1544 656 1724
rect 708 1544 718 1724
rect 838 1544 848 1724
rect 900 1544 910 1724
rect 1030 1544 1040 1724
rect 1092 1544 1102 1724
rect -32 1496 956 1504
rect -32 1396 52 1496
rect 640 1424 956 1496
rect 640 1396 700 1424
rect -32 1384 700 1396
rect -56 1124 1048 1260
rect -56 652 40 1124
rect 162 912 172 1092
rect 224 912 234 1092
rect 354 912 364 1092
rect 416 912 426 1092
rect 546 912 556 1092
rect 608 912 618 1092
rect 738 912 748 1092
rect 800 912 810 1092
rect 930 912 940 1092
rect 992 912 1002 1092
rect 70 688 80 868
rect 132 688 142 868
rect 258 688 268 868
rect 320 688 330 868
rect 450 688 460 868
rect 512 688 522 868
rect 642 688 652 868
rect 704 688 714 868
rect 834 688 844 868
rect 896 688 906 868
rect 1026 688 1036 868
rect 1088 688 1098 868
rect -56 504 956 652
rect -56 32 40 504
rect 166 292 176 472
rect 228 292 238 472
rect 358 292 368 472
rect 420 292 430 472
rect 550 292 560 472
rect 612 292 622 472
rect 742 292 752 472
rect 804 292 814 472
rect 934 292 944 472
rect 996 292 1006 472
rect 74 68 84 248
rect 136 68 146 248
rect 262 68 272 248
rect 324 68 334 248
rect 454 68 464 248
rect 516 68 526 248
rect 646 68 656 248
rect 708 68 718 248
rect 838 68 848 248
rect 900 68 910 248
rect 1030 68 1040 248
rect 1092 68 1102 248
rect -56 -96 1092 32
rect -56 -208 40 -96
rect -56 -364 1368 -208
rect -56 -828 40 -364
rect 330 -572 340 -392
rect 392 -572 402 -392
rect 846 -572 856 -392
rect 908 -572 918 -392
rect 1362 -572 1372 -392
rect 1424 -572 1434 -392
rect 70 -796 80 -616
rect 132 -796 142 -616
rect 586 -796 596 -616
rect 648 -796 658 -616
rect 1102 -796 1112 -616
rect 1164 -796 1174 -616
rect -56 -984 1368 -828
rect -56 -1444 40 -984
rect 330 -1192 340 -1012
rect 392 -1192 402 -1012
rect 846 -1192 856 -1012
rect 908 -1192 918 -1012
rect 1362 -1192 1372 -1012
rect 1424 -1192 1434 -1012
rect 70 -1416 80 -1236
rect 132 -1416 142 -1236
rect 586 -1416 596 -1236
rect 648 -1416 658 -1236
rect 1102 -1416 1112 -1236
rect 1164 -1416 1174 -1236
rect -56 -1600 1368 -1444
rect -56 -2064 40 -1600
rect 330 -1808 340 -1628
rect 392 -1808 402 -1628
rect 846 -1808 856 -1628
rect 908 -1808 918 -1628
rect 1362 -1808 1372 -1628
rect 1424 -1808 1434 -1628
rect 70 -2032 80 -1852
rect 132 -2032 142 -1852
rect 586 -2032 596 -1852
rect 648 -2032 658 -1852
rect 1102 -2032 1112 -1852
rect 1164 -2032 1174 -1852
rect -56 -2220 1368 -2064
rect -56 -2680 40 -2220
rect 330 -2428 340 -2248
rect 392 -2428 402 -2248
rect 846 -2428 856 -2248
rect 908 -2428 918 -2248
rect 1362 -2428 1372 -2248
rect 1424 -2428 1434 -2248
rect 70 -2652 80 -2472
rect 132 -2652 142 -2472
rect 586 -2652 596 -2472
rect 648 -2652 658 -2472
rect 1102 -2652 1112 -2472
rect 1164 -2652 1174 -2472
rect -56 -2836 1368 -2680
rect 248 -2920 472 -2914
rect 248 -3020 260 -2920
rect 460 -3020 472 -2920
rect 248 -3026 472 -3020
<< via1 >>
rect 108 2344 468 2776
rect 824 2288 1012 2372
rect 176 1768 228 1948
rect 368 1768 420 1948
rect 560 1768 612 1948
rect 752 1768 804 1948
rect 944 1768 996 1948
rect 80 1544 132 1724
rect 272 1544 324 1724
rect 464 1544 516 1724
rect 656 1544 708 1724
rect 848 1544 900 1724
rect 1040 1544 1092 1724
rect 52 1396 640 1496
rect 172 912 224 1092
rect 364 912 416 1092
rect 556 912 608 1092
rect 748 912 800 1092
rect 940 912 992 1092
rect 80 688 132 868
rect 268 688 320 868
rect 460 688 512 868
rect 652 688 704 868
rect 844 688 896 868
rect 1036 688 1088 868
rect 176 292 228 472
rect 368 292 420 472
rect 560 292 612 472
rect 752 292 804 472
rect 944 292 996 472
rect 84 68 136 248
rect 272 68 324 248
rect 464 68 516 248
rect 656 68 708 248
rect 848 68 900 248
rect 1040 68 1092 248
rect 340 -572 392 -392
rect 856 -572 908 -392
rect 1372 -572 1424 -392
rect 80 -796 132 -616
rect 596 -796 648 -616
rect 1112 -796 1164 -616
rect 340 -1192 392 -1012
rect 856 -1192 908 -1012
rect 1372 -1192 1424 -1012
rect 80 -1416 132 -1236
rect 596 -1416 648 -1236
rect 1112 -1416 1164 -1236
rect 340 -1808 392 -1628
rect 856 -1808 908 -1628
rect 1372 -1808 1424 -1628
rect 80 -2032 132 -1852
rect 596 -2032 648 -1852
rect 1112 -2032 1164 -1852
rect 340 -2428 392 -2248
rect 856 -2428 908 -2248
rect 1372 -2428 1424 -2248
rect 80 -2652 132 -2472
rect 596 -2652 648 -2472
rect 1112 -2652 1164 -2472
rect 260 -3020 460 -2920
<< metal2 >>
rect 108 2776 468 2786
rect 468 2344 480 2776
rect 108 2334 480 2344
rect 116 2080 480 2334
rect 824 2372 1012 2382
rect 824 2278 1012 2288
rect 116 1948 1188 2080
rect 116 1772 176 1948
rect 228 1772 368 1948
rect 176 1758 228 1768
rect 420 1772 560 1948
rect 368 1758 420 1768
rect 612 1772 752 1948
rect 560 1758 612 1768
rect 804 1772 944 1948
rect 752 1758 804 1768
rect 996 1772 1188 1948
rect 944 1758 996 1768
rect 80 1724 132 1734
rect 52 1708 80 1718
rect 272 1724 324 1734
rect 132 1708 272 1720
rect 464 1724 516 1734
rect 324 1708 464 1720
rect 656 1724 708 1734
rect 516 1708 656 1720
rect 640 1544 656 1708
rect 848 1724 900 1734
rect 708 1544 848 1720
rect 1040 1724 1092 1734
rect 900 1544 1040 1720
rect 640 1412 1092 1544
rect 52 1386 640 1396
rect 172 1162 992 1260
rect 64 1152 992 1162
rect 644 1092 992 1152
rect 644 920 748 1092
rect 64 912 172 920
rect 224 912 364 920
rect 416 912 556 920
rect 608 916 748 920
rect 608 912 644 916
rect 64 910 644 912
rect 800 916 940 1092
rect 172 902 224 910
rect 364 902 416 910
rect 556 902 608 910
rect 748 902 800 912
rect 940 902 992 912
rect 80 868 132 878
rect 268 868 320 878
rect 132 688 268 864
rect 460 868 512 878
rect 320 688 460 864
rect 652 868 704 878
rect 512 688 652 864
rect 844 868 896 878
rect 704 840 844 864
rect 1036 868 1088 878
rect 896 840 1036 864
rect 1088 850 1092 864
rect 1088 840 1408 850
rect 704 688 776 840
rect 80 612 776 688
rect 80 602 1408 612
rect 80 600 1092 602
rect 64 540 996 564
rect 644 472 996 540
rect 644 308 752 472
rect 64 298 176 308
rect 228 296 368 308
rect 176 282 228 292
rect 420 296 560 308
rect 368 282 420 292
rect 612 296 752 308
rect 560 282 612 292
rect 804 296 944 472
rect 752 282 804 292
rect 944 282 996 292
rect 84 252 136 258
rect 272 252 324 258
rect 464 252 516 258
rect 656 252 708 258
rect 848 254 900 258
rect 1040 254 1092 258
rect 780 252 1412 254
rect 84 248 1416 252
rect 136 68 272 248
rect 324 68 464 248
rect 516 68 656 248
rect 708 244 848 248
rect 900 244 1040 248
rect 1092 244 1416 248
rect 708 68 780 244
rect 84 16 780 68
rect 1412 16 1416 244
rect 84 4 1416 16
rect 776 -324 1408 -314
rect 340 -392 776 -324
rect 1408 -392 1424 -324
rect 392 -552 776 -392
rect 392 -568 856 -552
rect 340 -582 392 -572
rect 908 -568 1372 -552
rect 856 -582 908 -572
rect 1372 -582 1424 -572
rect 80 -616 132 -606
rect 596 -616 648 -606
rect 132 -628 596 -618
rect 1112 -616 1164 -606
rect 648 -620 668 -618
rect 648 -628 1112 -620
rect 668 -796 1112 -628
rect 80 -856 88 -796
rect 668 -856 1164 -796
rect 80 -864 1164 -856
rect 88 -866 668 -864
rect 776 -944 1408 -938
rect 340 -948 1424 -944
rect 340 -1012 776 -948
rect 1408 -1012 1424 -948
rect 392 -1176 776 -1012
rect 392 -1188 856 -1176
rect 340 -1202 392 -1192
rect 908 -1188 1372 -1176
rect 856 -1202 908 -1192
rect 1372 -1202 1424 -1192
rect 80 -1236 132 -1226
rect 596 -1236 648 -1226
rect 132 -1248 596 -1238
rect 1112 -1236 1164 -1226
rect 648 -1240 668 -1238
rect 648 -1248 1112 -1240
rect 668 -1416 1112 -1248
rect 80 -1476 88 -1416
rect 668 -1476 1164 -1416
rect 80 -1484 1164 -1476
rect 88 -1486 668 -1484
rect 776 -1560 1408 -1554
rect 340 -1564 1424 -1560
rect 340 -1628 776 -1564
rect 1408 -1628 1424 -1564
rect 392 -1792 776 -1628
rect 392 -1804 856 -1792
rect 340 -1818 392 -1808
rect 908 -1804 1372 -1792
rect 856 -1818 908 -1808
rect 1372 -1818 1424 -1808
rect 80 -1852 132 -1842
rect 596 -1852 648 -1842
rect 132 -1864 596 -1854
rect 1112 -1852 1164 -1842
rect 648 -1856 668 -1854
rect 648 -1864 1112 -1856
rect 668 -2032 1112 -1864
rect 80 -2092 88 -2032
rect 668 -2092 1164 -2032
rect 80 -2100 1164 -2092
rect 88 -2102 668 -2100
rect 780 -2160 1412 -2150
rect 340 -2248 780 -2180
rect 1412 -2248 1424 -2180
rect 392 -2388 780 -2248
rect 392 -2424 856 -2388
rect 340 -2438 392 -2428
rect 908 -2424 1372 -2388
rect 856 -2438 908 -2428
rect 1372 -2438 1424 -2428
rect 80 -2472 132 -2462
rect 596 -2472 648 -2462
rect 132 -2484 596 -2474
rect 1112 -2472 1164 -2462
rect 648 -2476 668 -2474
rect 648 -2484 1112 -2476
rect 668 -2652 1112 -2484
rect 80 -2712 88 -2652
rect 668 -2712 1164 -2652
rect 80 -2720 1164 -2712
rect 88 -2722 668 -2720
rect 260 -2920 460 -2910
rect 260 -3030 460 -3020
<< via2 >>
rect 824 2288 1012 2372
rect 52 1544 80 1708
rect 80 1544 132 1708
rect 132 1544 272 1708
rect 272 1544 324 1708
rect 324 1544 464 1708
rect 464 1544 516 1708
rect 516 1544 640 1708
rect 52 1496 640 1544
rect 52 1408 640 1496
rect 64 1092 644 1152
rect 64 920 172 1092
rect 172 920 224 1092
rect 224 920 364 1092
rect 364 920 416 1092
rect 416 920 556 1092
rect 556 920 608 1092
rect 608 920 644 1092
rect 776 688 844 840
rect 844 688 896 840
rect 896 688 1036 840
rect 1036 688 1088 840
rect 1088 688 1408 840
rect 776 612 1408 688
rect 64 472 644 540
rect 64 308 176 472
rect 176 308 228 472
rect 228 308 368 472
rect 368 308 420 472
rect 420 308 560 472
rect 560 308 612 472
rect 612 308 644 472
rect 780 68 848 244
rect 848 68 900 244
rect 900 68 1040 244
rect 1040 68 1092 244
rect 1092 68 1412 244
rect 780 16 1412 68
rect 776 -392 1408 -324
rect 776 -552 856 -392
rect 856 -552 908 -392
rect 908 -552 1372 -392
rect 1372 -552 1408 -392
rect 88 -796 132 -628
rect 132 -796 596 -628
rect 596 -796 648 -628
rect 648 -796 668 -628
rect 88 -856 668 -796
rect 776 -1012 1408 -948
rect 776 -1176 856 -1012
rect 856 -1176 908 -1012
rect 908 -1176 1372 -1012
rect 1372 -1176 1408 -1012
rect 88 -1416 132 -1248
rect 132 -1416 596 -1248
rect 596 -1416 648 -1248
rect 648 -1416 668 -1248
rect 88 -1476 668 -1416
rect 776 -1628 1408 -1564
rect 776 -1792 856 -1628
rect 856 -1792 908 -1628
rect 908 -1792 1372 -1628
rect 1372 -1792 1408 -1628
rect 88 -2032 132 -1864
rect 132 -2032 596 -1864
rect 596 -2032 648 -1864
rect 648 -2032 668 -1864
rect 88 -2092 668 -2032
rect 780 -2248 1412 -2160
rect 780 -2388 856 -2248
rect 856 -2388 908 -2248
rect 908 -2388 1372 -2248
rect 1372 -2388 1412 -2248
rect 88 -2652 132 -2484
rect 132 -2652 596 -2484
rect 596 -2652 648 -2484
rect 648 -2652 668 -2484
rect 88 -2712 668 -2652
rect 260 -3020 460 -2920
<< metal3 >>
rect 800 2372 1900 2460
rect 800 2288 824 2372
rect 1012 2288 1900 2372
rect 800 2240 1900 2288
rect 42 1708 650 1713
rect 42 1408 52 1708
rect 640 1408 650 1708
rect 42 1403 650 1408
rect 52 1157 640 1403
rect 52 1152 654 1157
rect 52 920 64 1152
rect 644 920 654 1152
rect 1640 1140 1900 2120
rect 52 915 654 920
rect 52 545 640 915
rect 764 840 1420 856
rect 764 612 776 840
rect 1408 612 1420 840
rect 52 540 654 545
rect 52 308 64 540
rect 644 308 654 540
rect 52 303 654 308
rect 52 300 640 303
rect 764 249 1420 612
rect 764 244 1422 249
rect 764 16 780 244
rect 1412 16 1422 244
rect 764 11 1422 16
rect 764 -324 1420 11
rect 764 -552 776 -324
rect 1408 -552 1420 -324
rect 80 -623 676 -620
rect 78 -628 678 -623
rect 78 -856 88 -628
rect 668 -856 678 -628
rect 78 -861 678 -856
rect 80 -1243 676 -861
rect 764 -948 1420 -552
rect 764 -1176 776 -948
rect 1408 -1176 1420 -948
rect 78 -1248 678 -1243
rect 78 -1476 88 -1248
rect 668 -1476 678 -1248
rect 78 -1481 678 -1476
rect 80 -1859 676 -1481
rect 764 -1564 1420 -1176
rect 764 -1792 776 -1564
rect 1408 -1792 1420 -1564
rect 78 -1864 678 -1859
rect 78 -2092 88 -1864
rect 668 -2092 678 -1864
rect 78 -2097 678 -2092
rect 80 -2479 676 -2097
rect 764 -2155 1420 -1792
rect 764 -2160 1422 -2155
rect 764 -2388 780 -2160
rect 1412 -2388 1422 -2160
rect 764 -2393 1422 -2388
rect 764 -2400 1420 -2393
rect 78 -2484 678 -2479
rect 78 -2712 88 -2484
rect 668 -2712 678 -2484
rect 78 -2717 678 -2712
rect 80 -2920 676 -2717
rect 80 -2976 260 -2920
rect 250 -3020 260 -2976
rect 460 -2976 676 -2920
rect 460 -3020 470 -2976
rect 250 -3025 470 -3020
<< metal4 >>
rect 1720 1080 1940 2120
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_0
timestamp 1684252655
transform 1 0 3826 0 1 4020
box -2186 -2040 2186 2040
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  sky130_fd_pr__cap_mim_m3_1_WXTTNJ_1
timestamp 1684252655
transform 1 0 3826 0 1 -820
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_lvt_9U3MKJ  sky130_fd_pr__nfet_01v8_lvt_9U3MKJ_1
timestamp 1683627527
transform -1 0 587 0 -1 579
box -647 -719 647 719
use sky130_fd_pr__nfet_01v8_lvt_67XT6R  sky130_fd_pr__nfet_01v8_lvt_67XT6R_1
timestamp 1683557511
transform 1 0 752 0 1 -1523
box -812 -1337 812 1337
use sky130_fd_pr__pfet_01v8_G3L97A  sky130_fd_pr__pfet_01v8_G3L97A_0
timestamp 1683713379
transform 0 -1 919 1 0 3160
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_VCB84W  sky130_fd_pr__pfet_01v8_VCB84W_0
timestamp 1683563853
transform 1 0 587 0 1 1747
box -647 -419 647 419
use sky130_fd_pr__res_xhigh_po_1p41_E28PWF  sky130_fd_pr__res_xhigh_po_1p41_E28PWF_0
timestamp 1683558843
transform 1 0 247 0 1 3178
box -307 -998 307 998
<< end >>
