magic
tech sky130A
magscale 1 2
timestamp 1683540360
<< metal3 >>
rect -2186 1012 2186 1040
rect -2186 -1012 2102 1012
rect 2166 -1012 2186 1012
rect -2186 -1040 2186 -1012
<< via3 >>
rect 2102 -1012 2166 1012
<< mimcap >>
rect -2146 960 1854 1000
rect -2146 -960 -2106 960
rect 1814 -960 1854 960
rect -2146 -1000 1854 -960
<< mimcapcontact >>
rect -2106 -960 1814 960
<< metal4 >>
rect 2086 1012 2182 1028
rect -2107 960 1815 961
rect -2107 -960 -2106 960
rect 1814 -960 1815 960
rect -2107 -961 1815 -960
rect 2086 -1012 2102 1012
rect 2166 -1012 2182 1012
rect 2086 -1028 2182 -1012
<< properties >>
string FIXED_BBOX -2186 -1040 1894 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20.0 l 10 val 411.4 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
