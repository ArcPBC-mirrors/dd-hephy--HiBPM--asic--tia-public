magic
tech sky130A
magscale 1 2
timestamp 1683557511
<< error_p >>
rect -461 1235 -403 1241
rect -269 1235 -211 1241
rect -77 1235 -19 1241
rect 115 1235 173 1241
rect 307 1235 365 1241
rect -461 1201 -449 1235
rect -269 1201 -257 1235
rect -77 1201 -65 1235
rect 115 1201 127 1235
rect 307 1201 319 1235
rect -461 1195 -403 1201
rect -269 1195 -211 1201
rect -77 1195 -19 1201
rect 115 1195 173 1201
rect 307 1195 365 1201
rect -365 707 -307 713
rect -173 707 -115 713
rect 19 707 77 713
rect 211 707 269 713
rect 403 707 461 713
rect -365 673 -353 707
rect -173 673 -161 707
rect 19 673 31 707
rect 211 673 223 707
rect 403 673 415 707
rect -365 667 -307 673
rect -173 667 -115 673
rect 19 667 77 673
rect 211 667 269 673
rect 403 667 461 673
rect -365 599 -307 605
rect -173 599 -115 605
rect 19 599 77 605
rect 211 599 269 605
rect 403 599 461 605
rect -365 565 -353 599
rect -173 565 -161 599
rect 19 565 31 599
rect 211 565 223 599
rect 403 565 415 599
rect -365 559 -307 565
rect -173 559 -115 565
rect 19 559 77 565
rect 211 559 269 565
rect 403 559 461 565
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect -365 -565 -307 -559
rect -173 -565 -115 -559
rect 19 -565 77 -559
rect 211 -565 269 -559
rect 403 -565 461 -559
rect -365 -599 -353 -565
rect -173 -599 -161 -565
rect 19 -599 31 -565
rect 211 -599 223 -565
rect 403 -599 415 -565
rect -365 -605 -307 -599
rect -173 -605 -115 -599
rect 19 -605 77 -599
rect 211 -605 269 -599
rect 403 -605 461 -599
rect -365 -673 -307 -667
rect -173 -673 -115 -667
rect 19 -673 77 -667
rect 211 -673 269 -667
rect 403 -673 461 -667
rect -365 -707 -353 -673
rect -173 -707 -161 -673
rect 19 -707 31 -673
rect 211 -707 223 -673
rect 403 -707 415 -673
rect -365 -713 -307 -707
rect -173 -713 -115 -707
rect 19 -713 77 -707
rect 211 -713 269 -707
rect 403 -713 461 -707
rect -461 -1201 -403 -1195
rect -269 -1201 -211 -1195
rect -77 -1201 -19 -1195
rect 115 -1201 173 -1195
rect 307 -1201 365 -1195
rect -461 -1235 -449 -1201
rect -269 -1235 -257 -1201
rect -77 -1235 -65 -1201
rect 115 -1235 127 -1201
rect 307 -1235 319 -1201
rect -461 -1241 -403 -1235
rect -269 -1241 -211 -1235
rect -77 -1241 -19 -1235
rect 115 -1241 173 -1235
rect 307 -1241 365 -1235
<< nwell >>
rect -647 -1373 647 1373
<< pmos >>
rect -447 754 -417 1154
rect -351 754 -321 1154
rect -255 754 -225 1154
rect -159 754 -129 1154
rect -63 754 -33 1154
rect 33 754 63 1154
rect 129 754 159 1154
rect 225 754 255 1154
rect 321 754 351 1154
rect 417 754 447 1154
rect -447 118 -417 518
rect -351 118 -321 518
rect -255 118 -225 518
rect -159 118 -129 518
rect -63 118 -33 518
rect 33 118 63 518
rect 129 118 159 518
rect 225 118 255 518
rect 321 118 351 518
rect 417 118 447 518
rect -447 -518 -417 -118
rect -351 -518 -321 -118
rect -255 -518 -225 -118
rect -159 -518 -129 -118
rect -63 -518 -33 -118
rect 33 -518 63 -118
rect 129 -518 159 -118
rect 225 -518 255 -118
rect 321 -518 351 -118
rect 417 -518 447 -118
rect -447 -1154 -417 -754
rect -351 -1154 -321 -754
rect -255 -1154 -225 -754
rect -159 -1154 -129 -754
rect -63 -1154 -33 -754
rect 33 -1154 63 -754
rect 129 -1154 159 -754
rect 225 -1154 255 -754
rect 321 -1154 351 -754
rect 417 -1154 447 -754
<< pdiff >>
rect -509 1142 -447 1154
rect -509 766 -497 1142
rect -463 766 -447 1142
rect -509 754 -447 766
rect -417 1142 -351 1154
rect -417 766 -401 1142
rect -367 766 -351 1142
rect -417 754 -351 766
rect -321 1142 -255 1154
rect -321 766 -305 1142
rect -271 766 -255 1142
rect -321 754 -255 766
rect -225 1142 -159 1154
rect -225 766 -209 1142
rect -175 766 -159 1142
rect -225 754 -159 766
rect -129 1142 -63 1154
rect -129 766 -113 1142
rect -79 766 -63 1142
rect -129 754 -63 766
rect -33 1142 33 1154
rect -33 766 -17 1142
rect 17 766 33 1142
rect -33 754 33 766
rect 63 1142 129 1154
rect 63 766 79 1142
rect 113 766 129 1142
rect 63 754 129 766
rect 159 1142 225 1154
rect 159 766 175 1142
rect 209 766 225 1142
rect 159 754 225 766
rect 255 1142 321 1154
rect 255 766 271 1142
rect 305 766 321 1142
rect 255 754 321 766
rect 351 1142 417 1154
rect 351 766 367 1142
rect 401 766 417 1142
rect 351 754 417 766
rect 447 1142 509 1154
rect 447 766 463 1142
rect 497 766 509 1142
rect 447 754 509 766
rect -509 506 -447 518
rect -509 130 -497 506
rect -463 130 -447 506
rect -509 118 -447 130
rect -417 506 -351 518
rect -417 130 -401 506
rect -367 130 -351 506
rect -417 118 -351 130
rect -321 506 -255 518
rect -321 130 -305 506
rect -271 130 -255 506
rect -321 118 -255 130
rect -225 506 -159 518
rect -225 130 -209 506
rect -175 130 -159 506
rect -225 118 -159 130
rect -129 506 -63 518
rect -129 130 -113 506
rect -79 130 -63 506
rect -129 118 -63 130
rect -33 506 33 518
rect -33 130 -17 506
rect 17 130 33 506
rect -33 118 33 130
rect 63 506 129 518
rect 63 130 79 506
rect 113 130 129 506
rect 63 118 129 130
rect 159 506 225 518
rect 159 130 175 506
rect 209 130 225 506
rect 159 118 225 130
rect 255 506 321 518
rect 255 130 271 506
rect 305 130 321 506
rect 255 118 321 130
rect 351 506 417 518
rect 351 130 367 506
rect 401 130 417 506
rect 351 118 417 130
rect 447 506 509 518
rect 447 130 463 506
rect 497 130 509 506
rect 447 118 509 130
rect -509 -130 -447 -118
rect -509 -506 -497 -130
rect -463 -506 -447 -130
rect -509 -518 -447 -506
rect -417 -130 -351 -118
rect -417 -506 -401 -130
rect -367 -506 -351 -130
rect -417 -518 -351 -506
rect -321 -130 -255 -118
rect -321 -506 -305 -130
rect -271 -506 -255 -130
rect -321 -518 -255 -506
rect -225 -130 -159 -118
rect -225 -506 -209 -130
rect -175 -506 -159 -130
rect -225 -518 -159 -506
rect -129 -130 -63 -118
rect -129 -506 -113 -130
rect -79 -506 -63 -130
rect -129 -518 -63 -506
rect -33 -130 33 -118
rect -33 -506 -17 -130
rect 17 -506 33 -130
rect -33 -518 33 -506
rect 63 -130 129 -118
rect 63 -506 79 -130
rect 113 -506 129 -130
rect 63 -518 129 -506
rect 159 -130 225 -118
rect 159 -506 175 -130
rect 209 -506 225 -130
rect 159 -518 225 -506
rect 255 -130 321 -118
rect 255 -506 271 -130
rect 305 -506 321 -130
rect 255 -518 321 -506
rect 351 -130 417 -118
rect 351 -506 367 -130
rect 401 -506 417 -130
rect 351 -518 417 -506
rect 447 -130 509 -118
rect 447 -506 463 -130
rect 497 -506 509 -130
rect 447 -518 509 -506
rect -509 -766 -447 -754
rect -509 -1142 -497 -766
rect -463 -1142 -447 -766
rect -509 -1154 -447 -1142
rect -417 -766 -351 -754
rect -417 -1142 -401 -766
rect -367 -1142 -351 -766
rect -417 -1154 -351 -1142
rect -321 -766 -255 -754
rect -321 -1142 -305 -766
rect -271 -1142 -255 -766
rect -321 -1154 -255 -1142
rect -225 -766 -159 -754
rect -225 -1142 -209 -766
rect -175 -1142 -159 -766
rect -225 -1154 -159 -1142
rect -129 -766 -63 -754
rect -129 -1142 -113 -766
rect -79 -1142 -63 -766
rect -129 -1154 -63 -1142
rect -33 -766 33 -754
rect -33 -1142 -17 -766
rect 17 -1142 33 -766
rect -33 -1154 33 -1142
rect 63 -766 129 -754
rect 63 -1142 79 -766
rect 113 -1142 129 -766
rect 63 -1154 129 -1142
rect 159 -766 225 -754
rect 159 -1142 175 -766
rect 209 -1142 225 -766
rect 159 -1154 225 -1142
rect 255 -766 321 -754
rect 255 -1142 271 -766
rect 305 -1142 321 -766
rect 255 -1154 321 -1142
rect 351 -766 417 -754
rect 351 -1142 367 -766
rect 401 -1142 417 -766
rect 351 -1154 417 -1142
rect 447 -766 509 -754
rect 447 -1142 463 -766
rect 497 -1142 509 -766
rect 447 -1154 509 -1142
<< pdiffc >>
rect -497 766 -463 1142
rect -401 766 -367 1142
rect -305 766 -271 1142
rect -209 766 -175 1142
rect -113 766 -79 1142
rect -17 766 17 1142
rect 79 766 113 1142
rect 175 766 209 1142
rect 271 766 305 1142
rect 367 766 401 1142
rect 463 766 497 1142
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect -497 -1142 -463 -766
rect -401 -1142 -367 -766
rect -305 -1142 -271 -766
rect -209 -1142 -175 -766
rect -113 -1142 -79 -766
rect -17 -1142 17 -766
rect 79 -1142 113 -766
rect 175 -1142 209 -766
rect 271 -1142 305 -766
rect 367 -1142 401 -766
rect 463 -1142 497 -766
<< nsubdiff >>
rect -611 1303 -515 1337
rect 515 1303 611 1337
rect -611 1241 -577 1303
rect 577 1241 611 1303
rect -611 -1303 -577 -1241
rect 577 -1303 611 -1241
rect -611 -1337 -515 -1303
rect 515 -1337 611 -1303
<< nsubdiffcont >>
rect -515 1303 515 1337
rect -611 -1241 -577 1241
rect 577 -1241 611 1241
rect -515 -1337 515 -1303
<< poly >>
rect -465 1235 -399 1251
rect -465 1201 -449 1235
rect -415 1201 -399 1235
rect -465 1185 -399 1201
rect -273 1235 -207 1251
rect -273 1201 -257 1235
rect -223 1201 -207 1235
rect -273 1185 -207 1201
rect -81 1235 -15 1251
rect -81 1201 -65 1235
rect -31 1201 -15 1235
rect -81 1185 -15 1201
rect 111 1235 177 1251
rect 111 1201 127 1235
rect 161 1201 177 1235
rect 111 1185 177 1201
rect 303 1235 369 1251
rect 303 1201 319 1235
rect 353 1201 369 1235
rect 303 1185 369 1201
rect -447 1154 -417 1185
rect -351 1154 -321 1180
rect -255 1154 -225 1185
rect -159 1154 -129 1180
rect -63 1154 -33 1185
rect 33 1154 63 1180
rect 129 1154 159 1185
rect 225 1154 255 1180
rect 321 1154 351 1185
rect 417 1154 447 1180
rect -447 728 -417 754
rect -351 723 -321 754
rect -255 728 -225 754
rect -159 723 -129 754
rect -63 728 -33 754
rect 33 723 63 754
rect 129 728 159 754
rect 225 723 255 754
rect 321 728 351 754
rect 417 723 447 754
rect -369 707 -303 723
rect -369 673 -353 707
rect -319 673 -303 707
rect -369 657 -303 673
rect -177 707 -111 723
rect -177 673 -161 707
rect -127 673 -111 707
rect -177 657 -111 673
rect 15 707 81 723
rect 15 673 31 707
rect 65 673 81 707
rect 15 657 81 673
rect 207 707 273 723
rect 207 673 223 707
rect 257 673 273 707
rect 207 657 273 673
rect 399 707 465 723
rect 399 673 415 707
rect 449 673 465 707
rect 399 657 465 673
rect -369 599 -303 615
rect -369 565 -353 599
rect -319 565 -303 599
rect -369 549 -303 565
rect -177 599 -111 615
rect -177 565 -161 599
rect -127 565 -111 599
rect -177 549 -111 565
rect 15 599 81 615
rect 15 565 31 599
rect 65 565 81 599
rect 15 549 81 565
rect 207 599 273 615
rect 207 565 223 599
rect 257 565 273 599
rect 207 549 273 565
rect 399 599 465 615
rect 399 565 415 599
rect 449 565 465 599
rect 399 549 465 565
rect -447 518 -417 544
rect -351 518 -321 549
rect -255 518 -225 544
rect -159 518 -129 549
rect -63 518 -33 544
rect 33 518 63 549
rect 129 518 159 544
rect 225 518 255 549
rect 321 518 351 544
rect 417 518 447 549
rect -447 87 -417 118
rect -351 92 -321 118
rect -255 87 -225 118
rect -159 92 -129 118
rect -63 87 -33 118
rect 33 92 63 118
rect 129 87 159 118
rect 225 92 255 118
rect 321 87 351 118
rect 417 92 447 118
rect -465 71 -399 87
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 303 -87 369 -71
rect -447 -118 -417 -87
rect -351 -118 -321 -92
rect -255 -118 -225 -87
rect -159 -118 -129 -92
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect 129 -118 159 -87
rect 225 -118 255 -92
rect 321 -118 351 -87
rect 417 -118 447 -92
rect -447 -544 -417 -518
rect -351 -549 -321 -518
rect -255 -544 -225 -518
rect -159 -549 -129 -518
rect -63 -544 -33 -518
rect 33 -549 63 -518
rect 129 -544 159 -518
rect 225 -549 255 -518
rect 321 -544 351 -518
rect 417 -549 447 -518
rect -369 -565 -303 -549
rect -369 -599 -353 -565
rect -319 -599 -303 -565
rect -369 -615 -303 -599
rect -177 -565 -111 -549
rect -177 -599 -161 -565
rect -127 -599 -111 -565
rect -177 -615 -111 -599
rect 15 -565 81 -549
rect 15 -599 31 -565
rect 65 -599 81 -565
rect 15 -615 81 -599
rect 207 -565 273 -549
rect 207 -599 223 -565
rect 257 -599 273 -565
rect 207 -615 273 -599
rect 399 -565 465 -549
rect 399 -599 415 -565
rect 449 -599 465 -565
rect 399 -615 465 -599
rect -369 -673 -303 -657
rect -369 -707 -353 -673
rect -319 -707 -303 -673
rect -369 -723 -303 -707
rect -177 -673 -111 -657
rect -177 -707 -161 -673
rect -127 -707 -111 -673
rect -177 -723 -111 -707
rect 15 -673 81 -657
rect 15 -707 31 -673
rect 65 -707 81 -673
rect 15 -723 81 -707
rect 207 -673 273 -657
rect 207 -707 223 -673
rect 257 -707 273 -673
rect 207 -723 273 -707
rect 399 -673 465 -657
rect 399 -707 415 -673
rect 449 -707 465 -673
rect 399 -723 465 -707
rect -447 -754 -417 -728
rect -351 -754 -321 -723
rect -255 -754 -225 -728
rect -159 -754 -129 -723
rect -63 -754 -33 -728
rect 33 -754 63 -723
rect 129 -754 159 -728
rect 225 -754 255 -723
rect 321 -754 351 -728
rect 417 -754 447 -723
rect -447 -1185 -417 -1154
rect -351 -1180 -321 -1154
rect -255 -1185 -225 -1154
rect -159 -1180 -129 -1154
rect -63 -1185 -33 -1154
rect 33 -1180 63 -1154
rect 129 -1185 159 -1154
rect 225 -1180 255 -1154
rect 321 -1185 351 -1154
rect 417 -1180 447 -1154
rect -465 -1201 -399 -1185
rect -465 -1235 -449 -1201
rect -415 -1235 -399 -1201
rect -465 -1251 -399 -1235
rect -273 -1201 -207 -1185
rect -273 -1235 -257 -1201
rect -223 -1235 -207 -1201
rect -273 -1251 -207 -1235
rect -81 -1201 -15 -1185
rect -81 -1235 -65 -1201
rect -31 -1235 -15 -1201
rect -81 -1251 -15 -1235
rect 111 -1201 177 -1185
rect 111 -1235 127 -1201
rect 161 -1235 177 -1201
rect 111 -1251 177 -1235
rect 303 -1201 369 -1185
rect 303 -1235 319 -1201
rect 353 -1235 369 -1201
rect 303 -1251 369 -1235
<< polycont >>
rect -449 1201 -415 1235
rect -257 1201 -223 1235
rect -65 1201 -31 1235
rect 127 1201 161 1235
rect 319 1201 353 1235
rect -353 673 -319 707
rect -161 673 -127 707
rect 31 673 65 707
rect 223 673 257 707
rect 415 673 449 707
rect -353 565 -319 599
rect -161 565 -127 599
rect 31 565 65 599
rect 223 565 257 599
rect 415 565 449 599
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect -353 -599 -319 -565
rect -161 -599 -127 -565
rect 31 -599 65 -565
rect 223 -599 257 -565
rect 415 -599 449 -565
rect -353 -707 -319 -673
rect -161 -707 -127 -673
rect 31 -707 65 -673
rect 223 -707 257 -673
rect 415 -707 449 -673
rect -449 -1235 -415 -1201
rect -257 -1235 -223 -1201
rect -65 -1235 -31 -1201
rect 127 -1235 161 -1201
rect 319 -1235 353 -1201
<< locali >>
rect -611 1303 -515 1337
rect 515 1303 611 1337
rect -611 1241 -577 1303
rect 577 1241 611 1303
rect -465 1201 -449 1235
rect -415 1201 -399 1235
rect -273 1201 -257 1235
rect -223 1201 -207 1235
rect -81 1201 -65 1235
rect -31 1201 -15 1235
rect 111 1201 127 1235
rect 161 1201 177 1235
rect 303 1201 319 1235
rect 353 1201 369 1235
rect -497 1142 -463 1158
rect -497 750 -463 766
rect -401 1142 -367 1158
rect -401 750 -367 766
rect -305 1142 -271 1158
rect -305 750 -271 766
rect -209 1142 -175 1158
rect -209 750 -175 766
rect -113 1142 -79 1158
rect -113 750 -79 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 79 1142 113 1158
rect 79 750 113 766
rect 175 1142 209 1158
rect 175 750 209 766
rect 271 1142 305 1158
rect 271 750 305 766
rect 367 1142 401 1158
rect 367 750 401 766
rect 463 1142 497 1158
rect 463 750 497 766
rect -369 673 -353 707
rect -319 673 -303 707
rect -177 673 -161 707
rect -127 673 -111 707
rect 15 673 31 707
rect 65 673 81 707
rect 207 673 223 707
rect 257 673 273 707
rect 399 673 415 707
rect 449 673 465 707
rect -369 565 -353 599
rect -319 565 -303 599
rect -177 565 -161 599
rect -127 565 -111 599
rect 15 565 31 599
rect 65 565 81 599
rect 207 565 223 599
rect 257 565 273 599
rect 399 565 415 599
rect 449 565 465 599
rect -497 506 -463 522
rect -497 114 -463 130
rect -401 506 -367 522
rect -401 114 -367 130
rect -305 506 -271 522
rect -305 114 -271 130
rect -209 506 -175 522
rect -209 114 -175 130
rect -113 506 -79 522
rect -113 114 -79 130
rect -17 506 17 522
rect -17 114 17 130
rect 79 506 113 522
rect 79 114 113 130
rect 175 506 209 522
rect 175 114 209 130
rect 271 506 305 522
rect 271 114 305 130
rect 367 506 401 522
rect 367 114 401 130
rect 463 506 497 522
rect 463 114 497 130
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect -497 -130 -463 -114
rect -497 -522 -463 -506
rect -401 -130 -367 -114
rect -401 -522 -367 -506
rect -305 -130 -271 -114
rect -305 -522 -271 -506
rect -209 -130 -175 -114
rect -209 -522 -175 -506
rect -113 -130 -79 -114
rect -113 -522 -79 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 79 -130 113 -114
rect 79 -522 113 -506
rect 175 -130 209 -114
rect 175 -522 209 -506
rect 271 -130 305 -114
rect 271 -522 305 -506
rect 367 -130 401 -114
rect 367 -522 401 -506
rect 463 -130 497 -114
rect 463 -522 497 -506
rect -369 -599 -353 -565
rect -319 -599 -303 -565
rect -177 -599 -161 -565
rect -127 -599 -111 -565
rect 15 -599 31 -565
rect 65 -599 81 -565
rect 207 -599 223 -565
rect 257 -599 273 -565
rect 399 -599 415 -565
rect 449 -599 465 -565
rect -369 -707 -353 -673
rect -319 -707 -303 -673
rect -177 -707 -161 -673
rect -127 -707 -111 -673
rect 15 -707 31 -673
rect 65 -707 81 -673
rect 207 -707 223 -673
rect 257 -707 273 -673
rect 399 -707 415 -673
rect 449 -707 465 -673
rect -497 -766 -463 -750
rect -497 -1158 -463 -1142
rect -401 -766 -367 -750
rect -401 -1158 -367 -1142
rect -305 -766 -271 -750
rect -305 -1158 -271 -1142
rect -209 -766 -175 -750
rect -209 -1158 -175 -1142
rect -113 -766 -79 -750
rect -113 -1158 -79 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 79 -766 113 -750
rect 79 -1158 113 -1142
rect 175 -766 209 -750
rect 175 -1158 209 -1142
rect 271 -766 305 -750
rect 271 -1158 305 -1142
rect 367 -766 401 -750
rect 367 -1158 401 -1142
rect 463 -766 497 -750
rect 463 -1158 497 -1142
rect -465 -1235 -449 -1201
rect -415 -1235 -399 -1201
rect -273 -1235 -257 -1201
rect -223 -1235 -207 -1201
rect -81 -1235 -65 -1201
rect -31 -1235 -15 -1201
rect 111 -1235 127 -1201
rect 161 -1235 177 -1201
rect 303 -1235 319 -1201
rect 353 -1235 369 -1201
rect -611 -1303 -577 -1241
rect 577 -1303 611 -1241
rect -611 -1337 -515 -1303
rect 515 -1337 611 -1303
<< viali >>
rect -449 1201 -415 1235
rect -257 1201 -223 1235
rect -65 1201 -31 1235
rect 127 1201 161 1235
rect 319 1201 353 1235
rect -497 766 -463 1142
rect -401 766 -367 1142
rect -305 766 -271 1142
rect -209 766 -175 1142
rect -113 766 -79 1142
rect -17 766 17 1142
rect 79 766 113 1142
rect 175 766 209 1142
rect 271 766 305 1142
rect 367 766 401 1142
rect 463 766 497 1142
rect -353 673 -319 707
rect -161 673 -127 707
rect 31 673 65 707
rect 223 673 257 707
rect 415 673 449 707
rect -353 565 -319 599
rect -161 565 -127 599
rect 31 565 65 599
rect 223 565 257 599
rect 415 565 449 599
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect -353 -599 -319 -565
rect -161 -599 -127 -565
rect 31 -599 65 -565
rect 223 -599 257 -565
rect 415 -599 449 -565
rect -353 -707 -319 -673
rect -161 -707 -127 -673
rect 31 -707 65 -673
rect 223 -707 257 -673
rect 415 -707 449 -673
rect -497 -1142 -463 -766
rect -401 -1142 -367 -766
rect -305 -1142 -271 -766
rect -209 -1142 -175 -766
rect -113 -1142 -79 -766
rect -17 -1142 17 -766
rect 79 -1142 113 -766
rect 175 -1142 209 -766
rect 271 -1142 305 -766
rect 367 -1142 401 -766
rect 463 -1142 497 -766
rect -449 -1235 -415 -1201
rect -257 -1235 -223 -1201
rect -65 -1235 -31 -1201
rect 127 -1235 161 -1201
rect 319 -1235 353 -1201
<< metal1 >>
rect -461 1235 -403 1241
rect -461 1201 -449 1235
rect -415 1201 -403 1235
rect -461 1195 -403 1201
rect -269 1235 -211 1241
rect -269 1201 -257 1235
rect -223 1201 -211 1235
rect -269 1195 -211 1201
rect -77 1235 -19 1241
rect -77 1201 -65 1235
rect -31 1201 -19 1235
rect -77 1195 -19 1201
rect 115 1235 173 1241
rect 115 1201 127 1235
rect 161 1201 173 1235
rect 115 1195 173 1201
rect 307 1235 365 1241
rect 307 1201 319 1235
rect 353 1201 365 1235
rect 307 1195 365 1201
rect -503 1142 -457 1154
rect -503 766 -497 1142
rect -463 766 -457 1142
rect -503 754 -457 766
rect -407 1142 -361 1154
rect -407 766 -401 1142
rect -367 766 -361 1142
rect -407 754 -361 766
rect -311 1142 -265 1154
rect -311 766 -305 1142
rect -271 766 -265 1142
rect -311 754 -265 766
rect -215 1142 -169 1154
rect -215 766 -209 1142
rect -175 766 -169 1142
rect -215 754 -169 766
rect -119 1142 -73 1154
rect -119 766 -113 1142
rect -79 766 -73 1142
rect -119 754 -73 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 73 1142 119 1154
rect 73 766 79 1142
rect 113 766 119 1142
rect 73 754 119 766
rect 169 1142 215 1154
rect 169 766 175 1142
rect 209 766 215 1142
rect 169 754 215 766
rect 265 1142 311 1154
rect 265 766 271 1142
rect 305 766 311 1142
rect 265 754 311 766
rect 361 1142 407 1154
rect 361 766 367 1142
rect 401 766 407 1142
rect 361 754 407 766
rect 457 1142 503 1154
rect 457 766 463 1142
rect 497 766 503 1142
rect 457 754 503 766
rect -365 707 -307 713
rect -365 673 -353 707
rect -319 673 -307 707
rect -365 667 -307 673
rect -173 707 -115 713
rect -173 673 -161 707
rect -127 673 -115 707
rect -173 667 -115 673
rect 19 707 77 713
rect 19 673 31 707
rect 65 673 77 707
rect 19 667 77 673
rect 211 707 269 713
rect 211 673 223 707
rect 257 673 269 707
rect 211 667 269 673
rect 403 707 461 713
rect 403 673 415 707
rect 449 673 461 707
rect 403 667 461 673
rect -365 599 -307 605
rect -365 565 -353 599
rect -319 565 -307 599
rect -365 559 -307 565
rect -173 599 -115 605
rect -173 565 -161 599
rect -127 565 -115 599
rect -173 559 -115 565
rect 19 599 77 605
rect 19 565 31 599
rect 65 565 77 599
rect 19 559 77 565
rect 211 599 269 605
rect 211 565 223 599
rect 257 565 269 599
rect 211 559 269 565
rect 403 599 461 605
rect 403 565 415 599
rect 449 565 461 599
rect 403 559 461 565
rect -503 506 -457 518
rect -503 130 -497 506
rect -463 130 -457 506
rect -503 118 -457 130
rect -407 506 -361 518
rect -407 130 -401 506
rect -367 130 -361 506
rect -407 118 -361 130
rect -311 506 -265 518
rect -311 130 -305 506
rect -271 130 -265 506
rect -311 118 -265 130
rect -215 506 -169 518
rect -215 130 -209 506
rect -175 130 -169 506
rect -215 118 -169 130
rect -119 506 -73 518
rect -119 130 -113 506
rect -79 130 -73 506
rect -119 118 -73 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 73 506 119 518
rect 73 130 79 506
rect 113 130 119 506
rect 73 118 119 130
rect 169 506 215 518
rect 169 130 175 506
rect 209 130 215 506
rect 169 118 215 130
rect 265 506 311 518
rect 265 130 271 506
rect 305 130 311 506
rect 265 118 311 130
rect 361 506 407 518
rect 361 130 367 506
rect 401 130 407 506
rect 361 118 407 130
rect 457 506 503 518
rect 457 130 463 506
rect 497 130 503 506
rect 457 118 503 130
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect -503 -130 -457 -118
rect -503 -506 -497 -130
rect -463 -506 -457 -130
rect -503 -518 -457 -506
rect -407 -130 -361 -118
rect -407 -506 -401 -130
rect -367 -506 -361 -130
rect -407 -518 -361 -506
rect -311 -130 -265 -118
rect -311 -506 -305 -130
rect -271 -506 -265 -130
rect -311 -518 -265 -506
rect -215 -130 -169 -118
rect -215 -506 -209 -130
rect -175 -506 -169 -130
rect -215 -518 -169 -506
rect -119 -130 -73 -118
rect -119 -506 -113 -130
rect -79 -506 -73 -130
rect -119 -518 -73 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 73 -130 119 -118
rect 73 -506 79 -130
rect 113 -506 119 -130
rect 73 -518 119 -506
rect 169 -130 215 -118
rect 169 -506 175 -130
rect 209 -506 215 -130
rect 169 -518 215 -506
rect 265 -130 311 -118
rect 265 -506 271 -130
rect 305 -506 311 -130
rect 265 -518 311 -506
rect 361 -130 407 -118
rect 361 -506 367 -130
rect 401 -506 407 -130
rect 361 -518 407 -506
rect 457 -130 503 -118
rect 457 -506 463 -130
rect 497 -506 503 -130
rect 457 -518 503 -506
rect -365 -565 -307 -559
rect -365 -599 -353 -565
rect -319 -599 -307 -565
rect -365 -605 -307 -599
rect -173 -565 -115 -559
rect -173 -599 -161 -565
rect -127 -599 -115 -565
rect -173 -605 -115 -599
rect 19 -565 77 -559
rect 19 -599 31 -565
rect 65 -599 77 -565
rect 19 -605 77 -599
rect 211 -565 269 -559
rect 211 -599 223 -565
rect 257 -599 269 -565
rect 211 -605 269 -599
rect 403 -565 461 -559
rect 403 -599 415 -565
rect 449 -599 461 -565
rect 403 -605 461 -599
rect -365 -673 -307 -667
rect -365 -707 -353 -673
rect -319 -707 -307 -673
rect -365 -713 -307 -707
rect -173 -673 -115 -667
rect -173 -707 -161 -673
rect -127 -707 -115 -673
rect -173 -713 -115 -707
rect 19 -673 77 -667
rect 19 -707 31 -673
rect 65 -707 77 -673
rect 19 -713 77 -707
rect 211 -673 269 -667
rect 211 -707 223 -673
rect 257 -707 269 -673
rect 211 -713 269 -707
rect 403 -673 461 -667
rect 403 -707 415 -673
rect 449 -707 461 -673
rect 403 -713 461 -707
rect -503 -766 -457 -754
rect -503 -1142 -497 -766
rect -463 -1142 -457 -766
rect -503 -1154 -457 -1142
rect -407 -766 -361 -754
rect -407 -1142 -401 -766
rect -367 -1142 -361 -766
rect -407 -1154 -361 -1142
rect -311 -766 -265 -754
rect -311 -1142 -305 -766
rect -271 -1142 -265 -766
rect -311 -1154 -265 -1142
rect -215 -766 -169 -754
rect -215 -1142 -209 -766
rect -175 -1142 -169 -766
rect -215 -1154 -169 -1142
rect -119 -766 -73 -754
rect -119 -1142 -113 -766
rect -79 -1142 -73 -766
rect -119 -1154 -73 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 73 -766 119 -754
rect 73 -1142 79 -766
rect 113 -1142 119 -766
rect 73 -1154 119 -1142
rect 169 -766 215 -754
rect 169 -1142 175 -766
rect 209 -1142 215 -766
rect 169 -1154 215 -1142
rect 265 -766 311 -754
rect 265 -1142 271 -766
rect 305 -1142 311 -766
rect 265 -1154 311 -1142
rect 361 -766 407 -754
rect 361 -1142 367 -766
rect 401 -1142 407 -766
rect 361 -1154 407 -1142
rect 457 -766 503 -754
rect 457 -1142 463 -766
rect 497 -1142 503 -766
rect 457 -1154 503 -1142
rect -461 -1201 -403 -1195
rect -461 -1235 -449 -1201
rect -415 -1235 -403 -1201
rect -461 -1241 -403 -1235
rect -269 -1201 -211 -1195
rect -269 -1235 -257 -1201
rect -223 -1235 -211 -1201
rect -269 -1241 -211 -1235
rect -77 -1201 -19 -1195
rect -77 -1235 -65 -1201
rect -31 -1235 -19 -1201
rect -77 -1241 -19 -1235
rect 115 -1201 173 -1195
rect 115 -1235 127 -1201
rect 161 -1235 173 -1201
rect 115 -1241 173 -1235
rect 307 -1201 365 -1195
rect 307 -1235 319 -1201
rect 353 -1235 365 -1201
rect 307 -1241 365 -1235
<< properties >>
string FIXED_BBOX -594 -1320 594 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 4 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
