magic
tech sky130A
magscale 1 2
timestamp 1683564698
<< error_p >>
rect -6070 1945 -4010 1972
rect -3550 1945 -1490 1972
rect -1030 1945 1030 1972
rect 1490 1945 3550 1972
rect 4010 1945 6070 1972
rect -6070 1136 -4010 1163
rect -3550 1136 -1490 1163
rect -1030 1136 1030 1163
rect 1490 1136 3550 1163
rect 4010 1136 6070 1163
rect -6070 909 -4010 936
rect -3550 909 -1490 936
rect -1030 909 1030 936
rect 1490 909 3550 936
rect 4010 909 6070 936
rect -6070 100 -4010 127
rect -3550 100 -1490 127
rect -1030 100 1030 127
rect 1490 100 3550 127
rect 4010 100 6070 127
rect -6070 -127 -4010 -100
rect -3550 -127 -1490 -100
rect -1030 -127 1030 -100
rect 1490 -127 3550 -100
rect 4010 -127 6070 -100
rect -6070 -936 -4010 -909
rect -3550 -936 -1490 -909
rect -1030 -936 1030 -909
rect 1490 -936 3550 -909
rect 4010 -936 6070 -909
rect -6070 -1163 -4010 -1136
rect -3550 -1163 -1490 -1136
rect -1030 -1163 1030 -1136
rect 1490 -1163 3550 -1136
rect 4010 -1163 6070 -1136
rect -6070 -1972 -4010 -1945
rect -3550 -1972 -1490 -1945
rect -1030 -1972 1030 -1945
rect 1490 -1972 3550 -1945
rect 4010 -1972 6070 -1945
<< nwell >>
rect -6173 1163 -3907 1945
rect -3653 1163 -1387 1945
rect -1133 1163 1133 1945
rect 1387 1163 3653 1945
rect 3907 1163 6173 1945
rect -6173 127 -3907 909
rect -3653 127 -1387 909
rect -1133 127 1133 909
rect 1387 127 3653 909
rect 3907 127 6173 909
rect -6173 -909 -3907 -127
rect -3653 -909 -1387 -127
rect -1133 -909 1133 -127
rect 1387 -909 3653 -127
rect 3907 -909 6173 -127
rect -6173 -1945 -3907 -1163
rect -3653 -1945 -1387 -1163
rect -1133 -1945 1133 -1163
rect 1387 -1945 3653 -1163
rect 3907 -1945 6173 -1163
<< pwell >>
rect -6283 1945 6283 2055
rect -6283 1163 -6173 1945
rect -3907 1163 -3653 1945
rect -1387 1163 -1133 1945
rect 1133 1163 1387 1945
rect 3653 1163 3907 1945
rect 6173 1163 6283 1945
rect -6283 909 6283 1163
rect -6283 127 -6173 909
rect -3907 127 -3653 909
rect -1387 127 -1133 909
rect 1133 127 1387 909
rect 3653 127 3907 909
rect 6173 127 6283 909
rect -6283 -127 6283 127
rect -6283 -909 -6173 -127
rect -3907 -909 -3653 -127
rect -1387 -909 -1133 -127
rect 1133 -909 1387 -127
rect 3653 -909 3907 -127
rect 6173 -909 6283 -127
rect -6283 -1163 6283 -909
rect -6283 -1945 -6173 -1163
rect -3907 -1945 -3653 -1163
rect -1387 -1945 -1133 -1163
rect 1133 -1945 1387 -1163
rect 3653 -1945 3907 -1163
rect 6173 -1945 6283 -1163
rect -6283 -2055 6283 -1945
<< varactor >>
rect -6040 1254 -4040 1854
rect -3520 1254 -1520 1854
rect -1000 1254 1000 1854
rect 1520 1254 3520 1854
rect 4040 1254 6040 1854
rect -6040 218 -4040 818
rect -3520 218 -1520 818
rect -1000 218 1000 818
rect 1520 218 3520 818
rect 4040 218 6040 818
rect -6040 -818 -4040 -218
rect -3520 -818 -1520 -218
rect -1000 -818 1000 -218
rect 1520 -818 3520 -218
rect 4040 -818 6040 -218
rect -6040 -1854 -4040 -1254
rect -3520 -1854 -1520 -1254
rect -1000 -1854 1000 -1254
rect 1520 -1854 3520 -1254
rect 4040 -1854 6040 -1254
<< psubdiff >>
rect -6247 1985 -6151 2019
rect 6151 1985 6247 2019
rect -6247 1923 -6213 1985
rect 6213 1923 6247 1985
rect -6247 -1985 -6213 -1923
rect 6213 -1985 6247 -1923
rect -6247 -2019 -6151 -1985
rect 6151 -2019 6247 -1985
<< nsubdiff >>
rect -6137 1830 -6040 1854
rect -6137 1278 -6125 1830
rect -6091 1278 -6040 1830
rect -6137 1254 -6040 1278
rect -4040 1830 -3943 1854
rect -4040 1278 -3989 1830
rect -3955 1278 -3943 1830
rect -4040 1254 -3943 1278
rect -3617 1830 -3520 1854
rect -3617 1278 -3605 1830
rect -3571 1278 -3520 1830
rect -3617 1254 -3520 1278
rect -1520 1830 -1423 1854
rect -1520 1278 -1469 1830
rect -1435 1278 -1423 1830
rect -1520 1254 -1423 1278
rect -1097 1830 -1000 1854
rect -1097 1278 -1085 1830
rect -1051 1278 -1000 1830
rect -1097 1254 -1000 1278
rect 1000 1830 1097 1854
rect 1000 1278 1051 1830
rect 1085 1278 1097 1830
rect 1000 1254 1097 1278
rect 1423 1830 1520 1854
rect 1423 1278 1435 1830
rect 1469 1278 1520 1830
rect 1423 1254 1520 1278
rect 3520 1830 3617 1854
rect 3520 1278 3571 1830
rect 3605 1278 3617 1830
rect 3520 1254 3617 1278
rect 3943 1830 4040 1854
rect 3943 1278 3955 1830
rect 3989 1278 4040 1830
rect 3943 1254 4040 1278
rect 6040 1830 6137 1854
rect 6040 1278 6091 1830
rect 6125 1278 6137 1830
rect 6040 1254 6137 1278
rect -6137 794 -6040 818
rect -6137 242 -6125 794
rect -6091 242 -6040 794
rect -6137 218 -6040 242
rect -4040 794 -3943 818
rect -4040 242 -3989 794
rect -3955 242 -3943 794
rect -4040 218 -3943 242
rect -3617 794 -3520 818
rect -3617 242 -3605 794
rect -3571 242 -3520 794
rect -3617 218 -3520 242
rect -1520 794 -1423 818
rect -1520 242 -1469 794
rect -1435 242 -1423 794
rect -1520 218 -1423 242
rect -1097 794 -1000 818
rect -1097 242 -1085 794
rect -1051 242 -1000 794
rect -1097 218 -1000 242
rect 1000 794 1097 818
rect 1000 242 1051 794
rect 1085 242 1097 794
rect 1000 218 1097 242
rect 1423 794 1520 818
rect 1423 242 1435 794
rect 1469 242 1520 794
rect 1423 218 1520 242
rect 3520 794 3617 818
rect 3520 242 3571 794
rect 3605 242 3617 794
rect 3520 218 3617 242
rect 3943 794 4040 818
rect 3943 242 3955 794
rect 3989 242 4040 794
rect 3943 218 4040 242
rect 6040 794 6137 818
rect 6040 242 6091 794
rect 6125 242 6137 794
rect 6040 218 6137 242
rect -6137 -242 -6040 -218
rect -6137 -794 -6125 -242
rect -6091 -794 -6040 -242
rect -6137 -818 -6040 -794
rect -4040 -242 -3943 -218
rect -4040 -794 -3989 -242
rect -3955 -794 -3943 -242
rect -4040 -818 -3943 -794
rect -3617 -242 -3520 -218
rect -3617 -794 -3605 -242
rect -3571 -794 -3520 -242
rect -3617 -818 -3520 -794
rect -1520 -242 -1423 -218
rect -1520 -794 -1469 -242
rect -1435 -794 -1423 -242
rect -1520 -818 -1423 -794
rect -1097 -242 -1000 -218
rect -1097 -794 -1085 -242
rect -1051 -794 -1000 -242
rect -1097 -818 -1000 -794
rect 1000 -242 1097 -218
rect 1000 -794 1051 -242
rect 1085 -794 1097 -242
rect 1000 -818 1097 -794
rect 1423 -242 1520 -218
rect 1423 -794 1435 -242
rect 1469 -794 1520 -242
rect 1423 -818 1520 -794
rect 3520 -242 3617 -218
rect 3520 -794 3571 -242
rect 3605 -794 3617 -242
rect 3520 -818 3617 -794
rect 3943 -242 4040 -218
rect 3943 -794 3955 -242
rect 3989 -794 4040 -242
rect 3943 -818 4040 -794
rect 6040 -242 6137 -218
rect 6040 -794 6091 -242
rect 6125 -794 6137 -242
rect 6040 -818 6137 -794
rect -6137 -1278 -6040 -1254
rect -6137 -1830 -6125 -1278
rect -6091 -1830 -6040 -1278
rect -6137 -1854 -6040 -1830
rect -4040 -1278 -3943 -1254
rect -4040 -1830 -3989 -1278
rect -3955 -1830 -3943 -1278
rect -4040 -1854 -3943 -1830
rect -3617 -1278 -3520 -1254
rect -3617 -1830 -3605 -1278
rect -3571 -1830 -3520 -1278
rect -3617 -1854 -3520 -1830
rect -1520 -1278 -1423 -1254
rect -1520 -1830 -1469 -1278
rect -1435 -1830 -1423 -1278
rect -1520 -1854 -1423 -1830
rect -1097 -1278 -1000 -1254
rect -1097 -1830 -1085 -1278
rect -1051 -1830 -1000 -1278
rect -1097 -1854 -1000 -1830
rect 1000 -1278 1097 -1254
rect 1000 -1830 1051 -1278
rect 1085 -1830 1097 -1278
rect 1000 -1854 1097 -1830
rect 1423 -1278 1520 -1254
rect 1423 -1830 1435 -1278
rect 1469 -1830 1520 -1278
rect 1423 -1854 1520 -1830
rect 3520 -1278 3617 -1254
rect 3520 -1830 3571 -1278
rect 3605 -1830 3617 -1278
rect 3520 -1854 3617 -1830
rect 3943 -1278 4040 -1254
rect 3943 -1830 3955 -1278
rect 3989 -1830 4040 -1278
rect 3943 -1854 4040 -1830
rect 6040 -1278 6137 -1254
rect 6040 -1830 6091 -1278
rect 6125 -1830 6137 -1278
rect 6040 -1854 6137 -1830
<< psubdiffcont >>
rect -6151 1985 6151 2019
rect -6247 -1923 -6213 1923
rect 6213 -1923 6247 1923
rect -6151 -2019 6151 -1985
<< nsubdiffcont >>
rect -6125 1278 -6091 1830
rect -3989 1278 -3955 1830
rect -3605 1278 -3571 1830
rect -1469 1278 -1435 1830
rect -1085 1278 -1051 1830
rect 1051 1278 1085 1830
rect 1435 1278 1469 1830
rect 3571 1278 3605 1830
rect 3955 1278 3989 1830
rect 6091 1278 6125 1830
rect -6125 242 -6091 794
rect -3989 242 -3955 794
rect -3605 242 -3571 794
rect -1469 242 -1435 794
rect -1085 242 -1051 794
rect 1051 242 1085 794
rect 1435 242 1469 794
rect 3571 242 3605 794
rect 3955 242 3989 794
rect 6091 242 6125 794
rect -6125 -794 -6091 -242
rect -3989 -794 -3955 -242
rect -3605 -794 -3571 -242
rect -1469 -794 -1435 -242
rect -1085 -794 -1051 -242
rect 1051 -794 1085 -242
rect 1435 -794 1469 -242
rect 3571 -794 3605 -242
rect 3955 -794 3989 -242
rect 6091 -794 6125 -242
rect -6125 -1830 -6091 -1278
rect -3989 -1830 -3955 -1278
rect -3605 -1830 -3571 -1278
rect -1469 -1830 -1435 -1278
rect -1085 -1830 -1051 -1278
rect 1051 -1830 1085 -1278
rect 1435 -1830 1469 -1278
rect 3571 -1830 3605 -1278
rect 3955 -1830 3989 -1278
rect 6091 -1830 6125 -1278
<< poly >>
rect -6040 1926 -4040 1942
rect -6040 1892 -6024 1926
rect -4056 1892 -4040 1926
rect -6040 1854 -4040 1892
rect -3520 1926 -1520 1942
rect -3520 1892 -3504 1926
rect -1536 1892 -1520 1926
rect -3520 1854 -1520 1892
rect -1000 1926 1000 1942
rect -1000 1892 -984 1926
rect 984 1892 1000 1926
rect -1000 1854 1000 1892
rect 1520 1926 3520 1942
rect 1520 1892 1536 1926
rect 3504 1892 3520 1926
rect 1520 1854 3520 1892
rect 4040 1926 6040 1942
rect 4040 1892 4056 1926
rect 6024 1892 6040 1926
rect 4040 1854 6040 1892
rect -6040 1216 -4040 1254
rect -6040 1182 -6024 1216
rect -4056 1182 -4040 1216
rect -6040 1166 -4040 1182
rect -3520 1216 -1520 1254
rect -3520 1182 -3504 1216
rect -1536 1182 -1520 1216
rect -3520 1166 -1520 1182
rect -1000 1216 1000 1254
rect -1000 1182 -984 1216
rect 984 1182 1000 1216
rect -1000 1166 1000 1182
rect 1520 1216 3520 1254
rect 1520 1182 1536 1216
rect 3504 1182 3520 1216
rect 1520 1166 3520 1182
rect 4040 1216 6040 1254
rect 4040 1182 4056 1216
rect 6024 1182 6040 1216
rect 4040 1166 6040 1182
rect -6040 890 -4040 906
rect -6040 856 -6024 890
rect -4056 856 -4040 890
rect -6040 818 -4040 856
rect -3520 890 -1520 906
rect -3520 856 -3504 890
rect -1536 856 -1520 890
rect -3520 818 -1520 856
rect -1000 890 1000 906
rect -1000 856 -984 890
rect 984 856 1000 890
rect -1000 818 1000 856
rect 1520 890 3520 906
rect 1520 856 1536 890
rect 3504 856 3520 890
rect 1520 818 3520 856
rect 4040 890 6040 906
rect 4040 856 4056 890
rect 6024 856 6040 890
rect 4040 818 6040 856
rect -6040 180 -4040 218
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -6040 130 -4040 146
rect -3520 180 -1520 218
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -3520 130 -1520 146
rect -1000 180 1000 218
rect -1000 146 -984 180
rect 984 146 1000 180
rect -1000 130 1000 146
rect 1520 180 3520 218
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 1520 130 3520 146
rect 4040 180 6040 218
rect 4040 146 4056 180
rect 6024 146 6040 180
rect 4040 130 6040 146
rect -6040 -146 -4040 -130
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -6040 -218 -4040 -180
rect -3520 -146 -1520 -130
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -3520 -218 -1520 -180
rect -1000 -146 1000 -130
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect -1000 -218 1000 -180
rect 1520 -146 3520 -130
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 1520 -218 3520 -180
rect 4040 -146 6040 -130
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect 4040 -218 6040 -180
rect -6040 -856 -4040 -818
rect -6040 -890 -6024 -856
rect -4056 -890 -4040 -856
rect -6040 -906 -4040 -890
rect -3520 -856 -1520 -818
rect -3520 -890 -3504 -856
rect -1536 -890 -1520 -856
rect -3520 -906 -1520 -890
rect -1000 -856 1000 -818
rect -1000 -890 -984 -856
rect 984 -890 1000 -856
rect -1000 -906 1000 -890
rect 1520 -856 3520 -818
rect 1520 -890 1536 -856
rect 3504 -890 3520 -856
rect 1520 -906 3520 -890
rect 4040 -856 6040 -818
rect 4040 -890 4056 -856
rect 6024 -890 6040 -856
rect 4040 -906 6040 -890
rect -6040 -1182 -4040 -1166
rect -6040 -1216 -6024 -1182
rect -4056 -1216 -4040 -1182
rect -6040 -1254 -4040 -1216
rect -3520 -1182 -1520 -1166
rect -3520 -1216 -3504 -1182
rect -1536 -1216 -1520 -1182
rect -3520 -1254 -1520 -1216
rect -1000 -1182 1000 -1166
rect -1000 -1216 -984 -1182
rect 984 -1216 1000 -1182
rect -1000 -1254 1000 -1216
rect 1520 -1182 3520 -1166
rect 1520 -1216 1536 -1182
rect 3504 -1216 3520 -1182
rect 1520 -1254 3520 -1216
rect 4040 -1182 6040 -1166
rect 4040 -1216 4056 -1182
rect 6024 -1216 6040 -1182
rect 4040 -1254 6040 -1216
rect -6040 -1892 -4040 -1854
rect -6040 -1926 -6024 -1892
rect -4056 -1926 -4040 -1892
rect -6040 -1942 -4040 -1926
rect -3520 -1892 -1520 -1854
rect -3520 -1926 -3504 -1892
rect -1536 -1926 -1520 -1892
rect -3520 -1942 -1520 -1926
rect -1000 -1892 1000 -1854
rect -1000 -1926 -984 -1892
rect 984 -1926 1000 -1892
rect -1000 -1942 1000 -1926
rect 1520 -1892 3520 -1854
rect 1520 -1926 1536 -1892
rect 3504 -1926 3520 -1892
rect 1520 -1942 3520 -1926
rect 4040 -1892 6040 -1854
rect 4040 -1926 4056 -1892
rect 6024 -1926 6040 -1892
rect 4040 -1942 6040 -1926
<< polycont >>
rect -6024 1892 -4056 1926
rect -3504 1892 -1536 1926
rect -984 1892 984 1926
rect 1536 1892 3504 1926
rect 4056 1892 6024 1926
rect -6024 1182 -4056 1216
rect -3504 1182 -1536 1216
rect -984 1182 984 1216
rect 1536 1182 3504 1216
rect 4056 1182 6024 1216
rect -6024 856 -4056 890
rect -3504 856 -1536 890
rect -984 856 984 890
rect 1536 856 3504 890
rect 4056 856 6024 890
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6024 -890 -4056 -856
rect -3504 -890 -1536 -856
rect -984 -890 984 -856
rect 1536 -890 3504 -856
rect 4056 -890 6024 -856
rect -6024 -1216 -4056 -1182
rect -3504 -1216 -1536 -1182
rect -984 -1216 984 -1182
rect 1536 -1216 3504 -1182
rect 4056 -1216 6024 -1182
rect -6024 -1926 -4056 -1892
rect -3504 -1926 -1536 -1892
rect -984 -1926 984 -1892
rect 1536 -1926 3504 -1892
rect 4056 -1926 6024 -1892
<< locali >>
rect -6247 1985 -6151 2019
rect 6151 1985 6247 2019
rect -6247 1923 -6213 1985
rect -6040 1892 -6024 1926
rect -4056 1892 -4040 1926
rect -3520 1892 -3504 1926
rect -1536 1892 -1520 1926
rect -1000 1892 -984 1926
rect 984 1892 1000 1926
rect 1520 1892 1536 1926
rect 3504 1892 3520 1926
rect 4040 1892 4056 1926
rect 6024 1892 6040 1926
rect 6213 1923 6247 1985
rect -6125 1830 -6091 1846
rect -6125 1262 -6091 1278
rect -3989 1830 -3955 1846
rect -3989 1262 -3955 1278
rect -3605 1830 -3571 1846
rect -3605 1262 -3571 1278
rect -1469 1830 -1435 1846
rect -1469 1262 -1435 1278
rect -1085 1830 -1051 1846
rect -1085 1262 -1051 1278
rect 1051 1830 1085 1846
rect 1051 1262 1085 1278
rect 1435 1830 1469 1846
rect 1435 1262 1469 1278
rect 3571 1830 3605 1846
rect 3571 1262 3605 1278
rect 3955 1830 3989 1846
rect 3955 1262 3989 1278
rect 6091 1830 6125 1846
rect 6091 1262 6125 1278
rect -6040 1182 -6024 1216
rect -4056 1182 -4040 1216
rect -3520 1182 -3504 1216
rect -1536 1182 -1520 1216
rect -1000 1182 -984 1216
rect 984 1182 1000 1216
rect 1520 1182 1536 1216
rect 3504 1182 3520 1216
rect 4040 1182 4056 1216
rect 6024 1182 6040 1216
rect -6040 856 -6024 890
rect -4056 856 -4040 890
rect -3520 856 -3504 890
rect -1536 856 -1520 890
rect -1000 856 -984 890
rect 984 856 1000 890
rect 1520 856 1536 890
rect 3504 856 3520 890
rect 4040 856 4056 890
rect 6024 856 6040 890
rect -6125 794 -6091 810
rect -6125 226 -6091 242
rect -3989 794 -3955 810
rect -3989 226 -3955 242
rect -3605 794 -3571 810
rect -3605 226 -3571 242
rect -1469 794 -1435 810
rect -1469 226 -1435 242
rect -1085 794 -1051 810
rect -1085 226 -1051 242
rect 1051 794 1085 810
rect 1051 226 1085 242
rect 1435 794 1469 810
rect 1435 226 1469 242
rect 3571 794 3605 810
rect 3571 226 3605 242
rect 3955 794 3989 810
rect 3955 226 3989 242
rect 6091 794 6125 810
rect 6091 226 6125 242
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -1000 146 -984 180
rect 984 146 1000 180
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 4040 146 4056 180
rect 6024 146 6040 180
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect -6125 -242 -6091 -226
rect -6125 -810 -6091 -794
rect -3989 -242 -3955 -226
rect -3989 -810 -3955 -794
rect -3605 -242 -3571 -226
rect -3605 -810 -3571 -794
rect -1469 -242 -1435 -226
rect -1469 -810 -1435 -794
rect -1085 -242 -1051 -226
rect -1085 -810 -1051 -794
rect 1051 -242 1085 -226
rect 1051 -810 1085 -794
rect 1435 -242 1469 -226
rect 1435 -810 1469 -794
rect 3571 -242 3605 -226
rect 3571 -810 3605 -794
rect 3955 -242 3989 -226
rect 3955 -810 3989 -794
rect 6091 -242 6125 -226
rect 6091 -810 6125 -794
rect -6040 -890 -6024 -856
rect -4056 -890 -4040 -856
rect -3520 -890 -3504 -856
rect -1536 -890 -1520 -856
rect -1000 -890 -984 -856
rect 984 -890 1000 -856
rect 1520 -890 1536 -856
rect 3504 -890 3520 -856
rect 4040 -890 4056 -856
rect 6024 -890 6040 -856
rect -6040 -1216 -6024 -1182
rect -4056 -1216 -4040 -1182
rect -3520 -1216 -3504 -1182
rect -1536 -1216 -1520 -1182
rect -1000 -1216 -984 -1182
rect 984 -1216 1000 -1182
rect 1520 -1216 1536 -1182
rect 3504 -1216 3520 -1182
rect 4040 -1216 4056 -1182
rect 6024 -1216 6040 -1182
rect -6125 -1278 -6091 -1262
rect -6125 -1846 -6091 -1830
rect -3989 -1278 -3955 -1262
rect -3989 -1846 -3955 -1830
rect -3605 -1278 -3571 -1262
rect -3605 -1846 -3571 -1830
rect -1469 -1278 -1435 -1262
rect -1469 -1846 -1435 -1830
rect -1085 -1278 -1051 -1262
rect -1085 -1846 -1051 -1830
rect 1051 -1278 1085 -1262
rect 1051 -1846 1085 -1830
rect 1435 -1278 1469 -1262
rect 1435 -1846 1469 -1830
rect 3571 -1278 3605 -1262
rect 3571 -1846 3605 -1830
rect 3955 -1278 3989 -1262
rect 3955 -1846 3989 -1830
rect 6091 -1278 6125 -1262
rect 6091 -1846 6125 -1830
rect -6247 -1985 -6213 -1923
rect -6040 -1926 -6024 -1892
rect -4056 -1926 -4040 -1892
rect -3520 -1926 -3504 -1892
rect -1536 -1926 -1520 -1892
rect -1000 -1926 -984 -1892
rect 984 -1926 1000 -1892
rect 1520 -1926 1536 -1892
rect 3504 -1926 3520 -1892
rect 4040 -1926 4056 -1892
rect 6024 -1926 6040 -1892
rect 6213 -1985 6247 -1923
rect -6247 -2019 -6151 -1985
rect 6151 -2019 6247 -1985
<< viali >>
rect -6024 1892 -4056 1926
rect -3504 1892 -1536 1926
rect -984 1892 984 1926
rect 1536 1892 3504 1926
rect 4056 1892 6024 1926
rect -6125 1278 -6091 1830
rect -3989 1278 -3955 1830
rect -3605 1278 -3571 1830
rect -1469 1278 -1435 1830
rect -1085 1278 -1051 1830
rect 1051 1278 1085 1830
rect 1435 1278 1469 1830
rect 3571 1278 3605 1830
rect 3955 1278 3989 1830
rect 6091 1278 6125 1830
rect -6024 1182 -4056 1216
rect -3504 1182 -1536 1216
rect -984 1182 984 1216
rect 1536 1182 3504 1216
rect 4056 1182 6024 1216
rect -6024 856 -4056 890
rect -3504 856 -1536 890
rect -984 856 984 890
rect 1536 856 3504 890
rect 4056 856 6024 890
rect -6125 242 -6091 794
rect -3989 242 -3955 794
rect -3605 242 -3571 794
rect -1469 242 -1435 794
rect -1085 242 -1051 794
rect 1051 242 1085 794
rect 1435 242 1469 794
rect 3571 242 3605 794
rect 3955 242 3989 794
rect 6091 242 6125 794
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6125 -794 -6091 -242
rect -3989 -794 -3955 -242
rect -3605 -794 -3571 -242
rect -1469 -794 -1435 -242
rect -1085 -794 -1051 -242
rect 1051 -794 1085 -242
rect 1435 -794 1469 -242
rect 3571 -794 3605 -242
rect 3955 -794 3989 -242
rect 6091 -794 6125 -242
rect -6024 -890 -4056 -856
rect -3504 -890 -1536 -856
rect -984 -890 984 -856
rect 1536 -890 3504 -856
rect 4056 -890 6024 -856
rect -6024 -1216 -4056 -1182
rect -3504 -1216 -1536 -1182
rect -984 -1216 984 -1182
rect 1536 -1216 3504 -1182
rect 4056 -1216 6024 -1182
rect -6125 -1830 -6091 -1278
rect -3989 -1830 -3955 -1278
rect -3605 -1830 -3571 -1278
rect -1469 -1830 -1435 -1278
rect -1085 -1830 -1051 -1278
rect 1051 -1830 1085 -1278
rect 1435 -1830 1469 -1278
rect 3571 -1830 3605 -1278
rect 3955 -1830 3989 -1278
rect 6091 -1830 6125 -1278
rect -6024 -1926 -4056 -1892
rect -3504 -1926 -1536 -1892
rect -984 -1926 984 -1892
rect 1536 -1926 3504 -1892
rect 4056 -1926 6024 -1892
<< metal1 >>
rect -6036 1926 -4044 1932
rect -6036 1892 -6024 1926
rect -4056 1892 -4044 1926
rect -6036 1886 -4044 1892
rect -3516 1926 -1524 1932
rect -3516 1892 -3504 1926
rect -1536 1892 -1524 1926
rect -3516 1886 -1524 1892
rect -996 1926 996 1932
rect -996 1892 -984 1926
rect 984 1892 996 1926
rect -996 1886 996 1892
rect 1524 1926 3516 1932
rect 1524 1892 1536 1926
rect 3504 1892 3516 1926
rect 1524 1886 3516 1892
rect 4044 1926 6036 1932
rect 4044 1892 4056 1926
rect 6024 1892 6036 1926
rect 4044 1886 6036 1892
rect -6131 1830 -6085 1842
rect -3995 1830 -3949 1842
rect -6131 1278 -6125 1830
rect -6091 1278 -3989 1830
rect -3955 1278 -3949 1830
rect -6131 1266 -6085 1278
rect -3995 1266 -3949 1278
rect -3611 1830 -3565 1842
rect -1475 1830 -1429 1842
rect -3611 1278 -3605 1830
rect -3571 1278 -1469 1830
rect -1435 1278 -1429 1830
rect -3611 1266 -3565 1278
rect -1475 1266 -1429 1278
rect -1091 1830 -1045 1842
rect 1045 1830 1091 1842
rect -1091 1278 -1085 1830
rect -1051 1278 1051 1830
rect 1085 1278 1091 1830
rect -1091 1266 -1045 1278
rect 1045 1266 1091 1278
rect 1429 1830 1475 1842
rect 3565 1830 3611 1842
rect 1429 1278 1435 1830
rect 1469 1278 3571 1830
rect 3605 1278 3611 1830
rect 1429 1266 1475 1278
rect 3565 1266 3611 1278
rect 3949 1830 3995 1842
rect 6085 1830 6131 1842
rect 3949 1278 3955 1830
rect 3989 1278 6091 1830
rect 6125 1278 6131 1830
rect 3949 1266 3995 1278
rect 6085 1266 6131 1278
rect -6036 1216 -4044 1222
rect -6036 1182 -6024 1216
rect -4056 1182 -4044 1216
rect -6036 1176 -4044 1182
rect -3516 1216 -1524 1222
rect -3516 1182 -3504 1216
rect -1536 1182 -1524 1216
rect -3516 1176 -1524 1182
rect -996 1216 996 1222
rect -996 1182 -984 1216
rect 984 1182 996 1216
rect -996 1176 996 1182
rect 1524 1216 3516 1222
rect 1524 1182 1536 1216
rect 3504 1182 3516 1216
rect 1524 1176 3516 1182
rect 4044 1216 6036 1222
rect 4044 1182 4056 1216
rect 6024 1182 6036 1216
rect 4044 1176 6036 1182
rect -6036 890 -4044 896
rect -6036 856 -6024 890
rect -4056 856 -4044 890
rect -6036 850 -4044 856
rect -3516 890 -1524 896
rect -3516 856 -3504 890
rect -1536 856 -1524 890
rect -3516 850 -1524 856
rect -996 890 996 896
rect -996 856 -984 890
rect 984 856 996 890
rect -996 850 996 856
rect 1524 890 3516 896
rect 1524 856 1536 890
rect 3504 856 3516 890
rect 1524 850 3516 856
rect 4044 890 6036 896
rect 4044 856 4056 890
rect 6024 856 6036 890
rect 4044 850 6036 856
rect -6131 794 -6085 806
rect -3995 794 -3949 806
rect -6131 242 -6125 794
rect -6091 242 -3989 794
rect -3955 242 -3949 794
rect -6131 230 -6085 242
rect -3995 230 -3949 242
rect -3611 794 -3565 806
rect -1475 794 -1429 806
rect -3611 242 -3605 794
rect -3571 242 -1469 794
rect -1435 242 -1429 794
rect -3611 230 -3565 242
rect -1475 230 -1429 242
rect -1091 794 -1045 806
rect 1045 794 1091 806
rect -1091 242 -1085 794
rect -1051 242 1051 794
rect 1085 242 1091 794
rect -1091 230 -1045 242
rect 1045 230 1091 242
rect 1429 794 1475 806
rect 3565 794 3611 806
rect 1429 242 1435 794
rect 1469 242 3571 794
rect 3605 242 3611 794
rect 1429 230 1475 242
rect 3565 230 3611 242
rect 3949 794 3995 806
rect 6085 794 6131 806
rect 3949 242 3955 794
rect 3989 242 6091 794
rect 6125 242 6131 794
rect 3949 230 3995 242
rect 6085 230 6131 242
rect -6036 180 -4044 186
rect -6036 146 -6024 180
rect -4056 146 -4044 180
rect -6036 140 -4044 146
rect -3516 180 -1524 186
rect -3516 146 -3504 180
rect -1536 146 -1524 180
rect -3516 140 -1524 146
rect -996 180 996 186
rect -996 146 -984 180
rect 984 146 996 180
rect -996 140 996 146
rect 1524 180 3516 186
rect 1524 146 1536 180
rect 3504 146 3516 180
rect 1524 140 3516 146
rect 4044 180 6036 186
rect 4044 146 4056 180
rect 6024 146 6036 180
rect 4044 140 6036 146
rect -6036 -146 -4044 -140
rect -6036 -180 -6024 -146
rect -4056 -180 -4044 -146
rect -6036 -186 -4044 -180
rect -3516 -146 -1524 -140
rect -3516 -180 -3504 -146
rect -1536 -180 -1524 -146
rect -3516 -186 -1524 -180
rect -996 -146 996 -140
rect -996 -180 -984 -146
rect 984 -180 996 -146
rect -996 -186 996 -180
rect 1524 -146 3516 -140
rect 1524 -180 1536 -146
rect 3504 -180 3516 -146
rect 1524 -186 3516 -180
rect 4044 -146 6036 -140
rect 4044 -180 4056 -146
rect 6024 -180 6036 -146
rect 4044 -186 6036 -180
rect -6131 -242 -6085 -230
rect -3995 -242 -3949 -230
rect -6131 -794 -6125 -242
rect -6091 -794 -3989 -242
rect -3955 -794 -3949 -242
rect -6131 -806 -6085 -794
rect -3995 -806 -3949 -794
rect -3611 -242 -3565 -230
rect -1475 -242 -1429 -230
rect -3611 -794 -3605 -242
rect -3571 -794 -1469 -242
rect -1435 -794 -1429 -242
rect -3611 -806 -3565 -794
rect -1475 -806 -1429 -794
rect -1091 -242 -1045 -230
rect 1045 -242 1091 -230
rect -1091 -794 -1085 -242
rect -1051 -794 1051 -242
rect 1085 -794 1091 -242
rect -1091 -806 -1045 -794
rect 1045 -806 1091 -794
rect 1429 -242 1475 -230
rect 3565 -242 3611 -230
rect 1429 -794 1435 -242
rect 1469 -794 3571 -242
rect 3605 -794 3611 -242
rect 1429 -806 1475 -794
rect 3565 -806 3611 -794
rect 3949 -242 3995 -230
rect 6085 -242 6131 -230
rect 3949 -794 3955 -242
rect 3989 -794 6091 -242
rect 6125 -794 6131 -242
rect 3949 -806 3995 -794
rect 6085 -806 6131 -794
rect -6036 -856 -4044 -850
rect -6036 -890 -6024 -856
rect -4056 -890 -4044 -856
rect -6036 -896 -4044 -890
rect -3516 -856 -1524 -850
rect -3516 -890 -3504 -856
rect -1536 -890 -1524 -856
rect -3516 -896 -1524 -890
rect -996 -856 996 -850
rect -996 -890 -984 -856
rect 984 -890 996 -856
rect -996 -896 996 -890
rect 1524 -856 3516 -850
rect 1524 -890 1536 -856
rect 3504 -890 3516 -856
rect 1524 -896 3516 -890
rect 4044 -856 6036 -850
rect 4044 -890 4056 -856
rect 6024 -890 6036 -856
rect 4044 -896 6036 -890
rect -6036 -1182 -4044 -1176
rect -6036 -1216 -6024 -1182
rect -4056 -1216 -4044 -1182
rect -6036 -1222 -4044 -1216
rect -3516 -1182 -1524 -1176
rect -3516 -1216 -3504 -1182
rect -1536 -1216 -1524 -1182
rect -3516 -1222 -1524 -1216
rect -996 -1182 996 -1176
rect -996 -1216 -984 -1182
rect 984 -1216 996 -1182
rect -996 -1222 996 -1216
rect 1524 -1182 3516 -1176
rect 1524 -1216 1536 -1182
rect 3504 -1216 3516 -1182
rect 1524 -1222 3516 -1216
rect 4044 -1182 6036 -1176
rect 4044 -1216 4056 -1182
rect 6024 -1216 6036 -1182
rect 4044 -1222 6036 -1216
rect -6131 -1278 -6085 -1266
rect -3995 -1278 -3949 -1266
rect -6131 -1830 -6125 -1278
rect -6091 -1830 -3989 -1278
rect -3955 -1830 -3949 -1278
rect -6131 -1842 -6085 -1830
rect -3995 -1842 -3949 -1830
rect -3611 -1278 -3565 -1266
rect -1475 -1278 -1429 -1266
rect -3611 -1830 -3605 -1278
rect -3571 -1830 -1469 -1278
rect -1435 -1830 -1429 -1278
rect -3611 -1842 -3565 -1830
rect -1475 -1842 -1429 -1830
rect -1091 -1278 -1045 -1266
rect 1045 -1278 1091 -1266
rect -1091 -1830 -1085 -1278
rect -1051 -1830 1051 -1278
rect 1085 -1830 1091 -1278
rect -1091 -1842 -1045 -1830
rect 1045 -1842 1091 -1830
rect 1429 -1278 1475 -1266
rect 3565 -1278 3611 -1266
rect 1429 -1830 1435 -1278
rect 1469 -1830 3571 -1278
rect 3605 -1830 3611 -1278
rect 1429 -1842 1475 -1830
rect 3565 -1842 3611 -1830
rect 3949 -1278 3995 -1266
rect 6085 -1278 6131 -1266
rect 3949 -1830 3955 -1278
rect 3989 -1830 6091 -1278
rect 6125 -1830 6131 -1278
rect 3949 -1842 3995 -1830
rect 6085 -1842 6131 -1830
rect -6036 -1892 -4044 -1886
rect -6036 -1926 -6024 -1892
rect -4056 -1926 -4044 -1892
rect -6036 -1932 -4044 -1926
rect -3516 -1892 -1524 -1886
rect -3516 -1926 -3504 -1892
rect -1536 -1926 -1524 -1892
rect -3516 -1932 -1524 -1926
rect -996 -1892 996 -1886
rect -996 -1926 -984 -1892
rect 984 -1926 996 -1892
rect -996 -1932 996 -1926
rect 1524 -1892 3516 -1886
rect 1524 -1926 1536 -1892
rect 3504 -1926 3516 -1892
rect 1524 -1932 3516 -1926
rect 4044 -1892 6036 -1886
rect 4044 -1926 4056 -1892
rect 6024 -1926 6036 -1892
rect 4044 -1932 6036 -1926
<< properties >>
string FIXED_BBOX -6230 -2002 6230 2002
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 3 l 10 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
