magic
tech sky130A
magscale 1 2
timestamp 1683557511
<< error_p >>
rect -941 599 -883 605
rect -749 599 -691 605
rect -557 599 -499 605
rect -365 599 -307 605
rect -173 599 -115 605
rect 19 599 77 605
rect 211 599 269 605
rect 403 599 461 605
rect 595 599 653 605
rect 787 599 845 605
rect -941 565 -929 599
rect -749 565 -737 599
rect -557 565 -545 599
rect -365 565 -353 599
rect -173 565 -161 599
rect 19 565 31 599
rect 211 565 223 599
rect 403 565 415 599
rect 595 565 607 599
rect 787 565 799 599
rect -941 559 -883 565
rect -749 559 -691 565
rect -557 559 -499 565
rect -365 559 -307 565
rect -173 559 -115 565
rect 19 559 77 565
rect 211 559 269 565
rect 403 559 461 565
rect 595 559 653 565
rect 787 559 845 565
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect -941 -565 -883 -559
rect -749 -565 -691 -559
rect -557 -565 -499 -559
rect -365 -565 -307 -559
rect -173 -565 -115 -559
rect 19 -565 77 -559
rect 211 -565 269 -559
rect 403 -565 461 -559
rect 595 -565 653 -559
rect 787 -565 845 -559
rect -941 -599 -929 -565
rect -749 -599 -737 -565
rect -557 -599 -545 -565
rect -365 -599 -353 -565
rect -173 -599 -161 -565
rect 19 -599 31 -565
rect 211 -599 223 -565
rect 403 -599 415 -565
rect 595 -599 607 -565
rect 787 -599 799 -565
rect -941 -605 -883 -599
rect -749 -605 -691 -599
rect -557 -605 -499 -599
rect -365 -605 -307 -599
rect -173 -605 -115 -599
rect 19 -605 77 -599
rect 211 -605 269 -599
rect 403 -605 461 -599
rect 595 -605 653 -599
rect 787 -605 845 -599
<< nwell >>
rect -1127 -737 1127 737
<< pmos >>
rect -927 118 -897 518
rect -831 118 -801 518
rect -735 118 -705 518
rect -639 118 -609 518
rect -543 118 -513 518
rect -447 118 -417 518
rect -351 118 -321 518
rect -255 118 -225 518
rect -159 118 -129 518
rect -63 118 -33 518
rect 33 118 63 518
rect 129 118 159 518
rect 225 118 255 518
rect 321 118 351 518
rect 417 118 447 518
rect 513 118 543 518
rect 609 118 639 518
rect 705 118 735 518
rect 801 118 831 518
rect 897 118 927 518
rect -927 -518 -897 -118
rect -831 -518 -801 -118
rect -735 -518 -705 -118
rect -639 -518 -609 -118
rect -543 -518 -513 -118
rect -447 -518 -417 -118
rect -351 -518 -321 -118
rect -255 -518 -225 -118
rect -159 -518 -129 -118
rect -63 -518 -33 -118
rect 33 -518 63 -118
rect 129 -518 159 -118
rect 225 -518 255 -118
rect 321 -518 351 -118
rect 417 -518 447 -118
rect 513 -518 543 -118
rect 609 -518 639 -118
rect 705 -518 735 -118
rect 801 -518 831 -118
rect 897 -518 927 -118
<< pdiff >>
rect -989 506 -927 518
rect -989 130 -977 506
rect -943 130 -927 506
rect -989 118 -927 130
rect -897 506 -831 518
rect -897 130 -881 506
rect -847 130 -831 506
rect -897 118 -831 130
rect -801 506 -735 518
rect -801 130 -785 506
rect -751 130 -735 506
rect -801 118 -735 130
rect -705 506 -639 518
rect -705 130 -689 506
rect -655 130 -639 506
rect -705 118 -639 130
rect -609 506 -543 518
rect -609 130 -593 506
rect -559 130 -543 506
rect -609 118 -543 130
rect -513 506 -447 518
rect -513 130 -497 506
rect -463 130 -447 506
rect -513 118 -447 130
rect -417 506 -351 518
rect -417 130 -401 506
rect -367 130 -351 506
rect -417 118 -351 130
rect -321 506 -255 518
rect -321 130 -305 506
rect -271 130 -255 506
rect -321 118 -255 130
rect -225 506 -159 518
rect -225 130 -209 506
rect -175 130 -159 506
rect -225 118 -159 130
rect -129 506 -63 518
rect -129 130 -113 506
rect -79 130 -63 506
rect -129 118 -63 130
rect -33 506 33 518
rect -33 130 -17 506
rect 17 130 33 506
rect -33 118 33 130
rect 63 506 129 518
rect 63 130 79 506
rect 113 130 129 506
rect 63 118 129 130
rect 159 506 225 518
rect 159 130 175 506
rect 209 130 225 506
rect 159 118 225 130
rect 255 506 321 518
rect 255 130 271 506
rect 305 130 321 506
rect 255 118 321 130
rect 351 506 417 518
rect 351 130 367 506
rect 401 130 417 506
rect 351 118 417 130
rect 447 506 513 518
rect 447 130 463 506
rect 497 130 513 506
rect 447 118 513 130
rect 543 506 609 518
rect 543 130 559 506
rect 593 130 609 506
rect 543 118 609 130
rect 639 506 705 518
rect 639 130 655 506
rect 689 130 705 506
rect 639 118 705 130
rect 735 506 801 518
rect 735 130 751 506
rect 785 130 801 506
rect 735 118 801 130
rect 831 506 897 518
rect 831 130 847 506
rect 881 130 897 506
rect 831 118 897 130
rect 927 506 989 518
rect 927 130 943 506
rect 977 130 989 506
rect 927 118 989 130
rect -989 -130 -927 -118
rect -989 -506 -977 -130
rect -943 -506 -927 -130
rect -989 -518 -927 -506
rect -897 -130 -831 -118
rect -897 -506 -881 -130
rect -847 -506 -831 -130
rect -897 -518 -831 -506
rect -801 -130 -735 -118
rect -801 -506 -785 -130
rect -751 -506 -735 -130
rect -801 -518 -735 -506
rect -705 -130 -639 -118
rect -705 -506 -689 -130
rect -655 -506 -639 -130
rect -705 -518 -639 -506
rect -609 -130 -543 -118
rect -609 -506 -593 -130
rect -559 -506 -543 -130
rect -609 -518 -543 -506
rect -513 -130 -447 -118
rect -513 -506 -497 -130
rect -463 -506 -447 -130
rect -513 -518 -447 -506
rect -417 -130 -351 -118
rect -417 -506 -401 -130
rect -367 -506 -351 -130
rect -417 -518 -351 -506
rect -321 -130 -255 -118
rect -321 -506 -305 -130
rect -271 -506 -255 -130
rect -321 -518 -255 -506
rect -225 -130 -159 -118
rect -225 -506 -209 -130
rect -175 -506 -159 -130
rect -225 -518 -159 -506
rect -129 -130 -63 -118
rect -129 -506 -113 -130
rect -79 -506 -63 -130
rect -129 -518 -63 -506
rect -33 -130 33 -118
rect -33 -506 -17 -130
rect 17 -506 33 -130
rect -33 -518 33 -506
rect 63 -130 129 -118
rect 63 -506 79 -130
rect 113 -506 129 -130
rect 63 -518 129 -506
rect 159 -130 225 -118
rect 159 -506 175 -130
rect 209 -506 225 -130
rect 159 -518 225 -506
rect 255 -130 321 -118
rect 255 -506 271 -130
rect 305 -506 321 -130
rect 255 -518 321 -506
rect 351 -130 417 -118
rect 351 -506 367 -130
rect 401 -506 417 -130
rect 351 -518 417 -506
rect 447 -130 513 -118
rect 447 -506 463 -130
rect 497 -506 513 -130
rect 447 -518 513 -506
rect 543 -130 609 -118
rect 543 -506 559 -130
rect 593 -506 609 -130
rect 543 -518 609 -506
rect 639 -130 705 -118
rect 639 -506 655 -130
rect 689 -506 705 -130
rect 639 -518 705 -506
rect 735 -130 801 -118
rect 735 -506 751 -130
rect 785 -506 801 -130
rect 735 -518 801 -506
rect 831 -130 897 -118
rect 831 -506 847 -130
rect 881 -506 897 -130
rect 831 -518 897 -506
rect 927 -130 989 -118
rect 927 -506 943 -130
rect 977 -506 989 -130
rect 927 -518 989 -506
<< pdiffc >>
rect -977 130 -943 506
rect -881 130 -847 506
rect -785 130 -751 506
rect -689 130 -655 506
rect -593 130 -559 506
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect 559 130 593 506
rect 655 130 689 506
rect 751 130 785 506
rect 847 130 881 506
rect 943 130 977 506
rect -977 -506 -943 -130
rect -881 -506 -847 -130
rect -785 -506 -751 -130
rect -689 -506 -655 -130
rect -593 -506 -559 -130
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect 559 -506 593 -130
rect 655 -506 689 -130
rect 751 -506 785 -130
rect 847 -506 881 -130
rect 943 -506 977 -130
<< nsubdiff >>
rect -1091 667 -995 701
rect 995 667 1091 701
rect -1091 605 -1057 667
rect 1057 605 1091 667
rect -1091 -667 -1057 -605
rect 1057 -667 1091 -605
rect -1091 -701 -995 -667
rect 995 -701 1091 -667
<< nsubdiffcont >>
rect -995 667 995 701
rect -1091 -605 -1057 605
rect 1057 -605 1091 605
rect -995 -701 995 -667
<< poly >>
rect -945 599 -879 615
rect -945 565 -929 599
rect -895 565 -879 599
rect -945 549 -879 565
rect -753 599 -687 615
rect -753 565 -737 599
rect -703 565 -687 599
rect -753 549 -687 565
rect -561 599 -495 615
rect -561 565 -545 599
rect -511 565 -495 599
rect -561 549 -495 565
rect -369 599 -303 615
rect -369 565 -353 599
rect -319 565 -303 599
rect -369 549 -303 565
rect -177 599 -111 615
rect -177 565 -161 599
rect -127 565 -111 599
rect -177 549 -111 565
rect 15 599 81 615
rect 15 565 31 599
rect 65 565 81 599
rect 15 549 81 565
rect 207 599 273 615
rect 207 565 223 599
rect 257 565 273 599
rect 207 549 273 565
rect 399 599 465 615
rect 399 565 415 599
rect 449 565 465 599
rect 399 549 465 565
rect 591 599 657 615
rect 591 565 607 599
rect 641 565 657 599
rect 591 549 657 565
rect 783 599 849 615
rect 783 565 799 599
rect 833 565 849 599
rect 783 549 849 565
rect -927 518 -897 549
rect -831 518 -801 544
rect -735 518 -705 549
rect -639 518 -609 544
rect -543 518 -513 549
rect -447 518 -417 544
rect -351 518 -321 549
rect -255 518 -225 544
rect -159 518 -129 549
rect -63 518 -33 544
rect 33 518 63 549
rect 129 518 159 544
rect 225 518 255 549
rect 321 518 351 544
rect 417 518 447 549
rect 513 518 543 544
rect 609 518 639 549
rect 705 518 735 544
rect 801 518 831 549
rect 897 518 927 544
rect -927 92 -897 118
rect -831 87 -801 118
rect -735 92 -705 118
rect -639 87 -609 118
rect -543 92 -513 118
rect -447 87 -417 118
rect -351 92 -321 118
rect -255 87 -225 118
rect -159 92 -129 118
rect -63 87 -33 118
rect 33 92 63 118
rect 129 87 159 118
rect 225 92 255 118
rect 321 87 351 118
rect 417 92 447 118
rect 513 87 543 118
rect 609 92 639 118
rect 705 87 735 118
rect 801 92 831 118
rect 897 87 927 118
rect -849 71 -783 87
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 879 -87 945 -71
rect -927 -118 -897 -92
rect -831 -118 -801 -87
rect -735 -118 -705 -92
rect -639 -118 -609 -87
rect -543 -118 -513 -92
rect -447 -118 -417 -87
rect -351 -118 -321 -92
rect -255 -118 -225 -87
rect -159 -118 -129 -92
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect 129 -118 159 -87
rect 225 -118 255 -92
rect 321 -118 351 -87
rect 417 -118 447 -92
rect 513 -118 543 -87
rect 609 -118 639 -92
rect 705 -118 735 -87
rect 801 -118 831 -92
rect 897 -118 927 -87
rect -927 -549 -897 -518
rect -831 -544 -801 -518
rect -735 -549 -705 -518
rect -639 -544 -609 -518
rect -543 -549 -513 -518
rect -447 -544 -417 -518
rect -351 -549 -321 -518
rect -255 -544 -225 -518
rect -159 -549 -129 -518
rect -63 -544 -33 -518
rect 33 -549 63 -518
rect 129 -544 159 -518
rect 225 -549 255 -518
rect 321 -544 351 -518
rect 417 -549 447 -518
rect 513 -544 543 -518
rect 609 -549 639 -518
rect 705 -544 735 -518
rect 801 -549 831 -518
rect 897 -544 927 -518
rect -945 -565 -879 -549
rect -945 -599 -929 -565
rect -895 -599 -879 -565
rect -945 -615 -879 -599
rect -753 -565 -687 -549
rect -753 -599 -737 -565
rect -703 -599 -687 -565
rect -753 -615 -687 -599
rect -561 -565 -495 -549
rect -561 -599 -545 -565
rect -511 -599 -495 -565
rect -561 -615 -495 -599
rect -369 -565 -303 -549
rect -369 -599 -353 -565
rect -319 -599 -303 -565
rect -369 -615 -303 -599
rect -177 -565 -111 -549
rect -177 -599 -161 -565
rect -127 -599 -111 -565
rect -177 -615 -111 -599
rect 15 -565 81 -549
rect 15 -599 31 -565
rect 65 -599 81 -565
rect 15 -615 81 -599
rect 207 -565 273 -549
rect 207 -599 223 -565
rect 257 -599 273 -565
rect 207 -615 273 -599
rect 399 -565 465 -549
rect 399 -599 415 -565
rect 449 -599 465 -565
rect 399 -615 465 -599
rect 591 -565 657 -549
rect 591 -599 607 -565
rect 641 -599 657 -565
rect 591 -615 657 -599
rect 783 -565 849 -549
rect 783 -599 799 -565
rect 833 -599 849 -565
rect 783 -615 849 -599
<< polycont >>
rect -929 565 -895 599
rect -737 565 -703 599
rect -545 565 -511 599
rect -353 565 -319 599
rect -161 565 -127 599
rect 31 565 65 599
rect 223 565 257 599
rect 415 565 449 599
rect 607 565 641 599
rect 799 565 833 599
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -929 -599 -895 -565
rect -737 -599 -703 -565
rect -545 -599 -511 -565
rect -353 -599 -319 -565
rect -161 -599 -127 -565
rect 31 -599 65 -565
rect 223 -599 257 -565
rect 415 -599 449 -565
rect 607 -599 641 -565
rect 799 -599 833 -565
<< locali >>
rect -1091 667 -995 701
rect 995 667 1091 701
rect -1091 605 -1057 667
rect 1057 605 1091 667
rect -945 565 -929 599
rect -895 565 -879 599
rect -753 565 -737 599
rect -703 565 -687 599
rect -561 565 -545 599
rect -511 565 -495 599
rect -369 565 -353 599
rect -319 565 -303 599
rect -177 565 -161 599
rect -127 565 -111 599
rect 15 565 31 599
rect 65 565 81 599
rect 207 565 223 599
rect 257 565 273 599
rect 399 565 415 599
rect 449 565 465 599
rect 591 565 607 599
rect 641 565 657 599
rect 783 565 799 599
rect 833 565 849 599
rect -977 506 -943 522
rect -977 114 -943 130
rect -881 506 -847 522
rect -881 114 -847 130
rect -785 506 -751 522
rect -785 114 -751 130
rect -689 506 -655 522
rect -689 114 -655 130
rect -593 506 -559 522
rect -593 114 -559 130
rect -497 506 -463 522
rect -497 114 -463 130
rect -401 506 -367 522
rect -401 114 -367 130
rect -305 506 -271 522
rect -305 114 -271 130
rect -209 506 -175 522
rect -209 114 -175 130
rect -113 506 -79 522
rect -113 114 -79 130
rect -17 506 17 522
rect -17 114 17 130
rect 79 506 113 522
rect 79 114 113 130
rect 175 506 209 522
rect 175 114 209 130
rect 271 506 305 522
rect 271 114 305 130
rect 367 506 401 522
rect 367 114 401 130
rect 463 506 497 522
rect 463 114 497 130
rect 559 506 593 522
rect 559 114 593 130
rect 655 506 689 522
rect 655 114 689 130
rect 751 506 785 522
rect 751 114 785 130
rect 847 506 881 522
rect 847 114 881 130
rect 943 506 977 522
rect 943 114 977 130
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect -977 -130 -943 -114
rect -977 -522 -943 -506
rect -881 -130 -847 -114
rect -881 -522 -847 -506
rect -785 -130 -751 -114
rect -785 -522 -751 -506
rect -689 -130 -655 -114
rect -689 -522 -655 -506
rect -593 -130 -559 -114
rect -593 -522 -559 -506
rect -497 -130 -463 -114
rect -497 -522 -463 -506
rect -401 -130 -367 -114
rect -401 -522 -367 -506
rect -305 -130 -271 -114
rect -305 -522 -271 -506
rect -209 -130 -175 -114
rect -209 -522 -175 -506
rect -113 -130 -79 -114
rect -113 -522 -79 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 79 -130 113 -114
rect 79 -522 113 -506
rect 175 -130 209 -114
rect 175 -522 209 -506
rect 271 -130 305 -114
rect 271 -522 305 -506
rect 367 -130 401 -114
rect 367 -522 401 -506
rect 463 -130 497 -114
rect 463 -522 497 -506
rect 559 -130 593 -114
rect 559 -522 593 -506
rect 655 -130 689 -114
rect 655 -522 689 -506
rect 751 -130 785 -114
rect 751 -522 785 -506
rect 847 -130 881 -114
rect 847 -522 881 -506
rect 943 -130 977 -114
rect 943 -522 977 -506
rect -945 -599 -929 -565
rect -895 -599 -879 -565
rect -753 -599 -737 -565
rect -703 -599 -687 -565
rect -561 -599 -545 -565
rect -511 -599 -495 -565
rect -369 -599 -353 -565
rect -319 -599 -303 -565
rect -177 -599 -161 -565
rect -127 -599 -111 -565
rect 15 -599 31 -565
rect 65 -599 81 -565
rect 207 -599 223 -565
rect 257 -599 273 -565
rect 399 -599 415 -565
rect 449 -599 465 -565
rect 591 -599 607 -565
rect 641 -599 657 -565
rect 783 -599 799 -565
rect 833 -599 849 -565
rect -1091 -667 -1057 -605
rect 1057 -667 1091 -605
rect -1091 -701 -995 -667
rect 995 -701 1091 -667
<< viali >>
rect -929 565 -895 599
rect -737 565 -703 599
rect -545 565 -511 599
rect -353 565 -319 599
rect -161 565 -127 599
rect 31 565 65 599
rect 223 565 257 599
rect 415 565 449 599
rect 607 565 641 599
rect 799 565 833 599
rect -977 130 -943 506
rect -881 130 -847 506
rect -785 130 -751 506
rect -689 130 -655 506
rect -593 130 -559 506
rect -497 130 -463 506
rect -401 130 -367 506
rect -305 130 -271 506
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect 271 130 305 506
rect 367 130 401 506
rect 463 130 497 506
rect 559 130 593 506
rect 655 130 689 506
rect 751 130 785 506
rect 847 130 881 506
rect 943 130 977 506
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -977 -506 -943 -130
rect -881 -506 -847 -130
rect -785 -506 -751 -130
rect -689 -506 -655 -130
rect -593 -506 -559 -130
rect -497 -506 -463 -130
rect -401 -506 -367 -130
rect -305 -506 -271 -130
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect 271 -506 305 -130
rect 367 -506 401 -130
rect 463 -506 497 -130
rect 559 -506 593 -130
rect 655 -506 689 -130
rect 751 -506 785 -130
rect 847 -506 881 -130
rect 943 -506 977 -130
rect -929 -599 -895 -565
rect -737 -599 -703 -565
rect -545 -599 -511 -565
rect -353 -599 -319 -565
rect -161 -599 -127 -565
rect 31 -599 65 -565
rect 223 -599 257 -565
rect 415 -599 449 -565
rect 607 -599 641 -565
rect 799 -599 833 -565
<< metal1 >>
rect -941 599 -883 605
rect -941 565 -929 599
rect -895 565 -883 599
rect -941 559 -883 565
rect -749 599 -691 605
rect -749 565 -737 599
rect -703 565 -691 599
rect -749 559 -691 565
rect -557 599 -499 605
rect -557 565 -545 599
rect -511 565 -499 599
rect -557 559 -499 565
rect -365 599 -307 605
rect -365 565 -353 599
rect -319 565 -307 599
rect -365 559 -307 565
rect -173 599 -115 605
rect -173 565 -161 599
rect -127 565 -115 599
rect -173 559 -115 565
rect 19 599 77 605
rect 19 565 31 599
rect 65 565 77 599
rect 19 559 77 565
rect 211 599 269 605
rect 211 565 223 599
rect 257 565 269 599
rect 211 559 269 565
rect 403 599 461 605
rect 403 565 415 599
rect 449 565 461 599
rect 403 559 461 565
rect 595 599 653 605
rect 595 565 607 599
rect 641 565 653 599
rect 595 559 653 565
rect 787 599 845 605
rect 787 565 799 599
rect 833 565 845 599
rect 787 559 845 565
rect -983 506 -937 518
rect -983 130 -977 506
rect -943 130 -937 506
rect -983 118 -937 130
rect -887 506 -841 518
rect -887 130 -881 506
rect -847 130 -841 506
rect -887 118 -841 130
rect -791 506 -745 518
rect -791 130 -785 506
rect -751 130 -745 506
rect -791 118 -745 130
rect -695 506 -649 518
rect -695 130 -689 506
rect -655 130 -649 506
rect -695 118 -649 130
rect -599 506 -553 518
rect -599 130 -593 506
rect -559 130 -553 506
rect -599 118 -553 130
rect -503 506 -457 518
rect -503 130 -497 506
rect -463 130 -457 506
rect -503 118 -457 130
rect -407 506 -361 518
rect -407 130 -401 506
rect -367 130 -361 506
rect -407 118 -361 130
rect -311 506 -265 518
rect -311 130 -305 506
rect -271 130 -265 506
rect -311 118 -265 130
rect -215 506 -169 518
rect -215 130 -209 506
rect -175 130 -169 506
rect -215 118 -169 130
rect -119 506 -73 518
rect -119 130 -113 506
rect -79 130 -73 506
rect -119 118 -73 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 73 506 119 518
rect 73 130 79 506
rect 113 130 119 506
rect 73 118 119 130
rect 169 506 215 518
rect 169 130 175 506
rect 209 130 215 506
rect 169 118 215 130
rect 265 506 311 518
rect 265 130 271 506
rect 305 130 311 506
rect 265 118 311 130
rect 361 506 407 518
rect 361 130 367 506
rect 401 130 407 506
rect 361 118 407 130
rect 457 506 503 518
rect 457 130 463 506
rect 497 130 503 506
rect 457 118 503 130
rect 553 506 599 518
rect 553 130 559 506
rect 593 130 599 506
rect 553 118 599 130
rect 649 506 695 518
rect 649 130 655 506
rect 689 130 695 506
rect 649 118 695 130
rect 745 506 791 518
rect 745 130 751 506
rect 785 130 791 506
rect 745 118 791 130
rect 841 506 887 518
rect 841 130 847 506
rect 881 130 887 506
rect 841 118 887 130
rect 937 506 983 518
rect 937 130 943 506
rect 977 130 983 506
rect 937 118 983 130
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect -983 -130 -937 -118
rect -983 -506 -977 -130
rect -943 -506 -937 -130
rect -983 -518 -937 -506
rect -887 -130 -841 -118
rect -887 -506 -881 -130
rect -847 -506 -841 -130
rect -887 -518 -841 -506
rect -791 -130 -745 -118
rect -791 -506 -785 -130
rect -751 -506 -745 -130
rect -791 -518 -745 -506
rect -695 -130 -649 -118
rect -695 -506 -689 -130
rect -655 -506 -649 -130
rect -695 -518 -649 -506
rect -599 -130 -553 -118
rect -599 -506 -593 -130
rect -559 -506 -553 -130
rect -599 -518 -553 -506
rect -503 -130 -457 -118
rect -503 -506 -497 -130
rect -463 -506 -457 -130
rect -503 -518 -457 -506
rect -407 -130 -361 -118
rect -407 -506 -401 -130
rect -367 -506 -361 -130
rect -407 -518 -361 -506
rect -311 -130 -265 -118
rect -311 -506 -305 -130
rect -271 -506 -265 -130
rect -311 -518 -265 -506
rect -215 -130 -169 -118
rect -215 -506 -209 -130
rect -175 -506 -169 -130
rect -215 -518 -169 -506
rect -119 -130 -73 -118
rect -119 -506 -113 -130
rect -79 -506 -73 -130
rect -119 -518 -73 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 73 -130 119 -118
rect 73 -506 79 -130
rect 113 -506 119 -130
rect 73 -518 119 -506
rect 169 -130 215 -118
rect 169 -506 175 -130
rect 209 -506 215 -130
rect 169 -518 215 -506
rect 265 -130 311 -118
rect 265 -506 271 -130
rect 305 -506 311 -130
rect 265 -518 311 -506
rect 361 -130 407 -118
rect 361 -506 367 -130
rect 401 -506 407 -130
rect 361 -518 407 -506
rect 457 -130 503 -118
rect 457 -506 463 -130
rect 497 -506 503 -130
rect 457 -518 503 -506
rect 553 -130 599 -118
rect 553 -506 559 -130
rect 593 -506 599 -130
rect 553 -518 599 -506
rect 649 -130 695 -118
rect 649 -506 655 -130
rect 689 -506 695 -130
rect 649 -518 695 -506
rect 745 -130 791 -118
rect 745 -506 751 -130
rect 785 -506 791 -130
rect 745 -518 791 -506
rect 841 -130 887 -118
rect 841 -506 847 -130
rect 881 -506 887 -130
rect 841 -518 887 -506
rect 937 -130 983 -118
rect 937 -506 943 -130
rect 977 -506 983 -130
rect 937 -518 983 -506
rect -941 -565 -883 -559
rect -941 -599 -929 -565
rect -895 -599 -883 -565
rect -941 -605 -883 -599
rect -749 -565 -691 -559
rect -749 -599 -737 -565
rect -703 -599 -691 -565
rect -749 -605 -691 -599
rect -557 -565 -499 -559
rect -557 -599 -545 -565
rect -511 -599 -499 -565
rect -557 -605 -499 -599
rect -365 -565 -307 -559
rect -365 -599 -353 -565
rect -319 -599 -307 -565
rect -365 -605 -307 -599
rect -173 -565 -115 -559
rect -173 -599 -161 -565
rect -127 -599 -115 -565
rect -173 -605 -115 -599
rect 19 -565 77 -559
rect 19 -599 31 -565
rect 65 -599 77 -565
rect 19 -605 77 -599
rect 211 -565 269 -559
rect 211 -599 223 -565
rect 257 -599 269 -565
rect 211 -605 269 -599
rect 403 -565 461 -559
rect 403 -599 415 -565
rect 449 -599 461 -565
rect 403 -605 461 -599
rect 595 -565 653 -559
rect 595 -599 607 -565
rect 641 -599 653 -565
rect 595 -605 653 -599
rect 787 -565 845 -559
rect 787 -599 799 -565
rect 833 -599 845 -565
rect 787 -605 845 -599
<< properties >>
string FIXED_BBOX -1074 -684 1074 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 2 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
