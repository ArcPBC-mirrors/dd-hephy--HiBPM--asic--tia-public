magic
tech sky130A
magscale 1 2
timestamp 1683544843
<< metal3 >>
rect -1686 2512 1686 2540
rect -1686 -2512 1602 2512
rect 1666 -2512 1686 2512
rect -1686 -2540 1686 -2512
<< via3 >>
rect 1602 -2512 1666 2512
<< mimcap >>
rect -1646 2460 1354 2500
rect -1646 -2460 -1606 2460
rect 1314 -2460 1354 2460
rect -1646 -2500 1354 -2460
<< mimcapcontact >>
rect -1606 -2460 1314 2460
<< metal4 >>
rect 1586 2512 1682 2528
rect -1607 2460 1315 2461
rect -1607 -2460 -1606 2460
rect 1314 -2460 1315 2460
rect -1607 -2461 1315 -2460
rect 1586 -2512 1602 2512
rect 1666 -2512 1682 2512
rect 1586 -2528 1682 -2512
<< properties >>
string FIXED_BBOX -1686 -2540 1394 2540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15 l 25 val 765.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
