magic
tech sky130A
magscale 1 2
timestamp 1683564698
<< error_p >>
rect -6070 2345 -4010 2372
rect -3550 2345 -1490 2372
rect -1030 2345 1030 2372
rect 1490 2345 3550 2372
rect 4010 2345 6070 2372
rect -6070 1336 -4010 1363
rect -3550 1336 -1490 1363
rect -1030 1336 1030 1363
rect 1490 1336 3550 1363
rect 4010 1336 6070 1363
rect -6070 1109 -4010 1136
rect -3550 1109 -1490 1136
rect -1030 1109 1030 1136
rect 1490 1109 3550 1136
rect 4010 1109 6070 1136
rect -6070 100 -4010 127
rect -3550 100 -1490 127
rect -1030 100 1030 127
rect 1490 100 3550 127
rect 4010 100 6070 127
rect -6070 -127 -4010 -100
rect -3550 -127 -1490 -100
rect -1030 -127 1030 -100
rect 1490 -127 3550 -100
rect 4010 -127 6070 -100
rect -6070 -1136 -4010 -1109
rect -3550 -1136 -1490 -1109
rect -1030 -1136 1030 -1109
rect 1490 -1136 3550 -1109
rect 4010 -1136 6070 -1109
rect -6070 -1363 -4010 -1336
rect -3550 -1363 -1490 -1336
rect -1030 -1363 1030 -1336
rect 1490 -1363 3550 -1336
rect 4010 -1363 6070 -1336
rect -6070 -2372 -4010 -2345
rect -3550 -2372 -1490 -2345
rect -1030 -2372 1030 -2345
rect 1490 -2372 3550 -2345
rect 4010 -2372 6070 -2345
<< nwell >>
rect -6173 1363 -3907 2345
rect -3653 1363 -1387 2345
rect -1133 1363 1133 2345
rect 1387 1363 3653 2345
rect 3907 1363 6173 2345
rect -6173 127 -3907 1109
rect -3653 127 -1387 1109
rect -1133 127 1133 1109
rect 1387 127 3653 1109
rect 3907 127 6173 1109
rect -6173 -1109 -3907 -127
rect -3653 -1109 -1387 -127
rect -1133 -1109 1133 -127
rect 1387 -1109 3653 -127
rect 3907 -1109 6173 -127
rect -6173 -2345 -3907 -1363
rect -3653 -2345 -1387 -1363
rect -1133 -2345 1133 -1363
rect 1387 -2345 3653 -1363
rect 3907 -2345 6173 -1363
<< pwell >>
rect -6283 2345 6283 2455
rect -6283 1363 -6173 2345
rect -3907 1363 -3653 2345
rect -1387 1363 -1133 2345
rect 1133 1363 1387 2345
rect 3653 1363 3907 2345
rect 6173 1363 6283 2345
rect -6283 1109 6283 1363
rect -6283 127 -6173 1109
rect -3907 127 -3653 1109
rect -1387 127 -1133 1109
rect 1133 127 1387 1109
rect 3653 127 3907 1109
rect 6173 127 6283 1109
rect -6283 -127 6283 127
rect -6283 -1109 -6173 -127
rect -3907 -1109 -3653 -127
rect -1387 -1109 -1133 -127
rect 1133 -1109 1387 -127
rect 3653 -1109 3907 -127
rect 6173 -1109 6283 -127
rect -6283 -1363 6283 -1109
rect -6283 -2345 -6173 -1363
rect -3907 -2345 -3653 -1363
rect -1387 -2345 -1133 -1363
rect 1133 -2345 1387 -1363
rect 3653 -2345 3907 -1363
rect 6173 -2345 6283 -1363
rect -6283 -2455 6283 -2345
<< varactor >>
rect -6040 1454 -4040 2254
rect -3520 1454 -1520 2254
rect -1000 1454 1000 2254
rect 1520 1454 3520 2254
rect 4040 1454 6040 2254
rect -6040 218 -4040 1018
rect -3520 218 -1520 1018
rect -1000 218 1000 1018
rect 1520 218 3520 1018
rect 4040 218 6040 1018
rect -6040 -1018 -4040 -218
rect -3520 -1018 -1520 -218
rect -1000 -1018 1000 -218
rect 1520 -1018 3520 -218
rect 4040 -1018 6040 -218
rect -6040 -2254 -4040 -1454
rect -3520 -2254 -1520 -1454
rect -1000 -2254 1000 -1454
rect 1520 -2254 3520 -1454
rect 4040 -2254 6040 -1454
<< psubdiff >>
rect -6247 2385 -6151 2419
rect 6151 2385 6247 2419
rect -6247 2323 -6213 2385
rect 6213 2323 6247 2385
rect -6247 -2385 -6213 -2323
rect 6213 -2385 6247 -2323
rect -6247 -2419 -6151 -2385
rect 6151 -2419 6247 -2385
<< nsubdiff >>
rect -6137 2230 -6040 2254
rect -6137 1478 -6125 2230
rect -6091 1478 -6040 2230
rect -6137 1454 -6040 1478
rect -4040 2230 -3943 2254
rect -4040 1478 -3989 2230
rect -3955 1478 -3943 2230
rect -4040 1454 -3943 1478
rect -3617 2230 -3520 2254
rect -3617 1478 -3605 2230
rect -3571 1478 -3520 2230
rect -3617 1454 -3520 1478
rect -1520 2230 -1423 2254
rect -1520 1478 -1469 2230
rect -1435 1478 -1423 2230
rect -1520 1454 -1423 1478
rect -1097 2230 -1000 2254
rect -1097 1478 -1085 2230
rect -1051 1478 -1000 2230
rect -1097 1454 -1000 1478
rect 1000 2230 1097 2254
rect 1000 1478 1051 2230
rect 1085 1478 1097 2230
rect 1000 1454 1097 1478
rect 1423 2230 1520 2254
rect 1423 1478 1435 2230
rect 1469 1478 1520 2230
rect 1423 1454 1520 1478
rect 3520 2230 3617 2254
rect 3520 1478 3571 2230
rect 3605 1478 3617 2230
rect 3520 1454 3617 1478
rect 3943 2230 4040 2254
rect 3943 1478 3955 2230
rect 3989 1478 4040 2230
rect 3943 1454 4040 1478
rect 6040 2230 6137 2254
rect 6040 1478 6091 2230
rect 6125 1478 6137 2230
rect 6040 1454 6137 1478
rect -6137 994 -6040 1018
rect -6137 242 -6125 994
rect -6091 242 -6040 994
rect -6137 218 -6040 242
rect -4040 994 -3943 1018
rect -4040 242 -3989 994
rect -3955 242 -3943 994
rect -4040 218 -3943 242
rect -3617 994 -3520 1018
rect -3617 242 -3605 994
rect -3571 242 -3520 994
rect -3617 218 -3520 242
rect -1520 994 -1423 1018
rect -1520 242 -1469 994
rect -1435 242 -1423 994
rect -1520 218 -1423 242
rect -1097 994 -1000 1018
rect -1097 242 -1085 994
rect -1051 242 -1000 994
rect -1097 218 -1000 242
rect 1000 994 1097 1018
rect 1000 242 1051 994
rect 1085 242 1097 994
rect 1000 218 1097 242
rect 1423 994 1520 1018
rect 1423 242 1435 994
rect 1469 242 1520 994
rect 1423 218 1520 242
rect 3520 994 3617 1018
rect 3520 242 3571 994
rect 3605 242 3617 994
rect 3520 218 3617 242
rect 3943 994 4040 1018
rect 3943 242 3955 994
rect 3989 242 4040 994
rect 3943 218 4040 242
rect 6040 994 6137 1018
rect 6040 242 6091 994
rect 6125 242 6137 994
rect 6040 218 6137 242
rect -6137 -242 -6040 -218
rect -6137 -994 -6125 -242
rect -6091 -994 -6040 -242
rect -6137 -1018 -6040 -994
rect -4040 -242 -3943 -218
rect -4040 -994 -3989 -242
rect -3955 -994 -3943 -242
rect -4040 -1018 -3943 -994
rect -3617 -242 -3520 -218
rect -3617 -994 -3605 -242
rect -3571 -994 -3520 -242
rect -3617 -1018 -3520 -994
rect -1520 -242 -1423 -218
rect -1520 -994 -1469 -242
rect -1435 -994 -1423 -242
rect -1520 -1018 -1423 -994
rect -1097 -242 -1000 -218
rect -1097 -994 -1085 -242
rect -1051 -994 -1000 -242
rect -1097 -1018 -1000 -994
rect 1000 -242 1097 -218
rect 1000 -994 1051 -242
rect 1085 -994 1097 -242
rect 1000 -1018 1097 -994
rect 1423 -242 1520 -218
rect 1423 -994 1435 -242
rect 1469 -994 1520 -242
rect 1423 -1018 1520 -994
rect 3520 -242 3617 -218
rect 3520 -994 3571 -242
rect 3605 -994 3617 -242
rect 3520 -1018 3617 -994
rect 3943 -242 4040 -218
rect 3943 -994 3955 -242
rect 3989 -994 4040 -242
rect 3943 -1018 4040 -994
rect 6040 -242 6137 -218
rect 6040 -994 6091 -242
rect 6125 -994 6137 -242
rect 6040 -1018 6137 -994
rect -6137 -1478 -6040 -1454
rect -6137 -2230 -6125 -1478
rect -6091 -2230 -6040 -1478
rect -6137 -2254 -6040 -2230
rect -4040 -1478 -3943 -1454
rect -4040 -2230 -3989 -1478
rect -3955 -2230 -3943 -1478
rect -4040 -2254 -3943 -2230
rect -3617 -1478 -3520 -1454
rect -3617 -2230 -3605 -1478
rect -3571 -2230 -3520 -1478
rect -3617 -2254 -3520 -2230
rect -1520 -1478 -1423 -1454
rect -1520 -2230 -1469 -1478
rect -1435 -2230 -1423 -1478
rect -1520 -2254 -1423 -2230
rect -1097 -1478 -1000 -1454
rect -1097 -2230 -1085 -1478
rect -1051 -2230 -1000 -1478
rect -1097 -2254 -1000 -2230
rect 1000 -1478 1097 -1454
rect 1000 -2230 1051 -1478
rect 1085 -2230 1097 -1478
rect 1000 -2254 1097 -2230
rect 1423 -1478 1520 -1454
rect 1423 -2230 1435 -1478
rect 1469 -2230 1520 -1478
rect 1423 -2254 1520 -2230
rect 3520 -1478 3617 -1454
rect 3520 -2230 3571 -1478
rect 3605 -2230 3617 -1478
rect 3520 -2254 3617 -2230
rect 3943 -1478 4040 -1454
rect 3943 -2230 3955 -1478
rect 3989 -2230 4040 -1478
rect 3943 -2254 4040 -2230
rect 6040 -1478 6137 -1454
rect 6040 -2230 6091 -1478
rect 6125 -2230 6137 -1478
rect 6040 -2254 6137 -2230
<< psubdiffcont >>
rect -6151 2385 6151 2419
rect -6247 -2323 -6213 2323
rect 6213 -2323 6247 2323
rect -6151 -2419 6151 -2385
<< nsubdiffcont >>
rect -6125 1478 -6091 2230
rect -3989 1478 -3955 2230
rect -3605 1478 -3571 2230
rect -1469 1478 -1435 2230
rect -1085 1478 -1051 2230
rect 1051 1478 1085 2230
rect 1435 1478 1469 2230
rect 3571 1478 3605 2230
rect 3955 1478 3989 2230
rect 6091 1478 6125 2230
rect -6125 242 -6091 994
rect -3989 242 -3955 994
rect -3605 242 -3571 994
rect -1469 242 -1435 994
rect -1085 242 -1051 994
rect 1051 242 1085 994
rect 1435 242 1469 994
rect 3571 242 3605 994
rect 3955 242 3989 994
rect 6091 242 6125 994
rect -6125 -994 -6091 -242
rect -3989 -994 -3955 -242
rect -3605 -994 -3571 -242
rect -1469 -994 -1435 -242
rect -1085 -994 -1051 -242
rect 1051 -994 1085 -242
rect 1435 -994 1469 -242
rect 3571 -994 3605 -242
rect 3955 -994 3989 -242
rect 6091 -994 6125 -242
rect -6125 -2230 -6091 -1478
rect -3989 -2230 -3955 -1478
rect -3605 -2230 -3571 -1478
rect -1469 -2230 -1435 -1478
rect -1085 -2230 -1051 -1478
rect 1051 -2230 1085 -1478
rect 1435 -2230 1469 -1478
rect 3571 -2230 3605 -1478
rect 3955 -2230 3989 -1478
rect 6091 -2230 6125 -1478
<< poly >>
rect -6040 2326 -4040 2342
rect -6040 2292 -6024 2326
rect -4056 2292 -4040 2326
rect -6040 2254 -4040 2292
rect -3520 2326 -1520 2342
rect -3520 2292 -3504 2326
rect -1536 2292 -1520 2326
rect -3520 2254 -1520 2292
rect -1000 2326 1000 2342
rect -1000 2292 -984 2326
rect 984 2292 1000 2326
rect -1000 2254 1000 2292
rect 1520 2326 3520 2342
rect 1520 2292 1536 2326
rect 3504 2292 3520 2326
rect 1520 2254 3520 2292
rect 4040 2326 6040 2342
rect 4040 2292 4056 2326
rect 6024 2292 6040 2326
rect 4040 2254 6040 2292
rect -6040 1416 -4040 1454
rect -6040 1382 -6024 1416
rect -4056 1382 -4040 1416
rect -6040 1366 -4040 1382
rect -3520 1416 -1520 1454
rect -3520 1382 -3504 1416
rect -1536 1382 -1520 1416
rect -3520 1366 -1520 1382
rect -1000 1416 1000 1454
rect -1000 1382 -984 1416
rect 984 1382 1000 1416
rect -1000 1366 1000 1382
rect 1520 1416 3520 1454
rect 1520 1382 1536 1416
rect 3504 1382 3520 1416
rect 1520 1366 3520 1382
rect 4040 1416 6040 1454
rect 4040 1382 4056 1416
rect 6024 1382 6040 1416
rect 4040 1366 6040 1382
rect -6040 1090 -4040 1106
rect -6040 1056 -6024 1090
rect -4056 1056 -4040 1090
rect -6040 1018 -4040 1056
rect -3520 1090 -1520 1106
rect -3520 1056 -3504 1090
rect -1536 1056 -1520 1090
rect -3520 1018 -1520 1056
rect -1000 1090 1000 1106
rect -1000 1056 -984 1090
rect 984 1056 1000 1090
rect -1000 1018 1000 1056
rect 1520 1090 3520 1106
rect 1520 1056 1536 1090
rect 3504 1056 3520 1090
rect 1520 1018 3520 1056
rect 4040 1090 6040 1106
rect 4040 1056 4056 1090
rect 6024 1056 6040 1090
rect 4040 1018 6040 1056
rect -6040 180 -4040 218
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -6040 130 -4040 146
rect -3520 180 -1520 218
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -3520 130 -1520 146
rect -1000 180 1000 218
rect -1000 146 -984 180
rect 984 146 1000 180
rect -1000 130 1000 146
rect 1520 180 3520 218
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 1520 130 3520 146
rect 4040 180 6040 218
rect 4040 146 4056 180
rect 6024 146 6040 180
rect 4040 130 6040 146
rect -6040 -146 -4040 -130
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -6040 -218 -4040 -180
rect -3520 -146 -1520 -130
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -3520 -218 -1520 -180
rect -1000 -146 1000 -130
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect -1000 -218 1000 -180
rect 1520 -146 3520 -130
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 1520 -218 3520 -180
rect 4040 -146 6040 -130
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect 4040 -218 6040 -180
rect -6040 -1056 -4040 -1018
rect -6040 -1090 -6024 -1056
rect -4056 -1090 -4040 -1056
rect -6040 -1106 -4040 -1090
rect -3520 -1056 -1520 -1018
rect -3520 -1090 -3504 -1056
rect -1536 -1090 -1520 -1056
rect -3520 -1106 -1520 -1090
rect -1000 -1056 1000 -1018
rect -1000 -1090 -984 -1056
rect 984 -1090 1000 -1056
rect -1000 -1106 1000 -1090
rect 1520 -1056 3520 -1018
rect 1520 -1090 1536 -1056
rect 3504 -1090 3520 -1056
rect 1520 -1106 3520 -1090
rect 4040 -1056 6040 -1018
rect 4040 -1090 4056 -1056
rect 6024 -1090 6040 -1056
rect 4040 -1106 6040 -1090
rect -6040 -1382 -4040 -1366
rect -6040 -1416 -6024 -1382
rect -4056 -1416 -4040 -1382
rect -6040 -1454 -4040 -1416
rect -3520 -1382 -1520 -1366
rect -3520 -1416 -3504 -1382
rect -1536 -1416 -1520 -1382
rect -3520 -1454 -1520 -1416
rect -1000 -1382 1000 -1366
rect -1000 -1416 -984 -1382
rect 984 -1416 1000 -1382
rect -1000 -1454 1000 -1416
rect 1520 -1382 3520 -1366
rect 1520 -1416 1536 -1382
rect 3504 -1416 3520 -1382
rect 1520 -1454 3520 -1416
rect 4040 -1382 6040 -1366
rect 4040 -1416 4056 -1382
rect 6024 -1416 6040 -1382
rect 4040 -1454 6040 -1416
rect -6040 -2292 -4040 -2254
rect -6040 -2326 -6024 -2292
rect -4056 -2326 -4040 -2292
rect -6040 -2342 -4040 -2326
rect -3520 -2292 -1520 -2254
rect -3520 -2326 -3504 -2292
rect -1536 -2326 -1520 -2292
rect -3520 -2342 -1520 -2326
rect -1000 -2292 1000 -2254
rect -1000 -2326 -984 -2292
rect 984 -2326 1000 -2292
rect -1000 -2342 1000 -2326
rect 1520 -2292 3520 -2254
rect 1520 -2326 1536 -2292
rect 3504 -2326 3520 -2292
rect 1520 -2342 3520 -2326
rect 4040 -2292 6040 -2254
rect 4040 -2326 4056 -2292
rect 6024 -2326 6040 -2292
rect 4040 -2342 6040 -2326
<< polycont >>
rect -6024 2292 -4056 2326
rect -3504 2292 -1536 2326
rect -984 2292 984 2326
rect 1536 2292 3504 2326
rect 4056 2292 6024 2326
rect -6024 1382 -4056 1416
rect -3504 1382 -1536 1416
rect -984 1382 984 1416
rect 1536 1382 3504 1416
rect 4056 1382 6024 1416
rect -6024 1056 -4056 1090
rect -3504 1056 -1536 1090
rect -984 1056 984 1090
rect 1536 1056 3504 1090
rect 4056 1056 6024 1090
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6024 -1090 -4056 -1056
rect -3504 -1090 -1536 -1056
rect -984 -1090 984 -1056
rect 1536 -1090 3504 -1056
rect 4056 -1090 6024 -1056
rect -6024 -1416 -4056 -1382
rect -3504 -1416 -1536 -1382
rect -984 -1416 984 -1382
rect 1536 -1416 3504 -1382
rect 4056 -1416 6024 -1382
rect -6024 -2326 -4056 -2292
rect -3504 -2326 -1536 -2292
rect -984 -2326 984 -2292
rect 1536 -2326 3504 -2292
rect 4056 -2326 6024 -2292
<< locali >>
rect -6247 2385 -6151 2419
rect 6151 2385 6247 2419
rect -6247 2323 -6213 2385
rect -6040 2292 -6024 2326
rect -4056 2292 -4040 2326
rect -3520 2292 -3504 2326
rect -1536 2292 -1520 2326
rect -1000 2292 -984 2326
rect 984 2292 1000 2326
rect 1520 2292 1536 2326
rect 3504 2292 3520 2326
rect 4040 2292 4056 2326
rect 6024 2292 6040 2326
rect 6213 2323 6247 2385
rect -6125 2230 -6091 2246
rect -6125 1462 -6091 1478
rect -3989 2230 -3955 2246
rect -3989 1462 -3955 1478
rect -3605 2230 -3571 2246
rect -3605 1462 -3571 1478
rect -1469 2230 -1435 2246
rect -1469 1462 -1435 1478
rect -1085 2230 -1051 2246
rect -1085 1462 -1051 1478
rect 1051 2230 1085 2246
rect 1051 1462 1085 1478
rect 1435 2230 1469 2246
rect 1435 1462 1469 1478
rect 3571 2230 3605 2246
rect 3571 1462 3605 1478
rect 3955 2230 3989 2246
rect 3955 1462 3989 1478
rect 6091 2230 6125 2246
rect 6091 1462 6125 1478
rect -6040 1382 -6024 1416
rect -4056 1382 -4040 1416
rect -3520 1382 -3504 1416
rect -1536 1382 -1520 1416
rect -1000 1382 -984 1416
rect 984 1382 1000 1416
rect 1520 1382 1536 1416
rect 3504 1382 3520 1416
rect 4040 1382 4056 1416
rect 6024 1382 6040 1416
rect -6040 1056 -6024 1090
rect -4056 1056 -4040 1090
rect -3520 1056 -3504 1090
rect -1536 1056 -1520 1090
rect -1000 1056 -984 1090
rect 984 1056 1000 1090
rect 1520 1056 1536 1090
rect 3504 1056 3520 1090
rect 4040 1056 4056 1090
rect 6024 1056 6040 1090
rect -6125 994 -6091 1010
rect -6125 226 -6091 242
rect -3989 994 -3955 1010
rect -3989 226 -3955 242
rect -3605 994 -3571 1010
rect -3605 226 -3571 242
rect -1469 994 -1435 1010
rect -1469 226 -1435 242
rect -1085 994 -1051 1010
rect -1085 226 -1051 242
rect 1051 994 1085 1010
rect 1051 226 1085 242
rect 1435 994 1469 1010
rect 1435 226 1469 242
rect 3571 994 3605 1010
rect 3571 226 3605 242
rect 3955 994 3989 1010
rect 3955 226 3989 242
rect 6091 994 6125 1010
rect 6091 226 6125 242
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -1000 146 -984 180
rect 984 146 1000 180
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 4040 146 4056 180
rect 6024 146 6040 180
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect -6125 -242 -6091 -226
rect -6125 -1010 -6091 -994
rect -3989 -242 -3955 -226
rect -3989 -1010 -3955 -994
rect -3605 -242 -3571 -226
rect -3605 -1010 -3571 -994
rect -1469 -242 -1435 -226
rect -1469 -1010 -1435 -994
rect -1085 -242 -1051 -226
rect -1085 -1010 -1051 -994
rect 1051 -242 1085 -226
rect 1051 -1010 1085 -994
rect 1435 -242 1469 -226
rect 1435 -1010 1469 -994
rect 3571 -242 3605 -226
rect 3571 -1010 3605 -994
rect 3955 -242 3989 -226
rect 3955 -1010 3989 -994
rect 6091 -242 6125 -226
rect 6091 -1010 6125 -994
rect -6040 -1090 -6024 -1056
rect -4056 -1090 -4040 -1056
rect -3520 -1090 -3504 -1056
rect -1536 -1090 -1520 -1056
rect -1000 -1090 -984 -1056
rect 984 -1090 1000 -1056
rect 1520 -1090 1536 -1056
rect 3504 -1090 3520 -1056
rect 4040 -1090 4056 -1056
rect 6024 -1090 6040 -1056
rect -6040 -1416 -6024 -1382
rect -4056 -1416 -4040 -1382
rect -3520 -1416 -3504 -1382
rect -1536 -1416 -1520 -1382
rect -1000 -1416 -984 -1382
rect 984 -1416 1000 -1382
rect 1520 -1416 1536 -1382
rect 3504 -1416 3520 -1382
rect 4040 -1416 4056 -1382
rect 6024 -1416 6040 -1382
rect -6125 -1478 -6091 -1462
rect -6125 -2246 -6091 -2230
rect -3989 -1478 -3955 -1462
rect -3989 -2246 -3955 -2230
rect -3605 -1478 -3571 -1462
rect -3605 -2246 -3571 -2230
rect -1469 -1478 -1435 -1462
rect -1469 -2246 -1435 -2230
rect -1085 -1478 -1051 -1462
rect -1085 -2246 -1051 -2230
rect 1051 -1478 1085 -1462
rect 1051 -2246 1085 -2230
rect 1435 -1478 1469 -1462
rect 1435 -2246 1469 -2230
rect 3571 -1478 3605 -1462
rect 3571 -2246 3605 -2230
rect 3955 -1478 3989 -1462
rect 3955 -2246 3989 -2230
rect 6091 -1478 6125 -1462
rect 6091 -2246 6125 -2230
rect -6247 -2385 -6213 -2323
rect -6040 -2326 -6024 -2292
rect -4056 -2326 -4040 -2292
rect -3520 -2326 -3504 -2292
rect -1536 -2326 -1520 -2292
rect -1000 -2326 -984 -2292
rect 984 -2326 1000 -2292
rect 1520 -2326 1536 -2292
rect 3504 -2326 3520 -2292
rect 4040 -2326 4056 -2292
rect 6024 -2326 6040 -2292
rect 6213 -2385 6247 -2323
rect -6247 -2419 -6151 -2385
rect 6151 -2419 6247 -2385
<< viali >>
rect -6024 2292 -4056 2326
rect -3504 2292 -1536 2326
rect -984 2292 984 2326
rect 1536 2292 3504 2326
rect 4056 2292 6024 2326
rect -6125 1478 -6091 2230
rect -3989 1478 -3955 2230
rect -3605 1478 -3571 2230
rect -1469 1478 -1435 2230
rect -1085 1478 -1051 2230
rect 1051 1478 1085 2230
rect 1435 1478 1469 2230
rect 3571 1478 3605 2230
rect 3955 1478 3989 2230
rect 6091 1478 6125 2230
rect -6024 1382 -4056 1416
rect -3504 1382 -1536 1416
rect -984 1382 984 1416
rect 1536 1382 3504 1416
rect 4056 1382 6024 1416
rect -6024 1056 -4056 1090
rect -3504 1056 -1536 1090
rect -984 1056 984 1090
rect 1536 1056 3504 1090
rect 4056 1056 6024 1090
rect -6125 242 -6091 994
rect -3989 242 -3955 994
rect -3605 242 -3571 994
rect -1469 242 -1435 994
rect -1085 242 -1051 994
rect 1051 242 1085 994
rect 1435 242 1469 994
rect 3571 242 3605 994
rect 3955 242 3989 994
rect 6091 242 6125 994
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6125 -994 -6091 -242
rect -3989 -994 -3955 -242
rect -3605 -994 -3571 -242
rect -1469 -994 -1435 -242
rect -1085 -994 -1051 -242
rect 1051 -994 1085 -242
rect 1435 -994 1469 -242
rect 3571 -994 3605 -242
rect 3955 -994 3989 -242
rect 6091 -994 6125 -242
rect -6024 -1090 -4056 -1056
rect -3504 -1090 -1536 -1056
rect -984 -1090 984 -1056
rect 1536 -1090 3504 -1056
rect 4056 -1090 6024 -1056
rect -6024 -1416 -4056 -1382
rect -3504 -1416 -1536 -1382
rect -984 -1416 984 -1382
rect 1536 -1416 3504 -1382
rect 4056 -1416 6024 -1382
rect -6125 -2230 -6091 -1478
rect -3989 -2230 -3955 -1478
rect -3605 -2230 -3571 -1478
rect -1469 -2230 -1435 -1478
rect -1085 -2230 -1051 -1478
rect 1051 -2230 1085 -1478
rect 1435 -2230 1469 -1478
rect 3571 -2230 3605 -1478
rect 3955 -2230 3989 -1478
rect 6091 -2230 6125 -1478
rect -6024 -2326 -4056 -2292
rect -3504 -2326 -1536 -2292
rect -984 -2326 984 -2292
rect 1536 -2326 3504 -2292
rect 4056 -2326 6024 -2292
<< metal1 >>
rect -6036 2326 -4044 2332
rect -6036 2292 -6024 2326
rect -4056 2292 -4044 2326
rect -6036 2286 -4044 2292
rect -3516 2326 -1524 2332
rect -3516 2292 -3504 2326
rect -1536 2292 -1524 2326
rect -3516 2286 -1524 2292
rect -996 2326 996 2332
rect -996 2292 -984 2326
rect 984 2292 996 2326
rect -996 2286 996 2292
rect 1524 2326 3516 2332
rect 1524 2292 1536 2326
rect 3504 2292 3516 2326
rect 1524 2286 3516 2292
rect 4044 2326 6036 2332
rect 4044 2292 4056 2326
rect 6024 2292 6036 2326
rect 4044 2286 6036 2292
rect -6131 2230 -6085 2242
rect -3995 2230 -3949 2242
rect -6131 1478 -6125 2230
rect -6091 1478 -3989 2230
rect -3955 1478 -3949 2230
rect -6131 1466 -6085 1478
rect -3995 1466 -3949 1478
rect -3611 2230 -3565 2242
rect -1475 2230 -1429 2242
rect -3611 1478 -3605 2230
rect -3571 1478 -1469 2230
rect -1435 1478 -1429 2230
rect -3611 1466 -3565 1478
rect -1475 1466 -1429 1478
rect -1091 2230 -1045 2242
rect 1045 2230 1091 2242
rect -1091 1478 -1085 2230
rect -1051 1478 1051 2230
rect 1085 1478 1091 2230
rect -1091 1466 -1045 1478
rect 1045 1466 1091 1478
rect 1429 2230 1475 2242
rect 3565 2230 3611 2242
rect 1429 1478 1435 2230
rect 1469 1478 3571 2230
rect 3605 1478 3611 2230
rect 1429 1466 1475 1478
rect 3565 1466 3611 1478
rect 3949 2230 3995 2242
rect 6085 2230 6131 2242
rect 3949 1478 3955 2230
rect 3989 1478 6091 2230
rect 6125 1478 6131 2230
rect 3949 1466 3995 1478
rect 6085 1466 6131 1478
rect -6036 1416 -4044 1422
rect -6036 1382 -6024 1416
rect -4056 1382 -4044 1416
rect -6036 1376 -4044 1382
rect -3516 1416 -1524 1422
rect -3516 1382 -3504 1416
rect -1536 1382 -1524 1416
rect -3516 1376 -1524 1382
rect -996 1416 996 1422
rect -996 1382 -984 1416
rect 984 1382 996 1416
rect -996 1376 996 1382
rect 1524 1416 3516 1422
rect 1524 1382 1536 1416
rect 3504 1382 3516 1416
rect 1524 1376 3516 1382
rect 4044 1416 6036 1422
rect 4044 1382 4056 1416
rect 6024 1382 6036 1416
rect 4044 1376 6036 1382
rect -6036 1090 -4044 1096
rect -6036 1056 -6024 1090
rect -4056 1056 -4044 1090
rect -6036 1050 -4044 1056
rect -3516 1090 -1524 1096
rect -3516 1056 -3504 1090
rect -1536 1056 -1524 1090
rect -3516 1050 -1524 1056
rect -996 1090 996 1096
rect -996 1056 -984 1090
rect 984 1056 996 1090
rect -996 1050 996 1056
rect 1524 1090 3516 1096
rect 1524 1056 1536 1090
rect 3504 1056 3516 1090
rect 1524 1050 3516 1056
rect 4044 1090 6036 1096
rect 4044 1056 4056 1090
rect 6024 1056 6036 1090
rect 4044 1050 6036 1056
rect -6131 994 -6085 1006
rect -3995 994 -3949 1006
rect -6131 242 -6125 994
rect -6091 242 -3989 994
rect -3955 242 -3949 994
rect -6131 230 -6085 242
rect -3995 230 -3949 242
rect -3611 994 -3565 1006
rect -1475 994 -1429 1006
rect -3611 242 -3605 994
rect -3571 242 -1469 994
rect -1435 242 -1429 994
rect -3611 230 -3565 242
rect -1475 230 -1429 242
rect -1091 994 -1045 1006
rect 1045 994 1091 1006
rect -1091 242 -1085 994
rect -1051 242 1051 994
rect 1085 242 1091 994
rect -1091 230 -1045 242
rect 1045 230 1091 242
rect 1429 994 1475 1006
rect 3565 994 3611 1006
rect 1429 242 1435 994
rect 1469 242 3571 994
rect 3605 242 3611 994
rect 1429 230 1475 242
rect 3565 230 3611 242
rect 3949 994 3995 1006
rect 6085 994 6131 1006
rect 3949 242 3955 994
rect 3989 242 6091 994
rect 6125 242 6131 994
rect 3949 230 3995 242
rect 6085 230 6131 242
rect -6036 180 -4044 186
rect -6036 146 -6024 180
rect -4056 146 -4044 180
rect -6036 140 -4044 146
rect -3516 180 -1524 186
rect -3516 146 -3504 180
rect -1536 146 -1524 180
rect -3516 140 -1524 146
rect -996 180 996 186
rect -996 146 -984 180
rect 984 146 996 180
rect -996 140 996 146
rect 1524 180 3516 186
rect 1524 146 1536 180
rect 3504 146 3516 180
rect 1524 140 3516 146
rect 4044 180 6036 186
rect 4044 146 4056 180
rect 6024 146 6036 180
rect 4044 140 6036 146
rect -6036 -146 -4044 -140
rect -6036 -180 -6024 -146
rect -4056 -180 -4044 -146
rect -6036 -186 -4044 -180
rect -3516 -146 -1524 -140
rect -3516 -180 -3504 -146
rect -1536 -180 -1524 -146
rect -3516 -186 -1524 -180
rect -996 -146 996 -140
rect -996 -180 -984 -146
rect 984 -180 996 -146
rect -996 -186 996 -180
rect 1524 -146 3516 -140
rect 1524 -180 1536 -146
rect 3504 -180 3516 -146
rect 1524 -186 3516 -180
rect 4044 -146 6036 -140
rect 4044 -180 4056 -146
rect 6024 -180 6036 -146
rect 4044 -186 6036 -180
rect -6131 -242 -6085 -230
rect -3995 -242 -3949 -230
rect -6131 -994 -6125 -242
rect -6091 -994 -3989 -242
rect -3955 -994 -3949 -242
rect -6131 -1006 -6085 -994
rect -3995 -1006 -3949 -994
rect -3611 -242 -3565 -230
rect -1475 -242 -1429 -230
rect -3611 -994 -3605 -242
rect -3571 -994 -1469 -242
rect -1435 -994 -1429 -242
rect -3611 -1006 -3565 -994
rect -1475 -1006 -1429 -994
rect -1091 -242 -1045 -230
rect 1045 -242 1091 -230
rect -1091 -994 -1085 -242
rect -1051 -994 1051 -242
rect 1085 -994 1091 -242
rect -1091 -1006 -1045 -994
rect 1045 -1006 1091 -994
rect 1429 -242 1475 -230
rect 3565 -242 3611 -230
rect 1429 -994 1435 -242
rect 1469 -994 3571 -242
rect 3605 -994 3611 -242
rect 1429 -1006 1475 -994
rect 3565 -1006 3611 -994
rect 3949 -242 3995 -230
rect 6085 -242 6131 -230
rect 3949 -994 3955 -242
rect 3989 -994 6091 -242
rect 6125 -994 6131 -242
rect 3949 -1006 3995 -994
rect 6085 -1006 6131 -994
rect -6036 -1056 -4044 -1050
rect -6036 -1090 -6024 -1056
rect -4056 -1090 -4044 -1056
rect -6036 -1096 -4044 -1090
rect -3516 -1056 -1524 -1050
rect -3516 -1090 -3504 -1056
rect -1536 -1090 -1524 -1056
rect -3516 -1096 -1524 -1090
rect -996 -1056 996 -1050
rect -996 -1090 -984 -1056
rect 984 -1090 996 -1056
rect -996 -1096 996 -1090
rect 1524 -1056 3516 -1050
rect 1524 -1090 1536 -1056
rect 3504 -1090 3516 -1056
rect 1524 -1096 3516 -1090
rect 4044 -1056 6036 -1050
rect 4044 -1090 4056 -1056
rect 6024 -1090 6036 -1056
rect 4044 -1096 6036 -1090
rect -6036 -1382 -4044 -1376
rect -6036 -1416 -6024 -1382
rect -4056 -1416 -4044 -1382
rect -6036 -1422 -4044 -1416
rect -3516 -1382 -1524 -1376
rect -3516 -1416 -3504 -1382
rect -1536 -1416 -1524 -1382
rect -3516 -1422 -1524 -1416
rect -996 -1382 996 -1376
rect -996 -1416 -984 -1382
rect 984 -1416 996 -1382
rect -996 -1422 996 -1416
rect 1524 -1382 3516 -1376
rect 1524 -1416 1536 -1382
rect 3504 -1416 3516 -1382
rect 1524 -1422 3516 -1416
rect 4044 -1382 6036 -1376
rect 4044 -1416 4056 -1382
rect 6024 -1416 6036 -1382
rect 4044 -1422 6036 -1416
rect -6131 -1478 -6085 -1466
rect -3995 -1478 -3949 -1466
rect -6131 -2230 -6125 -1478
rect -6091 -2230 -3989 -1478
rect -3955 -2230 -3949 -1478
rect -6131 -2242 -6085 -2230
rect -3995 -2242 -3949 -2230
rect -3611 -1478 -3565 -1466
rect -1475 -1478 -1429 -1466
rect -3611 -2230 -3605 -1478
rect -3571 -2230 -1469 -1478
rect -1435 -2230 -1429 -1478
rect -3611 -2242 -3565 -2230
rect -1475 -2242 -1429 -2230
rect -1091 -1478 -1045 -1466
rect 1045 -1478 1091 -1466
rect -1091 -2230 -1085 -1478
rect -1051 -2230 1051 -1478
rect 1085 -2230 1091 -1478
rect -1091 -2242 -1045 -2230
rect 1045 -2242 1091 -2230
rect 1429 -1478 1475 -1466
rect 3565 -1478 3611 -1466
rect 1429 -2230 1435 -1478
rect 1469 -2230 3571 -1478
rect 3605 -2230 3611 -1478
rect 1429 -2242 1475 -2230
rect 3565 -2242 3611 -2230
rect 3949 -1478 3995 -1466
rect 6085 -1478 6131 -1466
rect 3949 -2230 3955 -1478
rect 3989 -2230 6091 -1478
rect 6125 -2230 6131 -1478
rect 3949 -2242 3995 -2230
rect 6085 -2242 6131 -2230
rect -6036 -2292 -4044 -2286
rect -6036 -2326 -6024 -2292
rect -4056 -2326 -4044 -2292
rect -6036 -2332 -4044 -2326
rect -3516 -2292 -1524 -2286
rect -3516 -2326 -3504 -2292
rect -1536 -2326 -1524 -2292
rect -3516 -2332 -1524 -2326
rect -996 -2292 996 -2286
rect -996 -2326 -984 -2292
rect 984 -2326 996 -2292
rect -996 -2332 996 -2326
rect 1524 -2292 3516 -2286
rect 1524 -2326 1536 -2292
rect 3504 -2326 3516 -2292
rect 1524 -2332 3516 -2326
rect 4044 -2292 6036 -2286
rect 4044 -2326 4056 -2292
rect 6024 -2326 6036 -2292
rect 4044 -2332 6036 -2326
<< properties >>
string FIXED_BBOX -6230 -2402 6230 2402
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 4 l 10 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
