magic
tech sky130A
magscale 1 2
timestamp 1689672086
<< psubdiff >>
rect -8900 -4720 -8160 -4696
rect -8900 -5604 -8160 -5580
rect -4500 -5160 -4100 -5136
rect -4500 -5584 -4100 -5560
rect -2420 -5160 -2020 -5136
rect -2420 -5584 -2020 -5560
rect -340 -5160 60 -5136
rect -340 -5584 60 -5560
rect 1740 -5160 2140 -5136
rect 1740 -5584 2140 -5560
<< psubdiffcont >>
rect -8900 -5580 -8160 -4720
rect -4500 -5560 -4100 -5160
rect -2420 -5560 -2020 -5160
rect -340 -5560 60 -5160
rect 1740 -5560 2140 -5160
<< locali >>
rect -10240 4380 -7200 4500
rect -10280 3604 -9380 3680
rect -8460 3604 -7240 3680
rect -10280 3560 -7240 3604
rect -10380 1320 -7340 1440
rect -9560 -100 -9420 1320
rect -6900 1220 -6680 1300
rect -9560 -2320 -9420 -800
rect -8900 -4720 -8160 -4704
rect -4500 -5160 -4100 -5144
rect -4500 -5576 -4100 -5560
rect -2420 -5160 -2020 -5144
rect -2420 -5576 -2020 -5560
rect -340 -5160 60 -5144
rect -340 -5576 60 -5560
rect 1740 -5160 2140 -5144
rect 1740 -5576 2140 -5560
rect -8900 -5596 -8160 -5580
<< viali >>
rect -6680 1220 -6600 1320
rect -10140 -3340 -9860 -3060
rect -8900 -5580 -8160 -4720
rect -4500 -5560 -4100 -5160
rect -2420 -5560 -2020 -5160
rect -340 -5560 60 -5160
rect 1740 -5560 2140 -5160
<< metal1 >>
rect -10520 7300 -6940 8440
rect -10520 7100 -6400 7300
rect -10520 6760 -6940 7100
rect -10340 4260 -9896 4376
rect -7676 4360 -7052 4376
rect -7676 4260 -7100 4360
rect -10340 3800 -10180 4260
rect -7152 3800 -7100 4260
rect -10340 3684 -10024 3800
rect -7720 3684 -7100 3800
rect -7110 3680 -7100 3684
rect -6980 3680 -6970 4360
rect -10228 1418 -7336 1558
rect -9480 -716 -9264 1418
rect -7520 1100 -7360 1418
rect -6680 1332 -6480 7100
rect -5324 4776 -2176 4812
rect -5498 4504 -5488 4776
rect -5204 4688 -2176 4776
rect -148 4688 3000 4812
rect -5204 4504 -5168 4688
rect -148 4668 -28 4688
rect -5324 4228 -5168 4504
rect -254 4432 -244 4668
rect -60 4432 -28 4668
rect -148 4228 -28 4432
rect -5324 4104 -2176 4228
rect -148 4104 3000 4228
rect -6686 1320 -6480 1332
rect -6686 1220 -6680 1320
rect -6600 1220 -6480 1320
rect -6686 1208 -6594 1220
rect -7520 920 -6060 1100
rect -7450 740 -7440 820
rect -7260 740 -7250 820
rect -6220 -300 -6060 920
rect -6220 -560 -5180 -300
rect -9480 -2990 -9262 -716
rect -6220 -800 -6060 -560
rect -6230 -940 -6220 -800
rect -6060 -940 -6050 -800
rect -6220 -1040 -6060 -940
rect -6220 -1160 -5904 -1040
rect -10152 -3060 -9848 -3054
rect -10152 -3340 -10140 -3060
rect -9860 -3340 -9848 -3060
rect -10152 -3346 -9848 -3340
rect -8906 -4720 -8154 -4708
rect -8910 -5580 -8900 -4720
rect -8160 -5580 -8150 -4720
rect -4512 -5160 -4088 -5154
rect -4512 -5560 -4500 -5160
rect -4100 -5560 -4088 -5160
rect -4512 -5566 -4088 -5560
rect -2432 -5160 -2008 -5154
rect -2432 -5560 -2420 -5160
rect -2020 -5560 -2008 -5160
rect -2432 -5566 -2008 -5560
rect -352 -5160 72 -5154
rect -352 -5560 -340 -5160
rect 60 -5560 72 -5160
rect -352 -5566 72 -5560
rect 1728 -5160 2152 -5154
rect 1728 -5560 1740 -5160
rect 2140 -5560 2152 -5160
rect 1728 -5566 2152 -5560
rect -8906 -5592 -8154 -5580
<< via1 >>
rect -7100 3680 -6980 4360
rect -5488 4504 -5204 4776
rect -244 4432 -60 4668
rect -7440 740 -7260 820
rect -6220 -940 -6060 -800
rect -10140 -3340 -9860 -3060
rect -8900 -5580 -8160 -4720
rect -4500 -5560 -4100 -5160
rect -2420 -5560 -2020 -5160
rect -340 -5560 60 -5160
rect 1740 -5560 2140 -5160
<< metal2 >>
rect -10520 6760 -6940 8440
rect -5488 4776 -5204 4786
rect -5488 4494 -5204 4504
rect -244 4668 -60 4678
rect -244 4422 -60 4432
rect -7100 4360 -6980 4370
rect -8448 3938 -7680 3942
rect -10132 3928 -9364 3938
rect -10132 3658 -9364 3668
rect -8460 3932 -7208 3938
rect -8460 3672 -8448 3932
rect -7680 3928 -7208 3932
rect -8460 3662 -8080 3672
rect -8460 3660 -8342 3662
rect -7610 3662 -7208 3672
rect -7100 3670 -6980 3680
rect -8080 3650 -7610 3660
rect -10156 3172 -9754 3182
rect -10156 2640 -9754 2650
rect -9116 3172 -8714 3182
rect -9116 2640 -8714 2650
rect -8084 3168 -7682 3178
rect -8084 2636 -7682 2646
rect -10418 1078 -10330 2402
rect -9552 2288 -8202 2364
rect -10280 1704 -7440 1742
rect -10280 1452 -9520 1704
rect -9134 1452 -8012 1704
rect -9520 1322 -9134 1374
rect -7636 1452 -7440 1704
rect -7636 1336 -7446 1452
rect -8012 1326 -7446 1336
rect -10168 928 -9766 938
rect -10168 396 -9766 406
rect -10420 -1078 -10330 116
rect -9484 0 -9134 1322
rect -7880 1324 -7446 1326
rect -7880 1270 -7520 1324
rect -7440 820 -7260 830
rect -7440 738 -7438 740
rect -7262 738 -7260 740
rect -7440 730 -7260 738
rect -7438 728 -7262 730
rect -9520 -488 -9134 0
rect -9660 -498 -9130 -488
rect -9660 -892 -9130 -882
rect -6220 -800 -6060 -790
rect -9520 -972 -9134 -892
rect -6220 -950 -6060 -940
rect -10174 -1320 -9772 -1310
rect -10174 -1852 -9772 -1842
rect -9476 -2252 -9134 -972
rect -9520 -2694 -9134 -2252
rect -9526 -2724 -9134 -2694
rect -9554 -2740 -9134 -2724
rect -9672 -2750 -9134 -2740
rect -10140 -3060 -9860 -3050
rect -9142 -3132 -9134 -2750
rect -9672 -3142 -9134 -3132
rect -10140 -3350 -9860 -3340
rect -9520 -4316 -9134 -3142
rect -8860 -3420 -8120 -3410
rect -8320 -3690 -8120 -3420
rect -8860 -3710 -8320 -3700
rect -9684 -4326 -9124 -4316
rect -10160 -5420 -9684 -5180
rect -10180 -5512 -9684 -5420
rect -8900 -4720 -8160 -4710
rect -9124 -5512 -8900 -5180
rect -10180 -5580 -8900 -5512
rect -4500 -5160 -4100 -5150
rect -8160 -5580 -5464 -5180
rect -4500 -5570 -4100 -5560
rect -2420 -5160 -2020 -5150
rect -2420 -5570 -2020 -5560
rect -340 -5160 60 -5150
rect -340 -5570 60 -5560
rect 1740 -5160 2140 -5150
rect 1740 -5570 2140 -5560
rect -10180 -5900 -5464 -5580
rect -10180 -7600 -8980 -5900
rect -6180 -7600 -5464 -5900
rect -10180 -7820 -5464 -7600
<< via2 >>
rect -5488 4504 -5204 4776
rect -244 4432 -60 4668
rect -10132 3668 -9364 3928
rect -8448 3928 -7680 3932
rect -8448 3672 -7208 3928
rect -8080 3660 -7610 3672
rect -7100 3860 -6980 4360
rect -10156 2650 -9754 3172
rect -9116 2650 -8714 3172
rect -8084 2646 -7682 3168
rect -9520 1374 -9134 1704
rect -8012 1336 -7636 1704
rect -10168 406 -9766 928
rect -7438 740 -7262 810
rect -7438 738 -7262 740
rect -9660 -882 -9130 -498
rect -6220 -940 -6060 -800
rect -10174 -1842 -9772 -1320
rect -10140 -3340 -9860 -3060
rect -9672 -3132 -9142 -2750
rect -8860 -3700 -8320 -3420
rect -9684 -5512 -9124 -4326
rect -8900 -5580 -8160 -4720
rect -4500 -5560 -4100 -5160
rect -2420 -5560 -2020 -5160
rect -340 -5560 60 -5160
rect 1740 -5560 2140 -5160
rect -8980 -7600 -6180 -5900
<< metal3 >>
rect -10520 8860 9360 8920
rect -10520 8780 4560 8860
rect -10520 8040 -5120 8780
rect 3900 8040 4560 8780
rect -10520 7496 4560 8040
rect -10522 7360 4560 7496
rect -10522 6800 -10400 7360
rect -6980 7000 -5380 7360
rect 4340 7040 4560 7360
rect 5740 7040 8120 8860
rect 9300 7040 9360 8860
rect -6980 6800 -6940 7000
rect 4340 6980 9360 7040
rect -10522 6762 -6940 6800
rect -10520 6760 -6940 6762
rect -4630 5880 -4620 6740
rect -4380 5880 -4370 6740
rect -3870 5880 -3860 6740
rect -3620 5880 -3610 6740
rect -3110 5900 -3100 6740
rect -2860 5900 -2850 6740
rect -2350 5900 -2340 6740
rect -2100 5900 -2090 6740
rect -1590 5900 -1580 6740
rect -1340 5900 -1330 6740
rect 570 5460 580 5640
rect 820 5460 830 5640
rect 1330 5460 1340 5640
rect 1580 5460 1590 5640
rect 2090 5460 2100 5640
rect 2340 5460 2350 5640
rect -9130 4600 -9120 5060
rect -8820 4600 -8810 5060
rect 550 5040 560 5460
rect 840 5040 850 5460
rect 1310 5040 1320 5460
rect 1600 5040 1610 5460
rect 2070 5040 2080 5460
rect 2360 5040 2370 5460
rect -7390 4580 -7380 5040
rect -7080 4580 -7070 5040
rect -5498 4776 -5194 4781
rect 570 4780 580 5040
rect 820 4780 830 5040
rect 1330 4780 1340 5040
rect 1580 4780 1590 5040
rect 2090 4780 2100 5040
rect 2340 4780 2350 5040
rect 2830 4780 2840 5640
rect 3080 5460 3090 5640
rect 3590 5460 3600 5640
rect 3840 5460 3850 5640
rect 3120 5040 3130 5460
rect 3570 5040 3580 5460
rect 3860 5040 3870 5460
rect 3080 4780 3090 5040
rect 3590 4780 3600 5040
rect 3840 4780 3850 5040
rect -5498 4504 -5488 4776
rect -5204 4504 -5194 4776
rect -5498 4499 -5194 4504
rect -254 4668 -50 4673
rect -254 4432 -244 4668
rect -60 4432 -50 4668
rect -254 4427 -50 4432
rect -7110 4360 -6970 4365
rect -10172 3976 -9748 3980
rect -8080 3976 -7680 3978
rect -10172 3937 -7680 3976
rect -10172 3933 -7670 3937
rect -10172 3932 -7198 3933
rect -10172 3928 -8448 3932
rect -7680 3928 -7198 3932
rect -10172 3668 -10132 3928
rect -9364 3672 -8448 3928
rect -7208 3672 -7198 3928
rect -7110 3860 -7100 4360
rect -6980 3860 -6760 4360
rect -7110 3855 -6760 3860
rect -9364 3668 -8080 3672
rect -10172 3660 -8080 3668
rect -7610 3667 -7198 3672
rect -7610 3660 -7600 3667
rect -10172 3656 -7600 3660
rect -10172 3177 -9748 3656
rect -8090 3655 -7600 3656
rect -10172 3172 -9744 3177
rect -10174 2650 -10156 3172
rect -9754 3170 -9744 3172
rect -9126 3172 -8704 3177
rect -8080 3173 -7680 3655
rect -7100 3460 -6760 3855
rect -9126 3170 -9116 3172
rect -9754 2650 -9116 3170
rect -8714 3170 -8704 3172
rect -8094 3170 -7672 3173
rect -8714 3168 -7672 3170
rect -8714 2650 -8084 3168
rect -10174 2645 -9744 2650
rect -9126 2645 -8704 2650
rect -8094 2646 -8084 2650
rect -7682 2646 -7672 3168
rect -10174 933 -9750 2645
rect -8094 2641 -7672 2646
rect 4520 2440 5820 6980
rect 8060 2320 9360 6980
rect -9682 1709 -7636 1728
rect -9682 1708 -7626 1709
rect -9684 1704 -7626 1708
rect -9684 1700 -9520 1704
rect -9690 1320 -9680 1700
rect -9134 1374 -8012 1704
rect -9140 1336 -8012 1374
rect -7636 1336 -7626 1704
rect -9140 1332 -7626 1336
rect -9140 1320 -9124 1332
rect -8022 1331 -7626 1332
rect -10178 928 -9750 933
rect -10178 406 -10168 928
rect -9766 406 -9750 928
rect -10178 401 -9750 406
rect -10174 -1315 -9750 401
rect -10184 -1320 -9750 -1315
rect -10184 -1842 -10174 -1320
rect -9772 -1842 -9750 -1320
rect -9684 -493 -9124 1320
rect -7448 810 -6728 882
rect -7448 738 -7438 810
rect -7262 802 -6728 810
rect -7262 738 -7252 802
rect -7448 733 -7252 738
rect -8492 384 -8124 510
rect -9684 -498 -9120 -493
rect -9684 -882 -9660 -498
rect -9130 -500 -9120 -498
rect -9120 -880 -9110 -500
rect -9130 -882 -9120 -880
rect -9684 -887 -9120 -882
rect -10184 -1847 -9762 -1842
rect -9684 -2750 -9124 -887
rect -6862 -1220 -6730 802
rect -6230 -800 -6050 -795
rect -6230 -940 -6220 -800
rect -6060 -940 -6050 -800
rect -6230 -945 -6050 -940
rect -6220 -1220 -6060 -945
rect -6862 -1340 -6060 -1220
rect -8840 -1440 -8700 -1380
rect -6862 -1400 -6140 -1340
rect -6862 -1926 -6730 -1400
rect -10150 -3060 -9850 -3055
rect -10150 -3340 -10140 -3060
rect -9860 -3340 -9850 -3060
rect -10150 -3345 -9850 -3340
rect -9684 -3132 -9672 -2750
rect -9142 -3132 -9124 -2750
rect -9684 -4321 -9124 -3132
rect -8870 -3420 -8310 -3415
rect -8870 -4040 -8860 -3420
rect -8320 -4040 -8310 -3420
rect 5040 -3820 6500 -2000
rect -9694 -4326 -9114 -4321
rect -9694 -5000 -9684 -4326
rect -10180 -5512 -9684 -5000
rect -9124 -5000 -9114 -4326
rect -4940 -4600 3220 -3900
rect 8460 -4040 9920 -2220
rect -8910 -4720 -8150 -4715
rect -8910 -5000 -8900 -4720
rect -9124 -5512 -8900 -5000
rect -10180 -5580 -8900 -5512
rect -8160 -5000 -8150 -4720
rect -4940 -5000 3240 -4600
rect -8160 -5100 3240 -5000
rect -8160 -5580 -4940 -5100
rect -10180 -5900 -4940 -5580
rect -10180 -7600 -8980 -5900
rect -6180 -6180 -4940 -5900
rect 3240 -6180 3250 -5100
rect -6180 -7600 3240 -6180
rect -10180 -7820 3240 -7600
<< via3 >>
rect -5120 8040 3900 8780
rect -10400 6800 -6980 7360
rect 4560 7040 5740 8860
rect 8120 7040 9300 8860
rect -4620 5880 -4380 6740
rect -3860 5880 -3620 6740
rect -3100 5900 -2860 6740
rect -2340 5900 -2100 6740
rect -1580 5900 -1340 6740
rect 580 5460 820 5640
rect 1340 5460 1580 5640
rect 2100 5460 2340 5640
rect -9120 4600 -8820 5060
rect 560 5040 840 5460
rect 1320 5040 1600 5460
rect 2080 5040 2360 5460
rect -7380 4580 -7080 5040
rect 580 4780 820 5040
rect 1340 4780 1580 5040
rect 2100 4780 2340 5040
rect 2840 5460 3080 5640
rect 3600 5460 3840 5640
rect 2840 5040 3120 5460
rect 3580 5040 3860 5460
rect 2840 4780 3080 5040
rect 3600 4780 3840 5040
rect -5488 4504 -5204 4776
rect -244 4432 -60 4668
rect -9680 1374 -9520 1700
rect -9520 1374 -9140 1700
rect -9680 1320 -9140 1374
rect -8012 1336 -7636 1704
rect -9660 -880 -9130 -500
rect -9130 -880 -9120 -500
rect -10140 -3340 -9860 -3060
rect -9660 -3120 -9160 -2760
rect -8860 -3700 -8320 -3420
rect -8860 -4040 -8320 -3700
rect -9684 -5512 -9124 -4326
rect -8900 -5580 -8160 -4720
rect -4940 -5160 3240 -5100
rect -4940 -5560 -4500 -5160
rect -4500 -5560 -4100 -5160
rect -4100 -5560 -2420 -5160
rect -2420 -5560 -2020 -5160
rect -2020 -5560 -340 -5160
rect -340 -5560 60 -5160
rect 60 -5560 1740 -5160
rect 1740 -5560 2140 -5160
rect 2140 -5560 3240 -5160
rect -8980 -7600 -6180 -5900
rect -4940 -6180 3240 -5560
<< metal4 >>
rect -2480 8900 9360 8920
rect -10520 8860 9360 8900
rect -10520 8780 4560 8860
rect -10520 8040 -5120 8780
rect 3900 8040 4560 8780
rect -10520 7360 4560 8040
rect -10520 6800 -10400 7360
rect -6980 7040 4560 7360
rect 5740 7040 8120 8860
rect 9300 7040 9360 8860
rect -6980 6980 9360 7040
rect -6980 6800 -6940 6980
rect -10520 6760 -6940 6800
rect -4660 6740 6840 6760
rect -4660 5880 -4620 6740
rect -4380 5880 -3860 6740
rect -3620 5900 -3100 6740
rect -2860 5900 -2340 6740
rect -2100 5900 -1580 6740
rect -1340 5900 6840 6740
rect -3620 5880 6840 5900
rect -4660 5860 6840 5880
rect -9120 5320 -5520 5740
rect -9120 5061 -8760 5320
rect -9121 5060 -8760 5061
rect -9121 4600 -9120 5060
rect -8820 4600 -8760 5060
rect -7381 5040 -7079 5041
rect -9121 4599 -8819 4600
rect -7381 4580 -7380 5040
rect -7080 4580 -6000 5040
rect -7381 4579 -7079 4580
rect -6320 4360 -6000 4580
rect -5840 4800 -5520 5320
rect -440 5640 6820 5660
rect -440 5460 580 5640
rect 820 5460 1340 5640
rect 1580 5460 2100 5640
rect 2340 5460 2840 5640
rect 3080 5460 3600 5640
rect 3840 5460 6820 5640
rect -440 5040 560 5460
rect 840 5040 1320 5460
rect 1600 5040 2080 5460
rect 2360 5040 2840 5460
rect 3120 5040 3580 5460
rect 3860 5040 6820 5460
rect -5840 4777 -5260 4800
rect -440 4780 580 5040
rect 820 4780 1340 5040
rect 1580 4780 2100 5040
rect 2340 4780 2840 5040
rect 3080 4780 3600 5040
rect 3840 4780 6820 5040
rect -5840 4776 -5203 4777
rect -5840 4504 -5488 4776
rect -5204 4504 -5203 4776
rect -440 4760 6820 4780
rect -5840 4503 -5203 4504
rect -1720 4669 -180 4680
rect -1720 4668 -59 4669
rect -5840 4480 -5260 4503
rect -1720 4432 -244 4668
rect -60 4432 -59 4668
rect -1720 4431 -59 4432
rect -1720 4420 -180 4431
rect -1720 4360 -1420 4420
rect -6320 4040 -1420 4360
rect -10200 1701 -9140 1720
rect -8013 1704 -7635 1705
rect -10200 1700 -9139 1701
rect -10200 1320 -9680 1700
rect -9140 1320 -8994 1700
rect -8013 1336 -8012 1704
rect -7636 1700 -7635 1704
rect -7636 1336 -6100 1700
rect -8013 1335 -6100 1336
rect -10200 840 -8994 1320
rect -8012 840 -6100 1335
rect -10200 -499 -9140 840
rect -10200 -500 -9119 -499
rect -10200 -880 -9660 -500
rect -9120 -880 -9119 -500
rect -10200 -881 -9119 -880
rect -10200 -2760 -9140 -881
rect -6760 -1960 -6100 840
rect -10200 -3060 -9660 -2760
rect -10200 -3340 -10140 -3060
rect -9860 -3120 -9660 -3060
rect -9160 -3120 -9140 -2760
rect -9860 -3340 -9140 -3120
rect -10200 -3380 -9140 -3340
rect -10200 -3419 -8320 -3380
rect -10200 -3420 -8319 -3419
rect -10200 -4040 -8860 -3420
rect -8320 -4040 -8319 -3420
rect 5140 -3620 6600 -2060
rect -10200 -4041 -8319 -4040
rect -10200 -4100 -8320 -4041
rect -10200 -4325 -9140 -4100
rect -10200 -4326 -9123 -4325
rect -10200 -5512 -9684 -4326
rect -9124 -4598 -9123 -4326
rect -7100 -4598 -6380 -4280
rect -9124 -4600 -6020 -4598
rect -4940 -4600 7320 -3620
rect 8580 -4020 10040 -2200
rect -9124 -4720 7320 -4600
rect -9124 -5512 -8900 -4720
rect -10200 -5580 -8900 -5512
rect -8160 -5100 7320 -4720
rect -8160 -5580 -4940 -5100
rect -10200 -5900 -4940 -5580
rect -10200 -7600 -8980 -5900
rect -6180 -6180 -4940 -5900
rect 3240 -6040 7320 -5100
rect 3240 -6180 3860 -6040
rect -6180 -7600 3860 -6180
rect -10200 -7800 3860 -7600
rect -10180 -7820 3860 -7800
use outd_curm  outd_curm_1
timestamp 1683888831
transform 1 0 -9340 0 1 464
box -40 916 1002 3158
use outd_curm  outd_curm_2
timestamp 1683888831
transform 1 0 -8300 0 1 464
box -40 916 1002 3158
use outd_curm  outd_curm_3
timestamp 1683888831
transform 1 0 -10380 0 1 -1776
box -40 916 1002 3158
use outd_curm  outd_curm_4
timestamp 1683888831
transform 1 0 -10382 0 1 -4020
box -40 916 1002 3158
use outd_curm  outd_curm_9
timestamp 1683888831
transform 1 0 -10380 0 1 464
box -40 916 1002 3158
use outd_diffamp_6  outd_diffamp_6_0
timestamp 1689672086
transform 1 0 -10340 0 1 3600
box -80 20 1668 3804
use outd_diffamp_6  outd_diffamp_6_1
timestamp 1689672086
transform 1 0 -8600 0 1 3600
box -80 20 1668 3804
use outd_diffamp_50ohm_top_lg  outd_diffamp_50ohm_top_lg_0
timestamp 1687119368
transform 1 0 -12060 0 1 2188
box 6740 -7100 16178 6720
use outd_filter  outd_filter_0
timestamp 1684930430
transform 1 0 -12000 0 1 -4650
box 2696 870 5300 5940
use sky130_fd_pr__cap_mim_m3_1_2YC3NK  sky130_fd_pr__cap_mim_m3_1_2YC3NK_0
timestamp 1685108691
transform 0 1 7280 -1 0 -4934
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_2YC3NK  sky130_fd_pr__cap_mim_m3_1_2YC3NK_1
timestamp 1685108691
transform -1 0 9786 0 -1 240
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_2YC3NK  sky130_fd_pr__cap_mim_m3_1_2YC3NK_2
timestamp 1685108691
transform 1 0 5986 0 1 240
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_5F7Q4P  sky130_fd_pr__cap_mim_m3_1_5F7Q4P_0
timestamp 1684833579
transform 0 -1 -6652 1 0 2380
box -1186 -640 1186 640
use sky130_fd_pr__cap_mim_m3_1_5KPPX9  sky130_fd_pr__cap_mim_m3_1_5KPPX9_0
timestamp 1684929745
transform 1 0 -6834 0 1 -2880
box -1186 -1640 1186 1640
<< labels >>
rlabel metal4 -9960 -6980 -9240 -4660 1 VN
port 4 n
rlabel metal1 -10318 3778 -10268 4194 1 InputSignal
port 5 n
rlabel metal3 -7068 3922 -6994 4080 1 InputRef
port 6 n
rlabel metal3 -10306 7624 -9980 7986 1 VP
port 7 n
rlabel metal3 -8412 406 -8214 500 1 I_Bias
port 8 n
rlabel metal3 -8840 -1440 -8700 -1380 1 VM18D
rlabel metal1 -6040 -1140 -5920 -1060 1 VM6D
rlabel metal4 -5800 4520 -5580 4760 1 V_da2_P
rlabel metal4 -5800 4100 -5580 4340 1 V_da2_N
rlabel metal4 6000 6000 6800 6600 1 outP
port 10 n
rlabel metal4 6000 4800 6800 5600 1 outN
<< end >>
