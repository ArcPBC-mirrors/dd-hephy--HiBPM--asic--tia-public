magic
tech sky130A
magscale 1 2
timestamp 1684165924
<< metal3 >>
rect -2686 6172 2686 6200
rect -2686 148 2602 6172
rect 2666 148 2686 6172
rect -2686 120 2686 148
rect -2686 -148 2686 -120
rect -2686 -6172 2602 -148
rect 2666 -6172 2686 -148
rect -2686 -6200 2686 -6172
<< via3 >>
rect 2602 148 2666 6172
rect 2602 -6172 2666 -148
<< mimcap >>
rect -2646 6120 2354 6160
rect -2646 200 -2606 6120
rect 2314 200 2354 6120
rect -2646 160 2354 200
rect -2646 -200 2354 -160
rect -2646 -6120 -2606 -200
rect 2314 -6120 2354 -200
rect -2646 -6160 2354 -6120
<< mimcapcontact >>
rect -2606 200 2314 6120
rect -2606 -6120 2314 -200
<< metal4 >>
rect 2586 6172 2682 6188
rect -2607 6120 2315 6121
rect -2607 200 -2606 6120
rect 2314 200 2315 6120
rect -2607 199 2315 200
rect 2586 148 2602 6172
rect 2666 148 2682 6172
rect 2586 132 2682 148
rect 2586 -148 2682 -132
rect -2607 -200 2315 -199
rect -2607 -6120 -2606 -200
rect 2314 -6120 2315 -200
rect -2607 -6121 2315 -6120
rect 2586 -6172 2602 -148
rect 2666 -6172 2682 -148
rect 2586 -6188 2682 -6172
<< properties >>
string FIXED_BBOX -2686 120 2394 6200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25 l 30 val 1.52k carea 2.00 cperi 0.19 nx 1 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
