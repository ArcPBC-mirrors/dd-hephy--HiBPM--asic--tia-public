magic
tech sky130A
magscale 1 2
timestamp 1687117224
<< error_p >>
rect -29 9233 29 9239
rect -29 9199 -17 9233
rect -29 9193 29 9199
rect -29 8723 29 8729
rect -29 8689 -17 8723
rect -29 8683 29 8689
rect -29 8615 29 8621
rect -29 8581 -17 8615
rect -29 8575 29 8581
rect -29 8105 29 8111
rect -29 8071 -17 8105
rect -29 8065 29 8071
rect -29 7997 29 8003
rect -29 7963 -17 7997
rect -29 7957 29 7963
rect -29 7487 29 7493
rect -29 7453 -17 7487
rect -29 7447 29 7453
rect -29 7379 29 7385
rect -29 7345 -17 7379
rect -29 7339 29 7345
rect -29 6869 29 6875
rect -29 6835 -17 6869
rect -29 6829 29 6835
rect -29 6761 29 6767
rect -29 6727 -17 6761
rect -29 6721 29 6727
rect -29 6251 29 6257
rect -29 6217 -17 6251
rect -29 6211 29 6217
rect -29 6143 29 6149
rect -29 6109 -17 6143
rect -29 6103 29 6109
rect -29 5633 29 5639
rect -29 5599 -17 5633
rect -29 5593 29 5599
rect -29 5525 29 5531
rect -29 5491 -17 5525
rect -29 5485 29 5491
rect -29 5015 29 5021
rect -29 4981 -17 5015
rect -29 4975 29 4981
rect -29 4907 29 4913
rect -29 4873 -17 4907
rect -29 4867 29 4873
rect -29 4397 29 4403
rect -29 4363 -17 4397
rect -29 4357 29 4363
rect -29 4289 29 4295
rect -29 4255 -17 4289
rect -29 4249 29 4255
rect -29 3779 29 3785
rect -29 3745 -17 3779
rect -29 3739 29 3745
rect -29 3671 29 3677
rect -29 3637 -17 3671
rect -29 3631 29 3637
rect -29 3161 29 3167
rect -29 3127 -17 3161
rect -29 3121 29 3127
rect -29 3053 29 3059
rect -29 3019 -17 3053
rect -29 3013 29 3019
rect -29 2543 29 2549
rect -29 2509 -17 2543
rect -29 2503 29 2509
rect -29 2435 29 2441
rect -29 2401 -17 2435
rect -29 2395 29 2401
rect -29 1925 29 1931
rect -29 1891 -17 1925
rect -29 1885 29 1891
rect -29 1817 29 1823
rect -29 1783 -17 1817
rect -29 1777 29 1783
rect -29 1307 29 1313
rect -29 1273 -17 1307
rect -29 1267 29 1273
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect -29 1159 29 1165
rect -29 689 29 695
rect -29 655 -17 689
rect -29 649 29 655
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
rect -29 -655 29 -649
rect -29 -689 -17 -655
rect -29 -695 29 -689
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect -29 -1205 29 -1199
rect -29 -1273 29 -1267
rect -29 -1307 -17 -1273
rect -29 -1313 29 -1307
rect -29 -1783 29 -1777
rect -29 -1817 -17 -1783
rect -29 -1823 29 -1817
rect -29 -1891 29 -1885
rect -29 -1925 -17 -1891
rect -29 -1931 29 -1925
rect -29 -2401 29 -2395
rect -29 -2435 -17 -2401
rect -29 -2441 29 -2435
rect -29 -2509 29 -2503
rect -29 -2543 -17 -2509
rect -29 -2549 29 -2543
rect -29 -3019 29 -3013
rect -29 -3053 -17 -3019
rect -29 -3059 29 -3053
rect -29 -3127 29 -3121
rect -29 -3161 -17 -3127
rect -29 -3167 29 -3161
rect -29 -3637 29 -3631
rect -29 -3671 -17 -3637
rect -29 -3677 29 -3671
rect -29 -3745 29 -3739
rect -29 -3779 -17 -3745
rect -29 -3785 29 -3779
rect -29 -4255 29 -4249
rect -29 -4289 -17 -4255
rect -29 -4295 29 -4289
rect -29 -4363 29 -4357
rect -29 -4397 -17 -4363
rect -29 -4403 29 -4397
rect -29 -4873 29 -4867
rect -29 -4907 -17 -4873
rect -29 -4913 29 -4907
rect -29 -4981 29 -4975
rect -29 -5015 -17 -4981
rect -29 -5021 29 -5015
rect -29 -5491 29 -5485
rect -29 -5525 -17 -5491
rect -29 -5531 29 -5525
rect -29 -5599 29 -5593
rect -29 -5633 -17 -5599
rect -29 -5639 29 -5633
rect -29 -6109 29 -6103
rect -29 -6143 -17 -6109
rect -29 -6149 29 -6143
rect -29 -6217 29 -6211
rect -29 -6251 -17 -6217
rect -29 -6257 29 -6251
rect -29 -6727 29 -6721
rect -29 -6761 -17 -6727
rect -29 -6767 29 -6761
rect -29 -6835 29 -6829
rect -29 -6869 -17 -6835
rect -29 -6875 29 -6869
rect -29 -7345 29 -7339
rect -29 -7379 -17 -7345
rect -29 -7385 29 -7379
rect -29 -7453 29 -7447
rect -29 -7487 -17 -7453
rect -29 -7493 29 -7487
rect -29 -7963 29 -7957
rect -29 -7997 -17 -7963
rect -29 -8003 29 -7997
rect -29 -8071 29 -8065
rect -29 -8105 -17 -8071
rect -29 -8111 29 -8105
rect -29 -8581 29 -8575
rect -29 -8615 -17 -8581
rect -29 -8621 29 -8615
rect -29 -8689 29 -8683
rect -29 -8723 -17 -8689
rect -29 -8729 29 -8723
rect -29 -9199 29 -9193
rect -29 -9233 -17 -9199
rect -29 -9239 29 -9233
<< pwell >>
rect -211 -9371 211 9371
<< nmoslvt >>
rect -15 8761 15 9161
rect -15 8143 15 8543
rect -15 7525 15 7925
rect -15 6907 15 7307
rect -15 6289 15 6689
rect -15 5671 15 6071
rect -15 5053 15 5453
rect -15 4435 15 4835
rect -15 3817 15 4217
rect -15 3199 15 3599
rect -15 2581 15 2981
rect -15 1963 15 2363
rect -15 1345 15 1745
rect -15 727 15 1127
rect -15 109 15 509
rect -15 -509 15 -109
rect -15 -1127 15 -727
rect -15 -1745 15 -1345
rect -15 -2363 15 -1963
rect -15 -2981 15 -2581
rect -15 -3599 15 -3199
rect -15 -4217 15 -3817
rect -15 -4835 15 -4435
rect -15 -5453 15 -5053
rect -15 -6071 15 -5671
rect -15 -6689 15 -6289
rect -15 -7307 15 -6907
rect -15 -7925 15 -7525
rect -15 -8543 15 -8143
rect -15 -9161 15 -8761
<< ndiff >>
rect -73 9149 -15 9161
rect -73 8773 -61 9149
rect -27 8773 -15 9149
rect -73 8761 -15 8773
rect 15 9149 73 9161
rect 15 8773 27 9149
rect 61 8773 73 9149
rect 15 8761 73 8773
rect -73 8531 -15 8543
rect -73 8155 -61 8531
rect -27 8155 -15 8531
rect -73 8143 -15 8155
rect 15 8531 73 8543
rect 15 8155 27 8531
rect 61 8155 73 8531
rect 15 8143 73 8155
rect -73 7913 -15 7925
rect -73 7537 -61 7913
rect -27 7537 -15 7913
rect -73 7525 -15 7537
rect 15 7913 73 7925
rect 15 7537 27 7913
rect 61 7537 73 7913
rect 15 7525 73 7537
rect -73 7295 -15 7307
rect -73 6919 -61 7295
rect -27 6919 -15 7295
rect -73 6907 -15 6919
rect 15 7295 73 7307
rect 15 6919 27 7295
rect 61 6919 73 7295
rect 15 6907 73 6919
rect -73 6677 -15 6689
rect -73 6301 -61 6677
rect -27 6301 -15 6677
rect -73 6289 -15 6301
rect 15 6677 73 6689
rect 15 6301 27 6677
rect 61 6301 73 6677
rect 15 6289 73 6301
rect -73 6059 -15 6071
rect -73 5683 -61 6059
rect -27 5683 -15 6059
rect -73 5671 -15 5683
rect 15 6059 73 6071
rect 15 5683 27 6059
rect 61 5683 73 6059
rect 15 5671 73 5683
rect -73 5441 -15 5453
rect -73 5065 -61 5441
rect -27 5065 -15 5441
rect -73 5053 -15 5065
rect 15 5441 73 5453
rect 15 5065 27 5441
rect 61 5065 73 5441
rect 15 5053 73 5065
rect -73 4823 -15 4835
rect -73 4447 -61 4823
rect -27 4447 -15 4823
rect -73 4435 -15 4447
rect 15 4823 73 4835
rect 15 4447 27 4823
rect 61 4447 73 4823
rect 15 4435 73 4447
rect -73 4205 -15 4217
rect -73 3829 -61 4205
rect -27 3829 -15 4205
rect -73 3817 -15 3829
rect 15 4205 73 4217
rect 15 3829 27 4205
rect 61 3829 73 4205
rect 15 3817 73 3829
rect -73 3587 -15 3599
rect -73 3211 -61 3587
rect -27 3211 -15 3587
rect -73 3199 -15 3211
rect 15 3587 73 3599
rect 15 3211 27 3587
rect 61 3211 73 3587
rect 15 3199 73 3211
rect -73 2969 -15 2981
rect -73 2593 -61 2969
rect -27 2593 -15 2969
rect -73 2581 -15 2593
rect 15 2969 73 2981
rect 15 2593 27 2969
rect 61 2593 73 2969
rect 15 2581 73 2593
rect -73 2351 -15 2363
rect -73 1975 -61 2351
rect -27 1975 -15 2351
rect -73 1963 -15 1975
rect 15 2351 73 2363
rect 15 1975 27 2351
rect 61 1975 73 2351
rect 15 1963 73 1975
rect -73 1733 -15 1745
rect -73 1357 -61 1733
rect -27 1357 -15 1733
rect -73 1345 -15 1357
rect 15 1733 73 1745
rect 15 1357 27 1733
rect 61 1357 73 1733
rect 15 1345 73 1357
rect -73 1115 -15 1127
rect -73 739 -61 1115
rect -27 739 -15 1115
rect -73 727 -15 739
rect 15 1115 73 1127
rect 15 739 27 1115
rect 61 739 73 1115
rect 15 727 73 739
rect -73 497 -15 509
rect -73 121 -61 497
rect -27 121 -15 497
rect -73 109 -15 121
rect 15 497 73 509
rect 15 121 27 497
rect 61 121 73 497
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -497 -61 -121
rect -27 -497 -15 -121
rect -73 -509 -15 -497
rect 15 -121 73 -109
rect 15 -497 27 -121
rect 61 -497 73 -121
rect 15 -509 73 -497
rect -73 -739 -15 -727
rect -73 -1115 -61 -739
rect -27 -1115 -15 -739
rect -73 -1127 -15 -1115
rect 15 -739 73 -727
rect 15 -1115 27 -739
rect 61 -1115 73 -739
rect 15 -1127 73 -1115
rect -73 -1357 -15 -1345
rect -73 -1733 -61 -1357
rect -27 -1733 -15 -1357
rect -73 -1745 -15 -1733
rect 15 -1357 73 -1345
rect 15 -1733 27 -1357
rect 61 -1733 73 -1357
rect 15 -1745 73 -1733
rect -73 -1975 -15 -1963
rect -73 -2351 -61 -1975
rect -27 -2351 -15 -1975
rect -73 -2363 -15 -2351
rect 15 -1975 73 -1963
rect 15 -2351 27 -1975
rect 61 -2351 73 -1975
rect 15 -2363 73 -2351
rect -73 -2593 -15 -2581
rect -73 -2969 -61 -2593
rect -27 -2969 -15 -2593
rect -73 -2981 -15 -2969
rect 15 -2593 73 -2581
rect 15 -2969 27 -2593
rect 61 -2969 73 -2593
rect 15 -2981 73 -2969
rect -73 -3211 -15 -3199
rect -73 -3587 -61 -3211
rect -27 -3587 -15 -3211
rect -73 -3599 -15 -3587
rect 15 -3211 73 -3199
rect 15 -3587 27 -3211
rect 61 -3587 73 -3211
rect 15 -3599 73 -3587
rect -73 -3829 -15 -3817
rect -73 -4205 -61 -3829
rect -27 -4205 -15 -3829
rect -73 -4217 -15 -4205
rect 15 -3829 73 -3817
rect 15 -4205 27 -3829
rect 61 -4205 73 -3829
rect 15 -4217 73 -4205
rect -73 -4447 -15 -4435
rect -73 -4823 -61 -4447
rect -27 -4823 -15 -4447
rect -73 -4835 -15 -4823
rect 15 -4447 73 -4435
rect 15 -4823 27 -4447
rect 61 -4823 73 -4447
rect 15 -4835 73 -4823
rect -73 -5065 -15 -5053
rect -73 -5441 -61 -5065
rect -27 -5441 -15 -5065
rect -73 -5453 -15 -5441
rect 15 -5065 73 -5053
rect 15 -5441 27 -5065
rect 61 -5441 73 -5065
rect 15 -5453 73 -5441
rect -73 -5683 -15 -5671
rect -73 -6059 -61 -5683
rect -27 -6059 -15 -5683
rect -73 -6071 -15 -6059
rect 15 -5683 73 -5671
rect 15 -6059 27 -5683
rect 61 -6059 73 -5683
rect 15 -6071 73 -6059
rect -73 -6301 -15 -6289
rect -73 -6677 -61 -6301
rect -27 -6677 -15 -6301
rect -73 -6689 -15 -6677
rect 15 -6301 73 -6289
rect 15 -6677 27 -6301
rect 61 -6677 73 -6301
rect 15 -6689 73 -6677
rect -73 -6919 -15 -6907
rect -73 -7295 -61 -6919
rect -27 -7295 -15 -6919
rect -73 -7307 -15 -7295
rect 15 -6919 73 -6907
rect 15 -7295 27 -6919
rect 61 -7295 73 -6919
rect 15 -7307 73 -7295
rect -73 -7537 -15 -7525
rect -73 -7913 -61 -7537
rect -27 -7913 -15 -7537
rect -73 -7925 -15 -7913
rect 15 -7537 73 -7525
rect 15 -7913 27 -7537
rect 61 -7913 73 -7537
rect 15 -7925 73 -7913
rect -73 -8155 -15 -8143
rect -73 -8531 -61 -8155
rect -27 -8531 -15 -8155
rect -73 -8543 -15 -8531
rect 15 -8155 73 -8143
rect 15 -8531 27 -8155
rect 61 -8531 73 -8155
rect 15 -8543 73 -8531
rect -73 -8773 -15 -8761
rect -73 -9149 -61 -8773
rect -27 -9149 -15 -8773
rect -73 -9161 -15 -9149
rect 15 -8773 73 -8761
rect 15 -9149 27 -8773
rect 61 -9149 73 -8773
rect 15 -9161 73 -9149
<< ndiffc >>
rect -61 8773 -27 9149
rect 27 8773 61 9149
rect -61 8155 -27 8531
rect 27 8155 61 8531
rect -61 7537 -27 7913
rect 27 7537 61 7913
rect -61 6919 -27 7295
rect 27 6919 61 7295
rect -61 6301 -27 6677
rect 27 6301 61 6677
rect -61 5683 -27 6059
rect 27 5683 61 6059
rect -61 5065 -27 5441
rect 27 5065 61 5441
rect -61 4447 -27 4823
rect 27 4447 61 4823
rect -61 3829 -27 4205
rect 27 3829 61 4205
rect -61 3211 -27 3587
rect 27 3211 61 3587
rect -61 2593 -27 2969
rect 27 2593 61 2969
rect -61 1975 -27 2351
rect 27 1975 61 2351
rect -61 1357 -27 1733
rect 27 1357 61 1733
rect -61 739 -27 1115
rect 27 739 61 1115
rect -61 121 -27 497
rect 27 121 61 497
rect -61 -497 -27 -121
rect 27 -497 61 -121
rect -61 -1115 -27 -739
rect 27 -1115 61 -739
rect -61 -1733 -27 -1357
rect 27 -1733 61 -1357
rect -61 -2351 -27 -1975
rect 27 -2351 61 -1975
rect -61 -2969 -27 -2593
rect 27 -2969 61 -2593
rect -61 -3587 -27 -3211
rect 27 -3587 61 -3211
rect -61 -4205 -27 -3829
rect 27 -4205 61 -3829
rect -61 -4823 -27 -4447
rect 27 -4823 61 -4447
rect -61 -5441 -27 -5065
rect 27 -5441 61 -5065
rect -61 -6059 -27 -5683
rect 27 -6059 61 -5683
rect -61 -6677 -27 -6301
rect 27 -6677 61 -6301
rect -61 -7295 -27 -6919
rect 27 -7295 61 -6919
rect -61 -7913 -27 -7537
rect 27 -7913 61 -7537
rect -61 -8531 -27 -8155
rect 27 -8531 61 -8155
rect -61 -9149 -27 -8773
rect 27 -9149 61 -8773
<< psubdiff >>
rect -175 9301 -79 9335
rect 79 9301 175 9335
rect -175 9239 -141 9301
rect 141 9239 175 9301
rect -175 -9301 -141 -9239
rect 141 -9301 175 -9239
rect -175 -9335 -79 -9301
rect 79 -9335 175 -9301
<< psubdiffcont >>
rect -79 9301 79 9335
rect -175 -9239 -141 9239
rect 141 -9239 175 9239
rect -79 -9335 79 -9301
<< poly >>
rect -33 9233 33 9249
rect -33 9199 -17 9233
rect 17 9199 33 9233
rect -33 9183 33 9199
rect -15 9161 15 9183
rect -15 8739 15 8761
rect -33 8723 33 8739
rect -33 8689 -17 8723
rect 17 8689 33 8723
rect -33 8673 33 8689
rect -33 8615 33 8631
rect -33 8581 -17 8615
rect 17 8581 33 8615
rect -33 8565 33 8581
rect -15 8543 15 8565
rect -15 8121 15 8143
rect -33 8105 33 8121
rect -33 8071 -17 8105
rect 17 8071 33 8105
rect -33 8055 33 8071
rect -33 7997 33 8013
rect -33 7963 -17 7997
rect 17 7963 33 7997
rect -33 7947 33 7963
rect -15 7925 15 7947
rect -15 7503 15 7525
rect -33 7487 33 7503
rect -33 7453 -17 7487
rect 17 7453 33 7487
rect -33 7437 33 7453
rect -33 7379 33 7395
rect -33 7345 -17 7379
rect 17 7345 33 7379
rect -33 7329 33 7345
rect -15 7307 15 7329
rect -15 6885 15 6907
rect -33 6869 33 6885
rect -33 6835 -17 6869
rect 17 6835 33 6869
rect -33 6819 33 6835
rect -33 6761 33 6777
rect -33 6727 -17 6761
rect 17 6727 33 6761
rect -33 6711 33 6727
rect -15 6689 15 6711
rect -15 6267 15 6289
rect -33 6251 33 6267
rect -33 6217 -17 6251
rect 17 6217 33 6251
rect -33 6201 33 6217
rect -33 6143 33 6159
rect -33 6109 -17 6143
rect 17 6109 33 6143
rect -33 6093 33 6109
rect -15 6071 15 6093
rect -15 5649 15 5671
rect -33 5633 33 5649
rect -33 5599 -17 5633
rect 17 5599 33 5633
rect -33 5583 33 5599
rect -33 5525 33 5541
rect -33 5491 -17 5525
rect 17 5491 33 5525
rect -33 5475 33 5491
rect -15 5453 15 5475
rect -15 5031 15 5053
rect -33 5015 33 5031
rect -33 4981 -17 5015
rect 17 4981 33 5015
rect -33 4965 33 4981
rect -33 4907 33 4923
rect -33 4873 -17 4907
rect 17 4873 33 4907
rect -33 4857 33 4873
rect -15 4835 15 4857
rect -15 4413 15 4435
rect -33 4397 33 4413
rect -33 4363 -17 4397
rect 17 4363 33 4397
rect -33 4347 33 4363
rect -33 4289 33 4305
rect -33 4255 -17 4289
rect 17 4255 33 4289
rect -33 4239 33 4255
rect -15 4217 15 4239
rect -15 3795 15 3817
rect -33 3779 33 3795
rect -33 3745 -17 3779
rect 17 3745 33 3779
rect -33 3729 33 3745
rect -33 3671 33 3687
rect -33 3637 -17 3671
rect 17 3637 33 3671
rect -33 3621 33 3637
rect -15 3599 15 3621
rect -15 3177 15 3199
rect -33 3161 33 3177
rect -33 3127 -17 3161
rect 17 3127 33 3161
rect -33 3111 33 3127
rect -33 3053 33 3069
rect -33 3019 -17 3053
rect 17 3019 33 3053
rect -33 3003 33 3019
rect -15 2981 15 3003
rect -15 2559 15 2581
rect -33 2543 33 2559
rect -33 2509 -17 2543
rect 17 2509 33 2543
rect -33 2493 33 2509
rect -33 2435 33 2451
rect -33 2401 -17 2435
rect 17 2401 33 2435
rect -33 2385 33 2401
rect -15 2363 15 2385
rect -15 1941 15 1963
rect -33 1925 33 1941
rect -33 1891 -17 1925
rect 17 1891 33 1925
rect -33 1875 33 1891
rect -33 1817 33 1833
rect -33 1783 -17 1817
rect 17 1783 33 1817
rect -33 1767 33 1783
rect -15 1745 15 1767
rect -15 1323 15 1345
rect -33 1307 33 1323
rect -33 1273 -17 1307
rect 17 1273 33 1307
rect -33 1257 33 1273
rect -33 1199 33 1215
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -33 1149 33 1165
rect -15 1127 15 1149
rect -15 705 15 727
rect -33 689 33 705
rect -33 655 -17 689
rect 17 655 33 689
rect -33 639 33 655
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect -15 509 15 531
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -531 15 -509
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect -33 -655 33 -639
rect -33 -689 -17 -655
rect 17 -689 33 -655
rect -33 -705 33 -689
rect -15 -727 15 -705
rect -15 -1149 15 -1127
rect -33 -1165 33 -1149
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -33 -1215 33 -1199
rect -33 -1273 33 -1257
rect -33 -1307 -17 -1273
rect 17 -1307 33 -1273
rect -33 -1323 33 -1307
rect -15 -1345 15 -1323
rect -15 -1767 15 -1745
rect -33 -1783 33 -1767
rect -33 -1817 -17 -1783
rect 17 -1817 33 -1783
rect -33 -1833 33 -1817
rect -33 -1891 33 -1875
rect -33 -1925 -17 -1891
rect 17 -1925 33 -1891
rect -33 -1941 33 -1925
rect -15 -1963 15 -1941
rect -15 -2385 15 -2363
rect -33 -2401 33 -2385
rect -33 -2435 -17 -2401
rect 17 -2435 33 -2401
rect -33 -2451 33 -2435
rect -33 -2509 33 -2493
rect -33 -2543 -17 -2509
rect 17 -2543 33 -2509
rect -33 -2559 33 -2543
rect -15 -2581 15 -2559
rect -15 -3003 15 -2981
rect -33 -3019 33 -3003
rect -33 -3053 -17 -3019
rect 17 -3053 33 -3019
rect -33 -3069 33 -3053
rect -33 -3127 33 -3111
rect -33 -3161 -17 -3127
rect 17 -3161 33 -3127
rect -33 -3177 33 -3161
rect -15 -3199 15 -3177
rect -15 -3621 15 -3599
rect -33 -3637 33 -3621
rect -33 -3671 -17 -3637
rect 17 -3671 33 -3637
rect -33 -3687 33 -3671
rect -33 -3745 33 -3729
rect -33 -3779 -17 -3745
rect 17 -3779 33 -3745
rect -33 -3795 33 -3779
rect -15 -3817 15 -3795
rect -15 -4239 15 -4217
rect -33 -4255 33 -4239
rect -33 -4289 -17 -4255
rect 17 -4289 33 -4255
rect -33 -4305 33 -4289
rect -33 -4363 33 -4347
rect -33 -4397 -17 -4363
rect 17 -4397 33 -4363
rect -33 -4413 33 -4397
rect -15 -4435 15 -4413
rect -15 -4857 15 -4835
rect -33 -4873 33 -4857
rect -33 -4907 -17 -4873
rect 17 -4907 33 -4873
rect -33 -4923 33 -4907
rect -33 -4981 33 -4965
rect -33 -5015 -17 -4981
rect 17 -5015 33 -4981
rect -33 -5031 33 -5015
rect -15 -5053 15 -5031
rect -15 -5475 15 -5453
rect -33 -5491 33 -5475
rect -33 -5525 -17 -5491
rect 17 -5525 33 -5491
rect -33 -5541 33 -5525
rect -33 -5599 33 -5583
rect -33 -5633 -17 -5599
rect 17 -5633 33 -5599
rect -33 -5649 33 -5633
rect -15 -5671 15 -5649
rect -15 -6093 15 -6071
rect -33 -6109 33 -6093
rect -33 -6143 -17 -6109
rect 17 -6143 33 -6109
rect -33 -6159 33 -6143
rect -33 -6217 33 -6201
rect -33 -6251 -17 -6217
rect 17 -6251 33 -6217
rect -33 -6267 33 -6251
rect -15 -6289 15 -6267
rect -15 -6711 15 -6689
rect -33 -6727 33 -6711
rect -33 -6761 -17 -6727
rect 17 -6761 33 -6727
rect -33 -6777 33 -6761
rect -33 -6835 33 -6819
rect -33 -6869 -17 -6835
rect 17 -6869 33 -6835
rect -33 -6885 33 -6869
rect -15 -6907 15 -6885
rect -15 -7329 15 -7307
rect -33 -7345 33 -7329
rect -33 -7379 -17 -7345
rect 17 -7379 33 -7345
rect -33 -7395 33 -7379
rect -33 -7453 33 -7437
rect -33 -7487 -17 -7453
rect 17 -7487 33 -7453
rect -33 -7503 33 -7487
rect -15 -7525 15 -7503
rect -15 -7947 15 -7925
rect -33 -7963 33 -7947
rect -33 -7997 -17 -7963
rect 17 -7997 33 -7963
rect -33 -8013 33 -7997
rect -33 -8071 33 -8055
rect -33 -8105 -17 -8071
rect 17 -8105 33 -8071
rect -33 -8121 33 -8105
rect -15 -8143 15 -8121
rect -15 -8565 15 -8543
rect -33 -8581 33 -8565
rect -33 -8615 -17 -8581
rect 17 -8615 33 -8581
rect -33 -8631 33 -8615
rect -33 -8689 33 -8673
rect -33 -8723 -17 -8689
rect 17 -8723 33 -8689
rect -33 -8739 33 -8723
rect -15 -8761 15 -8739
rect -15 -9183 15 -9161
rect -33 -9199 33 -9183
rect -33 -9233 -17 -9199
rect 17 -9233 33 -9199
rect -33 -9249 33 -9233
<< polycont >>
rect -17 9199 17 9233
rect -17 8689 17 8723
rect -17 8581 17 8615
rect -17 8071 17 8105
rect -17 7963 17 7997
rect -17 7453 17 7487
rect -17 7345 17 7379
rect -17 6835 17 6869
rect -17 6727 17 6761
rect -17 6217 17 6251
rect -17 6109 17 6143
rect -17 5599 17 5633
rect -17 5491 17 5525
rect -17 4981 17 5015
rect -17 4873 17 4907
rect -17 4363 17 4397
rect -17 4255 17 4289
rect -17 3745 17 3779
rect -17 3637 17 3671
rect -17 3127 17 3161
rect -17 3019 17 3053
rect -17 2509 17 2543
rect -17 2401 17 2435
rect -17 1891 17 1925
rect -17 1783 17 1817
rect -17 1273 17 1307
rect -17 1165 17 1199
rect -17 655 17 689
rect -17 547 17 581
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -581 17 -547
rect -17 -689 17 -655
rect -17 -1199 17 -1165
rect -17 -1307 17 -1273
rect -17 -1817 17 -1783
rect -17 -1925 17 -1891
rect -17 -2435 17 -2401
rect -17 -2543 17 -2509
rect -17 -3053 17 -3019
rect -17 -3161 17 -3127
rect -17 -3671 17 -3637
rect -17 -3779 17 -3745
rect -17 -4289 17 -4255
rect -17 -4397 17 -4363
rect -17 -4907 17 -4873
rect -17 -5015 17 -4981
rect -17 -5525 17 -5491
rect -17 -5633 17 -5599
rect -17 -6143 17 -6109
rect -17 -6251 17 -6217
rect -17 -6761 17 -6727
rect -17 -6869 17 -6835
rect -17 -7379 17 -7345
rect -17 -7487 17 -7453
rect -17 -7997 17 -7963
rect -17 -8105 17 -8071
rect -17 -8615 17 -8581
rect -17 -8723 17 -8689
rect -17 -9233 17 -9199
<< locali >>
rect -175 9301 -79 9335
rect 79 9301 175 9335
rect -175 9239 -141 9301
rect 141 9239 175 9301
rect -33 9199 -17 9233
rect 17 9199 33 9233
rect -61 9149 -27 9165
rect -61 8757 -27 8773
rect 27 9149 61 9165
rect 27 8757 61 8773
rect -33 8689 -17 8723
rect 17 8689 33 8723
rect -33 8581 -17 8615
rect 17 8581 33 8615
rect -61 8531 -27 8547
rect -61 8139 -27 8155
rect 27 8531 61 8547
rect 27 8139 61 8155
rect -33 8071 -17 8105
rect 17 8071 33 8105
rect -33 7963 -17 7997
rect 17 7963 33 7997
rect -61 7913 -27 7929
rect -61 7521 -27 7537
rect 27 7913 61 7929
rect 27 7521 61 7537
rect -33 7453 -17 7487
rect 17 7453 33 7487
rect -33 7345 -17 7379
rect 17 7345 33 7379
rect -61 7295 -27 7311
rect -61 6903 -27 6919
rect 27 7295 61 7311
rect 27 6903 61 6919
rect -33 6835 -17 6869
rect 17 6835 33 6869
rect -33 6727 -17 6761
rect 17 6727 33 6761
rect -61 6677 -27 6693
rect -61 6285 -27 6301
rect 27 6677 61 6693
rect 27 6285 61 6301
rect -33 6217 -17 6251
rect 17 6217 33 6251
rect -33 6109 -17 6143
rect 17 6109 33 6143
rect -61 6059 -27 6075
rect -61 5667 -27 5683
rect 27 6059 61 6075
rect 27 5667 61 5683
rect -33 5599 -17 5633
rect 17 5599 33 5633
rect -33 5491 -17 5525
rect 17 5491 33 5525
rect -61 5441 -27 5457
rect -61 5049 -27 5065
rect 27 5441 61 5457
rect 27 5049 61 5065
rect -33 4981 -17 5015
rect 17 4981 33 5015
rect -33 4873 -17 4907
rect 17 4873 33 4907
rect -61 4823 -27 4839
rect -61 4431 -27 4447
rect 27 4823 61 4839
rect 27 4431 61 4447
rect -33 4363 -17 4397
rect 17 4363 33 4397
rect -33 4255 -17 4289
rect 17 4255 33 4289
rect -61 4205 -27 4221
rect -61 3813 -27 3829
rect 27 4205 61 4221
rect 27 3813 61 3829
rect -33 3745 -17 3779
rect 17 3745 33 3779
rect -33 3637 -17 3671
rect 17 3637 33 3671
rect -61 3587 -27 3603
rect -61 3195 -27 3211
rect 27 3587 61 3603
rect 27 3195 61 3211
rect -33 3127 -17 3161
rect 17 3127 33 3161
rect -33 3019 -17 3053
rect 17 3019 33 3053
rect -61 2969 -27 2985
rect -61 2577 -27 2593
rect 27 2969 61 2985
rect 27 2577 61 2593
rect -33 2509 -17 2543
rect 17 2509 33 2543
rect -33 2401 -17 2435
rect 17 2401 33 2435
rect -61 2351 -27 2367
rect -61 1959 -27 1975
rect 27 2351 61 2367
rect 27 1959 61 1975
rect -33 1891 -17 1925
rect 17 1891 33 1925
rect -33 1783 -17 1817
rect 17 1783 33 1817
rect -61 1733 -27 1749
rect -61 1341 -27 1357
rect 27 1733 61 1749
rect 27 1341 61 1357
rect -33 1273 -17 1307
rect 17 1273 33 1307
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -61 1115 -27 1131
rect -61 723 -27 739
rect 27 1115 61 1131
rect 27 723 61 739
rect -33 655 -17 689
rect 17 655 33 689
rect -33 547 -17 581
rect 17 547 33 581
rect -61 497 -27 513
rect -61 105 -27 121
rect 27 497 61 513
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -513 -27 -497
rect 27 -121 61 -105
rect 27 -513 61 -497
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -689 -17 -655
rect 17 -689 33 -655
rect -61 -739 -27 -723
rect -61 -1131 -27 -1115
rect 27 -739 61 -723
rect 27 -1131 61 -1115
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -33 -1307 -17 -1273
rect 17 -1307 33 -1273
rect -61 -1357 -27 -1341
rect -61 -1749 -27 -1733
rect 27 -1357 61 -1341
rect 27 -1749 61 -1733
rect -33 -1817 -17 -1783
rect 17 -1817 33 -1783
rect -33 -1925 -17 -1891
rect 17 -1925 33 -1891
rect -61 -1975 -27 -1959
rect -61 -2367 -27 -2351
rect 27 -1975 61 -1959
rect 27 -2367 61 -2351
rect -33 -2435 -17 -2401
rect 17 -2435 33 -2401
rect -33 -2543 -17 -2509
rect 17 -2543 33 -2509
rect -61 -2593 -27 -2577
rect -61 -2985 -27 -2969
rect 27 -2593 61 -2577
rect 27 -2985 61 -2969
rect -33 -3053 -17 -3019
rect 17 -3053 33 -3019
rect -33 -3161 -17 -3127
rect 17 -3161 33 -3127
rect -61 -3211 -27 -3195
rect -61 -3603 -27 -3587
rect 27 -3211 61 -3195
rect 27 -3603 61 -3587
rect -33 -3671 -17 -3637
rect 17 -3671 33 -3637
rect -33 -3779 -17 -3745
rect 17 -3779 33 -3745
rect -61 -3829 -27 -3813
rect -61 -4221 -27 -4205
rect 27 -3829 61 -3813
rect 27 -4221 61 -4205
rect -33 -4289 -17 -4255
rect 17 -4289 33 -4255
rect -33 -4397 -17 -4363
rect 17 -4397 33 -4363
rect -61 -4447 -27 -4431
rect -61 -4839 -27 -4823
rect 27 -4447 61 -4431
rect 27 -4839 61 -4823
rect -33 -4907 -17 -4873
rect 17 -4907 33 -4873
rect -33 -5015 -17 -4981
rect 17 -5015 33 -4981
rect -61 -5065 -27 -5049
rect -61 -5457 -27 -5441
rect 27 -5065 61 -5049
rect 27 -5457 61 -5441
rect -33 -5525 -17 -5491
rect 17 -5525 33 -5491
rect -33 -5633 -17 -5599
rect 17 -5633 33 -5599
rect -61 -5683 -27 -5667
rect -61 -6075 -27 -6059
rect 27 -5683 61 -5667
rect 27 -6075 61 -6059
rect -33 -6143 -17 -6109
rect 17 -6143 33 -6109
rect -33 -6251 -17 -6217
rect 17 -6251 33 -6217
rect -61 -6301 -27 -6285
rect -61 -6693 -27 -6677
rect 27 -6301 61 -6285
rect 27 -6693 61 -6677
rect -33 -6761 -17 -6727
rect 17 -6761 33 -6727
rect -33 -6869 -17 -6835
rect 17 -6869 33 -6835
rect -61 -6919 -27 -6903
rect -61 -7311 -27 -7295
rect 27 -6919 61 -6903
rect 27 -7311 61 -7295
rect -33 -7379 -17 -7345
rect 17 -7379 33 -7345
rect -33 -7487 -17 -7453
rect 17 -7487 33 -7453
rect -61 -7537 -27 -7521
rect -61 -7929 -27 -7913
rect 27 -7537 61 -7521
rect 27 -7929 61 -7913
rect -33 -7997 -17 -7963
rect 17 -7997 33 -7963
rect -33 -8105 -17 -8071
rect 17 -8105 33 -8071
rect -61 -8155 -27 -8139
rect -61 -8547 -27 -8531
rect 27 -8155 61 -8139
rect 27 -8547 61 -8531
rect -33 -8615 -17 -8581
rect 17 -8615 33 -8581
rect -33 -8723 -17 -8689
rect 17 -8723 33 -8689
rect -61 -8773 -27 -8757
rect -61 -9165 -27 -9149
rect 27 -8773 61 -8757
rect 27 -9165 61 -9149
rect -33 -9233 -17 -9199
rect 17 -9233 33 -9199
rect -175 -9301 -141 -9239
rect 141 -9301 175 -9239
rect -175 -9335 -79 -9301
rect 79 -9335 175 -9301
<< viali >>
rect -17 9199 17 9233
rect -61 8773 -27 9149
rect 27 8773 61 9149
rect -17 8689 17 8723
rect -17 8581 17 8615
rect -61 8155 -27 8531
rect 27 8155 61 8531
rect -17 8071 17 8105
rect -17 7963 17 7997
rect -61 7537 -27 7913
rect 27 7537 61 7913
rect -17 7453 17 7487
rect -17 7345 17 7379
rect -61 6919 -27 7295
rect 27 6919 61 7295
rect -17 6835 17 6869
rect -17 6727 17 6761
rect -61 6301 -27 6677
rect 27 6301 61 6677
rect -17 6217 17 6251
rect -17 6109 17 6143
rect -61 5683 -27 6059
rect 27 5683 61 6059
rect -17 5599 17 5633
rect -17 5491 17 5525
rect -61 5065 -27 5441
rect 27 5065 61 5441
rect -17 4981 17 5015
rect -17 4873 17 4907
rect -61 4447 -27 4823
rect 27 4447 61 4823
rect -17 4363 17 4397
rect -17 4255 17 4289
rect -61 3829 -27 4205
rect 27 3829 61 4205
rect -17 3745 17 3779
rect -17 3637 17 3671
rect -61 3211 -27 3587
rect 27 3211 61 3587
rect -17 3127 17 3161
rect -17 3019 17 3053
rect -61 2593 -27 2969
rect 27 2593 61 2969
rect -17 2509 17 2543
rect -17 2401 17 2435
rect -61 1975 -27 2351
rect 27 1975 61 2351
rect -17 1891 17 1925
rect -17 1783 17 1817
rect -61 1357 -27 1733
rect 27 1357 61 1733
rect -17 1273 17 1307
rect -17 1165 17 1199
rect -61 739 -27 1115
rect 27 739 61 1115
rect -17 655 17 689
rect -17 547 17 581
rect -61 121 -27 497
rect 27 121 61 497
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -497 -27 -121
rect 27 -497 61 -121
rect -17 -581 17 -547
rect -17 -689 17 -655
rect -61 -1115 -27 -739
rect 27 -1115 61 -739
rect -17 -1199 17 -1165
rect -17 -1307 17 -1273
rect -61 -1733 -27 -1357
rect 27 -1733 61 -1357
rect -17 -1817 17 -1783
rect -17 -1925 17 -1891
rect -61 -2351 -27 -1975
rect 27 -2351 61 -1975
rect -17 -2435 17 -2401
rect -17 -2543 17 -2509
rect -61 -2969 -27 -2593
rect 27 -2969 61 -2593
rect -17 -3053 17 -3019
rect -17 -3161 17 -3127
rect -61 -3587 -27 -3211
rect 27 -3587 61 -3211
rect -17 -3671 17 -3637
rect -17 -3779 17 -3745
rect -61 -4205 -27 -3829
rect 27 -4205 61 -3829
rect -17 -4289 17 -4255
rect -17 -4397 17 -4363
rect -61 -4823 -27 -4447
rect 27 -4823 61 -4447
rect -17 -4907 17 -4873
rect -17 -5015 17 -4981
rect -61 -5441 -27 -5065
rect 27 -5441 61 -5065
rect -17 -5525 17 -5491
rect -17 -5633 17 -5599
rect -61 -6059 -27 -5683
rect 27 -6059 61 -5683
rect -17 -6143 17 -6109
rect -17 -6251 17 -6217
rect -61 -6677 -27 -6301
rect 27 -6677 61 -6301
rect -17 -6761 17 -6727
rect -17 -6869 17 -6835
rect -61 -7295 -27 -6919
rect 27 -7295 61 -6919
rect -17 -7379 17 -7345
rect -17 -7487 17 -7453
rect -61 -7913 -27 -7537
rect 27 -7913 61 -7537
rect -17 -7997 17 -7963
rect -17 -8105 17 -8071
rect -61 -8531 -27 -8155
rect 27 -8531 61 -8155
rect -17 -8615 17 -8581
rect -17 -8723 17 -8689
rect -61 -9149 -27 -8773
rect 27 -9149 61 -8773
rect -17 -9233 17 -9199
<< metal1 >>
rect -29 9233 29 9239
rect -29 9199 -17 9233
rect 17 9199 29 9233
rect -29 9193 29 9199
rect -67 9149 -21 9161
rect -67 8773 -61 9149
rect -27 8773 -21 9149
rect -67 8761 -21 8773
rect 21 9149 67 9161
rect 21 8773 27 9149
rect 61 8773 67 9149
rect 21 8761 67 8773
rect -29 8723 29 8729
rect -29 8689 -17 8723
rect 17 8689 29 8723
rect -29 8683 29 8689
rect -29 8615 29 8621
rect -29 8581 -17 8615
rect 17 8581 29 8615
rect -29 8575 29 8581
rect -67 8531 -21 8543
rect -67 8155 -61 8531
rect -27 8155 -21 8531
rect -67 8143 -21 8155
rect 21 8531 67 8543
rect 21 8155 27 8531
rect 61 8155 67 8531
rect 21 8143 67 8155
rect -29 8105 29 8111
rect -29 8071 -17 8105
rect 17 8071 29 8105
rect -29 8065 29 8071
rect -29 7997 29 8003
rect -29 7963 -17 7997
rect 17 7963 29 7997
rect -29 7957 29 7963
rect -67 7913 -21 7925
rect -67 7537 -61 7913
rect -27 7537 -21 7913
rect -67 7525 -21 7537
rect 21 7913 67 7925
rect 21 7537 27 7913
rect 61 7537 67 7913
rect 21 7525 67 7537
rect -29 7487 29 7493
rect -29 7453 -17 7487
rect 17 7453 29 7487
rect -29 7447 29 7453
rect -29 7379 29 7385
rect -29 7345 -17 7379
rect 17 7345 29 7379
rect -29 7339 29 7345
rect -67 7295 -21 7307
rect -67 6919 -61 7295
rect -27 6919 -21 7295
rect -67 6907 -21 6919
rect 21 7295 67 7307
rect 21 6919 27 7295
rect 61 6919 67 7295
rect 21 6907 67 6919
rect -29 6869 29 6875
rect -29 6835 -17 6869
rect 17 6835 29 6869
rect -29 6829 29 6835
rect -29 6761 29 6767
rect -29 6727 -17 6761
rect 17 6727 29 6761
rect -29 6721 29 6727
rect -67 6677 -21 6689
rect -67 6301 -61 6677
rect -27 6301 -21 6677
rect -67 6289 -21 6301
rect 21 6677 67 6689
rect 21 6301 27 6677
rect 61 6301 67 6677
rect 21 6289 67 6301
rect -29 6251 29 6257
rect -29 6217 -17 6251
rect 17 6217 29 6251
rect -29 6211 29 6217
rect -29 6143 29 6149
rect -29 6109 -17 6143
rect 17 6109 29 6143
rect -29 6103 29 6109
rect -67 6059 -21 6071
rect -67 5683 -61 6059
rect -27 5683 -21 6059
rect -67 5671 -21 5683
rect 21 6059 67 6071
rect 21 5683 27 6059
rect 61 5683 67 6059
rect 21 5671 67 5683
rect -29 5633 29 5639
rect -29 5599 -17 5633
rect 17 5599 29 5633
rect -29 5593 29 5599
rect -29 5525 29 5531
rect -29 5491 -17 5525
rect 17 5491 29 5525
rect -29 5485 29 5491
rect -67 5441 -21 5453
rect -67 5065 -61 5441
rect -27 5065 -21 5441
rect -67 5053 -21 5065
rect 21 5441 67 5453
rect 21 5065 27 5441
rect 61 5065 67 5441
rect 21 5053 67 5065
rect -29 5015 29 5021
rect -29 4981 -17 5015
rect 17 4981 29 5015
rect -29 4975 29 4981
rect -29 4907 29 4913
rect -29 4873 -17 4907
rect 17 4873 29 4907
rect -29 4867 29 4873
rect -67 4823 -21 4835
rect -67 4447 -61 4823
rect -27 4447 -21 4823
rect -67 4435 -21 4447
rect 21 4823 67 4835
rect 21 4447 27 4823
rect 61 4447 67 4823
rect 21 4435 67 4447
rect -29 4397 29 4403
rect -29 4363 -17 4397
rect 17 4363 29 4397
rect -29 4357 29 4363
rect -29 4289 29 4295
rect -29 4255 -17 4289
rect 17 4255 29 4289
rect -29 4249 29 4255
rect -67 4205 -21 4217
rect -67 3829 -61 4205
rect -27 3829 -21 4205
rect -67 3817 -21 3829
rect 21 4205 67 4217
rect 21 3829 27 4205
rect 61 3829 67 4205
rect 21 3817 67 3829
rect -29 3779 29 3785
rect -29 3745 -17 3779
rect 17 3745 29 3779
rect -29 3739 29 3745
rect -29 3671 29 3677
rect -29 3637 -17 3671
rect 17 3637 29 3671
rect -29 3631 29 3637
rect -67 3587 -21 3599
rect -67 3211 -61 3587
rect -27 3211 -21 3587
rect -67 3199 -21 3211
rect 21 3587 67 3599
rect 21 3211 27 3587
rect 61 3211 67 3587
rect 21 3199 67 3211
rect -29 3161 29 3167
rect -29 3127 -17 3161
rect 17 3127 29 3161
rect -29 3121 29 3127
rect -29 3053 29 3059
rect -29 3019 -17 3053
rect 17 3019 29 3053
rect -29 3013 29 3019
rect -67 2969 -21 2981
rect -67 2593 -61 2969
rect -27 2593 -21 2969
rect -67 2581 -21 2593
rect 21 2969 67 2981
rect 21 2593 27 2969
rect 61 2593 67 2969
rect 21 2581 67 2593
rect -29 2543 29 2549
rect -29 2509 -17 2543
rect 17 2509 29 2543
rect -29 2503 29 2509
rect -29 2435 29 2441
rect -29 2401 -17 2435
rect 17 2401 29 2435
rect -29 2395 29 2401
rect -67 2351 -21 2363
rect -67 1975 -61 2351
rect -27 1975 -21 2351
rect -67 1963 -21 1975
rect 21 2351 67 2363
rect 21 1975 27 2351
rect 61 1975 67 2351
rect 21 1963 67 1975
rect -29 1925 29 1931
rect -29 1891 -17 1925
rect 17 1891 29 1925
rect -29 1885 29 1891
rect -29 1817 29 1823
rect -29 1783 -17 1817
rect 17 1783 29 1817
rect -29 1777 29 1783
rect -67 1733 -21 1745
rect -67 1357 -61 1733
rect -27 1357 -21 1733
rect -67 1345 -21 1357
rect 21 1733 67 1745
rect 21 1357 27 1733
rect 61 1357 67 1733
rect 21 1345 67 1357
rect -29 1307 29 1313
rect -29 1273 -17 1307
rect 17 1273 29 1307
rect -29 1267 29 1273
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect 17 1165 29 1199
rect -29 1159 29 1165
rect -67 1115 -21 1127
rect -67 739 -61 1115
rect -27 739 -21 1115
rect -67 727 -21 739
rect 21 1115 67 1127
rect 21 739 27 1115
rect 61 739 67 1115
rect 21 727 67 739
rect -29 689 29 695
rect -29 655 -17 689
rect 17 655 29 689
rect -29 649 29 655
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -67 497 -21 509
rect -67 121 -61 497
rect -27 121 -21 497
rect -67 109 -21 121
rect 21 497 67 509
rect 21 121 27 497
rect 61 121 67 497
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -497 -61 -121
rect -27 -497 -21 -121
rect -67 -509 -21 -497
rect 21 -121 67 -109
rect 21 -497 27 -121
rect 61 -497 67 -121
rect 21 -509 67 -497
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect -29 -655 29 -649
rect -29 -689 -17 -655
rect 17 -689 29 -655
rect -29 -695 29 -689
rect -67 -739 -21 -727
rect -67 -1115 -61 -739
rect -27 -1115 -21 -739
rect -67 -1127 -21 -1115
rect 21 -739 67 -727
rect 21 -1115 27 -739
rect 61 -1115 67 -739
rect 21 -1127 67 -1115
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect 17 -1199 29 -1165
rect -29 -1205 29 -1199
rect -29 -1273 29 -1267
rect -29 -1307 -17 -1273
rect 17 -1307 29 -1273
rect -29 -1313 29 -1307
rect -67 -1357 -21 -1345
rect -67 -1733 -61 -1357
rect -27 -1733 -21 -1357
rect -67 -1745 -21 -1733
rect 21 -1357 67 -1345
rect 21 -1733 27 -1357
rect 61 -1733 67 -1357
rect 21 -1745 67 -1733
rect -29 -1783 29 -1777
rect -29 -1817 -17 -1783
rect 17 -1817 29 -1783
rect -29 -1823 29 -1817
rect -29 -1891 29 -1885
rect -29 -1925 -17 -1891
rect 17 -1925 29 -1891
rect -29 -1931 29 -1925
rect -67 -1975 -21 -1963
rect -67 -2351 -61 -1975
rect -27 -2351 -21 -1975
rect -67 -2363 -21 -2351
rect 21 -1975 67 -1963
rect 21 -2351 27 -1975
rect 61 -2351 67 -1975
rect 21 -2363 67 -2351
rect -29 -2401 29 -2395
rect -29 -2435 -17 -2401
rect 17 -2435 29 -2401
rect -29 -2441 29 -2435
rect -29 -2509 29 -2503
rect -29 -2543 -17 -2509
rect 17 -2543 29 -2509
rect -29 -2549 29 -2543
rect -67 -2593 -21 -2581
rect -67 -2969 -61 -2593
rect -27 -2969 -21 -2593
rect -67 -2981 -21 -2969
rect 21 -2593 67 -2581
rect 21 -2969 27 -2593
rect 61 -2969 67 -2593
rect 21 -2981 67 -2969
rect -29 -3019 29 -3013
rect -29 -3053 -17 -3019
rect 17 -3053 29 -3019
rect -29 -3059 29 -3053
rect -29 -3127 29 -3121
rect -29 -3161 -17 -3127
rect 17 -3161 29 -3127
rect -29 -3167 29 -3161
rect -67 -3211 -21 -3199
rect -67 -3587 -61 -3211
rect -27 -3587 -21 -3211
rect -67 -3599 -21 -3587
rect 21 -3211 67 -3199
rect 21 -3587 27 -3211
rect 61 -3587 67 -3211
rect 21 -3599 67 -3587
rect -29 -3637 29 -3631
rect -29 -3671 -17 -3637
rect 17 -3671 29 -3637
rect -29 -3677 29 -3671
rect -29 -3745 29 -3739
rect -29 -3779 -17 -3745
rect 17 -3779 29 -3745
rect -29 -3785 29 -3779
rect -67 -3829 -21 -3817
rect -67 -4205 -61 -3829
rect -27 -4205 -21 -3829
rect -67 -4217 -21 -4205
rect 21 -3829 67 -3817
rect 21 -4205 27 -3829
rect 61 -4205 67 -3829
rect 21 -4217 67 -4205
rect -29 -4255 29 -4249
rect -29 -4289 -17 -4255
rect 17 -4289 29 -4255
rect -29 -4295 29 -4289
rect -29 -4363 29 -4357
rect -29 -4397 -17 -4363
rect 17 -4397 29 -4363
rect -29 -4403 29 -4397
rect -67 -4447 -21 -4435
rect -67 -4823 -61 -4447
rect -27 -4823 -21 -4447
rect -67 -4835 -21 -4823
rect 21 -4447 67 -4435
rect 21 -4823 27 -4447
rect 61 -4823 67 -4447
rect 21 -4835 67 -4823
rect -29 -4873 29 -4867
rect -29 -4907 -17 -4873
rect 17 -4907 29 -4873
rect -29 -4913 29 -4907
rect -29 -4981 29 -4975
rect -29 -5015 -17 -4981
rect 17 -5015 29 -4981
rect -29 -5021 29 -5015
rect -67 -5065 -21 -5053
rect -67 -5441 -61 -5065
rect -27 -5441 -21 -5065
rect -67 -5453 -21 -5441
rect 21 -5065 67 -5053
rect 21 -5441 27 -5065
rect 61 -5441 67 -5065
rect 21 -5453 67 -5441
rect -29 -5491 29 -5485
rect -29 -5525 -17 -5491
rect 17 -5525 29 -5491
rect -29 -5531 29 -5525
rect -29 -5599 29 -5593
rect -29 -5633 -17 -5599
rect 17 -5633 29 -5599
rect -29 -5639 29 -5633
rect -67 -5683 -21 -5671
rect -67 -6059 -61 -5683
rect -27 -6059 -21 -5683
rect -67 -6071 -21 -6059
rect 21 -5683 67 -5671
rect 21 -6059 27 -5683
rect 61 -6059 67 -5683
rect 21 -6071 67 -6059
rect -29 -6109 29 -6103
rect -29 -6143 -17 -6109
rect 17 -6143 29 -6109
rect -29 -6149 29 -6143
rect -29 -6217 29 -6211
rect -29 -6251 -17 -6217
rect 17 -6251 29 -6217
rect -29 -6257 29 -6251
rect -67 -6301 -21 -6289
rect -67 -6677 -61 -6301
rect -27 -6677 -21 -6301
rect -67 -6689 -21 -6677
rect 21 -6301 67 -6289
rect 21 -6677 27 -6301
rect 61 -6677 67 -6301
rect 21 -6689 67 -6677
rect -29 -6727 29 -6721
rect -29 -6761 -17 -6727
rect 17 -6761 29 -6727
rect -29 -6767 29 -6761
rect -29 -6835 29 -6829
rect -29 -6869 -17 -6835
rect 17 -6869 29 -6835
rect -29 -6875 29 -6869
rect -67 -6919 -21 -6907
rect -67 -7295 -61 -6919
rect -27 -7295 -21 -6919
rect -67 -7307 -21 -7295
rect 21 -6919 67 -6907
rect 21 -7295 27 -6919
rect 61 -7295 67 -6919
rect 21 -7307 67 -7295
rect -29 -7345 29 -7339
rect -29 -7379 -17 -7345
rect 17 -7379 29 -7345
rect -29 -7385 29 -7379
rect -29 -7453 29 -7447
rect -29 -7487 -17 -7453
rect 17 -7487 29 -7453
rect -29 -7493 29 -7487
rect -67 -7537 -21 -7525
rect -67 -7913 -61 -7537
rect -27 -7913 -21 -7537
rect -67 -7925 -21 -7913
rect 21 -7537 67 -7525
rect 21 -7913 27 -7537
rect 61 -7913 67 -7537
rect 21 -7925 67 -7913
rect -29 -7963 29 -7957
rect -29 -7997 -17 -7963
rect 17 -7997 29 -7963
rect -29 -8003 29 -7997
rect -29 -8071 29 -8065
rect -29 -8105 -17 -8071
rect 17 -8105 29 -8071
rect -29 -8111 29 -8105
rect -67 -8155 -21 -8143
rect -67 -8531 -61 -8155
rect -27 -8531 -21 -8155
rect -67 -8543 -21 -8531
rect 21 -8155 67 -8143
rect 21 -8531 27 -8155
rect 61 -8531 67 -8155
rect 21 -8543 67 -8531
rect -29 -8581 29 -8575
rect -29 -8615 -17 -8581
rect 17 -8615 29 -8581
rect -29 -8621 29 -8615
rect -29 -8689 29 -8683
rect -29 -8723 -17 -8689
rect 17 -8723 29 -8689
rect -29 -8729 29 -8723
rect -67 -8773 -21 -8761
rect -67 -9149 -61 -8773
rect -27 -9149 -21 -8773
rect -67 -9161 -21 -9149
rect 21 -8773 67 -8761
rect 21 -9149 27 -8773
rect 61 -9149 67 -8773
rect 21 -9161 67 -9149
rect -29 -9199 29 -9193
rect -29 -9233 -17 -9199
rect 17 -9233 29 -9199
rect -29 -9239 29 -9233
<< properties >>
string FIXED_BBOX -158 -9318 158 9318
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 30 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
