magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< error_p >>
rect -701 599 -643 605
rect -509 599 -451 605
rect -317 599 -259 605
rect -125 599 -67 605
rect 67 599 125 605
rect 259 599 317 605
rect 451 599 509 605
rect 643 599 701 605
rect -701 565 -689 599
rect -509 565 -497 599
rect -317 565 -305 599
rect -125 565 -113 599
rect 67 565 79 599
rect 259 565 271 599
rect 451 565 463 599
rect 643 565 655 599
rect -701 559 -643 565
rect -509 559 -451 565
rect -317 559 -259 565
rect -125 559 -67 565
rect 67 559 125 565
rect 259 559 317 565
rect 451 559 509 565
rect 643 559 701 565
rect -605 71 -547 77
rect -413 71 -355 77
rect -221 71 -163 77
rect -29 71 29 77
rect 163 71 221 77
rect 355 71 413 77
rect 547 71 605 77
rect -605 37 -593 71
rect -413 37 -401 71
rect -221 37 -209 71
rect -29 37 -17 71
rect 163 37 175 71
rect 355 37 367 71
rect 547 37 559 71
rect -605 31 -547 37
rect -413 31 -355 37
rect -221 31 -163 37
rect -29 31 29 37
rect 163 31 221 37
rect 355 31 413 37
rect 547 31 605 37
rect -605 -37 -547 -31
rect -413 -37 -355 -31
rect -221 -37 -163 -31
rect -29 -37 29 -31
rect 163 -37 221 -31
rect 355 -37 413 -31
rect 547 -37 605 -31
rect -605 -71 -593 -37
rect -413 -71 -401 -37
rect -221 -71 -209 -37
rect -29 -71 -17 -37
rect 163 -71 175 -37
rect 355 -71 367 -37
rect 547 -71 559 -37
rect -605 -77 -547 -71
rect -413 -77 -355 -71
rect -221 -77 -163 -71
rect -29 -77 29 -71
rect 163 -77 221 -71
rect 355 -77 413 -71
rect 547 -77 605 -71
rect -701 -565 -643 -559
rect -509 -565 -451 -559
rect -317 -565 -259 -559
rect -125 -565 -67 -559
rect 67 -565 125 -559
rect 259 -565 317 -559
rect 451 -565 509 -559
rect 643 -565 701 -559
rect -701 -599 -689 -565
rect -509 -599 -497 -565
rect -317 -599 -305 -565
rect -125 -599 -113 -565
rect 67 -599 79 -565
rect 259 -599 271 -565
rect 451 -599 463 -565
rect 643 -599 655 -565
rect -701 -605 -643 -599
rect -509 -605 -451 -599
rect -317 -605 -259 -599
rect -125 -605 -67 -599
rect 67 -605 125 -599
rect 259 -605 317 -599
rect 451 -605 509 -599
rect 643 -605 701 -599
<< nwell >>
rect -887 -737 887 737
<< pmos >>
rect -687 118 -657 518
rect -591 118 -561 518
rect -495 118 -465 518
rect -399 118 -369 518
rect -303 118 -273 518
rect -207 118 -177 518
rect -111 118 -81 518
rect -15 118 15 518
rect 81 118 111 518
rect 177 118 207 518
rect 273 118 303 518
rect 369 118 399 518
rect 465 118 495 518
rect 561 118 591 518
rect 657 118 687 518
rect -687 -518 -657 -118
rect -591 -518 -561 -118
rect -495 -518 -465 -118
rect -399 -518 -369 -118
rect -303 -518 -273 -118
rect -207 -518 -177 -118
rect -111 -518 -81 -118
rect -15 -518 15 -118
rect 81 -518 111 -118
rect 177 -518 207 -118
rect 273 -518 303 -118
rect 369 -518 399 -118
rect 465 -518 495 -118
rect 561 -518 591 -118
rect 657 -518 687 -118
<< pdiff >>
rect -749 506 -687 518
rect -749 130 -737 506
rect -703 130 -687 506
rect -749 118 -687 130
rect -657 506 -591 518
rect -657 130 -641 506
rect -607 130 -591 506
rect -657 118 -591 130
rect -561 506 -495 518
rect -561 130 -545 506
rect -511 130 -495 506
rect -561 118 -495 130
rect -465 506 -399 518
rect -465 130 -449 506
rect -415 130 -399 506
rect -465 118 -399 130
rect -369 506 -303 518
rect -369 130 -353 506
rect -319 130 -303 506
rect -369 118 -303 130
rect -273 506 -207 518
rect -273 130 -257 506
rect -223 130 -207 506
rect -273 118 -207 130
rect -177 506 -111 518
rect -177 130 -161 506
rect -127 130 -111 506
rect -177 118 -111 130
rect -81 506 -15 518
rect -81 130 -65 506
rect -31 130 -15 506
rect -81 118 -15 130
rect 15 506 81 518
rect 15 130 31 506
rect 65 130 81 506
rect 15 118 81 130
rect 111 506 177 518
rect 111 130 127 506
rect 161 130 177 506
rect 111 118 177 130
rect 207 506 273 518
rect 207 130 223 506
rect 257 130 273 506
rect 207 118 273 130
rect 303 506 369 518
rect 303 130 319 506
rect 353 130 369 506
rect 303 118 369 130
rect 399 506 465 518
rect 399 130 415 506
rect 449 130 465 506
rect 399 118 465 130
rect 495 506 561 518
rect 495 130 511 506
rect 545 130 561 506
rect 495 118 561 130
rect 591 506 657 518
rect 591 130 607 506
rect 641 130 657 506
rect 591 118 657 130
rect 687 506 749 518
rect 687 130 703 506
rect 737 130 749 506
rect 687 118 749 130
rect -749 -130 -687 -118
rect -749 -506 -737 -130
rect -703 -506 -687 -130
rect -749 -518 -687 -506
rect -657 -130 -591 -118
rect -657 -506 -641 -130
rect -607 -506 -591 -130
rect -657 -518 -591 -506
rect -561 -130 -495 -118
rect -561 -506 -545 -130
rect -511 -506 -495 -130
rect -561 -518 -495 -506
rect -465 -130 -399 -118
rect -465 -506 -449 -130
rect -415 -506 -399 -130
rect -465 -518 -399 -506
rect -369 -130 -303 -118
rect -369 -506 -353 -130
rect -319 -506 -303 -130
rect -369 -518 -303 -506
rect -273 -130 -207 -118
rect -273 -506 -257 -130
rect -223 -506 -207 -130
rect -273 -518 -207 -506
rect -177 -130 -111 -118
rect -177 -506 -161 -130
rect -127 -506 -111 -130
rect -177 -518 -111 -506
rect -81 -130 -15 -118
rect -81 -506 -65 -130
rect -31 -506 -15 -130
rect -81 -518 -15 -506
rect 15 -130 81 -118
rect 15 -506 31 -130
rect 65 -506 81 -130
rect 15 -518 81 -506
rect 111 -130 177 -118
rect 111 -506 127 -130
rect 161 -506 177 -130
rect 111 -518 177 -506
rect 207 -130 273 -118
rect 207 -506 223 -130
rect 257 -506 273 -130
rect 207 -518 273 -506
rect 303 -130 369 -118
rect 303 -506 319 -130
rect 353 -506 369 -130
rect 303 -518 369 -506
rect 399 -130 465 -118
rect 399 -506 415 -130
rect 449 -506 465 -130
rect 399 -518 465 -506
rect 495 -130 561 -118
rect 495 -506 511 -130
rect 545 -506 561 -130
rect 495 -518 561 -506
rect 591 -130 657 -118
rect 591 -506 607 -130
rect 641 -506 657 -130
rect 591 -518 657 -506
rect 687 -130 749 -118
rect 687 -506 703 -130
rect 737 -506 749 -130
rect 687 -518 749 -506
<< pdiffc >>
rect -737 130 -703 506
rect -641 130 -607 506
rect -545 130 -511 506
rect -449 130 -415 506
rect -353 130 -319 506
rect -257 130 -223 506
rect -161 130 -127 506
rect -65 130 -31 506
rect 31 130 65 506
rect 127 130 161 506
rect 223 130 257 506
rect 319 130 353 506
rect 415 130 449 506
rect 511 130 545 506
rect 607 130 641 506
rect 703 130 737 506
rect -737 -506 -703 -130
rect -641 -506 -607 -130
rect -545 -506 -511 -130
rect -449 -506 -415 -130
rect -353 -506 -319 -130
rect -257 -506 -223 -130
rect -161 -506 -127 -130
rect -65 -506 -31 -130
rect 31 -506 65 -130
rect 127 -506 161 -130
rect 223 -506 257 -130
rect 319 -506 353 -130
rect 415 -506 449 -130
rect 511 -506 545 -130
rect 607 -506 641 -130
rect 703 -506 737 -130
<< nsubdiff >>
rect -851 667 -755 701
rect 755 667 851 701
rect -851 605 -817 667
rect 817 605 851 667
rect -851 -667 -817 -605
rect 817 -667 851 -605
rect -851 -701 -755 -667
rect 755 -701 851 -667
<< nsubdiffcont >>
rect -755 667 755 701
rect -851 -605 -817 605
rect 817 -605 851 605
rect -755 -701 755 -667
<< poly >>
rect -705 599 -639 615
rect -705 565 -689 599
rect -655 565 -639 599
rect -705 549 -639 565
rect -513 599 -447 615
rect -513 565 -497 599
rect -463 565 -447 599
rect -513 549 -447 565
rect -321 599 -255 615
rect -321 565 -305 599
rect -271 565 -255 599
rect -321 549 -255 565
rect -129 599 -63 615
rect -129 565 -113 599
rect -79 565 -63 599
rect -129 549 -63 565
rect 63 599 129 615
rect 63 565 79 599
rect 113 565 129 599
rect 63 549 129 565
rect 255 599 321 615
rect 255 565 271 599
rect 305 565 321 599
rect 255 549 321 565
rect 447 599 513 615
rect 447 565 463 599
rect 497 565 513 599
rect 447 549 513 565
rect 639 599 705 615
rect 639 565 655 599
rect 689 565 705 599
rect 639 549 705 565
rect -687 518 -657 549
rect -591 518 -561 544
rect -495 518 -465 549
rect -399 518 -369 544
rect -303 518 -273 549
rect -207 518 -177 544
rect -111 518 -81 549
rect -15 518 15 544
rect 81 518 111 549
rect 177 518 207 544
rect 273 518 303 549
rect 369 518 399 544
rect 465 518 495 549
rect 561 518 591 544
rect 657 518 687 549
rect -687 92 -657 118
rect -591 87 -561 118
rect -495 92 -465 118
rect -399 87 -369 118
rect -303 92 -273 118
rect -207 87 -177 118
rect -111 92 -81 118
rect -15 87 15 118
rect 81 92 111 118
rect 177 87 207 118
rect 273 92 303 118
rect 369 87 399 118
rect 465 92 495 118
rect 561 87 591 118
rect 657 92 687 118
rect -609 71 -543 87
rect -609 37 -593 71
rect -559 37 -543 71
rect -609 21 -543 37
rect -417 71 -351 87
rect -417 37 -401 71
rect -367 37 -351 71
rect -417 21 -351 37
rect -225 71 -159 87
rect -225 37 -209 71
rect -175 37 -159 71
rect -225 21 -159 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 159 71 225 87
rect 159 37 175 71
rect 209 37 225 71
rect 159 21 225 37
rect 351 71 417 87
rect 351 37 367 71
rect 401 37 417 71
rect 351 21 417 37
rect 543 71 609 87
rect 543 37 559 71
rect 593 37 609 71
rect 543 21 609 37
rect -609 -37 -543 -21
rect -609 -71 -593 -37
rect -559 -71 -543 -37
rect -609 -87 -543 -71
rect -417 -37 -351 -21
rect -417 -71 -401 -37
rect -367 -71 -351 -37
rect -417 -87 -351 -71
rect -225 -37 -159 -21
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -225 -87 -159 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 159 -37 225 -21
rect 159 -71 175 -37
rect 209 -71 225 -37
rect 159 -87 225 -71
rect 351 -37 417 -21
rect 351 -71 367 -37
rect 401 -71 417 -37
rect 351 -87 417 -71
rect 543 -37 609 -21
rect 543 -71 559 -37
rect 593 -71 609 -37
rect 543 -87 609 -71
rect -687 -118 -657 -92
rect -591 -118 -561 -87
rect -495 -118 -465 -92
rect -399 -118 -369 -87
rect -303 -118 -273 -92
rect -207 -118 -177 -87
rect -111 -118 -81 -92
rect -15 -118 15 -87
rect 81 -118 111 -92
rect 177 -118 207 -87
rect 273 -118 303 -92
rect 369 -118 399 -87
rect 465 -118 495 -92
rect 561 -118 591 -87
rect 657 -118 687 -92
rect -687 -549 -657 -518
rect -591 -544 -561 -518
rect -495 -549 -465 -518
rect -399 -544 -369 -518
rect -303 -549 -273 -518
rect -207 -544 -177 -518
rect -111 -549 -81 -518
rect -15 -544 15 -518
rect 81 -549 111 -518
rect 177 -544 207 -518
rect 273 -549 303 -518
rect 369 -544 399 -518
rect 465 -549 495 -518
rect 561 -544 591 -518
rect 657 -549 687 -518
rect -705 -565 -639 -549
rect -705 -599 -689 -565
rect -655 -599 -639 -565
rect -705 -615 -639 -599
rect -513 -565 -447 -549
rect -513 -599 -497 -565
rect -463 -599 -447 -565
rect -513 -615 -447 -599
rect -321 -565 -255 -549
rect -321 -599 -305 -565
rect -271 -599 -255 -565
rect -321 -615 -255 -599
rect -129 -565 -63 -549
rect -129 -599 -113 -565
rect -79 -599 -63 -565
rect -129 -615 -63 -599
rect 63 -565 129 -549
rect 63 -599 79 -565
rect 113 -599 129 -565
rect 63 -615 129 -599
rect 255 -565 321 -549
rect 255 -599 271 -565
rect 305 -599 321 -565
rect 255 -615 321 -599
rect 447 -565 513 -549
rect 447 -599 463 -565
rect 497 -599 513 -565
rect 447 -615 513 -599
rect 639 -565 705 -549
rect 639 -599 655 -565
rect 689 -599 705 -565
rect 639 -615 705 -599
<< polycont >>
rect -689 565 -655 599
rect -497 565 -463 599
rect -305 565 -271 599
rect -113 565 -79 599
rect 79 565 113 599
rect 271 565 305 599
rect 463 565 497 599
rect 655 565 689 599
rect -593 37 -559 71
rect -401 37 -367 71
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect 367 37 401 71
rect 559 37 593 71
rect -593 -71 -559 -37
rect -401 -71 -367 -37
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect 367 -71 401 -37
rect 559 -71 593 -37
rect -689 -599 -655 -565
rect -497 -599 -463 -565
rect -305 -599 -271 -565
rect -113 -599 -79 -565
rect 79 -599 113 -565
rect 271 -599 305 -565
rect 463 -599 497 -565
rect 655 -599 689 -565
<< locali >>
rect -851 667 -755 701
rect 755 667 851 701
rect -851 605 -817 667
rect 817 605 851 667
rect -705 565 -689 599
rect -655 565 -639 599
rect -513 565 -497 599
rect -463 565 -447 599
rect -321 565 -305 599
rect -271 565 -255 599
rect -129 565 -113 599
rect -79 565 -63 599
rect 63 565 79 599
rect 113 565 129 599
rect 255 565 271 599
rect 305 565 321 599
rect 447 565 463 599
rect 497 565 513 599
rect 639 565 655 599
rect 689 565 705 599
rect -737 506 -703 522
rect -737 114 -703 130
rect -641 506 -607 522
rect -641 114 -607 130
rect -545 506 -511 522
rect -545 114 -511 130
rect -449 506 -415 522
rect -449 114 -415 130
rect -353 506 -319 522
rect -353 114 -319 130
rect -257 506 -223 522
rect -257 114 -223 130
rect -161 506 -127 522
rect -161 114 -127 130
rect -65 506 -31 522
rect -65 114 -31 130
rect 31 506 65 522
rect 31 114 65 130
rect 127 506 161 522
rect 127 114 161 130
rect 223 506 257 522
rect 223 114 257 130
rect 319 506 353 522
rect 319 114 353 130
rect 415 506 449 522
rect 415 114 449 130
rect 511 506 545 522
rect 511 114 545 130
rect 607 506 641 522
rect 607 114 641 130
rect 703 506 737 522
rect 703 114 737 130
rect -609 37 -593 71
rect -559 37 -543 71
rect -417 37 -401 71
rect -367 37 -351 71
rect -225 37 -209 71
rect -175 37 -159 71
rect -33 37 -17 71
rect 17 37 33 71
rect 159 37 175 71
rect 209 37 225 71
rect 351 37 367 71
rect 401 37 417 71
rect 543 37 559 71
rect 593 37 609 71
rect -609 -71 -593 -37
rect -559 -71 -543 -37
rect -417 -71 -401 -37
rect -367 -71 -351 -37
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 159 -71 175 -37
rect 209 -71 225 -37
rect 351 -71 367 -37
rect 401 -71 417 -37
rect 543 -71 559 -37
rect 593 -71 609 -37
rect -737 -130 -703 -114
rect -737 -522 -703 -506
rect -641 -130 -607 -114
rect -641 -522 -607 -506
rect -545 -130 -511 -114
rect -545 -522 -511 -506
rect -449 -130 -415 -114
rect -449 -522 -415 -506
rect -353 -130 -319 -114
rect -353 -522 -319 -506
rect -257 -130 -223 -114
rect -257 -522 -223 -506
rect -161 -130 -127 -114
rect -161 -522 -127 -506
rect -65 -130 -31 -114
rect -65 -522 -31 -506
rect 31 -130 65 -114
rect 31 -522 65 -506
rect 127 -130 161 -114
rect 127 -522 161 -506
rect 223 -130 257 -114
rect 223 -522 257 -506
rect 319 -130 353 -114
rect 319 -522 353 -506
rect 415 -130 449 -114
rect 415 -522 449 -506
rect 511 -130 545 -114
rect 511 -522 545 -506
rect 607 -130 641 -114
rect 607 -522 641 -506
rect 703 -130 737 -114
rect 703 -522 737 -506
rect -705 -599 -689 -565
rect -655 -599 -639 -565
rect -513 -599 -497 -565
rect -463 -599 -447 -565
rect -321 -599 -305 -565
rect -271 -599 -255 -565
rect -129 -599 -113 -565
rect -79 -599 -63 -565
rect 63 -599 79 -565
rect 113 -599 129 -565
rect 255 -599 271 -565
rect 305 -599 321 -565
rect 447 -599 463 -565
rect 497 -599 513 -565
rect 639 -599 655 -565
rect 689 -599 705 -565
rect -851 -667 -817 -605
rect 817 -667 851 -605
rect -851 -701 -755 -667
rect 755 -701 851 -667
<< viali >>
rect -689 565 -655 599
rect -497 565 -463 599
rect -305 565 -271 599
rect -113 565 -79 599
rect 79 565 113 599
rect 271 565 305 599
rect 463 565 497 599
rect 655 565 689 599
rect -737 130 -703 506
rect -641 130 -607 506
rect -545 130 -511 506
rect -449 130 -415 506
rect -353 130 -319 506
rect -257 130 -223 506
rect -161 130 -127 506
rect -65 130 -31 506
rect 31 130 65 506
rect 127 130 161 506
rect 223 130 257 506
rect 319 130 353 506
rect 415 130 449 506
rect 511 130 545 506
rect 607 130 641 506
rect 703 130 737 506
rect -593 37 -559 71
rect -401 37 -367 71
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect 367 37 401 71
rect 559 37 593 71
rect -593 -71 -559 -37
rect -401 -71 -367 -37
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect 367 -71 401 -37
rect 559 -71 593 -37
rect -737 -506 -703 -130
rect -641 -506 -607 -130
rect -545 -506 -511 -130
rect -449 -506 -415 -130
rect -353 -506 -319 -130
rect -257 -506 -223 -130
rect -161 -506 -127 -130
rect -65 -506 -31 -130
rect 31 -506 65 -130
rect 127 -506 161 -130
rect 223 -506 257 -130
rect 319 -506 353 -130
rect 415 -506 449 -130
rect 511 -506 545 -130
rect 607 -506 641 -130
rect 703 -506 737 -130
rect -689 -599 -655 -565
rect -497 -599 -463 -565
rect -305 -599 -271 -565
rect -113 -599 -79 -565
rect 79 -599 113 -565
rect 271 -599 305 -565
rect 463 -599 497 -565
rect 655 -599 689 -565
<< metal1 >>
rect -701 599 -643 605
rect -701 565 -689 599
rect -655 565 -643 599
rect -701 559 -643 565
rect -509 599 -451 605
rect -509 565 -497 599
rect -463 565 -451 599
rect -509 559 -451 565
rect -317 599 -259 605
rect -317 565 -305 599
rect -271 565 -259 599
rect -317 559 -259 565
rect -125 599 -67 605
rect -125 565 -113 599
rect -79 565 -67 599
rect -125 559 -67 565
rect 67 599 125 605
rect 67 565 79 599
rect 113 565 125 599
rect 67 559 125 565
rect 259 599 317 605
rect 259 565 271 599
rect 305 565 317 599
rect 259 559 317 565
rect 451 599 509 605
rect 451 565 463 599
rect 497 565 509 599
rect 451 559 509 565
rect 643 599 701 605
rect 643 565 655 599
rect 689 565 701 599
rect 643 559 701 565
rect -743 506 -697 518
rect -743 130 -737 506
rect -703 130 -697 506
rect -743 118 -697 130
rect -647 506 -601 518
rect -647 130 -641 506
rect -607 130 -601 506
rect -647 118 -601 130
rect -551 506 -505 518
rect -551 130 -545 506
rect -511 130 -505 506
rect -551 118 -505 130
rect -455 506 -409 518
rect -455 130 -449 506
rect -415 130 -409 506
rect -455 118 -409 130
rect -359 506 -313 518
rect -359 130 -353 506
rect -319 130 -313 506
rect -359 118 -313 130
rect -263 506 -217 518
rect -263 130 -257 506
rect -223 130 -217 506
rect -263 118 -217 130
rect -167 506 -121 518
rect -167 130 -161 506
rect -127 130 -121 506
rect -167 118 -121 130
rect -71 506 -25 518
rect -71 130 -65 506
rect -31 130 -25 506
rect -71 118 -25 130
rect 25 506 71 518
rect 25 130 31 506
rect 65 130 71 506
rect 25 118 71 130
rect 121 506 167 518
rect 121 130 127 506
rect 161 130 167 506
rect 121 118 167 130
rect 217 506 263 518
rect 217 130 223 506
rect 257 130 263 506
rect 217 118 263 130
rect 313 506 359 518
rect 313 130 319 506
rect 353 130 359 506
rect 313 118 359 130
rect 409 506 455 518
rect 409 130 415 506
rect 449 130 455 506
rect 409 118 455 130
rect 505 506 551 518
rect 505 130 511 506
rect 545 130 551 506
rect 505 118 551 130
rect 601 506 647 518
rect 601 130 607 506
rect 641 130 647 506
rect 601 118 647 130
rect 697 506 743 518
rect 697 130 703 506
rect 737 130 743 506
rect 697 118 743 130
rect -605 71 -547 77
rect -605 37 -593 71
rect -559 37 -547 71
rect -605 31 -547 37
rect -413 71 -355 77
rect -413 37 -401 71
rect -367 37 -355 71
rect -413 31 -355 37
rect -221 71 -163 77
rect -221 37 -209 71
rect -175 37 -163 71
rect -221 31 -163 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 163 71 221 77
rect 163 37 175 71
rect 209 37 221 71
rect 163 31 221 37
rect 355 71 413 77
rect 355 37 367 71
rect 401 37 413 71
rect 355 31 413 37
rect 547 71 605 77
rect 547 37 559 71
rect 593 37 605 71
rect 547 31 605 37
rect -605 -37 -547 -31
rect -605 -71 -593 -37
rect -559 -71 -547 -37
rect -605 -77 -547 -71
rect -413 -37 -355 -31
rect -413 -71 -401 -37
rect -367 -71 -355 -37
rect -413 -77 -355 -71
rect -221 -37 -163 -31
rect -221 -71 -209 -37
rect -175 -71 -163 -37
rect -221 -77 -163 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 163 -37 221 -31
rect 163 -71 175 -37
rect 209 -71 221 -37
rect 163 -77 221 -71
rect 355 -37 413 -31
rect 355 -71 367 -37
rect 401 -71 413 -37
rect 355 -77 413 -71
rect 547 -37 605 -31
rect 547 -71 559 -37
rect 593 -71 605 -37
rect 547 -77 605 -71
rect -743 -130 -697 -118
rect -743 -506 -737 -130
rect -703 -506 -697 -130
rect -743 -518 -697 -506
rect -647 -130 -601 -118
rect -647 -506 -641 -130
rect -607 -506 -601 -130
rect -647 -518 -601 -506
rect -551 -130 -505 -118
rect -551 -506 -545 -130
rect -511 -506 -505 -130
rect -551 -518 -505 -506
rect -455 -130 -409 -118
rect -455 -506 -449 -130
rect -415 -506 -409 -130
rect -455 -518 -409 -506
rect -359 -130 -313 -118
rect -359 -506 -353 -130
rect -319 -506 -313 -130
rect -359 -518 -313 -506
rect -263 -130 -217 -118
rect -263 -506 -257 -130
rect -223 -506 -217 -130
rect -263 -518 -217 -506
rect -167 -130 -121 -118
rect -167 -506 -161 -130
rect -127 -506 -121 -130
rect -167 -518 -121 -506
rect -71 -130 -25 -118
rect -71 -506 -65 -130
rect -31 -506 -25 -130
rect -71 -518 -25 -506
rect 25 -130 71 -118
rect 25 -506 31 -130
rect 65 -506 71 -130
rect 25 -518 71 -506
rect 121 -130 167 -118
rect 121 -506 127 -130
rect 161 -506 167 -130
rect 121 -518 167 -506
rect 217 -130 263 -118
rect 217 -506 223 -130
rect 257 -506 263 -130
rect 217 -518 263 -506
rect 313 -130 359 -118
rect 313 -506 319 -130
rect 353 -506 359 -130
rect 313 -518 359 -506
rect 409 -130 455 -118
rect 409 -506 415 -130
rect 449 -506 455 -130
rect 409 -518 455 -506
rect 505 -130 551 -118
rect 505 -506 511 -130
rect 545 -506 551 -130
rect 505 -518 551 -506
rect 601 -130 647 -118
rect 601 -506 607 -130
rect 641 -506 647 -130
rect 601 -518 647 -506
rect 697 -130 743 -118
rect 697 -506 703 -130
rect 737 -506 743 -130
rect 697 -518 743 -506
rect -701 -565 -643 -559
rect -701 -599 -689 -565
rect -655 -599 -643 -565
rect -701 -605 -643 -599
rect -509 -565 -451 -559
rect -509 -599 -497 -565
rect -463 -599 -451 -565
rect -509 -605 -451 -599
rect -317 -565 -259 -559
rect -317 -599 -305 -565
rect -271 -599 -259 -565
rect -317 -605 -259 -599
rect -125 -565 -67 -559
rect -125 -599 -113 -565
rect -79 -599 -67 -565
rect -125 -605 -67 -599
rect 67 -565 125 -559
rect 67 -599 79 -565
rect 113 -599 125 -565
rect 67 -605 125 -599
rect 259 -565 317 -559
rect 259 -599 271 -565
rect 305 -599 317 -565
rect 259 -605 317 -599
rect 451 -565 509 -559
rect 451 -599 463 -565
rect 497 -599 509 -565
rect 451 -605 509 -599
rect 643 -565 701 -559
rect 643 -599 655 -565
rect 689 -599 701 -565
rect 643 -605 701 -599
<< properties >>
string FIXED_BBOX -834 -684 834 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 2 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
