magic
tech sky130A
magscale 1 2
timestamp 1683737876
<< error_p >>
rect -5741 581 -5683 587
rect -5549 581 -5491 587
rect -5357 581 -5299 587
rect -5165 581 -5107 587
rect -4973 581 -4915 587
rect -4781 581 -4723 587
rect -4589 581 -4531 587
rect -4397 581 -4339 587
rect -4205 581 -4147 587
rect -4013 581 -3955 587
rect -3821 581 -3763 587
rect -3629 581 -3571 587
rect -3437 581 -3379 587
rect -3245 581 -3187 587
rect -3053 581 -2995 587
rect -2861 581 -2803 587
rect -2669 581 -2611 587
rect -2477 581 -2419 587
rect -2285 581 -2227 587
rect -2093 581 -2035 587
rect -1901 581 -1843 587
rect -1709 581 -1651 587
rect -1517 581 -1459 587
rect -1325 581 -1267 587
rect -1133 581 -1075 587
rect -941 581 -883 587
rect -749 581 -691 587
rect -557 581 -499 587
rect -365 581 -307 587
rect -173 581 -115 587
rect 19 581 77 587
rect 211 581 269 587
rect 403 581 461 587
rect 595 581 653 587
rect 787 581 845 587
rect 979 581 1037 587
rect 1171 581 1229 587
rect 1363 581 1421 587
rect 1555 581 1613 587
rect 1747 581 1805 587
rect 1939 581 1997 587
rect 2131 581 2189 587
rect 2323 581 2381 587
rect 2515 581 2573 587
rect 2707 581 2765 587
rect 2899 581 2957 587
rect 3091 581 3149 587
rect 3283 581 3341 587
rect 3475 581 3533 587
rect 3667 581 3725 587
rect 3859 581 3917 587
rect 4051 581 4109 587
rect 4243 581 4301 587
rect 4435 581 4493 587
rect 4627 581 4685 587
rect 4819 581 4877 587
rect 5011 581 5069 587
rect 5203 581 5261 587
rect 5395 581 5453 587
rect 5587 581 5645 587
rect -5741 547 -5729 581
rect -5549 547 -5537 581
rect -5357 547 -5345 581
rect -5165 547 -5153 581
rect -4973 547 -4961 581
rect -4781 547 -4769 581
rect -4589 547 -4577 581
rect -4397 547 -4385 581
rect -4205 547 -4193 581
rect -4013 547 -4001 581
rect -3821 547 -3809 581
rect -3629 547 -3617 581
rect -3437 547 -3425 581
rect -3245 547 -3233 581
rect -3053 547 -3041 581
rect -2861 547 -2849 581
rect -2669 547 -2657 581
rect -2477 547 -2465 581
rect -2285 547 -2273 581
rect -2093 547 -2081 581
rect -1901 547 -1889 581
rect -1709 547 -1697 581
rect -1517 547 -1505 581
rect -1325 547 -1313 581
rect -1133 547 -1121 581
rect -941 547 -929 581
rect -749 547 -737 581
rect -557 547 -545 581
rect -365 547 -353 581
rect -173 547 -161 581
rect 19 547 31 581
rect 211 547 223 581
rect 403 547 415 581
rect 595 547 607 581
rect 787 547 799 581
rect 979 547 991 581
rect 1171 547 1183 581
rect 1363 547 1375 581
rect 1555 547 1567 581
rect 1747 547 1759 581
rect 1939 547 1951 581
rect 2131 547 2143 581
rect 2323 547 2335 581
rect 2515 547 2527 581
rect 2707 547 2719 581
rect 2899 547 2911 581
rect 3091 547 3103 581
rect 3283 547 3295 581
rect 3475 547 3487 581
rect 3667 547 3679 581
rect 3859 547 3871 581
rect 4051 547 4063 581
rect 4243 547 4255 581
rect 4435 547 4447 581
rect 4627 547 4639 581
rect 4819 547 4831 581
rect 5011 547 5023 581
rect 5203 547 5215 581
rect 5395 547 5407 581
rect 5587 547 5599 581
rect -5741 541 -5683 547
rect -5549 541 -5491 547
rect -5357 541 -5299 547
rect -5165 541 -5107 547
rect -4973 541 -4915 547
rect -4781 541 -4723 547
rect -4589 541 -4531 547
rect -4397 541 -4339 547
rect -4205 541 -4147 547
rect -4013 541 -3955 547
rect -3821 541 -3763 547
rect -3629 541 -3571 547
rect -3437 541 -3379 547
rect -3245 541 -3187 547
rect -3053 541 -2995 547
rect -2861 541 -2803 547
rect -2669 541 -2611 547
rect -2477 541 -2419 547
rect -2285 541 -2227 547
rect -2093 541 -2035 547
rect -1901 541 -1843 547
rect -1709 541 -1651 547
rect -1517 541 -1459 547
rect -1325 541 -1267 547
rect -1133 541 -1075 547
rect -941 541 -883 547
rect -749 541 -691 547
rect -557 541 -499 547
rect -365 541 -307 547
rect -173 541 -115 547
rect 19 541 77 547
rect 211 541 269 547
rect 403 541 461 547
rect 595 541 653 547
rect 787 541 845 547
rect 979 541 1037 547
rect 1171 541 1229 547
rect 1363 541 1421 547
rect 1555 541 1613 547
rect 1747 541 1805 547
rect 1939 541 1997 547
rect 2131 541 2189 547
rect 2323 541 2381 547
rect 2515 541 2573 547
rect 2707 541 2765 547
rect 2899 541 2957 547
rect 3091 541 3149 547
rect 3283 541 3341 547
rect 3475 541 3533 547
rect 3667 541 3725 547
rect 3859 541 3917 547
rect 4051 541 4109 547
rect 4243 541 4301 547
rect 4435 541 4493 547
rect 4627 541 4685 547
rect 4819 541 4877 547
rect 5011 541 5069 547
rect 5203 541 5261 547
rect 5395 541 5453 547
rect 5587 541 5645 547
rect -5645 71 -5587 77
rect -5453 71 -5395 77
rect -5261 71 -5203 77
rect -5069 71 -5011 77
rect -4877 71 -4819 77
rect -4685 71 -4627 77
rect -4493 71 -4435 77
rect -4301 71 -4243 77
rect -4109 71 -4051 77
rect -3917 71 -3859 77
rect -3725 71 -3667 77
rect -3533 71 -3475 77
rect -3341 71 -3283 77
rect -3149 71 -3091 77
rect -2957 71 -2899 77
rect -2765 71 -2707 77
rect -2573 71 -2515 77
rect -2381 71 -2323 77
rect -2189 71 -2131 77
rect -1997 71 -1939 77
rect -1805 71 -1747 77
rect -1613 71 -1555 77
rect -1421 71 -1363 77
rect -1229 71 -1171 77
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect 1267 71 1325 77
rect 1459 71 1517 77
rect 1651 71 1709 77
rect 1843 71 1901 77
rect 2035 71 2093 77
rect 2227 71 2285 77
rect 2419 71 2477 77
rect 2611 71 2669 77
rect 2803 71 2861 77
rect 2995 71 3053 77
rect 3187 71 3245 77
rect 3379 71 3437 77
rect 3571 71 3629 77
rect 3763 71 3821 77
rect 3955 71 4013 77
rect 4147 71 4205 77
rect 4339 71 4397 77
rect 4531 71 4589 77
rect 4723 71 4781 77
rect 4915 71 4973 77
rect 5107 71 5165 77
rect 5299 71 5357 77
rect 5491 71 5549 77
rect 5683 71 5741 77
rect -5645 37 -5633 71
rect -5453 37 -5441 71
rect -5261 37 -5249 71
rect -5069 37 -5057 71
rect -4877 37 -4865 71
rect -4685 37 -4673 71
rect -4493 37 -4481 71
rect -4301 37 -4289 71
rect -4109 37 -4097 71
rect -3917 37 -3905 71
rect -3725 37 -3713 71
rect -3533 37 -3521 71
rect -3341 37 -3329 71
rect -3149 37 -3137 71
rect -2957 37 -2945 71
rect -2765 37 -2753 71
rect -2573 37 -2561 71
rect -2381 37 -2369 71
rect -2189 37 -2177 71
rect -1997 37 -1985 71
rect -1805 37 -1793 71
rect -1613 37 -1601 71
rect -1421 37 -1409 71
rect -1229 37 -1217 71
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect 1267 37 1279 71
rect 1459 37 1471 71
rect 1651 37 1663 71
rect 1843 37 1855 71
rect 2035 37 2047 71
rect 2227 37 2239 71
rect 2419 37 2431 71
rect 2611 37 2623 71
rect 2803 37 2815 71
rect 2995 37 3007 71
rect 3187 37 3199 71
rect 3379 37 3391 71
rect 3571 37 3583 71
rect 3763 37 3775 71
rect 3955 37 3967 71
rect 4147 37 4159 71
rect 4339 37 4351 71
rect 4531 37 4543 71
rect 4723 37 4735 71
rect 4915 37 4927 71
rect 5107 37 5119 71
rect 5299 37 5311 71
rect 5491 37 5503 71
rect 5683 37 5695 71
rect -5645 31 -5587 37
rect -5453 31 -5395 37
rect -5261 31 -5203 37
rect -5069 31 -5011 37
rect -4877 31 -4819 37
rect -4685 31 -4627 37
rect -4493 31 -4435 37
rect -4301 31 -4243 37
rect -4109 31 -4051 37
rect -3917 31 -3859 37
rect -3725 31 -3667 37
rect -3533 31 -3475 37
rect -3341 31 -3283 37
rect -3149 31 -3091 37
rect -2957 31 -2899 37
rect -2765 31 -2707 37
rect -2573 31 -2515 37
rect -2381 31 -2323 37
rect -2189 31 -2131 37
rect -1997 31 -1939 37
rect -1805 31 -1747 37
rect -1613 31 -1555 37
rect -1421 31 -1363 37
rect -1229 31 -1171 37
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect 1267 31 1325 37
rect 1459 31 1517 37
rect 1651 31 1709 37
rect 1843 31 1901 37
rect 2035 31 2093 37
rect 2227 31 2285 37
rect 2419 31 2477 37
rect 2611 31 2669 37
rect 2803 31 2861 37
rect 2995 31 3053 37
rect 3187 31 3245 37
rect 3379 31 3437 37
rect 3571 31 3629 37
rect 3763 31 3821 37
rect 3955 31 4013 37
rect 4147 31 4205 37
rect 4339 31 4397 37
rect 4531 31 4589 37
rect 4723 31 4781 37
rect 4915 31 4973 37
rect 5107 31 5165 37
rect 5299 31 5357 37
rect 5491 31 5549 37
rect 5683 31 5741 37
rect -5645 -37 -5587 -31
rect -5453 -37 -5395 -31
rect -5261 -37 -5203 -31
rect -5069 -37 -5011 -31
rect -4877 -37 -4819 -31
rect -4685 -37 -4627 -31
rect -4493 -37 -4435 -31
rect -4301 -37 -4243 -31
rect -4109 -37 -4051 -31
rect -3917 -37 -3859 -31
rect -3725 -37 -3667 -31
rect -3533 -37 -3475 -31
rect -3341 -37 -3283 -31
rect -3149 -37 -3091 -31
rect -2957 -37 -2899 -31
rect -2765 -37 -2707 -31
rect -2573 -37 -2515 -31
rect -2381 -37 -2323 -31
rect -2189 -37 -2131 -31
rect -1997 -37 -1939 -31
rect -1805 -37 -1747 -31
rect -1613 -37 -1555 -31
rect -1421 -37 -1363 -31
rect -1229 -37 -1171 -31
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect 1267 -37 1325 -31
rect 1459 -37 1517 -31
rect 1651 -37 1709 -31
rect 1843 -37 1901 -31
rect 2035 -37 2093 -31
rect 2227 -37 2285 -31
rect 2419 -37 2477 -31
rect 2611 -37 2669 -31
rect 2803 -37 2861 -31
rect 2995 -37 3053 -31
rect 3187 -37 3245 -31
rect 3379 -37 3437 -31
rect 3571 -37 3629 -31
rect 3763 -37 3821 -31
rect 3955 -37 4013 -31
rect 4147 -37 4205 -31
rect 4339 -37 4397 -31
rect 4531 -37 4589 -31
rect 4723 -37 4781 -31
rect 4915 -37 4973 -31
rect 5107 -37 5165 -31
rect 5299 -37 5357 -31
rect 5491 -37 5549 -31
rect 5683 -37 5741 -31
rect -5645 -71 -5633 -37
rect -5453 -71 -5441 -37
rect -5261 -71 -5249 -37
rect -5069 -71 -5057 -37
rect -4877 -71 -4865 -37
rect -4685 -71 -4673 -37
rect -4493 -71 -4481 -37
rect -4301 -71 -4289 -37
rect -4109 -71 -4097 -37
rect -3917 -71 -3905 -37
rect -3725 -71 -3713 -37
rect -3533 -71 -3521 -37
rect -3341 -71 -3329 -37
rect -3149 -71 -3137 -37
rect -2957 -71 -2945 -37
rect -2765 -71 -2753 -37
rect -2573 -71 -2561 -37
rect -2381 -71 -2369 -37
rect -2189 -71 -2177 -37
rect -1997 -71 -1985 -37
rect -1805 -71 -1793 -37
rect -1613 -71 -1601 -37
rect -1421 -71 -1409 -37
rect -1229 -71 -1217 -37
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect 1267 -71 1279 -37
rect 1459 -71 1471 -37
rect 1651 -71 1663 -37
rect 1843 -71 1855 -37
rect 2035 -71 2047 -37
rect 2227 -71 2239 -37
rect 2419 -71 2431 -37
rect 2611 -71 2623 -37
rect 2803 -71 2815 -37
rect 2995 -71 3007 -37
rect 3187 -71 3199 -37
rect 3379 -71 3391 -37
rect 3571 -71 3583 -37
rect 3763 -71 3775 -37
rect 3955 -71 3967 -37
rect 4147 -71 4159 -37
rect 4339 -71 4351 -37
rect 4531 -71 4543 -37
rect 4723 -71 4735 -37
rect 4915 -71 4927 -37
rect 5107 -71 5119 -37
rect 5299 -71 5311 -37
rect 5491 -71 5503 -37
rect 5683 -71 5695 -37
rect -5645 -77 -5587 -71
rect -5453 -77 -5395 -71
rect -5261 -77 -5203 -71
rect -5069 -77 -5011 -71
rect -4877 -77 -4819 -71
rect -4685 -77 -4627 -71
rect -4493 -77 -4435 -71
rect -4301 -77 -4243 -71
rect -4109 -77 -4051 -71
rect -3917 -77 -3859 -71
rect -3725 -77 -3667 -71
rect -3533 -77 -3475 -71
rect -3341 -77 -3283 -71
rect -3149 -77 -3091 -71
rect -2957 -77 -2899 -71
rect -2765 -77 -2707 -71
rect -2573 -77 -2515 -71
rect -2381 -77 -2323 -71
rect -2189 -77 -2131 -71
rect -1997 -77 -1939 -71
rect -1805 -77 -1747 -71
rect -1613 -77 -1555 -71
rect -1421 -77 -1363 -71
rect -1229 -77 -1171 -71
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect 1267 -77 1325 -71
rect 1459 -77 1517 -71
rect 1651 -77 1709 -71
rect 1843 -77 1901 -71
rect 2035 -77 2093 -71
rect 2227 -77 2285 -71
rect 2419 -77 2477 -71
rect 2611 -77 2669 -71
rect 2803 -77 2861 -71
rect 2995 -77 3053 -71
rect 3187 -77 3245 -71
rect 3379 -77 3437 -71
rect 3571 -77 3629 -71
rect 3763 -77 3821 -71
rect 3955 -77 4013 -71
rect 4147 -77 4205 -71
rect 4339 -77 4397 -71
rect 4531 -77 4589 -71
rect 4723 -77 4781 -71
rect 4915 -77 4973 -71
rect 5107 -77 5165 -71
rect 5299 -77 5357 -71
rect 5491 -77 5549 -71
rect 5683 -77 5741 -71
rect -5741 -547 -5683 -541
rect -5549 -547 -5491 -541
rect -5357 -547 -5299 -541
rect -5165 -547 -5107 -541
rect -4973 -547 -4915 -541
rect -4781 -547 -4723 -541
rect -4589 -547 -4531 -541
rect -4397 -547 -4339 -541
rect -4205 -547 -4147 -541
rect -4013 -547 -3955 -541
rect -3821 -547 -3763 -541
rect -3629 -547 -3571 -541
rect -3437 -547 -3379 -541
rect -3245 -547 -3187 -541
rect -3053 -547 -2995 -541
rect -2861 -547 -2803 -541
rect -2669 -547 -2611 -541
rect -2477 -547 -2419 -541
rect -2285 -547 -2227 -541
rect -2093 -547 -2035 -541
rect -1901 -547 -1843 -541
rect -1709 -547 -1651 -541
rect -1517 -547 -1459 -541
rect -1325 -547 -1267 -541
rect -1133 -547 -1075 -541
rect -941 -547 -883 -541
rect -749 -547 -691 -541
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect 595 -547 653 -541
rect 787 -547 845 -541
rect 979 -547 1037 -541
rect 1171 -547 1229 -541
rect 1363 -547 1421 -541
rect 1555 -547 1613 -541
rect 1747 -547 1805 -541
rect 1939 -547 1997 -541
rect 2131 -547 2189 -541
rect 2323 -547 2381 -541
rect 2515 -547 2573 -541
rect 2707 -547 2765 -541
rect 2899 -547 2957 -541
rect 3091 -547 3149 -541
rect 3283 -547 3341 -541
rect 3475 -547 3533 -541
rect 3667 -547 3725 -541
rect 3859 -547 3917 -541
rect 4051 -547 4109 -541
rect 4243 -547 4301 -541
rect 4435 -547 4493 -541
rect 4627 -547 4685 -541
rect 4819 -547 4877 -541
rect 5011 -547 5069 -541
rect 5203 -547 5261 -541
rect 5395 -547 5453 -541
rect 5587 -547 5645 -541
rect -5741 -581 -5729 -547
rect -5549 -581 -5537 -547
rect -5357 -581 -5345 -547
rect -5165 -581 -5153 -547
rect -4973 -581 -4961 -547
rect -4781 -581 -4769 -547
rect -4589 -581 -4577 -547
rect -4397 -581 -4385 -547
rect -4205 -581 -4193 -547
rect -4013 -581 -4001 -547
rect -3821 -581 -3809 -547
rect -3629 -581 -3617 -547
rect -3437 -581 -3425 -547
rect -3245 -581 -3233 -547
rect -3053 -581 -3041 -547
rect -2861 -581 -2849 -547
rect -2669 -581 -2657 -547
rect -2477 -581 -2465 -547
rect -2285 -581 -2273 -547
rect -2093 -581 -2081 -547
rect -1901 -581 -1889 -547
rect -1709 -581 -1697 -547
rect -1517 -581 -1505 -547
rect -1325 -581 -1313 -547
rect -1133 -581 -1121 -547
rect -941 -581 -929 -547
rect -749 -581 -737 -547
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect 595 -581 607 -547
rect 787 -581 799 -547
rect 979 -581 991 -547
rect 1171 -581 1183 -547
rect 1363 -581 1375 -547
rect 1555 -581 1567 -547
rect 1747 -581 1759 -547
rect 1939 -581 1951 -547
rect 2131 -581 2143 -547
rect 2323 -581 2335 -547
rect 2515 -581 2527 -547
rect 2707 -581 2719 -547
rect 2899 -581 2911 -547
rect 3091 -581 3103 -547
rect 3283 -581 3295 -547
rect 3475 -581 3487 -547
rect 3667 -581 3679 -547
rect 3859 -581 3871 -547
rect 4051 -581 4063 -547
rect 4243 -581 4255 -547
rect 4435 -581 4447 -547
rect 4627 -581 4639 -547
rect 4819 -581 4831 -547
rect 5011 -581 5023 -547
rect 5203 -581 5215 -547
rect 5395 -581 5407 -547
rect 5587 -581 5599 -547
rect -5741 -587 -5683 -581
rect -5549 -587 -5491 -581
rect -5357 -587 -5299 -581
rect -5165 -587 -5107 -581
rect -4973 -587 -4915 -581
rect -4781 -587 -4723 -581
rect -4589 -587 -4531 -581
rect -4397 -587 -4339 -581
rect -4205 -587 -4147 -581
rect -4013 -587 -3955 -581
rect -3821 -587 -3763 -581
rect -3629 -587 -3571 -581
rect -3437 -587 -3379 -581
rect -3245 -587 -3187 -581
rect -3053 -587 -2995 -581
rect -2861 -587 -2803 -581
rect -2669 -587 -2611 -581
rect -2477 -587 -2419 -581
rect -2285 -587 -2227 -581
rect -2093 -587 -2035 -581
rect -1901 -587 -1843 -581
rect -1709 -587 -1651 -581
rect -1517 -587 -1459 -581
rect -1325 -587 -1267 -581
rect -1133 -587 -1075 -581
rect -941 -587 -883 -581
rect -749 -587 -691 -581
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
rect 595 -587 653 -581
rect 787 -587 845 -581
rect 979 -587 1037 -581
rect 1171 -587 1229 -581
rect 1363 -587 1421 -581
rect 1555 -587 1613 -581
rect 1747 -587 1805 -581
rect 1939 -587 1997 -581
rect 2131 -587 2189 -581
rect 2323 -587 2381 -581
rect 2515 -587 2573 -581
rect 2707 -587 2765 -581
rect 2899 -587 2957 -581
rect 3091 -587 3149 -581
rect 3283 -587 3341 -581
rect 3475 -587 3533 -581
rect 3667 -587 3725 -581
rect 3859 -587 3917 -581
rect 4051 -587 4109 -581
rect 4243 -587 4301 -581
rect 4435 -587 4493 -581
rect 4627 -587 4685 -581
rect 4819 -587 4877 -581
rect 5011 -587 5069 -581
rect 5203 -587 5261 -581
rect 5395 -587 5453 -581
rect 5587 -587 5645 -581
<< pwell >>
rect -5927 -719 5927 719
<< nmoslvt >>
rect -5727 109 -5697 509
rect -5631 109 -5601 509
rect -5535 109 -5505 509
rect -5439 109 -5409 509
rect -5343 109 -5313 509
rect -5247 109 -5217 509
rect -5151 109 -5121 509
rect -5055 109 -5025 509
rect -4959 109 -4929 509
rect -4863 109 -4833 509
rect -4767 109 -4737 509
rect -4671 109 -4641 509
rect -4575 109 -4545 509
rect -4479 109 -4449 509
rect -4383 109 -4353 509
rect -4287 109 -4257 509
rect -4191 109 -4161 509
rect -4095 109 -4065 509
rect -3999 109 -3969 509
rect -3903 109 -3873 509
rect -3807 109 -3777 509
rect -3711 109 -3681 509
rect -3615 109 -3585 509
rect -3519 109 -3489 509
rect -3423 109 -3393 509
rect -3327 109 -3297 509
rect -3231 109 -3201 509
rect -3135 109 -3105 509
rect -3039 109 -3009 509
rect -2943 109 -2913 509
rect -2847 109 -2817 509
rect -2751 109 -2721 509
rect -2655 109 -2625 509
rect -2559 109 -2529 509
rect -2463 109 -2433 509
rect -2367 109 -2337 509
rect -2271 109 -2241 509
rect -2175 109 -2145 509
rect -2079 109 -2049 509
rect -1983 109 -1953 509
rect -1887 109 -1857 509
rect -1791 109 -1761 509
rect -1695 109 -1665 509
rect -1599 109 -1569 509
rect -1503 109 -1473 509
rect -1407 109 -1377 509
rect -1311 109 -1281 509
rect -1215 109 -1185 509
rect -1119 109 -1089 509
rect -1023 109 -993 509
rect -927 109 -897 509
rect -831 109 -801 509
rect -735 109 -705 509
rect -639 109 -609 509
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect 609 109 639 509
rect 705 109 735 509
rect 801 109 831 509
rect 897 109 927 509
rect 993 109 1023 509
rect 1089 109 1119 509
rect 1185 109 1215 509
rect 1281 109 1311 509
rect 1377 109 1407 509
rect 1473 109 1503 509
rect 1569 109 1599 509
rect 1665 109 1695 509
rect 1761 109 1791 509
rect 1857 109 1887 509
rect 1953 109 1983 509
rect 2049 109 2079 509
rect 2145 109 2175 509
rect 2241 109 2271 509
rect 2337 109 2367 509
rect 2433 109 2463 509
rect 2529 109 2559 509
rect 2625 109 2655 509
rect 2721 109 2751 509
rect 2817 109 2847 509
rect 2913 109 2943 509
rect 3009 109 3039 509
rect 3105 109 3135 509
rect 3201 109 3231 509
rect 3297 109 3327 509
rect 3393 109 3423 509
rect 3489 109 3519 509
rect 3585 109 3615 509
rect 3681 109 3711 509
rect 3777 109 3807 509
rect 3873 109 3903 509
rect 3969 109 3999 509
rect 4065 109 4095 509
rect 4161 109 4191 509
rect 4257 109 4287 509
rect 4353 109 4383 509
rect 4449 109 4479 509
rect 4545 109 4575 509
rect 4641 109 4671 509
rect 4737 109 4767 509
rect 4833 109 4863 509
rect 4929 109 4959 509
rect 5025 109 5055 509
rect 5121 109 5151 509
rect 5217 109 5247 509
rect 5313 109 5343 509
rect 5409 109 5439 509
rect 5505 109 5535 509
rect 5601 109 5631 509
rect 5697 109 5727 509
rect -5727 -509 -5697 -109
rect -5631 -509 -5601 -109
rect -5535 -509 -5505 -109
rect -5439 -509 -5409 -109
rect -5343 -509 -5313 -109
rect -5247 -509 -5217 -109
rect -5151 -509 -5121 -109
rect -5055 -509 -5025 -109
rect -4959 -509 -4929 -109
rect -4863 -509 -4833 -109
rect -4767 -509 -4737 -109
rect -4671 -509 -4641 -109
rect -4575 -509 -4545 -109
rect -4479 -509 -4449 -109
rect -4383 -509 -4353 -109
rect -4287 -509 -4257 -109
rect -4191 -509 -4161 -109
rect -4095 -509 -4065 -109
rect -3999 -509 -3969 -109
rect -3903 -509 -3873 -109
rect -3807 -509 -3777 -109
rect -3711 -509 -3681 -109
rect -3615 -509 -3585 -109
rect -3519 -509 -3489 -109
rect -3423 -509 -3393 -109
rect -3327 -509 -3297 -109
rect -3231 -509 -3201 -109
rect -3135 -509 -3105 -109
rect -3039 -509 -3009 -109
rect -2943 -509 -2913 -109
rect -2847 -509 -2817 -109
rect -2751 -509 -2721 -109
rect -2655 -509 -2625 -109
rect -2559 -509 -2529 -109
rect -2463 -509 -2433 -109
rect -2367 -509 -2337 -109
rect -2271 -509 -2241 -109
rect -2175 -509 -2145 -109
rect -2079 -509 -2049 -109
rect -1983 -509 -1953 -109
rect -1887 -509 -1857 -109
rect -1791 -509 -1761 -109
rect -1695 -509 -1665 -109
rect -1599 -509 -1569 -109
rect -1503 -509 -1473 -109
rect -1407 -509 -1377 -109
rect -1311 -509 -1281 -109
rect -1215 -509 -1185 -109
rect -1119 -509 -1089 -109
rect -1023 -509 -993 -109
rect -927 -509 -897 -109
rect -831 -509 -801 -109
rect -735 -509 -705 -109
rect -639 -509 -609 -109
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect 609 -509 639 -109
rect 705 -509 735 -109
rect 801 -509 831 -109
rect 897 -509 927 -109
rect 993 -509 1023 -109
rect 1089 -509 1119 -109
rect 1185 -509 1215 -109
rect 1281 -509 1311 -109
rect 1377 -509 1407 -109
rect 1473 -509 1503 -109
rect 1569 -509 1599 -109
rect 1665 -509 1695 -109
rect 1761 -509 1791 -109
rect 1857 -509 1887 -109
rect 1953 -509 1983 -109
rect 2049 -509 2079 -109
rect 2145 -509 2175 -109
rect 2241 -509 2271 -109
rect 2337 -509 2367 -109
rect 2433 -509 2463 -109
rect 2529 -509 2559 -109
rect 2625 -509 2655 -109
rect 2721 -509 2751 -109
rect 2817 -509 2847 -109
rect 2913 -509 2943 -109
rect 3009 -509 3039 -109
rect 3105 -509 3135 -109
rect 3201 -509 3231 -109
rect 3297 -509 3327 -109
rect 3393 -509 3423 -109
rect 3489 -509 3519 -109
rect 3585 -509 3615 -109
rect 3681 -509 3711 -109
rect 3777 -509 3807 -109
rect 3873 -509 3903 -109
rect 3969 -509 3999 -109
rect 4065 -509 4095 -109
rect 4161 -509 4191 -109
rect 4257 -509 4287 -109
rect 4353 -509 4383 -109
rect 4449 -509 4479 -109
rect 4545 -509 4575 -109
rect 4641 -509 4671 -109
rect 4737 -509 4767 -109
rect 4833 -509 4863 -109
rect 4929 -509 4959 -109
rect 5025 -509 5055 -109
rect 5121 -509 5151 -109
rect 5217 -509 5247 -109
rect 5313 -509 5343 -109
rect 5409 -509 5439 -109
rect 5505 -509 5535 -109
rect 5601 -509 5631 -109
rect 5697 -509 5727 -109
<< ndiff >>
rect -5789 497 -5727 509
rect -5789 121 -5777 497
rect -5743 121 -5727 497
rect -5789 109 -5727 121
rect -5697 497 -5631 509
rect -5697 121 -5681 497
rect -5647 121 -5631 497
rect -5697 109 -5631 121
rect -5601 497 -5535 509
rect -5601 121 -5585 497
rect -5551 121 -5535 497
rect -5601 109 -5535 121
rect -5505 497 -5439 509
rect -5505 121 -5489 497
rect -5455 121 -5439 497
rect -5505 109 -5439 121
rect -5409 497 -5343 509
rect -5409 121 -5393 497
rect -5359 121 -5343 497
rect -5409 109 -5343 121
rect -5313 497 -5247 509
rect -5313 121 -5297 497
rect -5263 121 -5247 497
rect -5313 109 -5247 121
rect -5217 497 -5151 509
rect -5217 121 -5201 497
rect -5167 121 -5151 497
rect -5217 109 -5151 121
rect -5121 497 -5055 509
rect -5121 121 -5105 497
rect -5071 121 -5055 497
rect -5121 109 -5055 121
rect -5025 497 -4959 509
rect -5025 121 -5009 497
rect -4975 121 -4959 497
rect -5025 109 -4959 121
rect -4929 497 -4863 509
rect -4929 121 -4913 497
rect -4879 121 -4863 497
rect -4929 109 -4863 121
rect -4833 497 -4767 509
rect -4833 121 -4817 497
rect -4783 121 -4767 497
rect -4833 109 -4767 121
rect -4737 497 -4671 509
rect -4737 121 -4721 497
rect -4687 121 -4671 497
rect -4737 109 -4671 121
rect -4641 497 -4575 509
rect -4641 121 -4625 497
rect -4591 121 -4575 497
rect -4641 109 -4575 121
rect -4545 497 -4479 509
rect -4545 121 -4529 497
rect -4495 121 -4479 497
rect -4545 109 -4479 121
rect -4449 497 -4383 509
rect -4449 121 -4433 497
rect -4399 121 -4383 497
rect -4449 109 -4383 121
rect -4353 497 -4287 509
rect -4353 121 -4337 497
rect -4303 121 -4287 497
rect -4353 109 -4287 121
rect -4257 497 -4191 509
rect -4257 121 -4241 497
rect -4207 121 -4191 497
rect -4257 109 -4191 121
rect -4161 497 -4095 509
rect -4161 121 -4145 497
rect -4111 121 -4095 497
rect -4161 109 -4095 121
rect -4065 497 -3999 509
rect -4065 121 -4049 497
rect -4015 121 -3999 497
rect -4065 109 -3999 121
rect -3969 497 -3903 509
rect -3969 121 -3953 497
rect -3919 121 -3903 497
rect -3969 109 -3903 121
rect -3873 497 -3807 509
rect -3873 121 -3857 497
rect -3823 121 -3807 497
rect -3873 109 -3807 121
rect -3777 497 -3711 509
rect -3777 121 -3761 497
rect -3727 121 -3711 497
rect -3777 109 -3711 121
rect -3681 497 -3615 509
rect -3681 121 -3665 497
rect -3631 121 -3615 497
rect -3681 109 -3615 121
rect -3585 497 -3519 509
rect -3585 121 -3569 497
rect -3535 121 -3519 497
rect -3585 109 -3519 121
rect -3489 497 -3423 509
rect -3489 121 -3473 497
rect -3439 121 -3423 497
rect -3489 109 -3423 121
rect -3393 497 -3327 509
rect -3393 121 -3377 497
rect -3343 121 -3327 497
rect -3393 109 -3327 121
rect -3297 497 -3231 509
rect -3297 121 -3281 497
rect -3247 121 -3231 497
rect -3297 109 -3231 121
rect -3201 497 -3135 509
rect -3201 121 -3185 497
rect -3151 121 -3135 497
rect -3201 109 -3135 121
rect -3105 497 -3039 509
rect -3105 121 -3089 497
rect -3055 121 -3039 497
rect -3105 109 -3039 121
rect -3009 497 -2943 509
rect -3009 121 -2993 497
rect -2959 121 -2943 497
rect -3009 109 -2943 121
rect -2913 497 -2847 509
rect -2913 121 -2897 497
rect -2863 121 -2847 497
rect -2913 109 -2847 121
rect -2817 497 -2751 509
rect -2817 121 -2801 497
rect -2767 121 -2751 497
rect -2817 109 -2751 121
rect -2721 497 -2655 509
rect -2721 121 -2705 497
rect -2671 121 -2655 497
rect -2721 109 -2655 121
rect -2625 497 -2559 509
rect -2625 121 -2609 497
rect -2575 121 -2559 497
rect -2625 109 -2559 121
rect -2529 497 -2463 509
rect -2529 121 -2513 497
rect -2479 121 -2463 497
rect -2529 109 -2463 121
rect -2433 497 -2367 509
rect -2433 121 -2417 497
rect -2383 121 -2367 497
rect -2433 109 -2367 121
rect -2337 497 -2271 509
rect -2337 121 -2321 497
rect -2287 121 -2271 497
rect -2337 109 -2271 121
rect -2241 497 -2175 509
rect -2241 121 -2225 497
rect -2191 121 -2175 497
rect -2241 109 -2175 121
rect -2145 497 -2079 509
rect -2145 121 -2129 497
rect -2095 121 -2079 497
rect -2145 109 -2079 121
rect -2049 497 -1983 509
rect -2049 121 -2033 497
rect -1999 121 -1983 497
rect -2049 109 -1983 121
rect -1953 497 -1887 509
rect -1953 121 -1937 497
rect -1903 121 -1887 497
rect -1953 109 -1887 121
rect -1857 497 -1791 509
rect -1857 121 -1841 497
rect -1807 121 -1791 497
rect -1857 109 -1791 121
rect -1761 497 -1695 509
rect -1761 121 -1745 497
rect -1711 121 -1695 497
rect -1761 109 -1695 121
rect -1665 497 -1599 509
rect -1665 121 -1649 497
rect -1615 121 -1599 497
rect -1665 109 -1599 121
rect -1569 497 -1503 509
rect -1569 121 -1553 497
rect -1519 121 -1503 497
rect -1569 109 -1503 121
rect -1473 497 -1407 509
rect -1473 121 -1457 497
rect -1423 121 -1407 497
rect -1473 109 -1407 121
rect -1377 497 -1311 509
rect -1377 121 -1361 497
rect -1327 121 -1311 497
rect -1377 109 -1311 121
rect -1281 497 -1215 509
rect -1281 121 -1265 497
rect -1231 121 -1215 497
rect -1281 109 -1215 121
rect -1185 497 -1119 509
rect -1185 121 -1169 497
rect -1135 121 -1119 497
rect -1185 109 -1119 121
rect -1089 497 -1023 509
rect -1089 121 -1073 497
rect -1039 121 -1023 497
rect -1089 109 -1023 121
rect -993 497 -927 509
rect -993 121 -977 497
rect -943 121 -927 497
rect -993 109 -927 121
rect -897 497 -831 509
rect -897 121 -881 497
rect -847 121 -831 497
rect -897 109 -831 121
rect -801 497 -735 509
rect -801 121 -785 497
rect -751 121 -735 497
rect -801 109 -735 121
rect -705 497 -639 509
rect -705 121 -689 497
rect -655 121 -639 497
rect -705 109 -639 121
rect -609 497 -543 509
rect -609 121 -593 497
rect -559 121 -543 497
rect -609 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 609 509
rect 543 121 559 497
rect 593 121 609 497
rect 543 109 609 121
rect 639 497 705 509
rect 639 121 655 497
rect 689 121 705 497
rect 639 109 705 121
rect 735 497 801 509
rect 735 121 751 497
rect 785 121 801 497
rect 735 109 801 121
rect 831 497 897 509
rect 831 121 847 497
rect 881 121 897 497
rect 831 109 897 121
rect 927 497 993 509
rect 927 121 943 497
rect 977 121 993 497
rect 927 109 993 121
rect 1023 497 1089 509
rect 1023 121 1039 497
rect 1073 121 1089 497
rect 1023 109 1089 121
rect 1119 497 1185 509
rect 1119 121 1135 497
rect 1169 121 1185 497
rect 1119 109 1185 121
rect 1215 497 1281 509
rect 1215 121 1231 497
rect 1265 121 1281 497
rect 1215 109 1281 121
rect 1311 497 1377 509
rect 1311 121 1327 497
rect 1361 121 1377 497
rect 1311 109 1377 121
rect 1407 497 1473 509
rect 1407 121 1423 497
rect 1457 121 1473 497
rect 1407 109 1473 121
rect 1503 497 1569 509
rect 1503 121 1519 497
rect 1553 121 1569 497
rect 1503 109 1569 121
rect 1599 497 1665 509
rect 1599 121 1615 497
rect 1649 121 1665 497
rect 1599 109 1665 121
rect 1695 497 1761 509
rect 1695 121 1711 497
rect 1745 121 1761 497
rect 1695 109 1761 121
rect 1791 497 1857 509
rect 1791 121 1807 497
rect 1841 121 1857 497
rect 1791 109 1857 121
rect 1887 497 1953 509
rect 1887 121 1903 497
rect 1937 121 1953 497
rect 1887 109 1953 121
rect 1983 497 2049 509
rect 1983 121 1999 497
rect 2033 121 2049 497
rect 1983 109 2049 121
rect 2079 497 2145 509
rect 2079 121 2095 497
rect 2129 121 2145 497
rect 2079 109 2145 121
rect 2175 497 2241 509
rect 2175 121 2191 497
rect 2225 121 2241 497
rect 2175 109 2241 121
rect 2271 497 2337 509
rect 2271 121 2287 497
rect 2321 121 2337 497
rect 2271 109 2337 121
rect 2367 497 2433 509
rect 2367 121 2383 497
rect 2417 121 2433 497
rect 2367 109 2433 121
rect 2463 497 2529 509
rect 2463 121 2479 497
rect 2513 121 2529 497
rect 2463 109 2529 121
rect 2559 497 2625 509
rect 2559 121 2575 497
rect 2609 121 2625 497
rect 2559 109 2625 121
rect 2655 497 2721 509
rect 2655 121 2671 497
rect 2705 121 2721 497
rect 2655 109 2721 121
rect 2751 497 2817 509
rect 2751 121 2767 497
rect 2801 121 2817 497
rect 2751 109 2817 121
rect 2847 497 2913 509
rect 2847 121 2863 497
rect 2897 121 2913 497
rect 2847 109 2913 121
rect 2943 497 3009 509
rect 2943 121 2959 497
rect 2993 121 3009 497
rect 2943 109 3009 121
rect 3039 497 3105 509
rect 3039 121 3055 497
rect 3089 121 3105 497
rect 3039 109 3105 121
rect 3135 497 3201 509
rect 3135 121 3151 497
rect 3185 121 3201 497
rect 3135 109 3201 121
rect 3231 497 3297 509
rect 3231 121 3247 497
rect 3281 121 3297 497
rect 3231 109 3297 121
rect 3327 497 3393 509
rect 3327 121 3343 497
rect 3377 121 3393 497
rect 3327 109 3393 121
rect 3423 497 3489 509
rect 3423 121 3439 497
rect 3473 121 3489 497
rect 3423 109 3489 121
rect 3519 497 3585 509
rect 3519 121 3535 497
rect 3569 121 3585 497
rect 3519 109 3585 121
rect 3615 497 3681 509
rect 3615 121 3631 497
rect 3665 121 3681 497
rect 3615 109 3681 121
rect 3711 497 3777 509
rect 3711 121 3727 497
rect 3761 121 3777 497
rect 3711 109 3777 121
rect 3807 497 3873 509
rect 3807 121 3823 497
rect 3857 121 3873 497
rect 3807 109 3873 121
rect 3903 497 3969 509
rect 3903 121 3919 497
rect 3953 121 3969 497
rect 3903 109 3969 121
rect 3999 497 4065 509
rect 3999 121 4015 497
rect 4049 121 4065 497
rect 3999 109 4065 121
rect 4095 497 4161 509
rect 4095 121 4111 497
rect 4145 121 4161 497
rect 4095 109 4161 121
rect 4191 497 4257 509
rect 4191 121 4207 497
rect 4241 121 4257 497
rect 4191 109 4257 121
rect 4287 497 4353 509
rect 4287 121 4303 497
rect 4337 121 4353 497
rect 4287 109 4353 121
rect 4383 497 4449 509
rect 4383 121 4399 497
rect 4433 121 4449 497
rect 4383 109 4449 121
rect 4479 497 4545 509
rect 4479 121 4495 497
rect 4529 121 4545 497
rect 4479 109 4545 121
rect 4575 497 4641 509
rect 4575 121 4591 497
rect 4625 121 4641 497
rect 4575 109 4641 121
rect 4671 497 4737 509
rect 4671 121 4687 497
rect 4721 121 4737 497
rect 4671 109 4737 121
rect 4767 497 4833 509
rect 4767 121 4783 497
rect 4817 121 4833 497
rect 4767 109 4833 121
rect 4863 497 4929 509
rect 4863 121 4879 497
rect 4913 121 4929 497
rect 4863 109 4929 121
rect 4959 497 5025 509
rect 4959 121 4975 497
rect 5009 121 5025 497
rect 4959 109 5025 121
rect 5055 497 5121 509
rect 5055 121 5071 497
rect 5105 121 5121 497
rect 5055 109 5121 121
rect 5151 497 5217 509
rect 5151 121 5167 497
rect 5201 121 5217 497
rect 5151 109 5217 121
rect 5247 497 5313 509
rect 5247 121 5263 497
rect 5297 121 5313 497
rect 5247 109 5313 121
rect 5343 497 5409 509
rect 5343 121 5359 497
rect 5393 121 5409 497
rect 5343 109 5409 121
rect 5439 497 5505 509
rect 5439 121 5455 497
rect 5489 121 5505 497
rect 5439 109 5505 121
rect 5535 497 5601 509
rect 5535 121 5551 497
rect 5585 121 5601 497
rect 5535 109 5601 121
rect 5631 497 5697 509
rect 5631 121 5647 497
rect 5681 121 5697 497
rect 5631 109 5697 121
rect 5727 497 5789 509
rect 5727 121 5743 497
rect 5777 121 5789 497
rect 5727 109 5789 121
rect -5789 -121 -5727 -109
rect -5789 -497 -5777 -121
rect -5743 -497 -5727 -121
rect -5789 -509 -5727 -497
rect -5697 -121 -5631 -109
rect -5697 -497 -5681 -121
rect -5647 -497 -5631 -121
rect -5697 -509 -5631 -497
rect -5601 -121 -5535 -109
rect -5601 -497 -5585 -121
rect -5551 -497 -5535 -121
rect -5601 -509 -5535 -497
rect -5505 -121 -5439 -109
rect -5505 -497 -5489 -121
rect -5455 -497 -5439 -121
rect -5505 -509 -5439 -497
rect -5409 -121 -5343 -109
rect -5409 -497 -5393 -121
rect -5359 -497 -5343 -121
rect -5409 -509 -5343 -497
rect -5313 -121 -5247 -109
rect -5313 -497 -5297 -121
rect -5263 -497 -5247 -121
rect -5313 -509 -5247 -497
rect -5217 -121 -5151 -109
rect -5217 -497 -5201 -121
rect -5167 -497 -5151 -121
rect -5217 -509 -5151 -497
rect -5121 -121 -5055 -109
rect -5121 -497 -5105 -121
rect -5071 -497 -5055 -121
rect -5121 -509 -5055 -497
rect -5025 -121 -4959 -109
rect -5025 -497 -5009 -121
rect -4975 -497 -4959 -121
rect -5025 -509 -4959 -497
rect -4929 -121 -4863 -109
rect -4929 -497 -4913 -121
rect -4879 -497 -4863 -121
rect -4929 -509 -4863 -497
rect -4833 -121 -4767 -109
rect -4833 -497 -4817 -121
rect -4783 -497 -4767 -121
rect -4833 -509 -4767 -497
rect -4737 -121 -4671 -109
rect -4737 -497 -4721 -121
rect -4687 -497 -4671 -121
rect -4737 -509 -4671 -497
rect -4641 -121 -4575 -109
rect -4641 -497 -4625 -121
rect -4591 -497 -4575 -121
rect -4641 -509 -4575 -497
rect -4545 -121 -4479 -109
rect -4545 -497 -4529 -121
rect -4495 -497 -4479 -121
rect -4545 -509 -4479 -497
rect -4449 -121 -4383 -109
rect -4449 -497 -4433 -121
rect -4399 -497 -4383 -121
rect -4449 -509 -4383 -497
rect -4353 -121 -4287 -109
rect -4353 -497 -4337 -121
rect -4303 -497 -4287 -121
rect -4353 -509 -4287 -497
rect -4257 -121 -4191 -109
rect -4257 -497 -4241 -121
rect -4207 -497 -4191 -121
rect -4257 -509 -4191 -497
rect -4161 -121 -4095 -109
rect -4161 -497 -4145 -121
rect -4111 -497 -4095 -121
rect -4161 -509 -4095 -497
rect -4065 -121 -3999 -109
rect -4065 -497 -4049 -121
rect -4015 -497 -3999 -121
rect -4065 -509 -3999 -497
rect -3969 -121 -3903 -109
rect -3969 -497 -3953 -121
rect -3919 -497 -3903 -121
rect -3969 -509 -3903 -497
rect -3873 -121 -3807 -109
rect -3873 -497 -3857 -121
rect -3823 -497 -3807 -121
rect -3873 -509 -3807 -497
rect -3777 -121 -3711 -109
rect -3777 -497 -3761 -121
rect -3727 -497 -3711 -121
rect -3777 -509 -3711 -497
rect -3681 -121 -3615 -109
rect -3681 -497 -3665 -121
rect -3631 -497 -3615 -121
rect -3681 -509 -3615 -497
rect -3585 -121 -3519 -109
rect -3585 -497 -3569 -121
rect -3535 -497 -3519 -121
rect -3585 -509 -3519 -497
rect -3489 -121 -3423 -109
rect -3489 -497 -3473 -121
rect -3439 -497 -3423 -121
rect -3489 -509 -3423 -497
rect -3393 -121 -3327 -109
rect -3393 -497 -3377 -121
rect -3343 -497 -3327 -121
rect -3393 -509 -3327 -497
rect -3297 -121 -3231 -109
rect -3297 -497 -3281 -121
rect -3247 -497 -3231 -121
rect -3297 -509 -3231 -497
rect -3201 -121 -3135 -109
rect -3201 -497 -3185 -121
rect -3151 -497 -3135 -121
rect -3201 -509 -3135 -497
rect -3105 -121 -3039 -109
rect -3105 -497 -3089 -121
rect -3055 -497 -3039 -121
rect -3105 -509 -3039 -497
rect -3009 -121 -2943 -109
rect -3009 -497 -2993 -121
rect -2959 -497 -2943 -121
rect -3009 -509 -2943 -497
rect -2913 -121 -2847 -109
rect -2913 -497 -2897 -121
rect -2863 -497 -2847 -121
rect -2913 -509 -2847 -497
rect -2817 -121 -2751 -109
rect -2817 -497 -2801 -121
rect -2767 -497 -2751 -121
rect -2817 -509 -2751 -497
rect -2721 -121 -2655 -109
rect -2721 -497 -2705 -121
rect -2671 -497 -2655 -121
rect -2721 -509 -2655 -497
rect -2625 -121 -2559 -109
rect -2625 -497 -2609 -121
rect -2575 -497 -2559 -121
rect -2625 -509 -2559 -497
rect -2529 -121 -2463 -109
rect -2529 -497 -2513 -121
rect -2479 -497 -2463 -121
rect -2529 -509 -2463 -497
rect -2433 -121 -2367 -109
rect -2433 -497 -2417 -121
rect -2383 -497 -2367 -121
rect -2433 -509 -2367 -497
rect -2337 -121 -2271 -109
rect -2337 -497 -2321 -121
rect -2287 -497 -2271 -121
rect -2337 -509 -2271 -497
rect -2241 -121 -2175 -109
rect -2241 -497 -2225 -121
rect -2191 -497 -2175 -121
rect -2241 -509 -2175 -497
rect -2145 -121 -2079 -109
rect -2145 -497 -2129 -121
rect -2095 -497 -2079 -121
rect -2145 -509 -2079 -497
rect -2049 -121 -1983 -109
rect -2049 -497 -2033 -121
rect -1999 -497 -1983 -121
rect -2049 -509 -1983 -497
rect -1953 -121 -1887 -109
rect -1953 -497 -1937 -121
rect -1903 -497 -1887 -121
rect -1953 -509 -1887 -497
rect -1857 -121 -1791 -109
rect -1857 -497 -1841 -121
rect -1807 -497 -1791 -121
rect -1857 -509 -1791 -497
rect -1761 -121 -1695 -109
rect -1761 -497 -1745 -121
rect -1711 -497 -1695 -121
rect -1761 -509 -1695 -497
rect -1665 -121 -1599 -109
rect -1665 -497 -1649 -121
rect -1615 -497 -1599 -121
rect -1665 -509 -1599 -497
rect -1569 -121 -1503 -109
rect -1569 -497 -1553 -121
rect -1519 -497 -1503 -121
rect -1569 -509 -1503 -497
rect -1473 -121 -1407 -109
rect -1473 -497 -1457 -121
rect -1423 -497 -1407 -121
rect -1473 -509 -1407 -497
rect -1377 -121 -1311 -109
rect -1377 -497 -1361 -121
rect -1327 -497 -1311 -121
rect -1377 -509 -1311 -497
rect -1281 -121 -1215 -109
rect -1281 -497 -1265 -121
rect -1231 -497 -1215 -121
rect -1281 -509 -1215 -497
rect -1185 -121 -1119 -109
rect -1185 -497 -1169 -121
rect -1135 -497 -1119 -121
rect -1185 -509 -1119 -497
rect -1089 -121 -1023 -109
rect -1089 -497 -1073 -121
rect -1039 -497 -1023 -121
rect -1089 -509 -1023 -497
rect -993 -121 -927 -109
rect -993 -497 -977 -121
rect -943 -497 -927 -121
rect -993 -509 -927 -497
rect -897 -121 -831 -109
rect -897 -497 -881 -121
rect -847 -497 -831 -121
rect -897 -509 -831 -497
rect -801 -121 -735 -109
rect -801 -497 -785 -121
rect -751 -497 -735 -121
rect -801 -509 -735 -497
rect -705 -121 -639 -109
rect -705 -497 -689 -121
rect -655 -497 -639 -121
rect -705 -509 -639 -497
rect -609 -121 -543 -109
rect -609 -497 -593 -121
rect -559 -497 -543 -121
rect -609 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 609 -109
rect 543 -497 559 -121
rect 593 -497 609 -121
rect 543 -509 609 -497
rect 639 -121 705 -109
rect 639 -497 655 -121
rect 689 -497 705 -121
rect 639 -509 705 -497
rect 735 -121 801 -109
rect 735 -497 751 -121
rect 785 -497 801 -121
rect 735 -509 801 -497
rect 831 -121 897 -109
rect 831 -497 847 -121
rect 881 -497 897 -121
rect 831 -509 897 -497
rect 927 -121 993 -109
rect 927 -497 943 -121
rect 977 -497 993 -121
rect 927 -509 993 -497
rect 1023 -121 1089 -109
rect 1023 -497 1039 -121
rect 1073 -497 1089 -121
rect 1023 -509 1089 -497
rect 1119 -121 1185 -109
rect 1119 -497 1135 -121
rect 1169 -497 1185 -121
rect 1119 -509 1185 -497
rect 1215 -121 1281 -109
rect 1215 -497 1231 -121
rect 1265 -497 1281 -121
rect 1215 -509 1281 -497
rect 1311 -121 1377 -109
rect 1311 -497 1327 -121
rect 1361 -497 1377 -121
rect 1311 -509 1377 -497
rect 1407 -121 1473 -109
rect 1407 -497 1423 -121
rect 1457 -497 1473 -121
rect 1407 -509 1473 -497
rect 1503 -121 1569 -109
rect 1503 -497 1519 -121
rect 1553 -497 1569 -121
rect 1503 -509 1569 -497
rect 1599 -121 1665 -109
rect 1599 -497 1615 -121
rect 1649 -497 1665 -121
rect 1599 -509 1665 -497
rect 1695 -121 1761 -109
rect 1695 -497 1711 -121
rect 1745 -497 1761 -121
rect 1695 -509 1761 -497
rect 1791 -121 1857 -109
rect 1791 -497 1807 -121
rect 1841 -497 1857 -121
rect 1791 -509 1857 -497
rect 1887 -121 1953 -109
rect 1887 -497 1903 -121
rect 1937 -497 1953 -121
rect 1887 -509 1953 -497
rect 1983 -121 2049 -109
rect 1983 -497 1999 -121
rect 2033 -497 2049 -121
rect 1983 -509 2049 -497
rect 2079 -121 2145 -109
rect 2079 -497 2095 -121
rect 2129 -497 2145 -121
rect 2079 -509 2145 -497
rect 2175 -121 2241 -109
rect 2175 -497 2191 -121
rect 2225 -497 2241 -121
rect 2175 -509 2241 -497
rect 2271 -121 2337 -109
rect 2271 -497 2287 -121
rect 2321 -497 2337 -121
rect 2271 -509 2337 -497
rect 2367 -121 2433 -109
rect 2367 -497 2383 -121
rect 2417 -497 2433 -121
rect 2367 -509 2433 -497
rect 2463 -121 2529 -109
rect 2463 -497 2479 -121
rect 2513 -497 2529 -121
rect 2463 -509 2529 -497
rect 2559 -121 2625 -109
rect 2559 -497 2575 -121
rect 2609 -497 2625 -121
rect 2559 -509 2625 -497
rect 2655 -121 2721 -109
rect 2655 -497 2671 -121
rect 2705 -497 2721 -121
rect 2655 -509 2721 -497
rect 2751 -121 2817 -109
rect 2751 -497 2767 -121
rect 2801 -497 2817 -121
rect 2751 -509 2817 -497
rect 2847 -121 2913 -109
rect 2847 -497 2863 -121
rect 2897 -497 2913 -121
rect 2847 -509 2913 -497
rect 2943 -121 3009 -109
rect 2943 -497 2959 -121
rect 2993 -497 3009 -121
rect 2943 -509 3009 -497
rect 3039 -121 3105 -109
rect 3039 -497 3055 -121
rect 3089 -497 3105 -121
rect 3039 -509 3105 -497
rect 3135 -121 3201 -109
rect 3135 -497 3151 -121
rect 3185 -497 3201 -121
rect 3135 -509 3201 -497
rect 3231 -121 3297 -109
rect 3231 -497 3247 -121
rect 3281 -497 3297 -121
rect 3231 -509 3297 -497
rect 3327 -121 3393 -109
rect 3327 -497 3343 -121
rect 3377 -497 3393 -121
rect 3327 -509 3393 -497
rect 3423 -121 3489 -109
rect 3423 -497 3439 -121
rect 3473 -497 3489 -121
rect 3423 -509 3489 -497
rect 3519 -121 3585 -109
rect 3519 -497 3535 -121
rect 3569 -497 3585 -121
rect 3519 -509 3585 -497
rect 3615 -121 3681 -109
rect 3615 -497 3631 -121
rect 3665 -497 3681 -121
rect 3615 -509 3681 -497
rect 3711 -121 3777 -109
rect 3711 -497 3727 -121
rect 3761 -497 3777 -121
rect 3711 -509 3777 -497
rect 3807 -121 3873 -109
rect 3807 -497 3823 -121
rect 3857 -497 3873 -121
rect 3807 -509 3873 -497
rect 3903 -121 3969 -109
rect 3903 -497 3919 -121
rect 3953 -497 3969 -121
rect 3903 -509 3969 -497
rect 3999 -121 4065 -109
rect 3999 -497 4015 -121
rect 4049 -497 4065 -121
rect 3999 -509 4065 -497
rect 4095 -121 4161 -109
rect 4095 -497 4111 -121
rect 4145 -497 4161 -121
rect 4095 -509 4161 -497
rect 4191 -121 4257 -109
rect 4191 -497 4207 -121
rect 4241 -497 4257 -121
rect 4191 -509 4257 -497
rect 4287 -121 4353 -109
rect 4287 -497 4303 -121
rect 4337 -497 4353 -121
rect 4287 -509 4353 -497
rect 4383 -121 4449 -109
rect 4383 -497 4399 -121
rect 4433 -497 4449 -121
rect 4383 -509 4449 -497
rect 4479 -121 4545 -109
rect 4479 -497 4495 -121
rect 4529 -497 4545 -121
rect 4479 -509 4545 -497
rect 4575 -121 4641 -109
rect 4575 -497 4591 -121
rect 4625 -497 4641 -121
rect 4575 -509 4641 -497
rect 4671 -121 4737 -109
rect 4671 -497 4687 -121
rect 4721 -497 4737 -121
rect 4671 -509 4737 -497
rect 4767 -121 4833 -109
rect 4767 -497 4783 -121
rect 4817 -497 4833 -121
rect 4767 -509 4833 -497
rect 4863 -121 4929 -109
rect 4863 -497 4879 -121
rect 4913 -497 4929 -121
rect 4863 -509 4929 -497
rect 4959 -121 5025 -109
rect 4959 -497 4975 -121
rect 5009 -497 5025 -121
rect 4959 -509 5025 -497
rect 5055 -121 5121 -109
rect 5055 -497 5071 -121
rect 5105 -497 5121 -121
rect 5055 -509 5121 -497
rect 5151 -121 5217 -109
rect 5151 -497 5167 -121
rect 5201 -497 5217 -121
rect 5151 -509 5217 -497
rect 5247 -121 5313 -109
rect 5247 -497 5263 -121
rect 5297 -497 5313 -121
rect 5247 -509 5313 -497
rect 5343 -121 5409 -109
rect 5343 -497 5359 -121
rect 5393 -497 5409 -121
rect 5343 -509 5409 -497
rect 5439 -121 5505 -109
rect 5439 -497 5455 -121
rect 5489 -497 5505 -121
rect 5439 -509 5505 -497
rect 5535 -121 5601 -109
rect 5535 -497 5551 -121
rect 5585 -497 5601 -121
rect 5535 -509 5601 -497
rect 5631 -121 5697 -109
rect 5631 -497 5647 -121
rect 5681 -497 5697 -121
rect 5631 -509 5697 -497
rect 5727 -121 5789 -109
rect 5727 -497 5743 -121
rect 5777 -497 5789 -121
rect 5727 -509 5789 -497
<< ndiffc >>
rect -5777 121 -5743 497
rect -5681 121 -5647 497
rect -5585 121 -5551 497
rect -5489 121 -5455 497
rect -5393 121 -5359 497
rect -5297 121 -5263 497
rect -5201 121 -5167 497
rect -5105 121 -5071 497
rect -5009 121 -4975 497
rect -4913 121 -4879 497
rect -4817 121 -4783 497
rect -4721 121 -4687 497
rect -4625 121 -4591 497
rect -4529 121 -4495 497
rect -4433 121 -4399 497
rect -4337 121 -4303 497
rect -4241 121 -4207 497
rect -4145 121 -4111 497
rect -4049 121 -4015 497
rect -3953 121 -3919 497
rect -3857 121 -3823 497
rect -3761 121 -3727 497
rect -3665 121 -3631 497
rect -3569 121 -3535 497
rect -3473 121 -3439 497
rect -3377 121 -3343 497
rect -3281 121 -3247 497
rect -3185 121 -3151 497
rect -3089 121 -3055 497
rect -2993 121 -2959 497
rect -2897 121 -2863 497
rect -2801 121 -2767 497
rect -2705 121 -2671 497
rect -2609 121 -2575 497
rect -2513 121 -2479 497
rect -2417 121 -2383 497
rect -2321 121 -2287 497
rect -2225 121 -2191 497
rect -2129 121 -2095 497
rect -2033 121 -1999 497
rect -1937 121 -1903 497
rect -1841 121 -1807 497
rect -1745 121 -1711 497
rect -1649 121 -1615 497
rect -1553 121 -1519 497
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect 1519 121 1553 497
rect 1615 121 1649 497
rect 1711 121 1745 497
rect 1807 121 1841 497
rect 1903 121 1937 497
rect 1999 121 2033 497
rect 2095 121 2129 497
rect 2191 121 2225 497
rect 2287 121 2321 497
rect 2383 121 2417 497
rect 2479 121 2513 497
rect 2575 121 2609 497
rect 2671 121 2705 497
rect 2767 121 2801 497
rect 2863 121 2897 497
rect 2959 121 2993 497
rect 3055 121 3089 497
rect 3151 121 3185 497
rect 3247 121 3281 497
rect 3343 121 3377 497
rect 3439 121 3473 497
rect 3535 121 3569 497
rect 3631 121 3665 497
rect 3727 121 3761 497
rect 3823 121 3857 497
rect 3919 121 3953 497
rect 4015 121 4049 497
rect 4111 121 4145 497
rect 4207 121 4241 497
rect 4303 121 4337 497
rect 4399 121 4433 497
rect 4495 121 4529 497
rect 4591 121 4625 497
rect 4687 121 4721 497
rect 4783 121 4817 497
rect 4879 121 4913 497
rect 4975 121 5009 497
rect 5071 121 5105 497
rect 5167 121 5201 497
rect 5263 121 5297 497
rect 5359 121 5393 497
rect 5455 121 5489 497
rect 5551 121 5585 497
rect 5647 121 5681 497
rect 5743 121 5777 497
rect -5777 -497 -5743 -121
rect -5681 -497 -5647 -121
rect -5585 -497 -5551 -121
rect -5489 -497 -5455 -121
rect -5393 -497 -5359 -121
rect -5297 -497 -5263 -121
rect -5201 -497 -5167 -121
rect -5105 -497 -5071 -121
rect -5009 -497 -4975 -121
rect -4913 -497 -4879 -121
rect -4817 -497 -4783 -121
rect -4721 -497 -4687 -121
rect -4625 -497 -4591 -121
rect -4529 -497 -4495 -121
rect -4433 -497 -4399 -121
rect -4337 -497 -4303 -121
rect -4241 -497 -4207 -121
rect -4145 -497 -4111 -121
rect -4049 -497 -4015 -121
rect -3953 -497 -3919 -121
rect -3857 -497 -3823 -121
rect -3761 -497 -3727 -121
rect -3665 -497 -3631 -121
rect -3569 -497 -3535 -121
rect -3473 -497 -3439 -121
rect -3377 -497 -3343 -121
rect -3281 -497 -3247 -121
rect -3185 -497 -3151 -121
rect -3089 -497 -3055 -121
rect -2993 -497 -2959 -121
rect -2897 -497 -2863 -121
rect -2801 -497 -2767 -121
rect -2705 -497 -2671 -121
rect -2609 -497 -2575 -121
rect -2513 -497 -2479 -121
rect -2417 -497 -2383 -121
rect -2321 -497 -2287 -121
rect -2225 -497 -2191 -121
rect -2129 -497 -2095 -121
rect -2033 -497 -1999 -121
rect -1937 -497 -1903 -121
rect -1841 -497 -1807 -121
rect -1745 -497 -1711 -121
rect -1649 -497 -1615 -121
rect -1553 -497 -1519 -121
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect 1519 -497 1553 -121
rect 1615 -497 1649 -121
rect 1711 -497 1745 -121
rect 1807 -497 1841 -121
rect 1903 -497 1937 -121
rect 1999 -497 2033 -121
rect 2095 -497 2129 -121
rect 2191 -497 2225 -121
rect 2287 -497 2321 -121
rect 2383 -497 2417 -121
rect 2479 -497 2513 -121
rect 2575 -497 2609 -121
rect 2671 -497 2705 -121
rect 2767 -497 2801 -121
rect 2863 -497 2897 -121
rect 2959 -497 2993 -121
rect 3055 -497 3089 -121
rect 3151 -497 3185 -121
rect 3247 -497 3281 -121
rect 3343 -497 3377 -121
rect 3439 -497 3473 -121
rect 3535 -497 3569 -121
rect 3631 -497 3665 -121
rect 3727 -497 3761 -121
rect 3823 -497 3857 -121
rect 3919 -497 3953 -121
rect 4015 -497 4049 -121
rect 4111 -497 4145 -121
rect 4207 -497 4241 -121
rect 4303 -497 4337 -121
rect 4399 -497 4433 -121
rect 4495 -497 4529 -121
rect 4591 -497 4625 -121
rect 4687 -497 4721 -121
rect 4783 -497 4817 -121
rect 4879 -497 4913 -121
rect 4975 -497 5009 -121
rect 5071 -497 5105 -121
rect 5167 -497 5201 -121
rect 5263 -497 5297 -121
rect 5359 -497 5393 -121
rect 5455 -497 5489 -121
rect 5551 -497 5585 -121
rect 5647 -497 5681 -121
rect 5743 -497 5777 -121
<< psubdiff >>
rect -5891 649 -5795 683
rect 5795 649 5891 683
rect -5891 587 -5857 649
rect 5857 587 5891 649
rect -5891 -649 -5857 -587
rect 5857 -649 5891 -587
rect -5891 -683 -5795 -649
rect 5795 -683 5891 -649
<< psubdiffcont >>
rect -5795 649 5795 683
rect -5891 -587 -5857 587
rect 5857 -587 5891 587
rect -5795 -683 5795 -649
<< poly >>
rect -5745 581 -5679 597
rect -5745 547 -5729 581
rect -5695 547 -5679 581
rect -5745 531 -5679 547
rect -5553 581 -5487 597
rect -5553 547 -5537 581
rect -5503 547 -5487 581
rect -5727 509 -5697 531
rect -5631 509 -5601 535
rect -5553 531 -5487 547
rect -5361 581 -5295 597
rect -5361 547 -5345 581
rect -5311 547 -5295 581
rect -5535 509 -5505 531
rect -5439 509 -5409 535
rect -5361 531 -5295 547
rect -5169 581 -5103 597
rect -5169 547 -5153 581
rect -5119 547 -5103 581
rect -5343 509 -5313 531
rect -5247 509 -5217 535
rect -5169 531 -5103 547
rect -4977 581 -4911 597
rect -4977 547 -4961 581
rect -4927 547 -4911 581
rect -5151 509 -5121 531
rect -5055 509 -5025 535
rect -4977 531 -4911 547
rect -4785 581 -4719 597
rect -4785 547 -4769 581
rect -4735 547 -4719 581
rect -4959 509 -4929 531
rect -4863 509 -4833 535
rect -4785 531 -4719 547
rect -4593 581 -4527 597
rect -4593 547 -4577 581
rect -4543 547 -4527 581
rect -4767 509 -4737 531
rect -4671 509 -4641 535
rect -4593 531 -4527 547
rect -4401 581 -4335 597
rect -4401 547 -4385 581
rect -4351 547 -4335 581
rect -4575 509 -4545 531
rect -4479 509 -4449 535
rect -4401 531 -4335 547
rect -4209 581 -4143 597
rect -4209 547 -4193 581
rect -4159 547 -4143 581
rect -4383 509 -4353 531
rect -4287 509 -4257 535
rect -4209 531 -4143 547
rect -4017 581 -3951 597
rect -4017 547 -4001 581
rect -3967 547 -3951 581
rect -4191 509 -4161 531
rect -4095 509 -4065 535
rect -4017 531 -3951 547
rect -3825 581 -3759 597
rect -3825 547 -3809 581
rect -3775 547 -3759 581
rect -3999 509 -3969 531
rect -3903 509 -3873 535
rect -3825 531 -3759 547
rect -3633 581 -3567 597
rect -3633 547 -3617 581
rect -3583 547 -3567 581
rect -3807 509 -3777 531
rect -3711 509 -3681 535
rect -3633 531 -3567 547
rect -3441 581 -3375 597
rect -3441 547 -3425 581
rect -3391 547 -3375 581
rect -3615 509 -3585 531
rect -3519 509 -3489 535
rect -3441 531 -3375 547
rect -3249 581 -3183 597
rect -3249 547 -3233 581
rect -3199 547 -3183 581
rect -3423 509 -3393 531
rect -3327 509 -3297 535
rect -3249 531 -3183 547
rect -3057 581 -2991 597
rect -3057 547 -3041 581
rect -3007 547 -2991 581
rect -3231 509 -3201 531
rect -3135 509 -3105 535
rect -3057 531 -2991 547
rect -2865 581 -2799 597
rect -2865 547 -2849 581
rect -2815 547 -2799 581
rect -3039 509 -3009 531
rect -2943 509 -2913 535
rect -2865 531 -2799 547
rect -2673 581 -2607 597
rect -2673 547 -2657 581
rect -2623 547 -2607 581
rect -2847 509 -2817 531
rect -2751 509 -2721 535
rect -2673 531 -2607 547
rect -2481 581 -2415 597
rect -2481 547 -2465 581
rect -2431 547 -2415 581
rect -2655 509 -2625 531
rect -2559 509 -2529 535
rect -2481 531 -2415 547
rect -2289 581 -2223 597
rect -2289 547 -2273 581
rect -2239 547 -2223 581
rect -2463 509 -2433 531
rect -2367 509 -2337 535
rect -2289 531 -2223 547
rect -2097 581 -2031 597
rect -2097 547 -2081 581
rect -2047 547 -2031 581
rect -2271 509 -2241 531
rect -2175 509 -2145 535
rect -2097 531 -2031 547
rect -1905 581 -1839 597
rect -1905 547 -1889 581
rect -1855 547 -1839 581
rect -2079 509 -2049 531
rect -1983 509 -1953 535
rect -1905 531 -1839 547
rect -1713 581 -1647 597
rect -1713 547 -1697 581
rect -1663 547 -1647 581
rect -1887 509 -1857 531
rect -1791 509 -1761 535
rect -1713 531 -1647 547
rect -1521 581 -1455 597
rect -1521 547 -1505 581
rect -1471 547 -1455 581
rect -1695 509 -1665 531
rect -1599 509 -1569 535
rect -1521 531 -1455 547
rect -1329 581 -1263 597
rect -1329 547 -1313 581
rect -1279 547 -1263 581
rect -1503 509 -1473 531
rect -1407 509 -1377 535
rect -1329 531 -1263 547
rect -1137 581 -1071 597
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -1311 509 -1281 531
rect -1215 509 -1185 535
rect -1137 531 -1071 547
rect -945 581 -879 597
rect -945 547 -929 581
rect -895 547 -879 581
rect -1119 509 -1089 531
rect -1023 509 -993 535
rect -945 531 -879 547
rect -753 581 -687 597
rect -753 547 -737 581
rect -703 547 -687 581
rect -927 509 -897 531
rect -831 509 -801 535
rect -753 531 -687 547
rect -561 581 -495 597
rect -561 547 -545 581
rect -511 547 -495 581
rect -735 509 -705 531
rect -639 509 -609 535
rect -561 531 -495 547
rect -369 581 -303 597
rect -369 547 -353 581
rect -319 547 -303 581
rect -543 509 -513 531
rect -447 509 -417 535
rect -369 531 -303 547
rect -177 581 -111 597
rect -177 547 -161 581
rect -127 547 -111 581
rect -351 509 -321 531
rect -255 509 -225 535
rect -177 531 -111 547
rect 15 581 81 597
rect 15 547 31 581
rect 65 547 81 581
rect -159 509 -129 531
rect -63 509 -33 535
rect 15 531 81 547
rect 207 581 273 597
rect 207 547 223 581
rect 257 547 273 581
rect 33 509 63 531
rect 129 509 159 535
rect 207 531 273 547
rect 399 581 465 597
rect 399 547 415 581
rect 449 547 465 581
rect 225 509 255 531
rect 321 509 351 535
rect 399 531 465 547
rect 591 581 657 597
rect 591 547 607 581
rect 641 547 657 581
rect 417 509 447 531
rect 513 509 543 535
rect 591 531 657 547
rect 783 581 849 597
rect 783 547 799 581
rect 833 547 849 581
rect 609 509 639 531
rect 705 509 735 535
rect 783 531 849 547
rect 975 581 1041 597
rect 975 547 991 581
rect 1025 547 1041 581
rect 801 509 831 531
rect 897 509 927 535
rect 975 531 1041 547
rect 1167 581 1233 597
rect 1167 547 1183 581
rect 1217 547 1233 581
rect 993 509 1023 531
rect 1089 509 1119 535
rect 1167 531 1233 547
rect 1359 581 1425 597
rect 1359 547 1375 581
rect 1409 547 1425 581
rect 1185 509 1215 531
rect 1281 509 1311 535
rect 1359 531 1425 547
rect 1551 581 1617 597
rect 1551 547 1567 581
rect 1601 547 1617 581
rect 1377 509 1407 531
rect 1473 509 1503 535
rect 1551 531 1617 547
rect 1743 581 1809 597
rect 1743 547 1759 581
rect 1793 547 1809 581
rect 1569 509 1599 531
rect 1665 509 1695 535
rect 1743 531 1809 547
rect 1935 581 2001 597
rect 1935 547 1951 581
rect 1985 547 2001 581
rect 1761 509 1791 531
rect 1857 509 1887 535
rect 1935 531 2001 547
rect 2127 581 2193 597
rect 2127 547 2143 581
rect 2177 547 2193 581
rect 1953 509 1983 531
rect 2049 509 2079 535
rect 2127 531 2193 547
rect 2319 581 2385 597
rect 2319 547 2335 581
rect 2369 547 2385 581
rect 2145 509 2175 531
rect 2241 509 2271 535
rect 2319 531 2385 547
rect 2511 581 2577 597
rect 2511 547 2527 581
rect 2561 547 2577 581
rect 2337 509 2367 531
rect 2433 509 2463 535
rect 2511 531 2577 547
rect 2703 581 2769 597
rect 2703 547 2719 581
rect 2753 547 2769 581
rect 2529 509 2559 531
rect 2625 509 2655 535
rect 2703 531 2769 547
rect 2895 581 2961 597
rect 2895 547 2911 581
rect 2945 547 2961 581
rect 2721 509 2751 531
rect 2817 509 2847 535
rect 2895 531 2961 547
rect 3087 581 3153 597
rect 3087 547 3103 581
rect 3137 547 3153 581
rect 2913 509 2943 531
rect 3009 509 3039 535
rect 3087 531 3153 547
rect 3279 581 3345 597
rect 3279 547 3295 581
rect 3329 547 3345 581
rect 3105 509 3135 531
rect 3201 509 3231 535
rect 3279 531 3345 547
rect 3471 581 3537 597
rect 3471 547 3487 581
rect 3521 547 3537 581
rect 3297 509 3327 531
rect 3393 509 3423 535
rect 3471 531 3537 547
rect 3663 581 3729 597
rect 3663 547 3679 581
rect 3713 547 3729 581
rect 3489 509 3519 531
rect 3585 509 3615 535
rect 3663 531 3729 547
rect 3855 581 3921 597
rect 3855 547 3871 581
rect 3905 547 3921 581
rect 3681 509 3711 531
rect 3777 509 3807 535
rect 3855 531 3921 547
rect 4047 581 4113 597
rect 4047 547 4063 581
rect 4097 547 4113 581
rect 3873 509 3903 531
rect 3969 509 3999 535
rect 4047 531 4113 547
rect 4239 581 4305 597
rect 4239 547 4255 581
rect 4289 547 4305 581
rect 4065 509 4095 531
rect 4161 509 4191 535
rect 4239 531 4305 547
rect 4431 581 4497 597
rect 4431 547 4447 581
rect 4481 547 4497 581
rect 4257 509 4287 531
rect 4353 509 4383 535
rect 4431 531 4497 547
rect 4623 581 4689 597
rect 4623 547 4639 581
rect 4673 547 4689 581
rect 4449 509 4479 531
rect 4545 509 4575 535
rect 4623 531 4689 547
rect 4815 581 4881 597
rect 4815 547 4831 581
rect 4865 547 4881 581
rect 4641 509 4671 531
rect 4737 509 4767 535
rect 4815 531 4881 547
rect 5007 581 5073 597
rect 5007 547 5023 581
rect 5057 547 5073 581
rect 4833 509 4863 531
rect 4929 509 4959 535
rect 5007 531 5073 547
rect 5199 581 5265 597
rect 5199 547 5215 581
rect 5249 547 5265 581
rect 5025 509 5055 531
rect 5121 509 5151 535
rect 5199 531 5265 547
rect 5391 581 5457 597
rect 5391 547 5407 581
rect 5441 547 5457 581
rect 5217 509 5247 531
rect 5313 509 5343 535
rect 5391 531 5457 547
rect 5583 581 5649 597
rect 5583 547 5599 581
rect 5633 547 5649 581
rect 5409 509 5439 531
rect 5505 509 5535 535
rect 5583 531 5649 547
rect 5601 509 5631 531
rect 5697 509 5727 535
rect -5727 83 -5697 109
rect -5631 87 -5601 109
rect -5649 71 -5583 87
rect -5535 83 -5505 109
rect -5439 87 -5409 109
rect -5649 37 -5633 71
rect -5599 37 -5583 71
rect -5649 21 -5583 37
rect -5457 71 -5391 87
rect -5343 83 -5313 109
rect -5247 87 -5217 109
rect -5457 37 -5441 71
rect -5407 37 -5391 71
rect -5457 21 -5391 37
rect -5265 71 -5199 87
rect -5151 83 -5121 109
rect -5055 87 -5025 109
rect -5265 37 -5249 71
rect -5215 37 -5199 71
rect -5265 21 -5199 37
rect -5073 71 -5007 87
rect -4959 83 -4929 109
rect -4863 87 -4833 109
rect -5073 37 -5057 71
rect -5023 37 -5007 71
rect -5073 21 -5007 37
rect -4881 71 -4815 87
rect -4767 83 -4737 109
rect -4671 87 -4641 109
rect -4881 37 -4865 71
rect -4831 37 -4815 71
rect -4881 21 -4815 37
rect -4689 71 -4623 87
rect -4575 83 -4545 109
rect -4479 87 -4449 109
rect -4689 37 -4673 71
rect -4639 37 -4623 71
rect -4689 21 -4623 37
rect -4497 71 -4431 87
rect -4383 83 -4353 109
rect -4287 87 -4257 109
rect -4497 37 -4481 71
rect -4447 37 -4431 71
rect -4497 21 -4431 37
rect -4305 71 -4239 87
rect -4191 83 -4161 109
rect -4095 87 -4065 109
rect -4305 37 -4289 71
rect -4255 37 -4239 71
rect -4305 21 -4239 37
rect -4113 71 -4047 87
rect -3999 83 -3969 109
rect -3903 87 -3873 109
rect -4113 37 -4097 71
rect -4063 37 -4047 71
rect -4113 21 -4047 37
rect -3921 71 -3855 87
rect -3807 83 -3777 109
rect -3711 87 -3681 109
rect -3921 37 -3905 71
rect -3871 37 -3855 71
rect -3921 21 -3855 37
rect -3729 71 -3663 87
rect -3615 83 -3585 109
rect -3519 87 -3489 109
rect -3729 37 -3713 71
rect -3679 37 -3663 71
rect -3729 21 -3663 37
rect -3537 71 -3471 87
rect -3423 83 -3393 109
rect -3327 87 -3297 109
rect -3537 37 -3521 71
rect -3487 37 -3471 71
rect -3537 21 -3471 37
rect -3345 71 -3279 87
rect -3231 83 -3201 109
rect -3135 87 -3105 109
rect -3345 37 -3329 71
rect -3295 37 -3279 71
rect -3345 21 -3279 37
rect -3153 71 -3087 87
rect -3039 83 -3009 109
rect -2943 87 -2913 109
rect -3153 37 -3137 71
rect -3103 37 -3087 71
rect -3153 21 -3087 37
rect -2961 71 -2895 87
rect -2847 83 -2817 109
rect -2751 87 -2721 109
rect -2961 37 -2945 71
rect -2911 37 -2895 71
rect -2961 21 -2895 37
rect -2769 71 -2703 87
rect -2655 83 -2625 109
rect -2559 87 -2529 109
rect -2769 37 -2753 71
rect -2719 37 -2703 71
rect -2769 21 -2703 37
rect -2577 71 -2511 87
rect -2463 83 -2433 109
rect -2367 87 -2337 109
rect -2577 37 -2561 71
rect -2527 37 -2511 71
rect -2577 21 -2511 37
rect -2385 71 -2319 87
rect -2271 83 -2241 109
rect -2175 87 -2145 109
rect -2385 37 -2369 71
rect -2335 37 -2319 71
rect -2385 21 -2319 37
rect -2193 71 -2127 87
rect -2079 83 -2049 109
rect -1983 87 -1953 109
rect -2193 37 -2177 71
rect -2143 37 -2127 71
rect -2193 21 -2127 37
rect -2001 71 -1935 87
rect -1887 83 -1857 109
rect -1791 87 -1761 109
rect -2001 37 -1985 71
rect -1951 37 -1935 71
rect -2001 21 -1935 37
rect -1809 71 -1743 87
rect -1695 83 -1665 109
rect -1599 87 -1569 109
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1809 21 -1743 37
rect -1617 71 -1551 87
rect -1503 83 -1473 109
rect -1407 87 -1377 109
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1617 21 -1551 37
rect -1425 71 -1359 87
rect -1311 83 -1281 109
rect -1215 87 -1185 109
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1425 21 -1359 37
rect -1233 71 -1167 87
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1233 21 -1167 37
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1185 83 1215 109
rect 1281 87 1311 109
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect 1263 71 1329 87
rect 1377 83 1407 109
rect 1473 87 1503 109
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1263 21 1329 37
rect 1455 71 1521 87
rect 1569 83 1599 109
rect 1665 87 1695 109
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1455 21 1521 37
rect 1647 71 1713 87
rect 1761 83 1791 109
rect 1857 87 1887 109
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1647 21 1713 37
rect 1839 71 1905 87
rect 1953 83 1983 109
rect 2049 87 2079 109
rect 1839 37 1855 71
rect 1889 37 1905 71
rect 1839 21 1905 37
rect 2031 71 2097 87
rect 2145 83 2175 109
rect 2241 87 2271 109
rect 2031 37 2047 71
rect 2081 37 2097 71
rect 2031 21 2097 37
rect 2223 71 2289 87
rect 2337 83 2367 109
rect 2433 87 2463 109
rect 2223 37 2239 71
rect 2273 37 2289 71
rect 2223 21 2289 37
rect 2415 71 2481 87
rect 2529 83 2559 109
rect 2625 87 2655 109
rect 2415 37 2431 71
rect 2465 37 2481 71
rect 2415 21 2481 37
rect 2607 71 2673 87
rect 2721 83 2751 109
rect 2817 87 2847 109
rect 2607 37 2623 71
rect 2657 37 2673 71
rect 2607 21 2673 37
rect 2799 71 2865 87
rect 2913 83 2943 109
rect 3009 87 3039 109
rect 2799 37 2815 71
rect 2849 37 2865 71
rect 2799 21 2865 37
rect 2991 71 3057 87
rect 3105 83 3135 109
rect 3201 87 3231 109
rect 2991 37 3007 71
rect 3041 37 3057 71
rect 2991 21 3057 37
rect 3183 71 3249 87
rect 3297 83 3327 109
rect 3393 87 3423 109
rect 3183 37 3199 71
rect 3233 37 3249 71
rect 3183 21 3249 37
rect 3375 71 3441 87
rect 3489 83 3519 109
rect 3585 87 3615 109
rect 3375 37 3391 71
rect 3425 37 3441 71
rect 3375 21 3441 37
rect 3567 71 3633 87
rect 3681 83 3711 109
rect 3777 87 3807 109
rect 3567 37 3583 71
rect 3617 37 3633 71
rect 3567 21 3633 37
rect 3759 71 3825 87
rect 3873 83 3903 109
rect 3969 87 3999 109
rect 3759 37 3775 71
rect 3809 37 3825 71
rect 3759 21 3825 37
rect 3951 71 4017 87
rect 4065 83 4095 109
rect 4161 87 4191 109
rect 3951 37 3967 71
rect 4001 37 4017 71
rect 3951 21 4017 37
rect 4143 71 4209 87
rect 4257 83 4287 109
rect 4353 87 4383 109
rect 4143 37 4159 71
rect 4193 37 4209 71
rect 4143 21 4209 37
rect 4335 71 4401 87
rect 4449 83 4479 109
rect 4545 87 4575 109
rect 4335 37 4351 71
rect 4385 37 4401 71
rect 4335 21 4401 37
rect 4527 71 4593 87
rect 4641 83 4671 109
rect 4737 87 4767 109
rect 4527 37 4543 71
rect 4577 37 4593 71
rect 4527 21 4593 37
rect 4719 71 4785 87
rect 4833 83 4863 109
rect 4929 87 4959 109
rect 4719 37 4735 71
rect 4769 37 4785 71
rect 4719 21 4785 37
rect 4911 71 4977 87
rect 5025 83 5055 109
rect 5121 87 5151 109
rect 4911 37 4927 71
rect 4961 37 4977 71
rect 4911 21 4977 37
rect 5103 71 5169 87
rect 5217 83 5247 109
rect 5313 87 5343 109
rect 5103 37 5119 71
rect 5153 37 5169 71
rect 5103 21 5169 37
rect 5295 71 5361 87
rect 5409 83 5439 109
rect 5505 87 5535 109
rect 5295 37 5311 71
rect 5345 37 5361 71
rect 5295 21 5361 37
rect 5487 71 5553 87
rect 5601 83 5631 109
rect 5697 87 5727 109
rect 5487 37 5503 71
rect 5537 37 5553 71
rect 5487 21 5553 37
rect 5679 71 5745 87
rect 5679 37 5695 71
rect 5729 37 5745 71
rect 5679 21 5745 37
rect -5649 -37 -5583 -21
rect -5649 -71 -5633 -37
rect -5599 -71 -5583 -37
rect -5727 -109 -5697 -83
rect -5649 -87 -5583 -71
rect -5457 -37 -5391 -21
rect -5457 -71 -5441 -37
rect -5407 -71 -5391 -37
rect -5631 -109 -5601 -87
rect -5535 -109 -5505 -83
rect -5457 -87 -5391 -71
rect -5265 -37 -5199 -21
rect -5265 -71 -5249 -37
rect -5215 -71 -5199 -37
rect -5439 -109 -5409 -87
rect -5343 -109 -5313 -83
rect -5265 -87 -5199 -71
rect -5073 -37 -5007 -21
rect -5073 -71 -5057 -37
rect -5023 -71 -5007 -37
rect -5247 -109 -5217 -87
rect -5151 -109 -5121 -83
rect -5073 -87 -5007 -71
rect -4881 -37 -4815 -21
rect -4881 -71 -4865 -37
rect -4831 -71 -4815 -37
rect -5055 -109 -5025 -87
rect -4959 -109 -4929 -83
rect -4881 -87 -4815 -71
rect -4689 -37 -4623 -21
rect -4689 -71 -4673 -37
rect -4639 -71 -4623 -37
rect -4863 -109 -4833 -87
rect -4767 -109 -4737 -83
rect -4689 -87 -4623 -71
rect -4497 -37 -4431 -21
rect -4497 -71 -4481 -37
rect -4447 -71 -4431 -37
rect -4671 -109 -4641 -87
rect -4575 -109 -4545 -83
rect -4497 -87 -4431 -71
rect -4305 -37 -4239 -21
rect -4305 -71 -4289 -37
rect -4255 -71 -4239 -37
rect -4479 -109 -4449 -87
rect -4383 -109 -4353 -83
rect -4305 -87 -4239 -71
rect -4113 -37 -4047 -21
rect -4113 -71 -4097 -37
rect -4063 -71 -4047 -37
rect -4287 -109 -4257 -87
rect -4191 -109 -4161 -83
rect -4113 -87 -4047 -71
rect -3921 -37 -3855 -21
rect -3921 -71 -3905 -37
rect -3871 -71 -3855 -37
rect -4095 -109 -4065 -87
rect -3999 -109 -3969 -83
rect -3921 -87 -3855 -71
rect -3729 -37 -3663 -21
rect -3729 -71 -3713 -37
rect -3679 -71 -3663 -37
rect -3903 -109 -3873 -87
rect -3807 -109 -3777 -83
rect -3729 -87 -3663 -71
rect -3537 -37 -3471 -21
rect -3537 -71 -3521 -37
rect -3487 -71 -3471 -37
rect -3711 -109 -3681 -87
rect -3615 -109 -3585 -83
rect -3537 -87 -3471 -71
rect -3345 -37 -3279 -21
rect -3345 -71 -3329 -37
rect -3295 -71 -3279 -37
rect -3519 -109 -3489 -87
rect -3423 -109 -3393 -83
rect -3345 -87 -3279 -71
rect -3153 -37 -3087 -21
rect -3153 -71 -3137 -37
rect -3103 -71 -3087 -37
rect -3327 -109 -3297 -87
rect -3231 -109 -3201 -83
rect -3153 -87 -3087 -71
rect -2961 -37 -2895 -21
rect -2961 -71 -2945 -37
rect -2911 -71 -2895 -37
rect -3135 -109 -3105 -87
rect -3039 -109 -3009 -83
rect -2961 -87 -2895 -71
rect -2769 -37 -2703 -21
rect -2769 -71 -2753 -37
rect -2719 -71 -2703 -37
rect -2943 -109 -2913 -87
rect -2847 -109 -2817 -83
rect -2769 -87 -2703 -71
rect -2577 -37 -2511 -21
rect -2577 -71 -2561 -37
rect -2527 -71 -2511 -37
rect -2751 -109 -2721 -87
rect -2655 -109 -2625 -83
rect -2577 -87 -2511 -71
rect -2385 -37 -2319 -21
rect -2385 -71 -2369 -37
rect -2335 -71 -2319 -37
rect -2559 -109 -2529 -87
rect -2463 -109 -2433 -83
rect -2385 -87 -2319 -71
rect -2193 -37 -2127 -21
rect -2193 -71 -2177 -37
rect -2143 -71 -2127 -37
rect -2367 -109 -2337 -87
rect -2271 -109 -2241 -83
rect -2193 -87 -2127 -71
rect -2001 -37 -1935 -21
rect -2001 -71 -1985 -37
rect -1951 -71 -1935 -37
rect -2175 -109 -2145 -87
rect -2079 -109 -2049 -83
rect -2001 -87 -1935 -71
rect -1809 -37 -1743 -21
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1983 -109 -1953 -87
rect -1887 -109 -1857 -83
rect -1809 -87 -1743 -71
rect -1617 -37 -1551 -21
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1791 -109 -1761 -87
rect -1695 -109 -1665 -83
rect -1617 -87 -1551 -71
rect -1425 -37 -1359 -21
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1599 -109 -1569 -87
rect -1503 -109 -1473 -83
rect -1425 -87 -1359 -71
rect -1233 -37 -1167 -21
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -83
rect -1233 -87 -1167 -71
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1263 -37 1329 -21
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1089 -109 1119 -87
rect 1185 -109 1215 -83
rect 1263 -87 1329 -71
rect 1455 -37 1521 -21
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1281 -109 1311 -87
rect 1377 -109 1407 -83
rect 1455 -87 1521 -71
rect 1647 -37 1713 -21
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1473 -109 1503 -87
rect 1569 -109 1599 -83
rect 1647 -87 1713 -71
rect 1839 -37 1905 -21
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect 1665 -109 1695 -87
rect 1761 -109 1791 -83
rect 1839 -87 1905 -71
rect 2031 -37 2097 -21
rect 2031 -71 2047 -37
rect 2081 -71 2097 -37
rect 1857 -109 1887 -87
rect 1953 -109 1983 -83
rect 2031 -87 2097 -71
rect 2223 -37 2289 -21
rect 2223 -71 2239 -37
rect 2273 -71 2289 -37
rect 2049 -109 2079 -87
rect 2145 -109 2175 -83
rect 2223 -87 2289 -71
rect 2415 -37 2481 -21
rect 2415 -71 2431 -37
rect 2465 -71 2481 -37
rect 2241 -109 2271 -87
rect 2337 -109 2367 -83
rect 2415 -87 2481 -71
rect 2607 -37 2673 -21
rect 2607 -71 2623 -37
rect 2657 -71 2673 -37
rect 2433 -109 2463 -87
rect 2529 -109 2559 -83
rect 2607 -87 2673 -71
rect 2799 -37 2865 -21
rect 2799 -71 2815 -37
rect 2849 -71 2865 -37
rect 2625 -109 2655 -87
rect 2721 -109 2751 -83
rect 2799 -87 2865 -71
rect 2991 -37 3057 -21
rect 2991 -71 3007 -37
rect 3041 -71 3057 -37
rect 2817 -109 2847 -87
rect 2913 -109 2943 -83
rect 2991 -87 3057 -71
rect 3183 -37 3249 -21
rect 3183 -71 3199 -37
rect 3233 -71 3249 -37
rect 3009 -109 3039 -87
rect 3105 -109 3135 -83
rect 3183 -87 3249 -71
rect 3375 -37 3441 -21
rect 3375 -71 3391 -37
rect 3425 -71 3441 -37
rect 3201 -109 3231 -87
rect 3297 -109 3327 -83
rect 3375 -87 3441 -71
rect 3567 -37 3633 -21
rect 3567 -71 3583 -37
rect 3617 -71 3633 -37
rect 3393 -109 3423 -87
rect 3489 -109 3519 -83
rect 3567 -87 3633 -71
rect 3759 -37 3825 -21
rect 3759 -71 3775 -37
rect 3809 -71 3825 -37
rect 3585 -109 3615 -87
rect 3681 -109 3711 -83
rect 3759 -87 3825 -71
rect 3951 -37 4017 -21
rect 3951 -71 3967 -37
rect 4001 -71 4017 -37
rect 3777 -109 3807 -87
rect 3873 -109 3903 -83
rect 3951 -87 4017 -71
rect 4143 -37 4209 -21
rect 4143 -71 4159 -37
rect 4193 -71 4209 -37
rect 3969 -109 3999 -87
rect 4065 -109 4095 -83
rect 4143 -87 4209 -71
rect 4335 -37 4401 -21
rect 4335 -71 4351 -37
rect 4385 -71 4401 -37
rect 4161 -109 4191 -87
rect 4257 -109 4287 -83
rect 4335 -87 4401 -71
rect 4527 -37 4593 -21
rect 4527 -71 4543 -37
rect 4577 -71 4593 -37
rect 4353 -109 4383 -87
rect 4449 -109 4479 -83
rect 4527 -87 4593 -71
rect 4719 -37 4785 -21
rect 4719 -71 4735 -37
rect 4769 -71 4785 -37
rect 4545 -109 4575 -87
rect 4641 -109 4671 -83
rect 4719 -87 4785 -71
rect 4911 -37 4977 -21
rect 4911 -71 4927 -37
rect 4961 -71 4977 -37
rect 4737 -109 4767 -87
rect 4833 -109 4863 -83
rect 4911 -87 4977 -71
rect 5103 -37 5169 -21
rect 5103 -71 5119 -37
rect 5153 -71 5169 -37
rect 4929 -109 4959 -87
rect 5025 -109 5055 -83
rect 5103 -87 5169 -71
rect 5295 -37 5361 -21
rect 5295 -71 5311 -37
rect 5345 -71 5361 -37
rect 5121 -109 5151 -87
rect 5217 -109 5247 -83
rect 5295 -87 5361 -71
rect 5487 -37 5553 -21
rect 5487 -71 5503 -37
rect 5537 -71 5553 -37
rect 5313 -109 5343 -87
rect 5409 -109 5439 -83
rect 5487 -87 5553 -71
rect 5679 -37 5745 -21
rect 5679 -71 5695 -37
rect 5729 -71 5745 -37
rect 5505 -109 5535 -87
rect 5601 -109 5631 -83
rect 5679 -87 5745 -71
rect 5697 -109 5727 -87
rect -5727 -531 -5697 -509
rect -5745 -547 -5679 -531
rect -5631 -535 -5601 -509
rect -5535 -531 -5505 -509
rect -5745 -581 -5729 -547
rect -5695 -581 -5679 -547
rect -5745 -597 -5679 -581
rect -5553 -547 -5487 -531
rect -5439 -535 -5409 -509
rect -5343 -531 -5313 -509
rect -5553 -581 -5537 -547
rect -5503 -581 -5487 -547
rect -5553 -597 -5487 -581
rect -5361 -547 -5295 -531
rect -5247 -535 -5217 -509
rect -5151 -531 -5121 -509
rect -5361 -581 -5345 -547
rect -5311 -581 -5295 -547
rect -5361 -597 -5295 -581
rect -5169 -547 -5103 -531
rect -5055 -535 -5025 -509
rect -4959 -531 -4929 -509
rect -5169 -581 -5153 -547
rect -5119 -581 -5103 -547
rect -5169 -597 -5103 -581
rect -4977 -547 -4911 -531
rect -4863 -535 -4833 -509
rect -4767 -531 -4737 -509
rect -4977 -581 -4961 -547
rect -4927 -581 -4911 -547
rect -4977 -597 -4911 -581
rect -4785 -547 -4719 -531
rect -4671 -535 -4641 -509
rect -4575 -531 -4545 -509
rect -4785 -581 -4769 -547
rect -4735 -581 -4719 -547
rect -4785 -597 -4719 -581
rect -4593 -547 -4527 -531
rect -4479 -535 -4449 -509
rect -4383 -531 -4353 -509
rect -4593 -581 -4577 -547
rect -4543 -581 -4527 -547
rect -4593 -597 -4527 -581
rect -4401 -547 -4335 -531
rect -4287 -535 -4257 -509
rect -4191 -531 -4161 -509
rect -4401 -581 -4385 -547
rect -4351 -581 -4335 -547
rect -4401 -597 -4335 -581
rect -4209 -547 -4143 -531
rect -4095 -535 -4065 -509
rect -3999 -531 -3969 -509
rect -4209 -581 -4193 -547
rect -4159 -581 -4143 -547
rect -4209 -597 -4143 -581
rect -4017 -547 -3951 -531
rect -3903 -535 -3873 -509
rect -3807 -531 -3777 -509
rect -4017 -581 -4001 -547
rect -3967 -581 -3951 -547
rect -4017 -597 -3951 -581
rect -3825 -547 -3759 -531
rect -3711 -535 -3681 -509
rect -3615 -531 -3585 -509
rect -3825 -581 -3809 -547
rect -3775 -581 -3759 -547
rect -3825 -597 -3759 -581
rect -3633 -547 -3567 -531
rect -3519 -535 -3489 -509
rect -3423 -531 -3393 -509
rect -3633 -581 -3617 -547
rect -3583 -581 -3567 -547
rect -3633 -597 -3567 -581
rect -3441 -547 -3375 -531
rect -3327 -535 -3297 -509
rect -3231 -531 -3201 -509
rect -3441 -581 -3425 -547
rect -3391 -581 -3375 -547
rect -3441 -597 -3375 -581
rect -3249 -547 -3183 -531
rect -3135 -535 -3105 -509
rect -3039 -531 -3009 -509
rect -3249 -581 -3233 -547
rect -3199 -581 -3183 -547
rect -3249 -597 -3183 -581
rect -3057 -547 -2991 -531
rect -2943 -535 -2913 -509
rect -2847 -531 -2817 -509
rect -3057 -581 -3041 -547
rect -3007 -581 -2991 -547
rect -3057 -597 -2991 -581
rect -2865 -547 -2799 -531
rect -2751 -535 -2721 -509
rect -2655 -531 -2625 -509
rect -2865 -581 -2849 -547
rect -2815 -581 -2799 -547
rect -2865 -597 -2799 -581
rect -2673 -547 -2607 -531
rect -2559 -535 -2529 -509
rect -2463 -531 -2433 -509
rect -2673 -581 -2657 -547
rect -2623 -581 -2607 -547
rect -2673 -597 -2607 -581
rect -2481 -547 -2415 -531
rect -2367 -535 -2337 -509
rect -2271 -531 -2241 -509
rect -2481 -581 -2465 -547
rect -2431 -581 -2415 -547
rect -2481 -597 -2415 -581
rect -2289 -547 -2223 -531
rect -2175 -535 -2145 -509
rect -2079 -531 -2049 -509
rect -2289 -581 -2273 -547
rect -2239 -581 -2223 -547
rect -2289 -597 -2223 -581
rect -2097 -547 -2031 -531
rect -1983 -535 -1953 -509
rect -1887 -531 -1857 -509
rect -2097 -581 -2081 -547
rect -2047 -581 -2031 -547
rect -2097 -597 -2031 -581
rect -1905 -547 -1839 -531
rect -1791 -535 -1761 -509
rect -1695 -531 -1665 -509
rect -1905 -581 -1889 -547
rect -1855 -581 -1839 -547
rect -1905 -597 -1839 -581
rect -1713 -547 -1647 -531
rect -1599 -535 -1569 -509
rect -1503 -531 -1473 -509
rect -1713 -581 -1697 -547
rect -1663 -581 -1647 -547
rect -1713 -597 -1647 -581
rect -1521 -547 -1455 -531
rect -1407 -535 -1377 -509
rect -1311 -531 -1281 -509
rect -1521 -581 -1505 -547
rect -1471 -581 -1455 -547
rect -1521 -597 -1455 -581
rect -1329 -547 -1263 -531
rect -1215 -535 -1185 -509
rect -1119 -531 -1089 -509
rect -1329 -581 -1313 -547
rect -1279 -581 -1263 -547
rect -1329 -597 -1263 -581
rect -1137 -547 -1071 -531
rect -1023 -535 -993 -509
rect -927 -531 -897 -509
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -1137 -597 -1071 -581
rect -945 -547 -879 -531
rect -831 -535 -801 -509
rect -735 -531 -705 -509
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -945 -597 -879 -581
rect -753 -547 -687 -531
rect -639 -535 -609 -509
rect -543 -531 -513 -509
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -753 -597 -687 -581
rect -561 -547 -495 -531
rect -447 -535 -417 -509
rect -351 -531 -321 -509
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -255 -535 -225 -509
rect -159 -531 -129 -509
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -63 -535 -33 -509
rect 33 -531 63 -509
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 129 -535 159 -509
rect 225 -531 255 -509
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 321 -535 351 -509
rect 417 -531 447 -509
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 513 -535 543 -509
rect 609 -531 639 -509
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
rect 591 -547 657 -531
rect 705 -535 735 -509
rect 801 -531 831 -509
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 591 -597 657 -581
rect 783 -547 849 -531
rect 897 -535 927 -509
rect 993 -531 1023 -509
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 783 -597 849 -581
rect 975 -547 1041 -531
rect 1089 -535 1119 -509
rect 1185 -531 1215 -509
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 975 -597 1041 -581
rect 1167 -547 1233 -531
rect 1281 -535 1311 -509
rect 1377 -531 1407 -509
rect 1167 -581 1183 -547
rect 1217 -581 1233 -547
rect 1167 -597 1233 -581
rect 1359 -547 1425 -531
rect 1473 -535 1503 -509
rect 1569 -531 1599 -509
rect 1359 -581 1375 -547
rect 1409 -581 1425 -547
rect 1359 -597 1425 -581
rect 1551 -547 1617 -531
rect 1665 -535 1695 -509
rect 1761 -531 1791 -509
rect 1551 -581 1567 -547
rect 1601 -581 1617 -547
rect 1551 -597 1617 -581
rect 1743 -547 1809 -531
rect 1857 -535 1887 -509
rect 1953 -531 1983 -509
rect 1743 -581 1759 -547
rect 1793 -581 1809 -547
rect 1743 -597 1809 -581
rect 1935 -547 2001 -531
rect 2049 -535 2079 -509
rect 2145 -531 2175 -509
rect 1935 -581 1951 -547
rect 1985 -581 2001 -547
rect 1935 -597 2001 -581
rect 2127 -547 2193 -531
rect 2241 -535 2271 -509
rect 2337 -531 2367 -509
rect 2127 -581 2143 -547
rect 2177 -581 2193 -547
rect 2127 -597 2193 -581
rect 2319 -547 2385 -531
rect 2433 -535 2463 -509
rect 2529 -531 2559 -509
rect 2319 -581 2335 -547
rect 2369 -581 2385 -547
rect 2319 -597 2385 -581
rect 2511 -547 2577 -531
rect 2625 -535 2655 -509
rect 2721 -531 2751 -509
rect 2511 -581 2527 -547
rect 2561 -581 2577 -547
rect 2511 -597 2577 -581
rect 2703 -547 2769 -531
rect 2817 -535 2847 -509
rect 2913 -531 2943 -509
rect 2703 -581 2719 -547
rect 2753 -581 2769 -547
rect 2703 -597 2769 -581
rect 2895 -547 2961 -531
rect 3009 -535 3039 -509
rect 3105 -531 3135 -509
rect 2895 -581 2911 -547
rect 2945 -581 2961 -547
rect 2895 -597 2961 -581
rect 3087 -547 3153 -531
rect 3201 -535 3231 -509
rect 3297 -531 3327 -509
rect 3087 -581 3103 -547
rect 3137 -581 3153 -547
rect 3087 -597 3153 -581
rect 3279 -547 3345 -531
rect 3393 -535 3423 -509
rect 3489 -531 3519 -509
rect 3279 -581 3295 -547
rect 3329 -581 3345 -547
rect 3279 -597 3345 -581
rect 3471 -547 3537 -531
rect 3585 -535 3615 -509
rect 3681 -531 3711 -509
rect 3471 -581 3487 -547
rect 3521 -581 3537 -547
rect 3471 -597 3537 -581
rect 3663 -547 3729 -531
rect 3777 -535 3807 -509
rect 3873 -531 3903 -509
rect 3663 -581 3679 -547
rect 3713 -581 3729 -547
rect 3663 -597 3729 -581
rect 3855 -547 3921 -531
rect 3969 -535 3999 -509
rect 4065 -531 4095 -509
rect 3855 -581 3871 -547
rect 3905 -581 3921 -547
rect 3855 -597 3921 -581
rect 4047 -547 4113 -531
rect 4161 -535 4191 -509
rect 4257 -531 4287 -509
rect 4047 -581 4063 -547
rect 4097 -581 4113 -547
rect 4047 -597 4113 -581
rect 4239 -547 4305 -531
rect 4353 -535 4383 -509
rect 4449 -531 4479 -509
rect 4239 -581 4255 -547
rect 4289 -581 4305 -547
rect 4239 -597 4305 -581
rect 4431 -547 4497 -531
rect 4545 -535 4575 -509
rect 4641 -531 4671 -509
rect 4431 -581 4447 -547
rect 4481 -581 4497 -547
rect 4431 -597 4497 -581
rect 4623 -547 4689 -531
rect 4737 -535 4767 -509
rect 4833 -531 4863 -509
rect 4623 -581 4639 -547
rect 4673 -581 4689 -547
rect 4623 -597 4689 -581
rect 4815 -547 4881 -531
rect 4929 -535 4959 -509
rect 5025 -531 5055 -509
rect 4815 -581 4831 -547
rect 4865 -581 4881 -547
rect 4815 -597 4881 -581
rect 5007 -547 5073 -531
rect 5121 -535 5151 -509
rect 5217 -531 5247 -509
rect 5007 -581 5023 -547
rect 5057 -581 5073 -547
rect 5007 -597 5073 -581
rect 5199 -547 5265 -531
rect 5313 -535 5343 -509
rect 5409 -531 5439 -509
rect 5199 -581 5215 -547
rect 5249 -581 5265 -547
rect 5199 -597 5265 -581
rect 5391 -547 5457 -531
rect 5505 -535 5535 -509
rect 5601 -531 5631 -509
rect 5391 -581 5407 -547
rect 5441 -581 5457 -547
rect 5391 -597 5457 -581
rect 5583 -547 5649 -531
rect 5697 -535 5727 -509
rect 5583 -581 5599 -547
rect 5633 -581 5649 -547
rect 5583 -597 5649 -581
<< polycont >>
rect -5729 547 -5695 581
rect -5537 547 -5503 581
rect -5345 547 -5311 581
rect -5153 547 -5119 581
rect -4961 547 -4927 581
rect -4769 547 -4735 581
rect -4577 547 -4543 581
rect -4385 547 -4351 581
rect -4193 547 -4159 581
rect -4001 547 -3967 581
rect -3809 547 -3775 581
rect -3617 547 -3583 581
rect -3425 547 -3391 581
rect -3233 547 -3199 581
rect -3041 547 -3007 581
rect -2849 547 -2815 581
rect -2657 547 -2623 581
rect -2465 547 -2431 581
rect -2273 547 -2239 581
rect -2081 547 -2047 581
rect -1889 547 -1855 581
rect -1697 547 -1663 581
rect -1505 547 -1471 581
rect -1313 547 -1279 581
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect 1183 547 1217 581
rect 1375 547 1409 581
rect 1567 547 1601 581
rect 1759 547 1793 581
rect 1951 547 1985 581
rect 2143 547 2177 581
rect 2335 547 2369 581
rect 2527 547 2561 581
rect 2719 547 2753 581
rect 2911 547 2945 581
rect 3103 547 3137 581
rect 3295 547 3329 581
rect 3487 547 3521 581
rect 3679 547 3713 581
rect 3871 547 3905 581
rect 4063 547 4097 581
rect 4255 547 4289 581
rect 4447 547 4481 581
rect 4639 547 4673 581
rect 4831 547 4865 581
rect 5023 547 5057 581
rect 5215 547 5249 581
rect 5407 547 5441 581
rect 5599 547 5633 581
rect -5633 37 -5599 71
rect -5441 37 -5407 71
rect -5249 37 -5215 71
rect -5057 37 -5023 71
rect -4865 37 -4831 71
rect -4673 37 -4639 71
rect -4481 37 -4447 71
rect -4289 37 -4255 71
rect -4097 37 -4063 71
rect -3905 37 -3871 71
rect -3713 37 -3679 71
rect -3521 37 -3487 71
rect -3329 37 -3295 71
rect -3137 37 -3103 71
rect -2945 37 -2911 71
rect -2753 37 -2719 71
rect -2561 37 -2527 71
rect -2369 37 -2335 71
rect -2177 37 -2143 71
rect -1985 37 -1951 71
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect 2047 37 2081 71
rect 2239 37 2273 71
rect 2431 37 2465 71
rect 2623 37 2657 71
rect 2815 37 2849 71
rect 3007 37 3041 71
rect 3199 37 3233 71
rect 3391 37 3425 71
rect 3583 37 3617 71
rect 3775 37 3809 71
rect 3967 37 4001 71
rect 4159 37 4193 71
rect 4351 37 4385 71
rect 4543 37 4577 71
rect 4735 37 4769 71
rect 4927 37 4961 71
rect 5119 37 5153 71
rect 5311 37 5345 71
rect 5503 37 5537 71
rect 5695 37 5729 71
rect -5633 -71 -5599 -37
rect -5441 -71 -5407 -37
rect -5249 -71 -5215 -37
rect -5057 -71 -5023 -37
rect -4865 -71 -4831 -37
rect -4673 -71 -4639 -37
rect -4481 -71 -4447 -37
rect -4289 -71 -4255 -37
rect -4097 -71 -4063 -37
rect -3905 -71 -3871 -37
rect -3713 -71 -3679 -37
rect -3521 -71 -3487 -37
rect -3329 -71 -3295 -37
rect -3137 -71 -3103 -37
rect -2945 -71 -2911 -37
rect -2753 -71 -2719 -37
rect -2561 -71 -2527 -37
rect -2369 -71 -2335 -37
rect -2177 -71 -2143 -37
rect -1985 -71 -1951 -37
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect 2047 -71 2081 -37
rect 2239 -71 2273 -37
rect 2431 -71 2465 -37
rect 2623 -71 2657 -37
rect 2815 -71 2849 -37
rect 3007 -71 3041 -37
rect 3199 -71 3233 -37
rect 3391 -71 3425 -37
rect 3583 -71 3617 -37
rect 3775 -71 3809 -37
rect 3967 -71 4001 -37
rect 4159 -71 4193 -37
rect 4351 -71 4385 -37
rect 4543 -71 4577 -37
rect 4735 -71 4769 -37
rect 4927 -71 4961 -37
rect 5119 -71 5153 -37
rect 5311 -71 5345 -37
rect 5503 -71 5537 -37
rect 5695 -71 5729 -37
rect -5729 -581 -5695 -547
rect -5537 -581 -5503 -547
rect -5345 -581 -5311 -547
rect -5153 -581 -5119 -547
rect -4961 -581 -4927 -547
rect -4769 -581 -4735 -547
rect -4577 -581 -4543 -547
rect -4385 -581 -4351 -547
rect -4193 -581 -4159 -547
rect -4001 -581 -3967 -547
rect -3809 -581 -3775 -547
rect -3617 -581 -3583 -547
rect -3425 -581 -3391 -547
rect -3233 -581 -3199 -547
rect -3041 -581 -3007 -547
rect -2849 -581 -2815 -547
rect -2657 -581 -2623 -547
rect -2465 -581 -2431 -547
rect -2273 -581 -2239 -547
rect -2081 -581 -2047 -547
rect -1889 -581 -1855 -547
rect -1697 -581 -1663 -547
rect -1505 -581 -1471 -547
rect -1313 -581 -1279 -547
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect 1183 -581 1217 -547
rect 1375 -581 1409 -547
rect 1567 -581 1601 -547
rect 1759 -581 1793 -547
rect 1951 -581 1985 -547
rect 2143 -581 2177 -547
rect 2335 -581 2369 -547
rect 2527 -581 2561 -547
rect 2719 -581 2753 -547
rect 2911 -581 2945 -547
rect 3103 -581 3137 -547
rect 3295 -581 3329 -547
rect 3487 -581 3521 -547
rect 3679 -581 3713 -547
rect 3871 -581 3905 -547
rect 4063 -581 4097 -547
rect 4255 -581 4289 -547
rect 4447 -581 4481 -547
rect 4639 -581 4673 -547
rect 4831 -581 4865 -547
rect 5023 -581 5057 -547
rect 5215 -581 5249 -547
rect 5407 -581 5441 -547
rect 5599 -581 5633 -547
<< locali >>
rect -5891 649 -5795 683
rect 5795 649 5891 683
rect -5891 587 -5857 649
rect 5857 587 5891 649
rect -5745 547 -5729 581
rect -5695 547 -5679 581
rect -5553 547 -5537 581
rect -5503 547 -5487 581
rect -5361 547 -5345 581
rect -5311 547 -5295 581
rect -5169 547 -5153 581
rect -5119 547 -5103 581
rect -4977 547 -4961 581
rect -4927 547 -4911 581
rect -4785 547 -4769 581
rect -4735 547 -4719 581
rect -4593 547 -4577 581
rect -4543 547 -4527 581
rect -4401 547 -4385 581
rect -4351 547 -4335 581
rect -4209 547 -4193 581
rect -4159 547 -4143 581
rect -4017 547 -4001 581
rect -3967 547 -3951 581
rect -3825 547 -3809 581
rect -3775 547 -3759 581
rect -3633 547 -3617 581
rect -3583 547 -3567 581
rect -3441 547 -3425 581
rect -3391 547 -3375 581
rect -3249 547 -3233 581
rect -3199 547 -3183 581
rect -3057 547 -3041 581
rect -3007 547 -2991 581
rect -2865 547 -2849 581
rect -2815 547 -2799 581
rect -2673 547 -2657 581
rect -2623 547 -2607 581
rect -2481 547 -2465 581
rect -2431 547 -2415 581
rect -2289 547 -2273 581
rect -2239 547 -2223 581
rect -2097 547 -2081 581
rect -2047 547 -2031 581
rect -1905 547 -1889 581
rect -1855 547 -1839 581
rect -1713 547 -1697 581
rect -1663 547 -1647 581
rect -1521 547 -1505 581
rect -1471 547 -1455 581
rect -1329 547 -1313 581
rect -1279 547 -1263 581
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -945 547 -929 581
rect -895 547 -879 581
rect -753 547 -737 581
rect -703 547 -687 581
rect -561 547 -545 581
rect -511 547 -495 581
rect -369 547 -353 581
rect -319 547 -303 581
rect -177 547 -161 581
rect -127 547 -111 581
rect 15 547 31 581
rect 65 547 81 581
rect 207 547 223 581
rect 257 547 273 581
rect 399 547 415 581
rect 449 547 465 581
rect 591 547 607 581
rect 641 547 657 581
rect 783 547 799 581
rect 833 547 849 581
rect 975 547 991 581
rect 1025 547 1041 581
rect 1167 547 1183 581
rect 1217 547 1233 581
rect 1359 547 1375 581
rect 1409 547 1425 581
rect 1551 547 1567 581
rect 1601 547 1617 581
rect 1743 547 1759 581
rect 1793 547 1809 581
rect 1935 547 1951 581
rect 1985 547 2001 581
rect 2127 547 2143 581
rect 2177 547 2193 581
rect 2319 547 2335 581
rect 2369 547 2385 581
rect 2511 547 2527 581
rect 2561 547 2577 581
rect 2703 547 2719 581
rect 2753 547 2769 581
rect 2895 547 2911 581
rect 2945 547 2961 581
rect 3087 547 3103 581
rect 3137 547 3153 581
rect 3279 547 3295 581
rect 3329 547 3345 581
rect 3471 547 3487 581
rect 3521 547 3537 581
rect 3663 547 3679 581
rect 3713 547 3729 581
rect 3855 547 3871 581
rect 3905 547 3921 581
rect 4047 547 4063 581
rect 4097 547 4113 581
rect 4239 547 4255 581
rect 4289 547 4305 581
rect 4431 547 4447 581
rect 4481 547 4497 581
rect 4623 547 4639 581
rect 4673 547 4689 581
rect 4815 547 4831 581
rect 4865 547 4881 581
rect 5007 547 5023 581
rect 5057 547 5073 581
rect 5199 547 5215 581
rect 5249 547 5265 581
rect 5391 547 5407 581
rect 5441 547 5457 581
rect 5583 547 5599 581
rect 5633 547 5649 581
rect -5777 497 -5743 513
rect -5777 105 -5743 121
rect -5681 497 -5647 513
rect -5681 105 -5647 121
rect -5585 497 -5551 513
rect -5585 105 -5551 121
rect -5489 497 -5455 513
rect -5489 105 -5455 121
rect -5393 497 -5359 513
rect -5393 105 -5359 121
rect -5297 497 -5263 513
rect -5297 105 -5263 121
rect -5201 497 -5167 513
rect -5201 105 -5167 121
rect -5105 497 -5071 513
rect -5105 105 -5071 121
rect -5009 497 -4975 513
rect -5009 105 -4975 121
rect -4913 497 -4879 513
rect -4913 105 -4879 121
rect -4817 497 -4783 513
rect -4817 105 -4783 121
rect -4721 497 -4687 513
rect -4721 105 -4687 121
rect -4625 497 -4591 513
rect -4625 105 -4591 121
rect -4529 497 -4495 513
rect -4529 105 -4495 121
rect -4433 497 -4399 513
rect -4433 105 -4399 121
rect -4337 497 -4303 513
rect -4337 105 -4303 121
rect -4241 497 -4207 513
rect -4241 105 -4207 121
rect -4145 497 -4111 513
rect -4145 105 -4111 121
rect -4049 497 -4015 513
rect -4049 105 -4015 121
rect -3953 497 -3919 513
rect -3953 105 -3919 121
rect -3857 497 -3823 513
rect -3857 105 -3823 121
rect -3761 497 -3727 513
rect -3761 105 -3727 121
rect -3665 497 -3631 513
rect -3665 105 -3631 121
rect -3569 497 -3535 513
rect -3569 105 -3535 121
rect -3473 497 -3439 513
rect -3473 105 -3439 121
rect -3377 497 -3343 513
rect -3377 105 -3343 121
rect -3281 497 -3247 513
rect -3281 105 -3247 121
rect -3185 497 -3151 513
rect -3185 105 -3151 121
rect -3089 497 -3055 513
rect -3089 105 -3055 121
rect -2993 497 -2959 513
rect -2993 105 -2959 121
rect -2897 497 -2863 513
rect -2897 105 -2863 121
rect -2801 497 -2767 513
rect -2801 105 -2767 121
rect -2705 497 -2671 513
rect -2705 105 -2671 121
rect -2609 497 -2575 513
rect -2609 105 -2575 121
rect -2513 497 -2479 513
rect -2513 105 -2479 121
rect -2417 497 -2383 513
rect -2417 105 -2383 121
rect -2321 497 -2287 513
rect -2321 105 -2287 121
rect -2225 497 -2191 513
rect -2225 105 -2191 121
rect -2129 497 -2095 513
rect -2129 105 -2095 121
rect -2033 497 -1999 513
rect -2033 105 -1999 121
rect -1937 497 -1903 513
rect -1937 105 -1903 121
rect -1841 497 -1807 513
rect -1841 105 -1807 121
rect -1745 497 -1711 513
rect -1745 105 -1711 121
rect -1649 497 -1615 513
rect -1649 105 -1615 121
rect -1553 497 -1519 513
rect -1553 105 -1519 121
rect -1457 497 -1423 513
rect -1457 105 -1423 121
rect -1361 497 -1327 513
rect -1361 105 -1327 121
rect -1265 497 -1231 513
rect -1265 105 -1231 121
rect -1169 497 -1135 513
rect -1169 105 -1135 121
rect -1073 497 -1039 513
rect -1073 105 -1039 121
rect -977 497 -943 513
rect -977 105 -943 121
rect -881 497 -847 513
rect -881 105 -847 121
rect -785 497 -751 513
rect -785 105 -751 121
rect -689 497 -655 513
rect -689 105 -655 121
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect 655 497 689 513
rect 655 105 689 121
rect 751 497 785 513
rect 751 105 785 121
rect 847 497 881 513
rect 847 105 881 121
rect 943 497 977 513
rect 943 105 977 121
rect 1039 497 1073 513
rect 1039 105 1073 121
rect 1135 497 1169 513
rect 1135 105 1169 121
rect 1231 497 1265 513
rect 1231 105 1265 121
rect 1327 497 1361 513
rect 1327 105 1361 121
rect 1423 497 1457 513
rect 1423 105 1457 121
rect 1519 497 1553 513
rect 1519 105 1553 121
rect 1615 497 1649 513
rect 1615 105 1649 121
rect 1711 497 1745 513
rect 1711 105 1745 121
rect 1807 497 1841 513
rect 1807 105 1841 121
rect 1903 497 1937 513
rect 1903 105 1937 121
rect 1999 497 2033 513
rect 1999 105 2033 121
rect 2095 497 2129 513
rect 2095 105 2129 121
rect 2191 497 2225 513
rect 2191 105 2225 121
rect 2287 497 2321 513
rect 2287 105 2321 121
rect 2383 497 2417 513
rect 2383 105 2417 121
rect 2479 497 2513 513
rect 2479 105 2513 121
rect 2575 497 2609 513
rect 2575 105 2609 121
rect 2671 497 2705 513
rect 2671 105 2705 121
rect 2767 497 2801 513
rect 2767 105 2801 121
rect 2863 497 2897 513
rect 2863 105 2897 121
rect 2959 497 2993 513
rect 2959 105 2993 121
rect 3055 497 3089 513
rect 3055 105 3089 121
rect 3151 497 3185 513
rect 3151 105 3185 121
rect 3247 497 3281 513
rect 3247 105 3281 121
rect 3343 497 3377 513
rect 3343 105 3377 121
rect 3439 497 3473 513
rect 3439 105 3473 121
rect 3535 497 3569 513
rect 3535 105 3569 121
rect 3631 497 3665 513
rect 3631 105 3665 121
rect 3727 497 3761 513
rect 3727 105 3761 121
rect 3823 497 3857 513
rect 3823 105 3857 121
rect 3919 497 3953 513
rect 3919 105 3953 121
rect 4015 497 4049 513
rect 4015 105 4049 121
rect 4111 497 4145 513
rect 4111 105 4145 121
rect 4207 497 4241 513
rect 4207 105 4241 121
rect 4303 497 4337 513
rect 4303 105 4337 121
rect 4399 497 4433 513
rect 4399 105 4433 121
rect 4495 497 4529 513
rect 4495 105 4529 121
rect 4591 497 4625 513
rect 4591 105 4625 121
rect 4687 497 4721 513
rect 4687 105 4721 121
rect 4783 497 4817 513
rect 4783 105 4817 121
rect 4879 497 4913 513
rect 4879 105 4913 121
rect 4975 497 5009 513
rect 4975 105 5009 121
rect 5071 497 5105 513
rect 5071 105 5105 121
rect 5167 497 5201 513
rect 5167 105 5201 121
rect 5263 497 5297 513
rect 5263 105 5297 121
rect 5359 497 5393 513
rect 5359 105 5393 121
rect 5455 497 5489 513
rect 5455 105 5489 121
rect 5551 497 5585 513
rect 5551 105 5585 121
rect 5647 497 5681 513
rect 5647 105 5681 121
rect 5743 497 5777 513
rect 5743 105 5777 121
rect -5649 37 -5633 71
rect -5599 37 -5583 71
rect -5457 37 -5441 71
rect -5407 37 -5391 71
rect -5265 37 -5249 71
rect -5215 37 -5199 71
rect -5073 37 -5057 71
rect -5023 37 -5007 71
rect -4881 37 -4865 71
rect -4831 37 -4815 71
rect -4689 37 -4673 71
rect -4639 37 -4623 71
rect -4497 37 -4481 71
rect -4447 37 -4431 71
rect -4305 37 -4289 71
rect -4255 37 -4239 71
rect -4113 37 -4097 71
rect -4063 37 -4047 71
rect -3921 37 -3905 71
rect -3871 37 -3855 71
rect -3729 37 -3713 71
rect -3679 37 -3663 71
rect -3537 37 -3521 71
rect -3487 37 -3471 71
rect -3345 37 -3329 71
rect -3295 37 -3279 71
rect -3153 37 -3137 71
rect -3103 37 -3087 71
rect -2961 37 -2945 71
rect -2911 37 -2895 71
rect -2769 37 -2753 71
rect -2719 37 -2703 71
rect -2577 37 -2561 71
rect -2527 37 -2511 71
rect -2385 37 -2369 71
rect -2335 37 -2319 71
rect -2193 37 -2177 71
rect -2143 37 -2127 71
rect -2001 37 -1985 71
rect -1951 37 -1935 71
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1839 37 1855 71
rect 1889 37 1905 71
rect 2031 37 2047 71
rect 2081 37 2097 71
rect 2223 37 2239 71
rect 2273 37 2289 71
rect 2415 37 2431 71
rect 2465 37 2481 71
rect 2607 37 2623 71
rect 2657 37 2673 71
rect 2799 37 2815 71
rect 2849 37 2865 71
rect 2991 37 3007 71
rect 3041 37 3057 71
rect 3183 37 3199 71
rect 3233 37 3249 71
rect 3375 37 3391 71
rect 3425 37 3441 71
rect 3567 37 3583 71
rect 3617 37 3633 71
rect 3759 37 3775 71
rect 3809 37 3825 71
rect 3951 37 3967 71
rect 4001 37 4017 71
rect 4143 37 4159 71
rect 4193 37 4209 71
rect 4335 37 4351 71
rect 4385 37 4401 71
rect 4527 37 4543 71
rect 4577 37 4593 71
rect 4719 37 4735 71
rect 4769 37 4785 71
rect 4911 37 4927 71
rect 4961 37 4977 71
rect 5103 37 5119 71
rect 5153 37 5169 71
rect 5295 37 5311 71
rect 5345 37 5361 71
rect 5487 37 5503 71
rect 5537 37 5553 71
rect 5679 37 5695 71
rect 5729 37 5745 71
rect -5649 -71 -5633 -37
rect -5599 -71 -5583 -37
rect -5457 -71 -5441 -37
rect -5407 -71 -5391 -37
rect -5265 -71 -5249 -37
rect -5215 -71 -5199 -37
rect -5073 -71 -5057 -37
rect -5023 -71 -5007 -37
rect -4881 -71 -4865 -37
rect -4831 -71 -4815 -37
rect -4689 -71 -4673 -37
rect -4639 -71 -4623 -37
rect -4497 -71 -4481 -37
rect -4447 -71 -4431 -37
rect -4305 -71 -4289 -37
rect -4255 -71 -4239 -37
rect -4113 -71 -4097 -37
rect -4063 -71 -4047 -37
rect -3921 -71 -3905 -37
rect -3871 -71 -3855 -37
rect -3729 -71 -3713 -37
rect -3679 -71 -3663 -37
rect -3537 -71 -3521 -37
rect -3487 -71 -3471 -37
rect -3345 -71 -3329 -37
rect -3295 -71 -3279 -37
rect -3153 -71 -3137 -37
rect -3103 -71 -3087 -37
rect -2961 -71 -2945 -37
rect -2911 -71 -2895 -37
rect -2769 -71 -2753 -37
rect -2719 -71 -2703 -37
rect -2577 -71 -2561 -37
rect -2527 -71 -2511 -37
rect -2385 -71 -2369 -37
rect -2335 -71 -2319 -37
rect -2193 -71 -2177 -37
rect -2143 -71 -2127 -37
rect -2001 -71 -1985 -37
rect -1951 -71 -1935 -37
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect 2031 -71 2047 -37
rect 2081 -71 2097 -37
rect 2223 -71 2239 -37
rect 2273 -71 2289 -37
rect 2415 -71 2431 -37
rect 2465 -71 2481 -37
rect 2607 -71 2623 -37
rect 2657 -71 2673 -37
rect 2799 -71 2815 -37
rect 2849 -71 2865 -37
rect 2991 -71 3007 -37
rect 3041 -71 3057 -37
rect 3183 -71 3199 -37
rect 3233 -71 3249 -37
rect 3375 -71 3391 -37
rect 3425 -71 3441 -37
rect 3567 -71 3583 -37
rect 3617 -71 3633 -37
rect 3759 -71 3775 -37
rect 3809 -71 3825 -37
rect 3951 -71 3967 -37
rect 4001 -71 4017 -37
rect 4143 -71 4159 -37
rect 4193 -71 4209 -37
rect 4335 -71 4351 -37
rect 4385 -71 4401 -37
rect 4527 -71 4543 -37
rect 4577 -71 4593 -37
rect 4719 -71 4735 -37
rect 4769 -71 4785 -37
rect 4911 -71 4927 -37
rect 4961 -71 4977 -37
rect 5103 -71 5119 -37
rect 5153 -71 5169 -37
rect 5295 -71 5311 -37
rect 5345 -71 5361 -37
rect 5487 -71 5503 -37
rect 5537 -71 5553 -37
rect 5679 -71 5695 -37
rect 5729 -71 5745 -37
rect -5777 -121 -5743 -105
rect -5777 -513 -5743 -497
rect -5681 -121 -5647 -105
rect -5681 -513 -5647 -497
rect -5585 -121 -5551 -105
rect -5585 -513 -5551 -497
rect -5489 -121 -5455 -105
rect -5489 -513 -5455 -497
rect -5393 -121 -5359 -105
rect -5393 -513 -5359 -497
rect -5297 -121 -5263 -105
rect -5297 -513 -5263 -497
rect -5201 -121 -5167 -105
rect -5201 -513 -5167 -497
rect -5105 -121 -5071 -105
rect -5105 -513 -5071 -497
rect -5009 -121 -4975 -105
rect -5009 -513 -4975 -497
rect -4913 -121 -4879 -105
rect -4913 -513 -4879 -497
rect -4817 -121 -4783 -105
rect -4817 -513 -4783 -497
rect -4721 -121 -4687 -105
rect -4721 -513 -4687 -497
rect -4625 -121 -4591 -105
rect -4625 -513 -4591 -497
rect -4529 -121 -4495 -105
rect -4529 -513 -4495 -497
rect -4433 -121 -4399 -105
rect -4433 -513 -4399 -497
rect -4337 -121 -4303 -105
rect -4337 -513 -4303 -497
rect -4241 -121 -4207 -105
rect -4241 -513 -4207 -497
rect -4145 -121 -4111 -105
rect -4145 -513 -4111 -497
rect -4049 -121 -4015 -105
rect -4049 -513 -4015 -497
rect -3953 -121 -3919 -105
rect -3953 -513 -3919 -497
rect -3857 -121 -3823 -105
rect -3857 -513 -3823 -497
rect -3761 -121 -3727 -105
rect -3761 -513 -3727 -497
rect -3665 -121 -3631 -105
rect -3665 -513 -3631 -497
rect -3569 -121 -3535 -105
rect -3569 -513 -3535 -497
rect -3473 -121 -3439 -105
rect -3473 -513 -3439 -497
rect -3377 -121 -3343 -105
rect -3377 -513 -3343 -497
rect -3281 -121 -3247 -105
rect -3281 -513 -3247 -497
rect -3185 -121 -3151 -105
rect -3185 -513 -3151 -497
rect -3089 -121 -3055 -105
rect -3089 -513 -3055 -497
rect -2993 -121 -2959 -105
rect -2993 -513 -2959 -497
rect -2897 -121 -2863 -105
rect -2897 -513 -2863 -497
rect -2801 -121 -2767 -105
rect -2801 -513 -2767 -497
rect -2705 -121 -2671 -105
rect -2705 -513 -2671 -497
rect -2609 -121 -2575 -105
rect -2609 -513 -2575 -497
rect -2513 -121 -2479 -105
rect -2513 -513 -2479 -497
rect -2417 -121 -2383 -105
rect -2417 -513 -2383 -497
rect -2321 -121 -2287 -105
rect -2321 -513 -2287 -497
rect -2225 -121 -2191 -105
rect -2225 -513 -2191 -497
rect -2129 -121 -2095 -105
rect -2129 -513 -2095 -497
rect -2033 -121 -1999 -105
rect -2033 -513 -1999 -497
rect -1937 -121 -1903 -105
rect -1937 -513 -1903 -497
rect -1841 -121 -1807 -105
rect -1841 -513 -1807 -497
rect -1745 -121 -1711 -105
rect -1745 -513 -1711 -497
rect -1649 -121 -1615 -105
rect -1649 -513 -1615 -497
rect -1553 -121 -1519 -105
rect -1553 -513 -1519 -497
rect -1457 -121 -1423 -105
rect -1457 -513 -1423 -497
rect -1361 -121 -1327 -105
rect -1361 -513 -1327 -497
rect -1265 -121 -1231 -105
rect -1265 -513 -1231 -497
rect -1169 -121 -1135 -105
rect -1169 -513 -1135 -497
rect -1073 -121 -1039 -105
rect -1073 -513 -1039 -497
rect -977 -121 -943 -105
rect -977 -513 -943 -497
rect -881 -121 -847 -105
rect -881 -513 -847 -497
rect -785 -121 -751 -105
rect -785 -513 -751 -497
rect -689 -121 -655 -105
rect -689 -513 -655 -497
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect 655 -121 689 -105
rect 655 -513 689 -497
rect 751 -121 785 -105
rect 751 -513 785 -497
rect 847 -121 881 -105
rect 847 -513 881 -497
rect 943 -121 977 -105
rect 943 -513 977 -497
rect 1039 -121 1073 -105
rect 1039 -513 1073 -497
rect 1135 -121 1169 -105
rect 1135 -513 1169 -497
rect 1231 -121 1265 -105
rect 1231 -513 1265 -497
rect 1327 -121 1361 -105
rect 1327 -513 1361 -497
rect 1423 -121 1457 -105
rect 1423 -513 1457 -497
rect 1519 -121 1553 -105
rect 1519 -513 1553 -497
rect 1615 -121 1649 -105
rect 1615 -513 1649 -497
rect 1711 -121 1745 -105
rect 1711 -513 1745 -497
rect 1807 -121 1841 -105
rect 1807 -513 1841 -497
rect 1903 -121 1937 -105
rect 1903 -513 1937 -497
rect 1999 -121 2033 -105
rect 1999 -513 2033 -497
rect 2095 -121 2129 -105
rect 2095 -513 2129 -497
rect 2191 -121 2225 -105
rect 2191 -513 2225 -497
rect 2287 -121 2321 -105
rect 2287 -513 2321 -497
rect 2383 -121 2417 -105
rect 2383 -513 2417 -497
rect 2479 -121 2513 -105
rect 2479 -513 2513 -497
rect 2575 -121 2609 -105
rect 2575 -513 2609 -497
rect 2671 -121 2705 -105
rect 2671 -513 2705 -497
rect 2767 -121 2801 -105
rect 2767 -513 2801 -497
rect 2863 -121 2897 -105
rect 2863 -513 2897 -497
rect 2959 -121 2993 -105
rect 2959 -513 2993 -497
rect 3055 -121 3089 -105
rect 3055 -513 3089 -497
rect 3151 -121 3185 -105
rect 3151 -513 3185 -497
rect 3247 -121 3281 -105
rect 3247 -513 3281 -497
rect 3343 -121 3377 -105
rect 3343 -513 3377 -497
rect 3439 -121 3473 -105
rect 3439 -513 3473 -497
rect 3535 -121 3569 -105
rect 3535 -513 3569 -497
rect 3631 -121 3665 -105
rect 3631 -513 3665 -497
rect 3727 -121 3761 -105
rect 3727 -513 3761 -497
rect 3823 -121 3857 -105
rect 3823 -513 3857 -497
rect 3919 -121 3953 -105
rect 3919 -513 3953 -497
rect 4015 -121 4049 -105
rect 4015 -513 4049 -497
rect 4111 -121 4145 -105
rect 4111 -513 4145 -497
rect 4207 -121 4241 -105
rect 4207 -513 4241 -497
rect 4303 -121 4337 -105
rect 4303 -513 4337 -497
rect 4399 -121 4433 -105
rect 4399 -513 4433 -497
rect 4495 -121 4529 -105
rect 4495 -513 4529 -497
rect 4591 -121 4625 -105
rect 4591 -513 4625 -497
rect 4687 -121 4721 -105
rect 4687 -513 4721 -497
rect 4783 -121 4817 -105
rect 4783 -513 4817 -497
rect 4879 -121 4913 -105
rect 4879 -513 4913 -497
rect 4975 -121 5009 -105
rect 4975 -513 5009 -497
rect 5071 -121 5105 -105
rect 5071 -513 5105 -497
rect 5167 -121 5201 -105
rect 5167 -513 5201 -497
rect 5263 -121 5297 -105
rect 5263 -513 5297 -497
rect 5359 -121 5393 -105
rect 5359 -513 5393 -497
rect 5455 -121 5489 -105
rect 5455 -513 5489 -497
rect 5551 -121 5585 -105
rect 5551 -513 5585 -497
rect 5647 -121 5681 -105
rect 5647 -513 5681 -497
rect 5743 -121 5777 -105
rect 5743 -513 5777 -497
rect -5745 -581 -5729 -547
rect -5695 -581 -5679 -547
rect -5553 -581 -5537 -547
rect -5503 -581 -5487 -547
rect -5361 -581 -5345 -547
rect -5311 -581 -5295 -547
rect -5169 -581 -5153 -547
rect -5119 -581 -5103 -547
rect -4977 -581 -4961 -547
rect -4927 -581 -4911 -547
rect -4785 -581 -4769 -547
rect -4735 -581 -4719 -547
rect -4593 -581 -4577 -547
rect -4543 -581 -4527 -547
rect -4401 -581 -4385 -547
rect -4351 -581 -4335 -547
rect -4209 -581 -4193 -547
rect -4159 -581 -4143 -547
rect -4017 -581 -4001 -547
rect -3967 -581 -3951 -547
rect -3825 -581 -3809 -547
rect -3775 -581 -3759 -547
rect -3633 -581 -3617 -547
rect -3583 -581 -3567 -547
rect -3441 -581 -3425 -547
rect -3391 -581 -3375 -547
rect -3249 -581 -3233 -547
rect -3199 -581 -3183 -547
rect -3057 -581 -3041 -547
rect -3007 -581 -2991 -547
rect -2865 -581 -2849 -547
rect -2815 -581 -2799 -547
rect -2673 -581 -2657 -547
rect -2623 -581 -2607 -547
rect -2481 -581 -2465 -547
rect -2431 -581 -2415 -547
rect -2289 -581 -2273 -547
rect -2239 -581 -2223 -547
rect -2097 -581 -2081 -547
rect -2047 -581 -2031 -547
rect -1905 -581 -1889 -547
rect -1855 -581 -1839 -547
rect -1713 -581 -1697 -547
rect -1663 -581 -1647 -547
rect -1521 -581 -1505 -547
rect -1471 -581 -1455 -547
rect -1329 -581 -1313 -547
rect -1279 -581 -1263 -547
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 1167 -581 1183 -547
rect 1217 -581 1233 -547
rect 1359 -581 1375 -547
rect 1409 -581 1425 -547
rect 1551 -581 1567 -547
rect 1601 -581 1617 -547
rect 1743 -581 1759 -547
rect 1793 -581 1809 -547
rect 1935 -581 1951 -547
rect 1985 -581 2001 -547
rect 2127 -581 2143 -547
rect 2177 -581 2193 -547
rect 2319 -581 2335 -547
rect 2369 -581 2385 -547
rect 2511 -581 2527 -547
rect 2561 -581 2577 -547
rect 2703 -581 2719 -547
rect 2753 -581 2769 -547
rect 2895 -581 2911 -547
rect 2945 -581 2961 -547
rect 3087 -581 3103 -547
rect 3137 -581 3153 -547
rect 3279 -581 3295 -547
rect 3329 -581 3345 -547
rect 3471 -581 3487 -547
rect 3521 -581 3537 -547
rect 3663 -581 3679 -547
rect 3713 -581 3729 -547
rect 3855 -581 3871 -547
rect 3905 -581 3921 -547
rect 4047 -581 4063 -547
rect 4097 -581 4113 -547
rect 4239 -581 4255 -547
rect 4289 -581 4305 -547
rect 4431 -581 4447 -547
rect 4481 -581 4497 -547
rect 4623 -581 4639 -547
rect 4673 -581 4689 -547
rect 4815 -581 4831 -547
rect 4865 -581 4881 -547
rect 5007 -581 5023 -547
rect 5057 -581 5073 -547
rect 5199 -581 5215 -547
rect 5249 -581 5265 -547
rect 5391 -581 5407 -547
rect 5441 -581 5457 -547
rect 5583 -581 5599 -547
rect 5633 -581 5649 -547
rect -5891 -649 -5857 -587
rect 5857 -649 5891 -587
rect -5891 -683 -5795 -649
rect 5795 -683 5891 -649
<< viali >>
rect -5729 547 -5695 581
rect -5537 547 -5503 581
rect -5345 547 -5311 581
rect -5153 547 -5119 581
rect -4961 547 -4927 581
rect -4769 547 -4735 581
rect -4577 547 -4543 581
rect -4385 547 -4351 581
rect -4193 547 -4159 581
rect -4001 547 -3967 581
rect -3809 547 -3775 581
rect -3617 547 -3583 581
rect -3425 547 -3391 581
rect -3233 547 -3199 581
rect -3041 547 -3007 581
rect -2849 547 -2815 581
rect -2657 547 -2623 581
rect -2465 547 -2431 581
rect -2273 547 -2239 581
rect -2081 547 -2047 581
rect -1889 547 -1855 581
rect -1697 547 -1663 581
rect -1505 547 -1471 581
rect -1313 547 -1279 581
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect 1183 547 1217 581
rect 1375 547 1409 581
rect 1567 547 1601 581
rect 1759 547 1793 581
rect 1951 547 1985 581
rect 2143 547 2177 581
rect 2335 547 2369 581
rect 2527 547 2561 581
rect 2719 547 2753 581
rect 2911 547 2945 581
rect 3103 547 3137 581
rect 3295 547 3329 581
rect 3487 547 3521 581
rect 3679 547 3713 581
rect 3871 547 3905 581
rect 4063 547 4097 581
rect 4255 547 4289 581
rect 4447 547 4481 581
rect 4639 547 4673 581
rect 4831 547 4865 581
rect 5023 547 5057 581
rect 5215 547 5249 581
rect 5407 547 5441 581
rect 5599 547 5633 581
rect -5777 121 -5743 497
rect -5681 121 -5647 497
rect -5585 121 -5551 497
rect -5489 121 -5455 497
rect -5393 121 -5359 497
rect -5297 121 -5263 497
rect -5201 121 -5167 497
rect -5105 121 -5071 497
rect -5009 121 -4975 497
rect -4913 121 -4879 497
rect -4817 121 -4783 497
rect -4721 121 -4687 497
rect -4625 121 -4591 497
rect -4529 121 -4495 497
rect -4433 121 -4399 497
rect -4337 121 -4303 497
rect -4241 121 -4207 497
rect -4145 121 -4111 497
rect -4049 121 -4015 497
rect -3953 121 -3919 497
rect -3857 121 -3823 497
rect -3761 121 -3727 497
rect -3665 121 -3631 497
rect -3569 121 -3535 497
rect -3473 121 -3439 497
rect -3377 121 -3343 497
rect -3281 121 -3247 497
rect -3185 121 -3151 497
rect -3089 121 -3055 497
rect -2993 121 -2959 497
rect -2897 121 -2863 497
rect -2801 121 -2767 497
rect -2705 121 -2671 497
rect -2609 121 -2575 497
rect -2513 121 -2479 497
rect -2417 121 -2383 497
rect -2321 121 -2287 497
rect -2225 121 -2191 497
rect -2129 121 -2095 497
rect -2033 121 -1999 497
rect -1937 121 -1903 497
rect -1841 121 -1807 497
rect -1745 121 -1711 497
rect -1649 121 -1615 497
rect -1553 121 -1519 497
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect 1519 121 1553 497
rect 1615 121 1649 497
rect 1711 121 1745 497
rect 1807 121 1841 497
rect 1903 121 1937 497
rect 1999 121 2033 497
rect 2095 121 2129 497
rect 2191 121 2225 497
rect 2287 121 2321 497
rect 2383 121 2417 497
rect 2479 121 2513 497
rect 2575 121 2609 497
rect 2671 121 2705 497
rect 2767 121 2801 497
rect 2863 121 2897 497
rect 2959 121 2993 497
rect 3055 121 3089 497
rect 3151 121 3185 497
rect 3247 121 3281 497
rect 3343 121 3377 497
rect 3439 121 3473 497
rect 3535 121 3569 497
rect 3631 121 3665 497
rect 3727 121 3761 497
rect 3823 121 3857 497
rect 3919 121 3953 497
rect 4015 121 4049 497
rect 4111 121 4145 497
rect 4207 121 4241 497
rect 4303 121 4337 497
rect 4399 121 4433 497
rect 4495 121 4529 497
rect 4591 121 4625 497
rect 4687 121 4721 497
rect 4783 121 4817 497
rect 4879 121 4913 497
rect 4975 121 5009 497
rect 5071 121 5105 497
rect 5167 121 5201 497
rect 5263 121 5297 497
rect 5359 121 5393 497
rect 5455 121 5489 497
rect 5551 121 5585 497
rect 5647 121 5681 497
rect 5743 121 5777 497
rect -5633 37 -5599 71
rect -5441 37 -5407 71
rect -5249 37 -5215 71
rect -5057 37 -5023 71
rect -4865 37 -4831 71
rect -4673 37 -4639 71
rect -4481 37 -4447 71
rect -4289 37 -4255 71
rect -4097 37 -4063 71
rect -3905 37 -3871 71
rect -3713 37 -3679 71
rect -3521 37 -3487 71
rect -3329 37 -3295 71
rect -3137 37 -3103 71
rect -2945 37 -2911 71
rect -2753 37 -2719 71
rect -2561 37 -2527 71
rect -2369 37 -2335 71
rect -2177 37 -2143 71
rect -1985 37 -1951 71
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect 2047 37 2081 71
rect 2239 37 2273 71
rect 2431 37 2465 71
rect 2623 37 2657 71
rect 2815 37 2849 71
rect 3007 37 3041 71
rect 3199 37 3233 71
rect 3391 37 3425 71
rect 3583 37 3617 71
rect 3775 37 3809 71
rect 3967 37 4001 71
rect 4159 37 4193 71
rect 4351 37 4385 71
rect 4543 37 4577 71
rect 4735 37 4769 71
rect 4927 37 4961 71
rect 5119 37 5153 71
rect 5311 37 5345 71
rect 5503 37 5537 71
rect 5695 37 5729 71
rect -5633 -71 -5599 -37
rect -5441 -71 -5407 -37
rect -5249 -71 -5215 -37
rect -5057 -71 -5023 -37
rect -4865 -71 -4831 -37
rect -4673 -71 -4639 -37
rect -4481 -71 -4447 -37
rect -4289 -71 -4255 -37
rect -4097 -71 -4063 -37
rect -3905 -71 -3871 -37
rect -3713 -71 -3679 -37
rect -3521 -71 -3487 -37
rect -3329 -71 -3295 -37
rect -3137 -71 -3103 -37
rect -2945 -71 -2911 -37
rect -2753 -71 -2719 -37
rect -2561 -71 -2527 -37
rect -2369 -71 -2335 -37
rect -2177 -71 -2143 -37
rect -1985 -71 -1951 -37
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect 2047 -71 2081 -37
rect 2239 -71 2273 -37
rect 2431 -71 2465 -37
rect 2623 -71 2657 -37
rect 2815 -71 2849 -37
rect 3007 -71 3041 -37
rect 3199 -71 3233 -37
rect 3391 -71 3425 -37
rect 3583 -71 3617 -37
rect 3775 -71 3809 -37
rect 3967 -71 4001 -37
rect 4159 -71 4193 -37
rect 4351 -71 4385 -37
rect 4543 -71 4577 -37
rect 4735 -71 4769 -37
rect 4927 -71 4961 -37
rect 5119 -71 5153 -37
rect 5311 -71 5345 -37
rect 5503 -71 5537 -37
rect 5695 -71 5729 -37
rect -5777 -497 -5743 -121
rect -5681 -497 -5647 -121
rect -5585 -497 -5551 -121
rect -5489 -497 -5455 -121
rect -5393 -497 -5359 -121
rect -5297 -497 -5263 -121
rect -5201 -497 -5167 -121
rect -5105 -497 -5071 -121
rect -5009 -497 -4975 -121
rect -4913 -497 -4879 -121
rect -4817 -497 -4783 -121
rect -4721 -497 -4687 -121
rect -4625 -497 -4591 -121
rect -4529 -497 -4495 -121
rect -4433 -497 -4399 -121
rect -4337 -497 -4303 -121
rect -4241 -497 -4207 -121
rect -4145 -497 -4111 -121
rect -4049 -497 -4015 -121
rect -3953 -497 -3919 -121
rect -3857 -497 -3823 -121
rect -3761 -497 -3727 -121
rect -3665 -497 -3631 -121
rect -3569 -497 -3535 -121
rect -3473 -497 -3439 -121
rect -3377 -497 -3343 -121
rect -3281 -497 -3247 -121
rect -3185 -497 -3151 -121
rect -3089 -497 -3055 -121
rect -2993 -497 -2959 -121
rect -2897 -497 -2863 -121
rect -2801 -497 -2767 -121
rect -2705 -497 -2671 -121
rect -2609 -497 -2575 -121
rect -2513 -497 -2479 -121
rect -2417 -497 -2383 -121
rect -2321 -497 -2287 -121
rect -2225 -497 -2191 -121
rect -2129 -497 -2095 -121
rect -2033 -497 -1999 -121
rect -1937 -497 -1903 -121
rect -1841 -497 -1807 -121
rect -1745 -497 -1711 -121
rect -1649 -497 -1615 -121
rect -1553 -497 -1519 -121
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect 1519 -497 1553 -121
rect 1615 -497 1649 -121
rect 1711 -497 1745 -121
rect 1807 -497 1841 -121
rect 1903 -497 1937 -121
rect 1999 -497 2033 -121
rect 2095 -497 2129 -121
rect 2191 -497 2225 -121
rect 2287 -497 2321 -121
rect 2383 -497 2417 -121
rect 2479 -497 2513 -121
rect 2575 -497 2609 -121
rect 2671 -497 2705 -121
rect 2767 -497 2801 -121
rect 2863 -497 2897 -121
rect 2959 -497 2993 -121
rect 3055 -497 3089 -121
rect 3151 -497 3185 -121
rect 3247 -497 3281 -121
rect 3343 -497 3377 -121
rect 3439 -497 3473 -121
rect 3535 -497 3569 -121
rect 3631 -497 3665 -121
rect 3727 -497 3761 -121
rect 3823 -497 3857 -121
rect 3919 -497 3953 -121
rect 4015 -497 4049 -121
rect 4111 -497 4145 -121
rect 4207 -497 4241 -121
rect 4303 -497 4337 -121
rect 4399 -497 4433 -121
rect 4495 -497 4529 -121
rect 4591 -497 4625 -121
rect 4687 -497 4721 -121
rect 4783 -497 4817 -121
rect 4879 -497 4913 -121
rect 4975 -497 5009 -121
rect 5071 -497 5105 -121
rect 5167 -497 5201 -121
rect 5263 -497 5297 -121
rect 5359 -497 5393 -121
rect 5455 -497 5489 -121
rect 5551 -497 5585 -121
rect 5647 -497 5681 -121
rect 5743 -497 5777 -121
rect -5729 -581 -5695 -547
rect -5537 -581 -5503 -547
rect -5345 -581 -5311 -547
rect -5153 -581 -5119 -547
rect -4961 -581 -4927 -547
rect -4769 -581 -4735 -547
rect -4577 -581 -4543 -547
rect -4385 -581 -4351 -547
rect -4193 -581 -4159 -547
rect -4001 -581 -3967 -547
rect -3809 -581 -3775 -547
rect -3617 -581 -3583 -547
rect -3425 -581 -3391 -547
rect -3233 -581 -3199 -547
rect -3041 -581 -3007 -547
rect -2849 -581 -2815 -547
rect -2657 -581 -2623 -547
rect -2465 -581 -2431 -547
rect -2273 -581 -2239 -547
rect -2081 -581 -2047 -547
rect -1889 -581 -1855 -547
rect -1697 -581 -1663 -547
rect -1505 -581 -1471 -547
rect -1313 -581 -1279 -547
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect 1183 -581 1217 -547
rect 1375 -581 1409 -547
rect 1567 -581 1601 -547
rect 1759 -581 1793 -547
rect 1951 -581 1985 -547
rect 2143 -581 2177 -547
rect 2335 -581 2369 -547
rect 2527 -581 2561 -547
rect 2719 -581 2753 -547
rect 2911 -581 2945 -547
rect 3103 -581 3137 -547
rect 3295 -581 3329 -547
rect 3487 -581 3521 -547
rect 3679 -581 3713 -547
rect 3871 -581 3905 -547
rect 4063 -581 4097 -547
rect 4255 -581 4289 -547
rect 4447 -581 4481 -547
rect 4639 -581 4673 -547
rect 4831 -581 4865 -547
rect 5023 -581 5057 -547
rect 5215 -581 5249 -547
rect 5407 -581 5441 -547
rect 5599 -581 5633 -547
<< metal1 >>
rect -5741 581 -5683 587
rect -5741 547 -5729 581
rect -5695 547 -5683 581
rect -5741 541 -5683 547
rect -5549 581 -5491 587
rect -5549 547 -5537 581
rect -5503 547 -5491 581
rect -5549 541 -5491 547
rect -5357 581 -5299 587
rect -5357 547 -5345 581
rect -5311 547 -5299 581
rect -5357 541 -5299 547
rect -5165 581 -5107 587
rect -5165 547 -5153 581
rect -5119 547 -5107 581
rect -5165 541 -5107 547
rect -4973 581 -4915 587
rect -4973 547 -4961 581
rect -4927 547 -4915 581
rect -4973 541 -4915 547
rect -4781 581 -4723 587
rect -4781 547 -4769 581
rect -4735 547 -4723 581
rect -4781 541 -4723 547
rect -4589 581 -4531 587
rect -4589 547 -4577 581
rect -4543 547 -4531 581
rect -4589 541 -4531 547
rect -4397 581 -4339 587
rect -4397 547 -4385 581
rect -4351 547 -4339 581
rect -4397 541 -4339 547
rect -4205 581 -4147 587
rect -4205 547 -4193 581
rect -4159 547 -4147 581
rect -4205 541 -4147 547
rect -4013 581 -3955 587
rect -4013 547 -4001 581
rect -3967 547 -3955 581
rect -4013 541 -3955 547
rect -3821 581 -3763 587
rect -3821 547 -3809 581
rect -3775 547 -3763 581
rect -3821 541 -3763 547
rect -3629 581 -3571 587
rect -3629 547 -3617 581
rect -3583 547 -3571 581
rect -3629 541 -3571 547
rect -3437 581 -3379 587
rect -3437 547 -3425 581
rect -3391 547 -3379 581
rect -3437 541 -3379 547
rect -3245 581 -3187 587
rect -3245 547 -3233 581
rect -3199 547 -3187 581
rect -3245 541 -3187 547
rect -3053 581 -2995 587
rect -3053 547 -3041 581
rect -3007 547 -2995 581
rect -3053 541 -2995 547
rect -2861 581 -2803 587
rect -2861 547 -2849 581
rect -2815 547 -2803 581
rect -2861 541 -2803 547
rect -2669 581 -2611 587
rect -2669 547 -2657 581
rect -2623 547 -2611 581
rect -2669 541 -2611 547
rect -2477 581 -2419 587
rect -2477 547 -2465 581
rect -2431 547 -2419 581
rect -2477 541 -2419 547
rect -2285 581 -2227 587
rect -2285 547 -2273 581
rect -2239 547 -2227 581
rect -2285 541 -2227 547
rect -2093 581 -2035 587
rect -2093 547 -2081 581
rect -2047 547 -2035 581
rect -2093 541 -2035 547
rect -1901 581 -1843 587
rect -1901 547 -1889 581
rect -1855 547 -1843 581
rect -1901 541 -1843 547
rect -1709 581 -1651 587
rect -1709 547 -1697 581
rect -1663 547 -1651 581
rect -1709 541 -1651 547
rect -1517 581 -1459 587
rect -1517 547 -1505 581
rect -1471 547 -1459 581
rect -1517 541 -1459 547
rect -1325 581 -1267 587
rect -1325 547 -1313 581
rect -1279 547 -1267 581
rect -1325 541 -1267 547
rect -1133 581 -1075 587
rect -1133 547 -1121 581
rect -1087 547 -1075 581
rect -1133 541 -1075 547
rect -941 581 -883 587
rect -941 547 -929 581
rect -895 547 -883 581
rect -941 541 -883 547
rect -749 581 -691 587
rect -749 547 -737 581
rect -703 547 -691 581
rect -749 541 -691 547
rect -557 581 -499 587
rect -557 547 -545 581
rect -511 547 -499 581
rect -557 541 -499 547
rect -365 581 -307 587
rect -365 547 -353 581
rect -319 547 -307 581
rect -365 541 -307 547
rect -173 581 -115 587
rect -173 547 -161 581
rect -127 547 -115 581
rect -173 541 -115 547
rect 19 581 77 587
rect 19 547 31 581
rect 65 547 77 581
rect 19 541 77 547
rect 211 581 269 587
rect 211 547 223 581
rect 257 547 269 581
rect 211 541 269 547
rect 403 581 461 587
rect 403 547 415 581
rect 449 547 461 581
rect 403 541 461 547
rect 595 581 653 587
rect 595 547 607 581
rect 641 547 653 581
rect 595 541 653 547
rect 787 581 845 587
rect 787 547 799 581
rect 833 547 845 581
rect 787 541 845 547
rect 979 581 1037 587
rect 979 547 991 581
rect 1025 547 1037 581
rect 979 541 1037 547
rect 1171 581 1229 587
rect 1171 547 1183 581
rect 1217 547 1229 581
rect 1171 541 1229 547
rect 1363 581 1421 587
rect 1363 547 1375 581
rect 1409 547 1421 581
rect 1363 541 1421 547
rect 1555 581 1613 587
rect 1555 547 1567 581
rect 1601 547 1613 581
rect 1555 541 1613 547
rect 1747 581 1805 587
rect 1747 547 1759 581
rect 1793 547 1805 581
rect 1747 541 1805 547
rect 1939 581 1997 587
rect 1939 547 1951 581
rect 1985 547 1997 581
rect 1939 541 1997 547
rect 2131 581 2189 587
rect 2131 547 2143 581
rect 2177 547 2189 581
rect 2131 541 2189 547
rect 2323 581 2381 587
rect 2323 547 2335 581
rect 2369 547 2381 581
rect 2323 541 2381 547
rect 2515 581 2573 587
rect 2515 547 2527 581
rect 2561 547 2573 581
rect 2515 541 2573 547
rect 2707 581 2765 587
rect 2707 547 2719 581
rect 2753 547 2765 581
rect 2707 541 2765 547
rect 2899 581 2957 587
rect 2899 547 2911 581
rect 2945 547 2957 581
rect 2899 541 2957 547
rect 3091 581 3149 587
rect 3091 547 3103 581
rect 3137 547 3149 581
rect 3091 541 3149 547
rect 3283 581 3341 587
rect 3283 547 3295 581
rect 3329 547 3341 581
rect 3283 541 3341 547
rect 3475 581 3533 587
rect 3475 547 3487 581
rect 3521 547 3533 581
rect 3475 541 3533 547
rect 3667 581 3725 587
rect 3667 547 3679 581
rect 3713 547 3725 581
rect 3667 541 3725 547
rect 3859 581 3917 587
rect 3859 547 3871 581
rect 3905 547 3917 581
rect 3859 541 3917 547
rect 4051 581 4109 587
rect 4051 547 4063 581
rect 4097 547 4109 581
rect 4051 541 4109 547
rect 4243 581 4301 587
rect 4243 547 4255 581
rect 4289 547 4301 581
rect 4243 541 4301 547
rect 4435 581 4493 587
rect 4435 547 4447 581
rect 4481 547 4493 581
rect 4435 541 4493 547
rect 4627 581 4685 587
rect 4627 547 4639 581
rect 4673 547 4685 581
rect 4627 541 4685 547
rect 4819 581 4877 587
rect 4819 547 4831 581
rect 4865 547 4877 581
rect 4819 541 4877 547
rect 5011 581 5069 587
rect 5011 547 5023 581
rect 5057 547 5069 581
rect 5011 541 5069 547
rect 5203 581 5261 587
rect 5203 547 5215 581
rect 5249 547 5261 581
rect 5203 541 5261 547
rect 5395 581 5453 587
rect 5395 547 5407 581
rect 5441 547 5453 581
rect 5395 541 5453 547
rect 5587 581 5645 587
rect 5587 547 5599 581
rect 5633 547 5645 581
rect 5587 541 5645 547
rect -5783 497 -5737 509
rect -5783 121 -5777 497
rect -5743 121 -5737 497
rect -5783 109 -5737 121
rect -5687 497 -5641 509
rect -5687 121 -5681 497
rect -5647 121 -5641 497
rect -5687 109 -5641 121
rect -5591 497 -5545 509
rect -5591 121 -5585 497
rect -5551 121 -5545 497
rect -5591 109 -5545 121
rect -5495 497 -5449 509
rect -5495 121 -5489 497
rect -5455 121 -5449 497
rect -5495 109 -5449 121
rect -5399 497 -5353 509
rect -5399 121 -5393 497
rect -5359 121 -5353 497
rect -5399 109 -5353 121
rect -5303 497 -5257 509
rect -5303 121 -5297 497
rect -5263 121 -5257 497
rect -5303 109 -5257 121
rect -5207 497 -5161 509
rect -5207 121 -5201 497
rect -5167 121 -5161 497
rect -5207 109 -5161 121
rect -5111 497 -5065 509
rect -5111 121 -5105 497
rect -5071 121 -5065 497
rect -5111 109 -5065 121
rect -5015 497 -4969 509
rect -5015 121 -5009 497
rect -4975 121 -4969 497
rect -5015 109 -4969 121
rect -4919 497 -4873 509
rect -4919 121 -4913 497
rect -4879 121 -4873 497
rect -4919 109 -4873 121
rect -4823 497 -4777 509
rect -4823 121 -4817 497
rect -4783 121 -4777 497
rect -4823 109 -4777 121
rect -4727 497 -4681 509
rect -4727 121 -4721 497
rect -4687 121 -4681 497
rect -4727 109 -4681 121
rect -4631 497 -4585 509
rect -4631 121 -4625 497
rect -4591 121 -4585 497
rect -4631 109 -4585 121
rect -4535 497 -4489 509
rect -4535 121 -4529 497
rect -4495 121 -4489 497
rect -4535 109 -4489 121
rect -4439 497 -4393 509
rect -4439 121 -4433 497
rect -4399 121 -4393 497
rect -4439 109 -4393 121
rect -4343 497 -4297 509
rect -4343 121 -4337 497
rect -4303 121 -4297 497
rect -4343 109 -4297 121
rect -4247 497 -4201 509
rect -4247 121 -4241 497
rect -4207 121 -4201 497
rect -4247 109 -4201 121
rect -4151 497 -4105 509
rect -4151 121 -4145 497
rect -4111 121 -4105 497
rect -4151 109 -4105 121
rect -4055 497 -4009 509
rect -4055 121 -4049 497
rect -4015 121 -4009 497
rect -4055 109 -4009 121
rect -3959 497 -3913 509
rect -3959 121 -3953 497
rect -3919 121 -3913 497
rect -3959 109 -3913 121
rect -3863 497 -3817 509
rect -3863 121 -3857 497
rect -3823 121 -3817 497
rect -3863 109 -3817 121
rect -3767 497 -3721 509
rect -3767 121 -3761 497
rect -3727 121 -3721 497
rect -3767 109 -3721 121
rect -3671 497 -3625 509
rect -3671 121 -3665 497
rect -3631 121 -3625 497
rect -3671 109 -3625 121
rect -3575 497 -3529 509
rect -3575 121 -3569 497
rect -3535 121 -3529 497
rect -3575 109 -3529 121
rect -3479 497 -3433 509
rect -3479 121 -3473 497
rect -3439 121 -3433 497
rect -3479 109 -3433 121
rect -3383 497 -3337 509
rect -3383 121 -3377 497
rect -3343 121 -3337 497
rect -3383 109 -3337 121
rect -3287 497 -3241 509
rect -3287 121 -3281 497
rect -3247 121 -3241 497
rect -3287 109 -3241 121
rect -3191 497 -3145 509
rect -3191 121 -3185 497
rect -3151 121 -3145 497
rect -3191 109 -3145 121
rect -3095 497 -3049 509
rect -3095 121 -3089 497
rect -3055 121 -3049 497
rect -3095 109 -3049 121
rect -2999 497 -2953 509
rect -2999 121 -2993 497
rect -2959 121 -2953 497
rect -2999 109 -2953 121
rect -2903 497 -2857 509
rect -2903 121 -2897 497
rect -2863 121 -2857 497
rect -2903 109 -2857 121
rect -2807 497 -2761 509
rect -2807 121 -2801 497
rect -2767 121 -2761 497
rect -2807 109 -2761 121
rect -2711 497 -2665 509
rect -2711 121 -2705 497
rect -2671 121 -2665 497
rect -2711 109 -2665 121
rect -2615 497 -2569 509
rect -2615 121 -2609 497
rect -2575 121 -2569 497
rect -2615 109 -2569 121
rect -2519 497 -2473 509
rect -2519 121 -2513 497
rect -2479 121 -2473 497
rect -2519 109 -2473 121
rect -2423 497 -2377 509
rect -2423 121 -2417 497
rect -2383 121 -2377 497
rect -2423 109 -2377 121
rect -2327 497 -2281 509
rect -2327 121 -2321 497
rect -2287 121 -2281 497
rect -2327 109 -2281 121
rect -2231 497 -2185 509
rect -2231 121 -2225 497
rect -2191 121 -2185 497
rect -2231 109 -2185 121
rect -2135 497 -2089 509
rect -2135 121 -2129 497
rect -2095 121 -2089 497
rect -2135 109 -2089 121
rect -2039 497 -1993 509
rect -2039 121 -2033 497
rect -1999 121 -1993 497
rect -2039 109 -1993 121
rect -1943 497 -1897 509
rect -1943 121 -1937 497
rect -1903 121 -1897 497
rect -1943 109 -1897 121
rect -1847 497 -1801 509
rect -1847 121 -1841 497
rect -1807 121 -1801 497
rect -1847 109 -1801 121
rect -1751 497 -1705 509
rect -1751 121 -1745 497
rect -1711 121 -1705 497
rect -1751 109 -1705 121
rect -1655 497 -1609 509
rect -1655 121 -1649 497
rect -1615 121 -1609 497
rect -1655 109 -1609 121
rect -1559 497 -1513 509
rect -1559 121 -1553 497
rect -1519 121 -1513 497
rect -1559 109 -1513 121
rect -1463 497 -1417 509
rect -1463 121 -1457 497
rect -1423 121 -1417 497
rect -1463 109 -1417 121
rect -1367 497 -1321 509
rect -1367 121 -1361 497
rect -1327 121 -1321 497
rect -1367 109 -1321 121
rect -1271 497 -1225 509
rect -1271 121 -1265 497
rect -1231 121 -1225 497
rect -1271 109 -1225 121
rect -1175 497 -1129 509
rect -1175 121 -1169 497
rect -1135 121 -1129 497
rect -1175 109 -1129 121
rect -1079 497 -1033 509
rect -1079 121 -1073 497
rect -1039 121 -1033 497
rect -1079 109 -1033 121
rect -983 497 -937 509
rect -983 121 -977 497
rect -943 121 -937 497
rect -983 109 -937 121
rect -887 497 -841 509
rect -887 121 -881 497
rect -847 121 -841 497
rect -887 109 -841 121
rect -791 497 -745 509
rect -791 121 -785 497
rect -751 121 -745 497
rect -791 109 -745 121
rect -695 497 -649 509
rect -695 121 -689 497
rect -655 121 -649 497
rect -695 109 -649 121
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect 649 497 695 509
rect 649 121 655 497
rect 689 121 695 497
rect 649 109 695 121
rect 745 497 791 509
rect 745 121 751 497
rect 785 121 791 497
rect 745 109 791 121
rect 841 497 887 509
rect 841 121 847 497
rect 881 121 887 497
rect 841 109 887 121
rect 937 497 983 509
rect 937 121 943 497
rect 977 121 983 497
rect 937 109 983 121
rect 1033 497 1079 509
rect 1033 121 1039 497
rect 1073 121 1079 497
rect 1033 109 1079 121
rect 1129 497 1175 509
rect 1129 121 1135 497
rect 1169 121 1175 497
rect 1129 109 1175 121
rect 1225 497 1271 509
rect 1225 121 1231 497
rect 1265 121 1271 497
rect 1225 109 1271 121
rect 1321 497 1367 509
rect 1321 121 1327 497
rect 1361 121 1367 497
rect 1321 109 1367 121
rect 1417 497 1463 509
rect 1417 121 1423 497
rect 1457 121 1463 497
rect 1417 109 1463 121
rect 1513 497 1559 509
rect 1513 121 1519 497
rect 1553 121 1559 497
rect 1513 109 1559 121
rect 1609 497 1655 509
rect 1609 121 1615 497
rect 1649 121 1655 497
rect 1609 109 1655 121
rect 1705 497 1751 509
rect 1705 121 1711 497
rect 1745 121 1751 497
rect 1705 109 1751 121
rect 1801 497 1847 509
rect 1801 121 1807 497
rect 1841 121 1847 497
rect 1801 109 1847 121
rect 1897 497 1943 509
rect 1897 121 1903 497
rect 1937 121 1943 497
rect 1897 109 1943 121
rect 1993 497 2039 509
rect 1993 121 1999 497
rect 2033 121 2039 497
rect 1993 109 2039 121
rect 2089 497 2135 509
rect 2089 121 2095 497
rect 2129 121 2135 497
rect 2089 109 2135 121
rect 2185 497 2231 509
rect 2185 121 2191 497
rect 2225 121 2231 497
rect 2185 109 2231 121
rect 2281 497 2327 509
rect 2281 121 2287 497
rect 2321 121 2327 497
rect 2281 109 2327 121
rect 2377 497 2423 509
rect 2377 121 2383 497
rect 2417 121 2423 497
rect 2377 109 2423 121
rect 2473 497 2519 509
rect 2473 121 2479 497
rect 2513 121 2519 497
rect 2473 109 2519 121
rect 2569 497 2615 509
rect 2569 121 2575 497
rect 2609 121 2615 497
rect 2569 109 2615 121
rect 2665 497 2711 509
rect 2665 121 2671 497
rect 2705 121 2711 497
rect 2665 109 2711 121
rect 2761 497 2807 509
rect 2761 121 2767 497
rect 2801 121 2807 497
rect 2761 109 2807 121
rect 2857 497 2903 509
rect 2857 121 2863 497
rect 2897 121 2903 497
rect 2857 109 2903 121
rect 2953 497 2999 509
rect 2953 121 2959 497
rect 2993 121 2999 497
rect 2953 109 2999 121
rect 3049 497 3095 509
rect 3049 121 3055 497
rect 3089 121 3095 497
rect 3049 109 3095 121
rect 3145 497 3191 509
rect 3145 121 3151 497
rect 3185 121 3191 497
rect 3145 109 3191 121
rect 3241 497 3287 509
rect 3241 121 3247 497
rect 3281 121 3287 497
rect 3241 109 3287 121
rect 3337 497 3383 509
rect 3337 121 3343 497
rect 3377 121 3383 497
rect 3337 109 3383 121
rect 3433 497 3479 509
rect 3433 121 3439 497
rect 3473 121 3479 497
rect 3433 109 3479 121
rect 3529 497 3575 509
rect 3529 121 3535 497
rect 3569 121 3575 497
rect 3529 109 3575 121
rect 3625 497 3671 509
rect 3625 121 3631 497
rect 3665 121 3671 497
rect 3625 109 3671 121
rect 3721 497 3767 509
rect 3721 121 3727 497
rect 3761 121 3767 497
rect 3721 109 3767 121
rect 3817 497 3863 509
rect 3817 121 3823 497
rect 3857 121 3863 497
rect 3817 109 3863 121
rect 3913 497 3959 509
rect 3913 121 3919 497
rect 3953 121 3959 497
rect 3913 109 3959 121
rect 4009 497 4055 509
rect 4009 121 4015 497
rect 4049 121 4055 497
rect 4009 109 4055 121
rect 4105 497 4151 509
rect 4105 121 4111 497
rect 4145 121 4151 497
rect 4105 109 4151 121
rect 4201 497 4247 509
rect 4201 121 4207 497
rect 4241 121 4247 497
rect 4201 109 4247 121
rect 4297 497 4343 509
rect 4297 121 4303 497
rect 4337 121 4343 497
rect 4297 109 4343 121
rect 4393 497 4439 509
rect 4393 121 4399 497
rect 4433 121 4439 497
rect 4393 109 4439 121
rect 4489 497 4535 509
rect 4489 121 4495 497
rect 4529 121 4535 497
rect 4489 109 4535 121
rect 4585 497 4631 509
rect 4585 121 4591 497
rect 4625 121 4631 497
rect 4585 109 4631 121
rect 4681 497 4727 509
rect 4681 121 4687 497
rect 4721 121 4727 497
rect 4681 109 4727 121
rect 4777 497 4823 509
rect 4777 121 4783 497
rect 4817 121 4823 497
rect 4777 109 4823 121
rect 4873 497 4919 509
rect 4873 121 4879 497
rect 4913 121 4919 497
rect 4873 109 4919 121
rect 4969 497 5015 509
rect 4969 121 4975 497
rect 5009 121 5015 497
rect 4969 109 5015 121
rect 5065 497 5111 509
rect 5065 121 5071 497
rect 5105 121 5111 497
rect 5065 109 5111 121
rect 5161 497 5207 509
rect 5161 121 5167 497
rect 5201 121 5207 497
rect 5161 109 5207 121
rect 5257 497 5303 509
rect 5257 121 5263 497
rect 5297 121 5303 497
rect 5257 109 5303 121
rect 5353 497 5399 509
rect 5353 121 5359 497
rect 5393 121 5399 497
rect 5353 109 5399 121
rect 5449 497 5495 509
rect 5449 121 5455 497
rect 5489 121 5495 497
rect 5449 109 5495 121
rect 5545 497 5591 509
rect 5545 121 5551 497
rect 5585 121 5591 497
rect 5545 109 5591 121
rect 5641 497 5687 509
rect 5641 121 5647 497
rect 5681 121 5687 497
rect 5641 109 5687 121
rect 5737 497 5783 509
rect 5737 121 5743 497
rect 5777 121 5783 497
rect 5737 109 5783 121
rect -5645 71 -5587 77
rect -5645 37 -5633 71
rect -5599 37 -5587 71
rect -5645 31 -5587 37
rect -5453 71 -5395 77
rect -5453 37 -5441 71
rect -5407 37 -5395 71
rect -5453 31 -5395 37
rect -5261 71 -5203 77
rect -5261 37 -5249 71
rect -5215 37 -5203 71
rect -5261 31 -5203 37
rect -5069 71 -5011 77
rect -5069 37 -5057 71
rect -5023 37 -5011 71
rect -5069 31 -5011 37
rect -4877 71 -4819 77
rect -4877 37 -4865 71
rect -4831 37 -4819 71
rect -4877 31 -4819 37
rect -4685 71 -4627 77
rect -4685 37 -4673 71
rect -4639 37 -4627 71
rect -4685 31 -4627 37
rect -4493 71 -4435 77
rect -4493 37 -4481 71
rect -4447 37 -4435 71
rect -4493 31 -4435 37
rect -4301 71 -4243 77
rect -4301 37 -4289 71
rect -4255 37 -4243 71
rect -4301 31 -4243 37
rect -4109 71 -4051 77
rect -4109 37 -4097 71
rect -4063 37 -4051 71
rect -4109 31 -4051 37
rect -3917 71 -3859 77
rect -3917 37 -3905 71
rect -3871 37 -3859 71
rect -3917 31 -3859 37
rect -3725 71 -3667 77
rect -3725 37 -3713 71
rect -3679 37 -3667 71
rect -3725 31 -3667 37
rect -3533 71 -3475 77
rect -3533 37 -3521 71
rect -3487 37 -3475 71
rect -3533 31 -3475 37
rect -3341 71 -3283 77
rect -3341 37 -3329 71
rect -3295 37 -3283 71
rect -3341 31 -3283 37
rect -3149 71 -3091 77
rect -3149 37 -3137 71
rect -3103 37 -3091 71
rect -3149 31 -3091 37
rect -2957 71 -2899 77
rect -2957 37 -2945 71
rect -2911 37 -2899 71
rect -2957 31 -2899 37
rect -2765 71 -2707 77
rect -2765 37 -2753 71
rect -2719 37 -2707 71
rect -2765 31 -2707 37
rect -2573 71 -2515 77
rect -2573 37 -2561 71
rect -2527 37 -2515 71
rect -2573 31 -2515 37
rect -2381 71 -2323 77
rect -2381 37 -2369 71
rect -2335 37 -2323 71
rect -2381 31 -2323 37
rect -2189 71 -2131 77
rect -2189 37 -2177 71
rect -2143 37 -2131 71
rect -2189 31 -2131 37
rect -1997 71 -1939 77
rect -1997 37 -1985 71
rect -1951 37 -1939 71
rect -1997 31 -1939 37
rect -1805 71 -1747 77
rect -1805 37 -1793 71
rect -1759 37 -1747 71
rect -1805 31 -1747 37
rect -1613 71 -1555 77
rect -1613 37 -1601 71
rect -1567 37 -1555 71
rect -1613 31 -1555 37
rect -1421 71 -1363 77
rect -1421 37 -1409 71
rect -1375 37 -1363 71
rect -1421 31 -1363 37
rect -1229 71 -1171 77
rect -1229 37 -1217 71
rect -1183 37 -1171 71
rect -1229 31 -1171 37
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect 1267 71 1325 77
rect 1267 37 1279 71
rect 1313 37 1325 71
rect 1267 31 1325 37
rect 1459 71 1517 77
rect 1459 37 1471 71
rect 1505 37 1517 71
rect 1459 31 1517 37
rect 1651 71 1709 77
rect 1651 37 1663 71
rect 1697 37 1709 71
rect 1651 31 1709 37
rect 1843 71 1901 77
rect 1843 37 1855 71
rect 1889 37 1901 71
rect 1843 31 1901 37
rect 2035 71 2093 77
rect 2035 37 2047 71
rect 2081 37 2093 71
rect 2035 31 2093 37
rect 2227 71 2285 77
rect 2227 37 2239 71
rect 2273 37 2285 71
rect 2227 31 2285 37
rect 2419 71 2477 77
rect 2419 37 2431 71
rect 2465 37 2477 71
rect 2419 31 2477 37
rect 2611 71 2669 77
rect 2611 37 2623 71
rect 2657 37 2669 71
rect 2611 31 2669 37
rect 2803 71 2861 77
rect 2803 37 2815 71
rect 2849 37 2861 71
rect 2803 31 2861 37
rect 2995 71 3053 77
rect 2995 37 3007 71
rect 3041 37 3053 71
rect 2995 31 3053 37
rect 3187 71 3245 77
rect 3187 37 3199 71
rect 3233 37 3245 71
rect 3187 31 3245 37
rect 3379 71 3437 77
rect 3379 37 3391 71
rect 3425 37 3437 71
rect 3379 31 3437 37
rect 3571 71 3629 77
rect 3571 37 3583 71
rect 3617 37 3629 71
rect 3571 31 3629 37
rect 3763 71 3821 77
rect 3763 37 3775 71
rect 3809 37 3821 71
rect 3763 31 3821 37
rect 3955 71 4013 77
rect 3955 37 3967 71
rect 4001 37 4013 71
rect 3955 31 4013 37
rect 4147 71 4205 77
rect 4147 37 4159 71
rect 4193 37 4205 71
rect 4147 31 4205 37
rect 4339 71 4397 77
rect 4339 37 4351 71
rect 4385 37 4397 71
rect 4339 31 4397 37
rect 4531 71 4589 77
rect 4531 37 4543 71
rect 4577 37 4589 71
rect 4531 31 4589 37
rect 4723 71 4781 77
rect 4723 37 4735 71
rect 4769 37 4781 71
rect 4723 31 4781 37
rect 4915 71 4973 77
rect 4915 37 4927 71
rect 4961 37 4973 71
rect 4915 31 4973 37
rect 5107 71 5165 77
rect 5107 37 5119 71
rect 5153 37 5165 71
rect 5107 31 5165 37
rect 5299 71 5357 77
rect 5299 37 5311 71
rect 5345 37 5357 71
rect 5299 31 5357 37
rect 5491 71 5549 77
rect 5491 37 5503 71
rect 5537 37 5549 71
rect 5491 31 5549 37
rect 5683 71 5741 77
rect 5683 37 5695 71
rect 5729 37 5741 71
rect 5683 31 5741 37
rect -5645 -37 -5587 -31
rect -5645 -71 -5633 -37
rect -5599 -71 -5587 -37
rect -5645 -77 -5587 -71
rect -5453 -37 -5395 -31
rect -5453 -71 -5441 -37
rect -5407 -71 -5395 -37
rect -5453 -77 -5395 -71
rect -5261 -37 -5203 -31
rect -5261 -71 -5249 -37
rect -5215 -71 -5203 -37
rect -5261 -77 -5203 -71
rect -5069 -37 -5011 -31
rect -5069 -71 -5057 -37
rect -5023 -71 -5011 -37
rect -5069 -77 -5011 -71
rect -4877 -37 -4819 -31
rect -4877 -71 -4865 -37
rect -4831 -71 -4819 -37
rect -4877 -77 -4819 -71
rect -4685 -37 -4627 -31
rect -4685 -71 -4673 -37
rect -4639 -71 -4627 -37
rect -4685 -77 -4627 -71
rect -4493 -37 -4435 -31
rect -4493 -71 -4481 -37
rect -4447 -71 -4435 -37
rect -4493 -77 -4435 -71
rect -4301 -37 -4243 -31
rect -4301 -71 -4289 -37
rect -4255 -71 -4243 -37
rect -4301 -77 -4243 -71
rect -4109 -37 -4051 -31
rect -4109 -71 -4097 -37
rect -4063 -71 -4051 -37
rect -4109 -77 -4051 -71
rect -3917 -37 -3859 -31
rect -3917 -71 -3905 -37
rect -3871 -71 -3859 -37
rect -3917 -77 -3859 -71
rect -3725 -37 -3667 -31
rect -3725 -71 -3713 -37
rect -3679 -71 -3667 -37
rect -3725 -77 -3667 -71
rect -3533 -37 -3475 -31
rect -3533 -71 -3521 -37
rect -3487 -71 -3475 -37
rect -3533 -77 -3475 -71
rect -3341 -37 -3283 -31
rect -3341 -71 -3329 -37
rect -3295 -71 -3283 -37
rect -3341 -77 -3283 -71
rect -3149 -37 -3091 -31
rect -3149 -71 -3137 -37
rect -3103 -71 -3091 -37
rect -3149 -77 -3091 -71
rect -2957 -37 -2899 -31
rect -2957 -71 -2945 -37
rect -2911 -71 -2899 -37
rect -2957 -77 -2899 -71
rect -2765 -37 -2707 -31
rect -2765 -71 -2753 -37
rect -2719 -71 -2707 -37
rect -2765 -77 -2707 -71
rect -2573 -37 -2515 -31
rect -2573 -71 -2561 -37
rect -2527 -71 -2515 -37
rect -2573 -77 -2515 -71
rect -2381 -37 -2323 -31
rect -2381 -71 -2369 -37
rect -2335 -71 -2323 -37
rect -2381 -77 -2323 -71
rect -2189 -37 -2131 -31
rect -2189 -71 -2177 -37
rect -2143 -71 -2131 -37
rect -2189 -77 -2131 -71
rect -1997 -37 -1939 -31
rect -1997 -71 -1985 -37
rect -1951 -71 -1939 -37
rect -1997 -77 -1939 -71
rect -1805 -37 -1747 -31
rect -1805 -71 -1793 -37
rect -1759 -71 -1747 -37
rect -1805 -77 -1747 -71
rect -1613 -37 -1555 -31
rect -1613 -71 -1601 -37
rect -1567 -71 -1555 -37
rect -1613 -77 -1555 -71
rect -1421 -37 -1363 -31
rect -1421 -71 -1409 -37
rect -1375 -71 -1363 -37
rect -1421 -77 -1363 -71
rect -1229 -37 -1171 -31
rect -1229 -71 -1217 -37
rect -1183 -71 -1171 -37
rect -1229 -77 -1171 -71
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect 1267 -37 1325 -31
rect 1267 -71 1279 -37
rect 1313 -71 1325 -37
rect 1267 -77 1325 -71
rect 1459 -37 1517 -31
rect 1459 -71 1471 -37
rect 1505 -71 1517 -37
rect 1459 -77 1517 -71
rect 1651 -37 1709 -31
rect 1651 -71 1663 -37
rect 1697 -71 1709 -37
rect 1651 -77 1709 -71
rect 1843 -37 1901 -31
rect 1843 -71 1855 -37
rect 1889 -71 1901 -37
rect 1843 -77 1901 -71
rect 2035 -37 2093 -31
rect 2035 -71 2047 -37
rect 2081 -71 2093 -37
rect 2035 -77 2093 -71
rect 2227 -37 2285 -31
rect 2227 -71 2239 -37
rect 2273 -71 2285 -37
rect 2227 -77 2285 -71
rect 2419 -37 2477 -31
rect 2419 -71 2431 -37
rect 2465 -71 2477 -37
rect 2419 -77 2477 -71
rect 2611 -37 2669 -31
rect 2611 -71 2623 -37
rect 2657 -71 2669 -37
rect 2611 -77 2669 -71
rect 2803 -37 2861 -31
rect 2803 -71 2815 -37
rect 2849 -71 2861 -37
rect 2803 -77 2861 -71
rect 2995 -37 3053 -31
rect 2995 -71 3007 -37
rect 3041 -71 3053 -37
rect 2995 -77 3053 -71
rect 3187 -37 3245 -31
rect 3187 -71 3199 -37
rect 3233 -71 3245 -37
rect 3187 -77 3245 -71
rect 3379 -37 3437 -31
rect 3379 -71 3391 -37
rect 3425 -71 3437 -37
rect 3379 -77 3437 -71
rect 3571 -37 3629 -31
rect 3571 -71 3583 -37
rect 3617 -71 3629 -37
rect 3571 -77 3629 -71
rect 3763 -37 3821 -31
rect 3763 -71 3775 -37
rect 3809 -71 3821 -37
rect 3763 -77 3821 -71
rect 3955 -37 4013 -31
rect 3955 -71 3967 -37
rect 4001 -71 4013 -37
rect 3955 -77 4013 -71
rect 4147 -37 4205 -31
rect 4147 -71 4159 -37
rect 4193 -71 4205 -37
rect 4147 -77 4205 -71
rect 4339 -37 4397 -31
rect 4339 -71 4351 -37
rect 4385 -71 4397 -37
rect 4339 -77 4397 -71
rect 4531 -37 4589 -31
rect 4531 -71 4543 -37
rect 4577 -71 4589 -37
rect 4531 -77 4589 -71
rect 4723 -37 4781 -31
rect 4723 -71 4735 -37
rect 4769 -71 4781 -37
rect 4723 -77 4781 -71
rect 4915 -37 4973 -31
rect 4915 -71 4927 -37
rect 4961 -71 4973 -37
rect 4915 -77 4973 -71
rect 5107 -37 5165 -31
rect 5107 -71 5119 -37
rect 5153 -71 5165 -37
rect 5107 -77 5165 -71
rect 5299 -37 5357 -31
rect 5299 -71 5311 -37
rect 5345 -71 5357 -37
rect 5299 -77 5357 -71
rect 5491 -37 5549 -31
rect 5491 -71 5503 -37
rect 5537 -71 5549 -37
rect 5491 -77 5549 -71
rect 5683 -37 5741 -31
rect 5683 -71 5695 -37
rect 5729 -71 5741 -37
rect 5683 -77 5741 -71
rect -5783 -121 -5737 -109
rect -5783 -497 -5777 -121
rect -5743 -497 -5737 -121
rect -5783 -509 -5737 -497
rect -5687 -121 -5641 -109
rect -5687 -497 -5681 -121
rect -5647 -497 -5641 -121
rect -5687 -509 -5641 -497
rect -5591 -121 -5545 -109
rect -5591 -497 -5585 -121
rect -5551 -497 -5545 -121
rect -5591 -509 -5545 -497
rect -5495 -121 -5449 -109
rect -5495 -497 -5489 -121
rect -5455 -497 -5449 -121
rect -5495 -509 -5449 -497
rect -5399 -121 -5353 -109
rect -5399 -497 -5393 -121
rect -5359 -497 -5353 -121
rect -5399 -509 -5353 -497
rect -5303 -121 -5257 -109
rect -5303 -497 -5297 -121
rect -5263 -497 -5257 -121
rect -5303 -509 -5257 -497
rect -5207 -121 -5161 -109
rect -5207 -497 -5201 -121
rect -5167 -497 -5161 -121
rect -5207 -509 -5161 -497
rect -5111 -121 -5065 -109
rect -5111 -497 -5105 -121
rect -5071 -497 -5065 -121
rect -5111 -509 -5065 -497
rect -5015 -121 -4969 -109
rect -5015 -497 -5009 -121
rect -4975 -497 -4969 -121
rect -5015 -509 -4969 -497
rect -4919 -121 -4873 -109
rect -4919 -497 -4913 -121
rect -4879 -497 -4873 -121
rect -4919 -509 -4873 -497
rect -4823 -121 -4777 -109
rect -4823 -497 -4817 -121
rect -4783 -497 -4777 -121
rect -4823 -509 -4777 -497
rect -4727 -121 -4681 -109
rect -4727 -497 -4721 -121
rect -4687 -497 -4681 -121
rect -4727 -509 -4681 -497
rect -4631 -121 -4585 -109
rect -4631 -497 -4625 -121
rect -4591 -497 -4585 -121
rect -4631 -509 -4585 -497
rect -4535 -121 -4489 -109
rect -4535 -497 -4529 -121
rect -4495 -497 -4489 -121
rect -4535 -509 -4489 -497
rect -4439 -121 -4393 -109
rect -4439 -497 -4433 -121
rect -4399 -497 -4393 -121
rect -4439 -509 -4393 -497
rect -4343 -121 -4297 -109
rect -4343 -497 -4337 -121
rect -4303 -497 -4297 -121
rect -4343 -509 -4297 -497
rect -4247 -121 -4201 -109
rect -4247 -497 -4241 -121
rect -4207 -497 -4201 -121
rect -4247 -509 -4201 -497
rect -4151 -121 -4105 -109
rect -4151 -497 -4145 -121
rect -4111 -497 -4105 -121
rect -4151 -509 -4105 -497
rect -4055 -121 -4009 -109
rect -4055 -497 -4049 -121
rect -4015 -497 -4009 -121
rect -4055 -509 -4009 -497
rect -3959 -121 -3913 -109
rect -3959 -497 -3953 -121
rect -3919 -497 -3913 -121
rect -3959 -509 -3913 -497
rect -3863 -121 -3817 -109
rect -3863 -497 -3857 -121
rect -3823 -497 -3817 -121
rect -3863 -509 -3817 -497
rect -3767 -121 -3721 -109
rect -3767 -497 -3761 -121
rect -3727 -497 -3721 -121
rect -3767 -509 -3721 -497
rect -3671 -121 -3625 -109
rect -3671 -497 -3665 -121
rect -3631 -497 -3625 -121
rect -3671 -509 -3625 -497
rect -3575 -121 -3529 -109
rect -3575 -497 -3569 -121
rect -3535 -497 -3529 -121
rect -3575 -509 -3529 -497
rect -3479 -121 -3433 -109
rect -3479 -497 -3473 -121
rect -3439 -497 -3433 -121
rect -3479 -509 -3433 -497
rect -3383 -121 -3337 -109
rect -3383 -497 -3377 -121
rect -3343 -497 -3337 -121
rect -3383 -509 -3337 -497
rect -3287 -121 -3241 -109
rect -3287 -497 -3281 -121
rect -3247 -497 -3241 -121
rect -3287 -509 -3241 -497
rect -3191 -121 -3145 -109
rect -3191 -497 -3185 -121
rect -3151 -497 -3145 -121
rect -3191 -509 -3145 -497
rect -3095 -121 -3049 -109
rect -3095 -497 -3089 -121
rect -3055 -497 -3049 -121
rect -3095 -509 -3049 -497
rect -2999 -121 -2953 -109
rect -2999 -497 -2993 -121
rect -2959 -497 -2953 -121
rect -2999 -509 -2953 -497
rect -2903 -121 -2857 -109
rect -2903 -497 -2897 -121
rect -2863 -497 -2857 -121
rect -2903 -509 -2857 -497
rect -2807 -121 -2761 -109
rect -2807 -497 -2801 -121
rect -2767 -497 -2761 -121
rect -2807 -509 -2761 -497
rect -2711 -121 -2665 -109
rect -2711 -497 -2705 -121
rect -2671 -497 -2665 -121
rect -2711 -509 -2665 -497
rect -2615 -121 -2569 -109
rect -2615 -497 -2609 -121
rect -2575 -497 -2569 -121
rect -2615 -509 -2569 -497
rect -2519 -121 -2473 -109
rect -2519 -497 -2513 -121
rect -2479 -497 -2473 -121
rect -2519 -509 -2473 -497
rect -2423 -121 -2377 -109
rect -2423 -497 -2417 -121
rect -2383 -497 -2377 -121
rect -2423 -509 -2377 -497
rect -2327 -121 -2281 -109
rect -2327 -497 -2321 -121
rect -2287 -497 -2281 -121
rect -2327 -509 -2281 -497
rect -2231 -121 -2185 -109
rect -2231 -497 -2225 -121
rect -2191 -497 -2185 -121
rect -2231 -509 -2185 -497
rect -2135 -121 -2089 -109
rect -2135 -497 -2129 -121
rect -2095 -497 -2089 -121
rect -2135 -509 -2089 -497
rect -2039 -121 -1993 -109
rect -2039 -497 -2033 -121
rect -1999 -497 -1993 -121
rect -2039 -509 -1993 -497
rect -1943 -121 -1897 -109
rect -1943 -497 -1937 -121
rect -1903 -497 -1897 -121
rect -1943 -509 -1897 -497
rect -1847 -121 -1801 -109
rect -1847 -497 -1841 -121
rect -1807 -497 -1801 -121
rect -1847 -509 -1801 -497
rect -1751 -121 -1705 -109
rect -1751 -497 -1745 -121
rect -1711 -497 -1705 -121
rect -1751 -509 -1705 -497
rect -1655 -121 -1609 -109
rect -1655 -497 -1649 -121
rect -1615 -497 -1609 -121
rect -1655 -509 -1609 -497
rect -1559 -121 -1513 -109
rect -1559 -497 -1553 -121
rect -1519 -497 -1513 -121
rect -1559 -509 -1513 -497
rect -1463 -121 -1417 -109
rect -1463 -497 -1457 -121
rect -1423 -497 -1417 -121
rect -1463 -509 -1417 -497
rect -1367 -121 -1321 -109
rect -1367 -497 -1361 -121
rect -1327 -497 -1321 -121
rect -1367 -509 -1321 -497
rect -1271 -121 -1225 -109
rect -1271 -497 -1265 -121
rect -1231 -497 -1225 -121
rect -1271 -509 -1225 -497
rect -1175 -121 -1129 -109
rect -1175 -497 -1169 -121
rect -1135 -497 -1129 -121
rect -1175 -509 -1129 -497
rect -1079 -121 -1033 -109
rect -1079 -497 -1073 -121
rect -1039 -497 -1033 -121
rect -1079 -509 -1033 -497
rect -983 -121 -937 -109
rect -983 -497 -977 -121
rect -943 -497 -937 -121
rect -983 -509 -937 -497
rect -887 -121 -841 -109
rect -887 -497 -881 -121
rect -847 -497 -841 -121
rect -887 -509 -841 -497
rect -791 -121 -745 -109
rect -791 -497 -785 -121
rect -751 -497 -745 -121
rect -791 -509 -745 -497
rect -695 -121 -649 -109
rect -695 -497 -689 -121
rect -655 -497 -649 -121
rect -695 -509 -649 -497
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect 649 -121 695 -109
rect 649 -497 655 -121
rect 689 -497 695 -121
rect 649 -509 695 -497
rect 745 -121 791 -109
rect 745 -497 751 -121
rect 785 -497 791 -121
rect 745 -509 791 -497
rect 841 -121 887 -109
rect 841 -497 847 -121
rect 881 -497 887 -121
rect 841 -509 887 -497
rect 937 -121 983 -109
rect 937 -497 943 -121
rect 977 -497 983 -121
rect 937 -509 983 -497
rect 1033 -121 1079 -109
rect 1033 -497 1039 -121
rect 1073 -497 1079 -121
rect 1033 -509 1079 -497
rect 1129 -121 1175 -109
rect 1129 -497 1135 -121
rect 1169 -497 1175 -121
rect 1129 -509 1175 -497
rect 1225 -121 1271 -109
rect 1225 -497 1231 -121
rect 1265 -497 1271 -121
rect 1225 -509 1271 -497
rect 1321 -121 1367 -109
rect 1321 -497 1327 -121
rect 1361 -497 1367 -121
rect 1321 -509 1367 -497
rect 1417 -121 1463 -109
rect 1417 -497 1423 -121
rect 1457 -497 1463 -121
rect 1417 -509 1463 -497
rect 1513 -121 1559 -109
rect 1513 -497 1519 -121
rect 1553 -497 1559 -121
rect 1513 -509 1559 -497
rect 1609 -121 1655 -109
rect 1609 -497 1615 -121
rect 1649 -497 1655 -121
rect 1609 -509 1655 -497
rect 1705 -121 1751 -109
rect 1705 -497 1711 -121
rect 1745 -497 1751 -121
rect 1705 -509 1751 -497
rect 1801 -121 1847 -109
rect 1801 -497 1807 -121
rect 1841 -497 1847 -121
rect 1801 -509 1847 -497
rect 1897 -121 1943 -109
rect 1897 -497 1903 -121
rect 1937 -497 1943 -121
rect 1897 -509 1943 -497
rect 1993 -121 2039 -109
rect 1993 -497 1999 -121
rect 2033 -497 2039 -121
rect 1993 -509 2039 -497
rect 2089 -121 2135 -109
rect 2089 -497 2095 -121
rect 2129 -497 2135 -121
rect 2089 -509 2135 -497
rect 2185 -121 2231 -109
rect 2185 -497 2191 -121
rect 2225 -497 2231 -121
rect 2185 -509 2231 -497
rect 2281 -121 2327 -109
rect 2281 -497 2287 -121
rect 2321 -497 2327 -121
rect 2281 -509 2327 -497
rect 2377 -121 2423 -109
rect 2377 -497 2383 -121
rect 2417 -497 2423 -121
rect 2377 -509 2423 -497
rect 2473 -121 2519 -109
rect 2473 -497 2479 -121
rect 2513 -497 2519 -121
rect 2473 -509 2519 -497
rect 2569 -121 2615 -109
rect 2569 -497 2575 -121
rect 2609 -497 2615 -121
rect 2569 -509 2615 -497
rect 2665 -121 2711 -109
rect 2665 -497 2671 -121
rect 2705 -497 2711 -121
rect 2665 -509 2711 -497
rect 2761 -121 2807 -109
rect 2761 -497 2767 -121
rect 2801 -497 2807 -121
rect 2761 -509 2807 -497
rect 2857 -121 2903 -109
rect 2857 -497 2863 -121
rect 2897 -497 2903 -121
rect 2857 -509 2903 -497
rect 2953 -121 2999 -109
rect 2953 -497 2959 -121
rect 2993 -497 2999 -121
rect 2953 -509 2999 -497
rect 3049 -121 3095 -109
rect 3049 -497 3055 -121
rect 3089 -497 3095 -121
rect 3049 -509 3095 -497
rect 3145 -121 3191 -109
rect 3145 -497 3151 -121
rect 3185 -497 3191 -121
rect 3145 -509 3191 -497
rect 3241 -121 3287 -109
rect 3241 -497 3247 -121
rect 3281 -497 3287 -121
rect 3241 -509 3287 -497
rect 3337 -121 3383 -109
rect 3337 -497 3343 -121
rect 3377 -497 3383 -121
rect 3337 -509 3383 -497
rect 3433 -121 3479 -109
rect 3433 -497 3439 -121
rect 3473 -497 3479 -121
rect 3433 -509 3479 -497
rect 3529 -121 3575 -109
rect 3529 -497 3535 -121
rect 3569 -497 3575 -121
rect 3529 -509 3575 -497
rect 3625 -121 3671 -109
rect 3625 -497 3631 -121
rect 3665 -497 3671 -121
rect 3625 -509 3671 -497
rect 3721 -121 3767 -109
rect 3721 -497 3727 -121
rect 3761 -497 3767 -121
rect 3721 -509 3767 -497
rect 3817 -121 3863 -109
rect 3817 -497 3823 -121
rect 3857 -497 3863 -121
rect 3817 -509 3863 -497
rect 3913 -121 3959 -109
rect 3913 -497 3919 -121
rect 3953 -497 3959 -121
rect 3913 -509 3959 -497
rect 4009 -121 4055 -109
rect 4009 -497 4015 -121
rect 4049 -497 4055 -121
rect 4009 -509 4055 -497
rect 4105 -121 4151 -109
rect 4105 -497 4111 -121
rect 4145 -497 4151 -121
rect 4105 -509 4151 -497
rect 4201 -121 4247 -109
rect 4201 -497 4207 -121
rect 4241 -497 4247 -121
rect 4201 -509 4247 -497
rect 4297 -121 4343 -109
rect 4297 -497 4303 -121
rect 4337 -497 4343 -121
rect 4297 -509 4343 -497
rect 4393 -121 4439 -109
rect 4393 -497 4399 -121
rect 4433 -497 4439 -121
rect 4393 -509 4439 -497
rect 4489 -121 4535 -109
rect 4489 -497 4495 -121
rect 4529 -497 4535 -121
rect 4489 -509 4535 -497
rect 4585 -121 4631 -109
rect 4585 -497 4591 -121
rect 4625 -497 4631 -121
rect 4585 -509 4631 -497
rect 4681 -121 4727 -109
rect 4681 -497 4687 -121
rect 4721 -497 4727 -121
rect 4681 -509 4727 -497
rect 4777 -121 4823 -109
rect 4777 -497 4783 -121
rect 4817 -497 4823 -121
rect 4777 -509 4823 -497
rect 4873 -121 4919 -109
rect 4873 -497 4879 -121
rect 4913 -497 4919 -121
rect 4873 -509 4919 -497
rect 4969 -121 5015 -109
rect 4969 -497 4975 -121
rect 5009 -497 5015 -121
rect 4969 -509 5015 -497
rect 5065 -121 5111 -109
rect 5065 -497 5071 -121
rect 5105 -497 5111 -121
rect 5065 -509 5111 -497
rect 5161 -121 5207 -109
rect 5161 -497 5167 -121
rect 5201 -497 5207 -121
rect 5161 -509 5207 -497
rect 5257 -121 5303 -109
rect 5257 -497 5263 -121
rect 5297 -497 5303 -121
rect 5257 -509 5303 -497
rect 5353 -121 5399 -109
rect 5353 -497 5359 -121
rect 5393 -497 5399 -121
rect 5353 -509 5399 -497
rect 5449 -121 5495 -109
rect 5449 -497 5455 -121
rect 5489 -497 5495 -121
rect 5449 -509 5495 -497
rect 5545 -121 5591 -109
rect 5545 -497 5551 -121
rect 5585 -497 5591 -121
rect 5545 -509 5591 -497
rect 5641 -121 5687 -109
rect 5641 -497 5647 -121
rect 5681 -497 5687 -121
rect 5641 -509 5687 -497
rect 5737 -121 5783 -109
rect 5737 -497 5743 -121
rect 5777 -497 5783 -121
rect 5737 -509 5783 -497
rect -5741 -547 -5683 -541
rect -5741 -581 -5729 -547
rect -5695 -581 -5683 -547
rect -5741 -587 -5683 -581
rect -5549 -547 -5491 -541
rect -5549 -581 -5537 -547
rect -5503 -581 -5491 -547
rect -5549 -587 -5491 -581
rect -5357 -547 -5299 -541
rect -5357 -581 -5345 -547
rect -5311 -581 -5299 -547
rect -5357 -587 -5299 -581
rect -5165 -547 -5107 -541
rect -5165 -581 -5153 -547
rect -5119 -581 -5107 -547
rect -5165 -587 -5107 -581
rect -4973 -547 -4915 -541
rect -4973 -581 -4961 -547
rect -4927 -581 -4915 -547
rect -4973 -587 -4915 -581
rect -4781 -547 -4723 -541
rect -4781 -581 -4769 -547
rect -4735 -581 -4723 -547
rect -4781 -587 -4723 -581
rect -4589 -547 -4531 -541
rect -4589 -581 -4577 -547
rect -4543 -581 -4531 -547
rect -4589 -587 -4531 -581
rect -4397 -547 -4339 -541
rect -4397 -581 -4385 -547
rect -4351 -581 -4339 -547
rect -4397 -587 -4339 -581
rect -4205 -547 -4147 -541
rect -4205 -581 -4193 -547
rect -4159 -581 -4147 -547
rect -4205 -587 -4147 -581
rect -4013 -547 -3955 -541
rect -4013 -581 -4001 -547
rect -3967 -581 -3955 -547
rect -4013 -587 -3955 -581
rect -3821 -547 -3763 -541
rect -3821 -581 -3809 -547
rect -3775 -581 -3763 -547
rect -3821 -587 -3763 -581
rect -3629 -547 -3571 -541
rect -3629 -581 -3617 -547
rect -3583 -581 -3571 -547
rect -3629 -587 -3571 -581
rect -3437 -547 -3379 -541
rect -3437 -581 -3425 -547
rect -3391 -581 -3379 -547
rect -3437 -587 -3379 -581
rect -3245 -547 -3187 -541
rect -3245 -581 -3233 -547
rect -3199 -581 -3187 -547
rect -3245 -587 -3187 -581
rect -3053 -547 -2995 -541
rect -3053 -581 -3041 -547
rect -3007 -581 -2995 -547
rect -3053 -587 -2995 -581
rect -2861 -547 -2803 -541
rect -2861 -581 -2849 -547
rect -2815 -581 -2803 -547
rect -2861 -587 -2803 -581
rect -2669 -547 -2611 -541
rect -2669 -581 -2657 -547
rect -2623 -581 -2611 -547
rect -2669 -587 -2611 -581
rect -2477 -547 -2419 -541
rect -2477 -581 -2465 -547
rect -2431 -581 -2419 -547
rect -2477 -587 -2419 -581
rect -2285 -547 -2227 -541
rect -2285 -581 -2273 -547
rect -2239 -581 -2227 -547
rect -2285 -587 -2227 -581
rect -2093 -547 -2035 -541
rect -2093 -581 -2081 -547
rect -2047 -581 -2035 -547
rect -2093 -587 -2035 -581
rect -1901 -547 -1843 -541
rect -1901 -581 -1889 -547
rect -1855 -581 -1843 -547
rect -1901 -587 -1843 -581
rect -1709 -547 -1651 -541
rect -1709 -581 -1697 -547
rect -1663 -581 -1651 -547
rect -1709 -587 -1651 -581
rect -1517 -547 -1459 -541
rect -1517 -581 -1505 -547
rect -1471 -581 -1459 -547
rect -1517 -587 -1459 -581
rect -1325 -547 -1267 -541
rect -1325 -581 -1313 -547
rect -1279 -581 -1267 -547
rect -1325 -587 -1267 -581
rect -1133 -547 -1075 -541
rect -1133 -581 -1121 -547
rect -1087 -581 -1075 -547
rect -1133 -587 -1075 -581
rect -941 -547 -883 -541
rect -941 -581 -929 -547
rect -895 -581 -883 -547
rect -941 -587 -883 -581
rect -749 -547 -691 -541
rect -749 -581 -737 -547
rect -703 -581 -691 -547
rect -749 -587 -691 -581
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
rect 595 -547 653 -541
rect 595 -581 607 -547
rect 641 -581 653 -547
rect 595 -587 653 -581
rect 787 -547 845 -541
rect 787 -581 799 -547
rect 833 -581 845 -547
rect 787 -587 845 -581
rect 979 -547 1037 -541
rect 979 -581 991 -547
rect 1025 -581 1037 -547
rect 979 -587 1037 -581
rect 1171 -547 1229 -541
rect 1171 -581 1183 -547
rect 1217 -581 1229 -547
rect 1171 -587 1229 -581
rect 1363 -547 1421 -541
rect 1363 -581 1375 -547
rect 1409 -581 1421 -547
rect 1363 -587 1421 -581
rect 1555 -547 1613 -541
rect 1555 -581 1567 -547
rect 1601 -581 1613 -547
rect 1555 -587 1613 -581
rect 1747 -547 1805 -541
rect 1747 -581 1759 -547
rect 1793 -581 1805 -547
rect 1747 -587 1805 -581
rect 1939 -547 1997 -541
rect 1939 -581 1951 -547
rect 1985 -581 1997 -547
rect 1939 -587 1997 -581
rect 2131 -547 2189 -541
rect 2131 -581 2143 -547
rect 2177 -581 2189 -547
rect 2131 -587 2189 -581
rect 2323 -547 2381 -541
rect 2323 -581 2335 -547
rect 2369 -581 2381 -547
rect 2323 -587 2381 -581
rect 2515 -547 2573 -541
rect 2515 -581 2527 -547
rect 2561 -581 2573 -547
rect 2515 -587 2573 -581
rect 2707 -547 2765 -541
rect 2707 -581 2719 -547
rect 2753 -581 2765 -547
rect 2707 -587 2765 -581
rect 2899 -547 2957 -541
rect 2899 -581 2911 -547
rect 2945 -581 2957 -547
rect 2899 -587 2957 -581
rect 3091 -547 3149 -541
rect 3091 -581 3103 -547
rect 3137 -581 3149 -547
rect 3091 -587 3149 -581
rect 3283 -547 3341 -541
rect 3283 -581 3295 -547
rect 3329 -581 3341 -547
rect 3283 -587 3341 -581
rect 3475 -547 3533 -541
rect 3475 -581 3487 -547
rect 3521 -581 3533 -547
rect 3475 -587 3533 -581
rect 3667 -547 3725 -541
rect 3667 -581 3679 -547
rect 3713 -581 3725 -547
rect 3667 -587 3725 -581
rect 3859 -547 3917 -541
rect 3859 -581 3871 -547
rect 3905 -581 3917 -547
rect 3859 -587 3917 -581
rect 4051 -547 4109 -541
rect 4051 -581 4063 -547
rect 4097 -581 4109 -547
rect 4051 -587 4109 -581
rect 4243 -547 4301 -541
rect 4243 -581 4255 -547
rect 4289 -581 4301 -547
rect 4243 -587 4301 -581
rect 4435 -547 4493 -541
rect 4435 -581 4447 -547
rect 4481 -581 4493 -547
rect 4435 -587 4493 -581
rect 4627 -547 4685 -541
rect 4627 -581 4639 -547
rect 4673 -581 4685 -547
rect 4627 -587 4685 -581
rect 4819 -547 4877 -541
rect 4819 -581 4831 -547
rect 4865 -581 4877 -547
rect 4819 -587 4877 -581
rect 5011 -547 5069 -541
rect 5011 -581 5023 -547
rect 5057 -581 5069 -547
rect 5011 -587 5069 -581
rect 5203 -547 5261 -541
rect 5203 -581 5215 -547
rect 5249 -581 5261 -547
rect 5203 -587 5261 -581
rect 5395 -547 5453 -541
rect 5395 -581 5407 -547
rect 5441 -581 5453 -547
rect 5395 -587 5453 -581
rect 5587 -547 5645 -541
rect 5587 -581 5599 -547
rect 5633 -581 5645 -547
rect 5587 -587 5645 -581
<< properties >>
string FIXED_BBOX -5874 -666 5874 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 2 nf 120 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
