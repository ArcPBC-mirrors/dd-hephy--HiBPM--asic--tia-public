magic
tech sky130A
magscale 1 2
timestamp 1683540360
<< metal3 >>
rect -986 1012 986 1040
rect -986 -1012 902 1012
rect 966 -1012 986 1012
rect -986 -1040 986 -1012
<< via3 >>
rect 902 -1012 966 1012
<< mimcap >>
rect -946 960 654 1000
rect -946 -960 -906 960
rect 614 -960 654 960
rect -946 -1000 654 -960
<< mimcapcontact >>
rect -906 -960 614 960
<< metal4 >>
rect 886 1012 982 1028
rect -907 960 615 961
rect -907 -960 -906 960
rect 614 -960 615 960
rect -907 -961 615 -960
rect 886 -1012 902 1012
rect 966 -1012 982 1012
rect 886 -1028 982 -1012
<< properties >>
string FIXED_BBOX -986 -1040 694 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 8 l 10 val 166.84 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
