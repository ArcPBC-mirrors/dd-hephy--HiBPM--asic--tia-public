magic
tech sky130A
magscale 1 2
timestamp 1685113734
<< metal1 >>
rect 280 2476 3200 2600
rect 326 2264 336 2448
rect 388 2264 398 2448
rect 518 2264 528 2448
rect 580 2264 590 2448
rect 710 2264 720 2448
rect 772 2264 782 2448
rect 902 2264 912 2448
rect 964 2264 974 2448
rect 1094 2264 1104 2448
rect 1156 2264 1166 2448
rect 1286 2264 1296 2448
rect 1348 2264 1358 2448
rect 1478 2264 1488 2448
rect 1540 2264 1550 2448
rect 1670 2264 1680 2448
rect 1732 2264 1742 2448
rect 1862 2264 1872 2448
rect 1924 2264 1934 2448
rect 2054 2264 2064 2448
rect 2116 2264 2126 2448
rect 2246 2264 2256 2448
rect 2308 2264 2318 2448
rect 2438 2264 2448 2448
rect 2500 2264 2510 2448
rect 2630 2264 2640 2448
rect 2692 2264 2702 2448
rect 2822 2264 2832 2448
rect 2884 2264 2894 2448
rect 3014 2264 3024 2448
rect 3076 2264 3086 2448
rect 230 2044 240 2228
rect 292 2044 302 2228
rect 422 2044 432 2228
rect 484 2044 494 2228
rect 614 2044 624 2228
rect 676 2044 686 2228
rect 806 2044 816 2228
rect 868 2044 878 2228
rect 998 2044 1008 2228
rect 1060 2044 1070 2228
rect 1190 2044 1200 2228
rect 1252 2044 1262 2228
rect 1382 2044 1392 2228
rect 1444 2044 1454 2228
rect 1574 2044 1584 2228
rect 1636 2044 1646 2228
rect 1766 2044 1776 2228
rect 1828 2044 1838 2228
rect 1958 2044 1968 2228
rect 2020 2044 2030 2228
rect 2150 2044 2160 2228
rect 2212 2044 2222 2228
rect 2342 2044 2352 2228
rect 2404 2044 2414 2228
rect 2534 2044 2544 2228
rect 2596 2044 2606 2228
rect 2726 2044 2736 2228
rect 2788 2044 2798 2228
rect 2918 2044 2928 2228
rect 2980 2044 2990 2228
rect 3110 2044 3120 2228
rect 3172 2044 3182 2228
rect 376 1856 3200 2012
rect 326 1644 336 1828
rect 388 1644 398 1828
rect 518 1644 528 1828
rect 580 1644 590 1828
rect 710 1644 720 1828
rect 772 1644 782 1828
rect 902 1644 912 1828
rect 964 1644 974 1828
rect 1094 1644 1104 1828
rect 1156 1644 1166 1828
rect 1286 1644 1296 1828
rect 1348 1644 1358 1828
rect 1478 1644 1488 1828
rect 1540 1644 1550 1828
rect 1670 1644 1680 1828
rect 1732 1644 1742 1828
rect 1862 1644 1872 1828
rect 1924 1644 1934 1828
rect 2054 1644 2064 1828
rect 2116 1644 2126 1828
rect 2246 1644 2256 1828
rect 2308 1644 2318 1828
rect 2438 1644 2448 1828
rect 2500 1644 2510 1828
rect 2630 1644 2640 1828
rect 2692 1644 2702 1828
rect 2822 1644 2832 1828
rect 2884 1644 2894 1828
rect 3014 1644 3024 1828
rect 3076 1644 3086 1828
rect 230 1424 240 1608
rect 292 1424 302 1608
rect 422 1424 432 1608
rect 484 1424 494 1608
rect 614 1424 624 1608
rect 676 1424 686 1608
rect 806 1424 816 1608
rect 868 1424 878 1608
rect 998 1424 1008 1608
rect 1060 1424 1070 1608
rect 1190 1424 1200 1608
rect 1252 1424 1262 1608
rect 1382 1424 1392 1608
rect 1444 1424 1454 1608
rect 1574 1424 1584 1608
rect 1636 1424 1646 1608
rect 1766 1424 1776 1608
rect 1828 1424 1838 1608
rect 1958 1424 1968 1608
rect 2020 1424 2030 1608
rect 2150 1424 2160 1608
rect 2212 1424 2222 1608
rect 2342 1424 2352 1608
rect 2404 1424 2414 1608
rect 2534 1424 2544 1608
rect 2596 1424 2606 1608
rect 2726 1424 2736 1608
rect 2788 1424 2798 1608
rect 2918 1424 2928 1608
rect 2980 1424 2990 1608
rect 3110 1424 3120 1608
rect 3172 1424 3182 1608
rect 280 1240 3200 1396
rect 326 1028 336 1212
rect 388 1028 398 1212
rect 518 1028 528 1212
rect 580 1028 590 1212
rect 710 1028 720 1212
rect 772 1028 782 1212
rect 902 1028 912 1212
rect 964 1028 974 1212
rect 1094 1028 1104 1212
rect 1156 1028 1166 1212
rect 1286 1028 1296 1212
rect 1348 1028 1358 1212
rect 1478 1028 1488 1212
rect 1540 1028 1550 1212
rect 1670 1028 1680 1212
rect 1732 1028 1742 1212
rect 1862 1028 1872 1212
rect 1924 1028 1934 1212
rect 2054 1028 2064 1212
rect 2116 1028 2126 1212
rect 2246 1028 2256 1212
rect 2308 1028 2318 1212
rect 2438 1028 2448 1212
rect 2500 1028 2510 1212
rect 2630 1028 2640 1212
rect 2692 1028 2702 1212
rect 2822 1028 2832 1212
rect 2884 1028 2894 1212
rect 3014 1028 3024 1212
rect 3076 1028 3086 1212
rect 230 808 240 992
rect 292 808 302 992
rect 422 808 432 992
rect 484 808 494 992
rect 614 808 624 992
rect 676 808 686 992
rect 806 808 816 992
rect 868 808 878 992
rect 998 808 1008 992
rect 1060 808 1070 992
rect 1190 808 1200 992
rect 1252 808 1262 992
rect 1382 808 1392 992
rect 1444 808 1454 992
rect 1574 808 1584 992
rect 1636 808 1646 992
rect 1766 808 1776 992
rect 1828 808 1838 992
rect 1958 808 1968 992
rect 2020 808 2030 992
rect 2150 808 2160 992
rect 2212 808 2222 992
rect 2342 808 2352 992
rect 2404 808 2414 992
rect 2534 808 2544 992
rect 2596 808 2606 992
rect 2726 808 2736 992
rect 2788 808 2798 992
rect 2918 808 2928 992
rect 2980 808 2990 992
rect 3110 808 3120 992
rect 3172 808 3182 992
rect 372 620 3200 776
rect 326 408 336 592
rect 388 408 398 592
rect 518 408 528 592
rect 580 408 590 592
rect 710 408 720 592
rect 772 408 782 592
rect 902 408 912 592
rect 964 408 974 592
rect 1094 408 1104 592
rect 1156 408 1166 592
rect 1286 408 1296 592
rect 1348 408 1358 592
rect 1478 408 1488 592
rect 1540 408 1550 592
rect 1670 408 1680 592
rect 1732 408 1742 592
rect 1862 408 1872 592
rect 1924 408 1934 592
rect 2054 408 2064 592
rect 2116 408 2126 592
rect 2246 408 2256 592
rect 2308 408 2318 592
rect 2438 408 2448 592
rect 2500 408 2510 592
rect 2630 408 2640 592
rect 2692 408 2702 592
rect 2822 408 2832 592
rect 2884 408 2894 592
rect 3014 408 3024 592
rect 3076 408 3086 592
rect 230 188 240 372
rect 292 188 302 372
rect 422 188 432 372
rect 484 188 494 372
rect 614 188 624 372
rect 676 188 686 372
rect 806 188 816 372
rect 868 188 878 372
rect 998 188 1008 372
rect 1060 188 1070 372
rect 1190 188 1200 372
rect 1252 188 1262 372
rect 1382 188 1392 372
rect 1444 188 1454 372
rect 1574 188 1584 372
rect 1636 188 1646 372
rect 1766 188 1776 372
rect 1828 188 1838 372
rect 1958 188 1968 372
rect 2020 188 2030 372
rect 2150 188 2160 372
rect 2212 188 2222 372
rect 2342 188 2352 372
rect 2404 188 2414 372
rect 2534 188 2544 372
rect 2596 188 2606 372
rect 2726 188 2736 372
rect 2788 188 2798 372
rect 2918 188 2928 372
rect 2980 188 2990 372
rect 3110 188 3120 372
rect 3172 188 3182 372
rect 260 20 3200 160
<< via1 >>
rect 336 2264 388 2448
rect 528 2264 580 2448
rect 720 2264 772 2448
rect 912 2264 964 2448
rect 1104 2264 1156 2448
rect 1296 2264 1348 2448
rect 1488 2264 1540 2448
rect 1680 2264 1732 2448
rect 1872 2264 1924 2448
rect 2064 2264 2116 2448
rect 2256 2264 2308 2448
rect 2448 2264 2500 2448
rect 2640 2264 2692 2448
rect 2832 2264 2884 2448
rect 3024 2264 3076 2448
rect 240 2044 292 2228
rect 432 2044 484 2228
rect 624 2044 676 2228
rect 816 2044 868 2228
rect 1008 2044 1060 2228
rect 1200 2044 1252 2228
rect 1392 2044 1444 2228
rect 1584 2044 1636 2228
rect 1776 2044 1828 2228
rect 1968 2044 2020 2228
rect 2160 2044 2212 2228
rect 2352 2044 2404 2228
rect 2544 2044 2596 2228
rect 2736 2044 2788 2228
rect 2928 2044 2980 2228
rect 3120 2044 3172 2228
rect 336 1644 388 1828
rect 528 1644 580 1828
rect 720 1644 772 1828
rect 912 1644 964 1828
rect 1104 1644 1156 1828
rect 1296 1644 1348 1828
rect 1488 1644 1540 1828
rect 1680 1644 1732 1828
rect 1872 1644 1924 1828
rect 2064 1644 2116 1828
rect 2256 1644 2308 1828
rect 2448 1644 2500 1828
rect 2640 1644 2692 1828
rect 2832 1644 2884 1828
rect 3024 1644 3076 1828
rect 240 1424 292 1608
rect 432 1424 484 1608
rect 624 1424 676 1608
rect 816 1424 868 1608
rect 1008 1424 1060 1608
rect 1200 1424 1252 1608
rect 1392 1424 1444 1608
rect 1584 1424 1636 1608
rect 1776 1424 1828 1608
rect 1968 1424 2020 1608
rect 2160 1424 2212 1608
rect 2352 1424 2404 1608
rect 2544 1424 2596 1608
rect 2736 1424 2788 1608
rect 2928 1424 2980 1608
rect 3120 1424 3172 1608
rect 336 1028 388 1212
rect 528 1028 580 1212
rect 720 1028 772 1212
rect 912 1028 964 1212
rect 1104 1028 1156 1212
rect 1296 1028 1348 1212
rect 1488 1028 1540 1212
rect 1680 1028 1732 1212
rect 1872 1028 1924 1212
rect 2064 1028 2116 1212
rect 2256 1028 2308 1212
rect 2448 1028 2500 1212
rect 2640 1028 2692 1212
rect 2832 1028 2884 1212
rect 3024 1028 3076 1212
rect 240 808 292 992
rect 432 808 484 992
rect 624 808 676 992
rect 816 808 868 992
rect 1008 808 1060 992
rect 1200 808 1252 992
rect 1392 808 1444 992
rect 1584 808 1636 992
rect 1776 808 1828 992
rect 1968 808 2020 992
rect 2160 808 2212 992
rect 2352 808 2404 992
rect 2544 808 2596 992
rect 2736 808 2788 992
rect 2928 808 2980 992
rect 3120 808 3172 992
rect 336 408 388 592
rect 528 408 580 592
rect 720 408 772 592
rect 912 408 964 592
rect 1104 408 1156 592
rect 1296 408 1348 592
rect 1488 408 1540 592
rect 1680 408 1732 592
rect 1872 408 1924 592
rect 2064 408 2116 592
rect 2256 408 2308 592
rect 2448 408 2500 592
rect 2640 408 2692 592
rect 2832 408 2884 592
rect 3024 408 3076 592
rect 240 188 292 372
rect 432 188 484 372
rect 624 188 676 372
rect 816 188 868 372
rect 1008 188 1060 372
rect 1200 188 1252 372
rect 1392 188 1444 372
rect 1584 188 1636 372
rect 1776 188 1828 372
rect 1968 188 2020 372
rect 2160 188 2212 372
rect 2352 188 2404 372
rect 2544 188 2596 372
rect 2736 188 2788 372
rect 2928 188 2980 372
rect 3120 188 3172 372
<< metal2 >>
rect 336 2448 3076 2540
rect 388 2272 528 2448
rect 336 2254 388 2264
rect 580 2272 720 2448
rect 528 2254 580 2264
rect 772 2272 912 2448
rect 720 2254 772 2264
rect 964 2272 1104 2448
rect 912 2254 964 2264
rect 1156 2272 1296 2448
rect 1104 2254 1156 2264
rect 1348 2272 1488 2448
rect 1296 2254 1348 2264
rect 1540 2272 1680 2448
rect 1488 2254 1540 2264
rect 1732 2272 1872 2448
rect 1680 2254 1732 2264
rect 1924 2272 2064 2448
rect 1872 2254 1924 2264
rect 2116 2272 2256 2448
rect 2064 2254 2116 2264
rect 2308 2272 2448 2448
rect 2256 2254 2308 2264
rect 2500 2272 2640 2448
rect 2448 2254 2500 2264
rect 2692 2272 2832 2448
rect 2640 2254 2692 2264
rect 2884 2272 3024 2448
rect 2832 2254 2884 2264
rect 3024 2254 3076 2264
rect 240 2228 292 2238
rect 236 2044 240 2220
rect 432 2228 484 2238
rect 292 2044 432 2220
rect 624 2228 676 2238
rect 484 2044 624 2220
rect 816 2228 868 2238
rect 676 2044 816 2220
rect 1008 2228 1060 2238
rect 868 2044 1008 2220
rect 1200 2228 1252 2238
rect 1060 2044 1200 2220
rect 1392 2228 1444 2238
rect 1252 2044 1392 2220
rect 1584 2228 1636 2238
rect 1444 2044 1584 2220
rect 1776 2228 1828 2238
rect 1636 2044 1776 2220
rect 1968 2228 2020 2238
rect 1828 2044 1968 2220
rect 2160 2228 2212 2238
rect 2020 2044 2160 2220
rect 2352 2228 2404 2238
rect 2212 2044 2352 2220
rect 2544 2228 2596 2238
rect 2404 2044 2544 2220
rect 2736 2228 2788 2238
rect 2596 2044 2736 2220
rect 2928 2228 2980 2238
rect 2788 2044 2928 2220
rect 3120 2228 3172 2238
rect 2980 2044 3120 2220
rect 3172 2044 3176 2220
rect 236 1952 3176 2044
rect 336 1828 3076 1920
rect 388 1652 528 1828
rect 336 1634 388 1644
rect 580 1652 720 1828
rect 528 1634 580 1644
rect 772 1652 912 1828
rect 720 1634 772 1644
rect 964 1652 1104 1828
rect 912 1634 964 1644
rect 1156 1652 1296 1828
rect 1104 1634 1156 1644
rect 1348 1652 1488 1828
rect 1296 1634 1348 1644
rect 1540 1652 1680 1828
rect 1488 1634 1540 1644
rect 1732 1652 1872 1828
rect 1680 1634 1732 1644
rect 1924 1652 2064 1828
rect 1872 1634 1924 1644
rect 2116 1652 2256 1828
rect 2064 1634 2116 1644
rect 2308 1652 2448 1828
rect 2256 1634 2308 1644
rect 2500 1652 2640 1828
rect 2448 1634 2500 1644
rect 2692 1652 2832 1828
rect 2640 1634 2692 1644
rect 2884 1652 3024 1828
rect 2832 1634 2884 1644
rect 3024 1634 3076 1644
rect 240 1608 292 1618
rect 432 1608 484 1618
rect 292 1424 432 1600
rect 624 1608 676 1618
rect 484 1424 624 1600
rect 816 1608 868 1618
rect 676 1424 816 1600
rect 1008 1608 1060 1618
rect 868 1424 1008 1600
rect 1200 1608 1252 1618
rect 1060 1424 1200 1600
rect 1392 1608 1444 1618
rect 1252 1424 1392 1600
rect 1584 1608 1636 1618
rect 1444 1424 1584 1600
rect 1776 1608 1828 1618
rect 1636 1424 1776 1600
rect 1968 1608 2020 1618
rect 1828 1424 1968 1600
rect 2160 1608 2212 1618
rect 2020 1424 2160 1600
rect 2352 1608 2404 1618
rect 2212 1424 2352 1600
rect 2544 1608 2596 1618
rect 2404 1424 2544 1600
rect 2736 1608 2788 1618
rect 2596 1424 2736 1600
rect 2928 1608 2980 1618
rect 2788 1424 2928 1600
rect 3120 1608 3172 1618
rect 2980 1424 3120 1600
rect 3172 1424 3180 1600
rect 240 1332 3180 1424
rect 336 1212 3076 1304
rect 388 1036 528 1212
rect 336 1018 388 1028
rect 580 1036 720 1212
rect 528 1018 580 1028
rect 772 1036 912 1212
rect 720 1018 772 1028
rect 964 1036 1104 1212
rect 912 1018 964 1028
rect 1156 1036 1296 1212
rect 1104 1018 1156 1028
rect 1348 1036 1488 1212
rect 1296 1018 1348 1028
rect 1540 1036 1680 1212
rect 1488 1018 1540 1028
rect 1732 1036 1872 1212
rect 1680 1018 1732 1028
rect 1924 1036 2064 1212
rect 1872 1018 1924 1028
rect 2116 1036 2256 1212
rect 2064 1018 2116 1028
rect 2308 1036 2448 1212
rect 2256 1018 2308 1028
rect 2500 1036 2640 1212
rect 2448 1018 2500 1028
rect 2692 1036 2832 1212
rect 2640 1018 2692 1028
rect 2884 1036 3024 1212
rect 2832 1018 2884 1028
rect 3024 1018 3076 1028
rect 240 992 292 1002
rect 432 992 484 1002
rect 292 808 432 988
rect 624 992 676 1002
rect 484 808 624 988
rect 816 992 868 1002
rect 676 808 816 988
rect 1008 992 1060 1002
rect 868 808 1008 988
rect 1200 992 1252 1002
rect 1060 808 1200 988
rect 1392 992 1444 1002
rect 1252 808 1392 988
rect 1584 992 1636 1002
rect 1444 808 1584 988
rect 1776 992 1828 1002
rect 1636 808 1776 988
rect 1968 992 2020 1002
rect 1828 808 1968 988
rect 2160 992 2212 1002
rect 2020 808 2160 988
rect 2352 992 2404 1002
rect 2212 808 2352 988
rect 2544 992 2596 1002
rect 2404 808 2544 988
rect 2736 992 2788 1002
rect 2596 808 2736 988
rect 2928 992 2980 1002
rect 2788 808 2928 988
rect 3120 992 3172 1002
rect 2980 808 3120 988
rect 3172 808 3180 988
rect 240 720 3180 808
rect 336 592 3076 684
rect 388 416 528 592
rect 336 398 388 408
rect 580 416 720 592
rect 528 398 580 408
rect 772 416 912 592
rect 720 398 772 408
rect 964 416 1104 592
rect 912 398 964 408
rect 1156 416 1296 592
rect 1104 398 1156 408
rect 1348 416 1488 592
rect 1296 398 1348 408
rect 1540 416 1680 592
rect 1488 398 1540 408
rect 1732 416 1872 592
rect 1680 398 1732 408
rect 1924 416 2064 592
rect 1872 398 1924 408
rect 2116 416 2256 592
rect 2064 398 2116 408
rect 2308 416 2448 592
rect 2256 398 2308 408
rect 2500 416 2640 592
rect 2448 398 2500 408
rect 2692 416 2832 592
rect 2640 398 2692 408
rect 2884 416 3024 592
rect 2832 398 2884 408
rect 3024 398 3076 408
rect 240 372 292 382
rect 432 372 484 382
rect 292 188 432 364
rect 624 372 676 382
rect 484 188 624 364
rect 816 372 868 382
rect 676 188 816 364
rect 1008 372 1060 382
rect 868 188 1008 364
rect 1200 372 1252 382
rect 1060 188 1200 364
rect 1392 372 1444 382
rect 1252 188 1392 364
rect 1584 372 1636 382
rect 1444 188 1584 364
rect 1776 372 1828 382
rect 1636 188 1776 364
rect 1968 372 2020 382
rect 1828 188 1968 364
rect 2160 372 2212 382
rect 2020 188 2160 364
rect 2352 372 2404 382
rect 2212 188 2352 364
rect 2544 372 2596 382
rect 2404 188 2544 364
rect 2736 372 2788 382
rect 2596 188 2736 364
rect 2928 372 2980 382
rect 2788 188 2928 364
rect 3120 372 3172 382
rect 2980 188 3120 364
rect 3172 188 3180 364
rect 240 96 3180 188
use outd_curm#0  outd_curm_0
timestamp 1685113734
transform 1 0 2020 0 1 -3176
box -40 916 1002 3158
use outd_curm#0  outd_curm_1
timestamp 1685113734
transform 1 0 3060 0 1 -3176
box -40 916 1002 3158
use outd_curm#0  outd_curm_4
timestamp 1685113734
transform 1 0 980 0 1 -3176
box -40 916 1002 3158
use outd_curm#0  outd_curm_5
timestamp 1685113734
transform 1 0 -60 0 1 -3176
box -40 916 1002 3158
use outd_curm#0  outd_curm_8
timestamp 1685113734
transform 1 0 980 0 1 -7656
box -40 916 1002 3158
use outd_curm#0  outd_curm_19
timestamp 1685113734
transform 1 0 2020 0 1 -7656
box -40 916 1002 3158
use outd_curm#0  outd_curm_21
timestamp 1685113734
transform 1 0 2020 0 1 -5416
box -40 916 1002 3158
use outd_curm#0  outd_curm_22
timestamp 1685113734
transform 1 0 980 0 1 -5416
box -40 916 1002 3158
use outd_curm#0  outd_curm_23
timestamp 1685113734
transform 1 0 -60 0 1 -5416
box -40 916 1002 3158
use outd_curm#0  outd_curm_25
timestamp 1685113734
transform 1 0 -60 0 1 -7656
box -40 916 1002 3158
use sky130_fd_pr__nfet_01v8_lvt_T6YALJ  sky130_fd_pr__nfet_01v8_lvt_T6YALJ_2
timestamp 1683809155
transform 1 0 1707 0 1 1317
box -1607 -1337 1607 1337
<< end >>
