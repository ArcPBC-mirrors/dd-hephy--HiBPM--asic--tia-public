magic
tech sky130A
magscale 1 2
timestamp 1684252655
<< psubdiff >>
rect 2840 810 3050 834
rect 2840 536 3050 560
<< psubdiffcont >>
rect 2840 560 3050 810
<< locali >>
rect 2380 6300 2520 6520
rect 1220 6160 1320 6300
rect 1200 4020 1300 4220
rect 2840 810 3050 826
rect 3050 560 3090 670
rect 2840 544 3090 560
rect 2900 360 3090 544
rect 2720 200 2840 360
rect 2980 250 3090 360
<< viali >>
rect 2840 200 2980 360
<< metal1 >>
rect 1412 8208 2456 8216
rect 1412 8132 2296 8208
rect 2436 8132 2456 8208
rect 1412 8116 2456 8132
rect 1366 7908 1376 8088
rect 1428 7908 1438 8088
rect 1558 7908 1568 8088
rect 1620 7908 1630 8088
rect 1750 7908 1760 8088
rect 1812 7908 1822 8088
rect 1942 7908 1952 8088
rect 2004 7908 2014 8088
rect 2134 7908 2144 8088
rect 2196 7908 2206 8088
rect 1270 7684 1280 7864
rect 1332 7684 1342 7864
rect 1462 7684 1472 7864
rect 1524 7684 1534 7864
rect 1654 7684 1664 7864
rect 1716 7684 1726 7864
rect 1846 7684 1856 7864
rect 1908 7684 1918 7864
rect 2038 7684 2048 7864
rect 2100 7684 2110 7864
rect 2230 7684 2240 7864
rect 2292 7684 2302 7864
rect 2336 7656 2456 8116
rect 2670 8048 2680 8148
rect 2860 8048 2870 8148
rect 1320 7500 2456 7656
rect 1366 7292 1376 7472
rect 1428 7292 1438 7472
rect 1558 7292 1568 7472
rect 1620 7292 1630 7472
rect 1750 7292 1760 7472
rect 1812 7292 1822 7472
rect 1942 7292 1952 7472
rect 2004 7292 2014 7472
rect 2134 7292 2144 7472
rect 2196 7292 2206 7472
rect 1270 7068 1280 7248
rect 1332 7068 1342 7248
rect 1462 7068 1472 7248
rect 1524 7068 1534 7248
rect 1654 7068 1664 7248
rect 1716 7068 1726 7248
rect 1846 7068 1856 7248
rect 1908 7068 1918 7248
rect 2038 7068 2048 7248
rect 2100 7068 2110 7248
rect 2230 7068 2240 7248
rect 2292 7068 2302 7248
rect 2336 7036 2456 7500
rect 1416 6880 2456 7036
rect 1366 6672 1376 6852
rect 1428 6672 1438 6852
rect 1558 6672 1568 6852
rect 1620 6672 1630 6852
rect 1750 6672 1760 6852
rect 1812 6672 1822 6852
rect 1942 6672 1952 6852
rect 2004 6672 2014 6852
rect 2134 6672 2144 6852
rect 2196 6672 2206 6852
rect 1270 6448 1280 6628
rect 1332 6448 1342 6628
rect 1462 6448 1472 6628
rect 1524 6448 1534 6628
rect 1654 6448 1664 6628
rect 1716 6448 1726 6628
rect 1846 6448 1856 6628
rect 1908 6448 1918 6628
rect 2038 6448 2048 6628
rect 2100 6448 2110 6628
rect 2230 6448 2240 6628
rect 2292 6448 2302 6628
rect 2336 6420 2456 6880
rect 2574 6680 2584 6892
rect 2660 6680 2670 6892
rect 2874 6684 2884 6896
rect 2960 6684 2970 6896
rect 1320 6320 2456 6420
rect 2670 6344 2680 6424
rect 2860 6344 2870 6424
rect 2338 5840 2348 6016
rect 2516 5840 2526 6016
rect 2834 360 2986 372
rect 2830 200 2840 360
rect 2980 200 2990 360
rect 2834 188 2986 200
<< via1 >>
rect 2296 8132 2436 8208
rect 1376 7908 1428 8088
rect 1568 7908 1620 8088
rect 1760 7908 1812 8088
rect 1952 7908 2004 8088
rect 2144 7908 2196 8088
rect 1280 7684 1332 7864
rect 1472 7684 1524 7864
rect 1664 7684 1716 7864
rect 1856 7684 1908 7864
rect 2048 7684 2100 7864
rect 2240 7684 2292 7864
rect 2680 8048 2860 8148
rect 1376 7292 1428 7472
rect 1568 7292 1620 7472
rect 1760 7292 1812 7472
rect 1952 7292 2004 7472
rect 2144 7292 2196 7472
rect 1280 7068 1332 7248
rect 1472 7068 1524 7248
rect 1664 7068 1716 7248
rect 1856 7068 1908 7248
rect 2048 7068 2100 7248
rect 2240 7068 2292 7248
rect 1376 6672 1428 6852
rect 1568 6672 1620 6852
rect 1760 6672 1812 6852
rect 1952 6672 2004 6852
rect 2144 6672 2196 6852
rect 1280 6448 1332 6628
rect 1472 6448 1524 6628
rect 1664 6448 1716 6628
rect 1856 6448 1908 6628
rect 2048 6448 2100 6628
rect 2240 6448 2292 6628
rect 2584 6680 2660 6892
rect 2884 6684 2960 6896
rect 2680 6344 2860 6424
rect 2348 5840 2516 6016
rect 2840 200 2980 360
<< metal2 >>
rect 1380 8212 1650 8460
rect 2296 8212 2436 8218
rect 1376 8208 2624 8212
rect 1376 8132 2296 8208
rect 2436 8132 2624 8208
rect 1376 8088 2624 8132
rect 1428 7912 1568 8088
rect 1376 7898 1428 7908
rect 1620 7912 1760 8088
rect 1568 7898 1620 7908
rect 1812 7912 1952 8088
rect 1760 7898 1812 7908
rect 2004 7912 2144 8088
rect 1952 7898 2004 7908
rect 2196 7912 2624 8088
rect 2680 8148 2860 8158
rect 2680 8038 2860 8048
rect 2144 7898 2196 7908
rect 1280 7864 1332 7874
rect 1472 7864 1524 7874
rect 1332 7704 1472 7860
rect 1664 7864 1716 7874
rect 1524 7704 1664 7860
rect 1856 7864 1908 7874
rect 1716 7704 1856 7860
rect 2048 7864 2100 7874
rect 1908 7704 2048 7860
rect 1332 7684 1372 7704
rect 2024 7684 2048 7704
rect 2240 7864 2292 7874
rect 2100 7684 2240 7860
rect 1280 7436 1372 7684
rect 2024 7472 2292 7684
rect 2024 7436 2144 7472
rect 1280 7300 1376 7436
rect 1428 7300 1568 7436
rect 1376 7282 1428 7292
rect 1620 7300 1760 7436
rect 1568 7282 1620 7292
rect 1812 7300 1952 7436
rect 1760 7282 1812 7292
rect 2004 7300 2144 7436
rect 1952 7282 2004 7292
rect 2196 7300 2292 7472
rect 2144 7282 2196 7292
rect 1280 7248 1332 7258
rect 1276 7068 1280 7244
rect 1472 7248 1524 7258
rect 1332 7068 1472 7244
rect 1664 7248 1716 7258
rect 1524 7068 1664 7244
rect 1856 7248 1908 7258
rect 1716 7068 1856 7244
rect 2048 7248 2100 7258
rect 1908 7068 2048 7244
rect 2240 7248 2292 7258
rect 2100 7068 2240 7244
rect 2344 7244 2624 7912
rect 2292 7068 2624 7244
rect 1276 6902 2624 7068
rect 1276 6892 2660 6902
rect 2884 6896 2960 6906
rect 1276 6852 2584 6892
rect 1276 6680 1376 6852
rect 1428 6680 1568 6852
rect 1376 6662 1428 6672
rect 1620 6680 1760 6852
rect 1568 6662 1620 6672
rect 1812 6680 1952 6852
rect 1760 6662 1812 6672
rect 2004 6680 2144 6852
rect 1952 6662 2004 6672
rect 2196 6680 2584 6852
rect 2660 6684 2884 6892
rect 2660 6680 2960 6684
rect 2144 6662 2196 6672
rect 2584 6670 2660 6680
rect 2884 6674 2960 6680
rect 1280 6628 1332 6638
rect 1472 6628 1524 6638
rect 1332 6592 1472 6624
rect 1664 6628 1716 6638
rect 1524 6592 1664 6624
rect 1856 6628 1908 6638
rect 1716 6592 1856 6624
rect 2048 6628 2100 6638
rect 1908 6592 2048 6624
rect 1332 6448 1372 6592
rect 2024 6448 2048 6592
rect 2240 6628 2292 6638
rect 2100 6448 2240 6624
rect 2292 6448 2320 6624
rect 1280 6360 1372 6448
rect 2024 6324 2320 6448
rect 2680 6428 2860 6434
rect 1372 6314 2320 6324
rect 2016 6108 2320 6314
rect 2620 6424 2880 6428
rect 2620 6344 2680 6424
rect 2860 6344 2880 6424
rect 2620 6108 2880 6344
rect 1368 6016 2880 6108
rect 1368 5840 2348 6016
rect 2516 5840 2880 6016
rect 2348 5830 2516 5840
rect 2840 360 2980 370
rect 2840 190 2980 200
<< via2 >>
rect 2680 8048 2860 8148
rect 1372 7684 1472 7704
rect 1472 7684 1524 7704
rect 1524 7684 1664 7704
rect 1664 7684 1716 7704
rect 1716 7684 1856 7704
rect 1856 7684 1908 7704
rect 1908 7684 2024 7704
rect 1372 7472 2024 7684
rect 1372 7436 1376 7472
rect 1376 7436 1428 7472
rect 1428 7436 1568 7472
rect 1568 7436 1620 7472
rect 1620 7436 1760 7472
rect 1760 7436 1812 7472
rect 1812 7436 1952 7472
rect 1952 7436 2004 7472
rect 2004 7436 2024 7472
rect 1372 6448 1472 6592
rect 1472 6448 1524 6592
rect 1524 6448 1664 6592
rect 1664 6448 1716 6592
rect 1716 6448 1856 6592
rect 1856 6448 1908 6592
rect 1908 6448 2024 6592
rect 1372 6324 2024 6448
rect 2840 200 2980 360
<< metal3 >>
rect 2680 8153 3248 8228
rect 2670 8148 3248 8153
rect 2670 8048 2680 8148
rect 2860 8048 3248 8148
rect 2670 8043 2870 8048
rect 1356 7704 2048 7728
rect 1356 7436 1372 7704
rect 2024 7436 2048 7704
rect 1356 6592 2048 7436
rect 1356 6324 1372 6592
rect 2024 6324 2048 6592
rect 1356 6296 2048 6324
rect 3180 4140 3348 4572
rect 2024 136 2624 860
rect 2830 360 2990 365
rect 2830 200 2840 360
rect 2980 200 2990 360
rect 2830 195 2990 200
rect 2014 -144 2024 136
rect 2624 -144 2634 136
<< via3 >>
rect 2840 200 2980 360
rect 2024 -144 2624 136
<< metal4 >>
rect 3264 4600 3432 4636
rect 3260 4060 3720 4600
rect 3264 4024 3432 4060
rect 2839 360 2981 361
rect 2839 200 2840 360
rect 2980 200 2981 360
rect 2839 199 2981 200
rect 2023 136 2625 137
rect 2840 136 2980 199
rect 3260 136 3720 392
rect 2023 -144 2024 136
rect 2624 -144 3720 136
rect 2023 -145 2625 -144
rect 3260 -148 3720 -144
use curr_m  curr_m_0
timestamp 1684252655
transform 1 0 1140 0 1 4560
box 0 -4400 1624 1656
use sky130_fd_pr__cap_mim_m3_1_BCLRNG  sky130_fd_pr__cap_mim_m3_1_BCLRNG_0
timestamp 1683624190
transform 1 0 5366 0 1 4340
box -2186 -4200 2186 4200
use sky130_fd_pr__nfet_01v8_lvt_L8NDKD  sky130_fd_pr__nfet_01v8_lvt_L8NDKD_0
timestamp 1683713379
transform 0 1 2770 -1 0 7236
box -996 -310 996 310
use sky130_fd_pr__nfet_01v8_lvt_R2KHEY  sky130_fd_pr__nfet_01v8_lvt_R2KHEY_1
timestamp 1684252655
transform 1 0 1787 0 1 7268
box -647 -1028 647 1028
<< labels >>
rlabel metal2 1390 8310 1630 8450 1 I_Bias1
port 1 n
rlabel metal3 3190 4310 3240 4410 1 Out
port 2 n
rlabel metal4 2760 -90 2960 30 1 Vn
port 3 n
<< end >>
