magic
tech sky130A
magscale 1 2
timestamp 1683553987
<< nwell >>
rect -957 -1055 957 1055
<< pmos >>
rect -761 436 -661 836
rect -603 436 -503 836
rect -445 436 -345 836
rect -287 436 -187 836
rect -129 436 -29 836
rect 29 436 129 836
rect 187 436 287 836
rect 345 436 445 836
rect 503 436 603 836
rect 661 436 761 836
rect -761 -200 -661 200
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
rect 661 -200 761 200
rect -761 -836 -661 -436
rect -603 -836 -503 -436
rect -445 -836 -345 -436
rect -287 -836 -187 -436
rect -129 -836 -29 -436
rect 29 -836 129 -436
rect 187 -836 287 -436
rect 345 -836 445 -436
rect 503 -836 603 -436
rect 661 -836 761 -436
<< pdiff >>
rect -819 824 -761 836
rect -819 448 -807 824
rect -773 448 -761 824
rect -819 436 -761 448
rect -661 824 -603 836
rect -661 448 -649 824
rect -615 448 -603 824
rect -661 436 -603 448
rect -503 824 -445 836
rect -503 448 -491 824
rect -457 448 -445 824
rect -503 436 -445 448
rect -345 824 -287 836
rect -345 448 -333 824
rect -299 448 -287 824
rect -345 436 -287 448
rect -187 824 -129 836
rect -187 448 -175 824
rect -141 448 -129 824
rect -187 436 -129 448
rect -29 824 29 836
rect -29 448 -17 824
rect 17 448 29 824
rect -29 436 29 448
rect 129 824 187 836
rect 129 448 141 824
rect 175 448 187 824
rect 129 436 187 448
rect 287 824 345 836
rect 287 448 299 824
rect 333 448 345 824
rect 287 436 345 448
rect 445 824 503 836
rect 445 448 457 824
rect 491 448 503 824
rect 445 436 503 448
rect 603 824 661 836
rect 603 448 615 824
rect 649 448 661 824
rect 603 436 661 448
rect 761 824 819 836
rect 761 448 773 824
rect 807 448 819 824
rect 761 436 819 448
rect -819 188 -761 200
rect -819 -188 -807 188
rect -773 -188 -761 188
rect -819 -200 -761 -188
rect -661 188 -603 200
rect -661 -188 -649 188
rect -615 -188 -603 188
rect -661 -200 -603 -188
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
rect 603 188 661 200
rect 603 -188 615 188
rect 649 -188 661 188
rect 603 -200 661 -188
rect 761 188 819 200
rect 761 -188 773 188
rect 807 -188 819 188
rect 761 -200 819 -188
rect -819 -448 -761 -436
rect -819 -824 -807 -448
rect -773 -824 -761 -448
rect -819 -836 -761 -824
rect -661 -448 -603 -436
rect -661 -824 -649 -448
rect -615 -824 -603 -448
rect -661 -836 -603 -824
rect -503 -448 -445 -436
rect -503 -824 -491 -448
rect -457 -824 -445 -448
rect -503 -836 -445 -824
rect -345 -448 -287 -436
rect -345 -824 -333 -448
rect -299 -824 -287 -448
rect -345 -836 -287 -824
rect -187 -448 -129 -436
rect -187 -824 -175 -448
rect -141 -824 -129 -448
rect -187 -836 -129 -824
rect -29 -448 29 -436
rect -29 -824 -17 -448
rect 17 -824 29 -448
rect -29 -836 29 -824
rect 129 -448 187 -436
rect 129 -824 141 -448
rect 175 -824 187 -448
rect 129 -836 187 -824
rect 287 -448 345 -436
rect 287 -824 299 -448
rect 333 -824 345 -448
rect 287 -836 345 -824
rect 445 -448 503 -436
rect 445 -824 457 -448
rect 491 -824 503 -448
rect 445 -836 503 -824
rect 603 -448 661 -436
rect 603 -824 615 -448
rect 649 -824 661 -448
rect 603 -836 661 -824
rect 761 -448 819 -436
rect 761 -824 773 -448
rect 807 -824 819 -448
rect 761 -836 819 -824
<< pdiffc >>
rect -807 448 -773 824
rect -649 448 -615 824
rect -491 448 -457 824
rect -333 448 -299 824
rect -175 448 -141 824
rect -17 448 17 824
rect 141 448 175 824
rect 299 448 333 824
rect 457 448 491 824
rect 615 448 649 824
rect 773 448 807 824
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect -807 -824 -773 -448
rect -649 -824 -615 -448
rect -491 -824 -457 -448
rect -333 -824 -299 -448
rect -175 -824 -141 -448
rect -17 -824 17 -448
rect 141 -824 175 -448
rect 299 -824 333 -448
rect 457 -824 491 -448
rect 615 -824 649 -448
rect 773 -824 807 -448
<< nsubdiff >>
rect -921 985 -825 1019
rect 825 985 921 1019
rect -921 923 -887 985
rect 887 923 921 985
rect -921 -985 -887 -923
rect 887 -985 921 -923
rect -921 -1019 -825 -985
rect 825 -1019 921 -985
<< nsubdiffcont >>
rect -825 985 825 1019
rect -921 -923 -887 923
rect 887 -923 921 923
rect -825 -1019 825 -985
<< poly >>
rect -761 917 -661 933
rect -761 883 -745 917
rect -677 883 -661 917
rect -761 836 -661 883
rect -603 917 -503 933
rect -603 883 -587 917
rect -519 883 -503 917
rect -603 836 -503 883
rect -445 917 -345 933
rect -445 883 -429 917
rect -361 883 -345 917
rect -445 836 -345 883
rect -287 917 -187 933
rect -287 883 -271 917
rect -203 883 -187 917
rect -287 836 -187 883
rect -129 917 -29 933
rect -129 883 -113 917
rect -45 883 -29 917
rect -129 836 -29 883
rect 29 917 129 933
rect 29 883 45 917
rect 113 883 129 917
rect 29 836 129 883
rect 187 917 287 933
rect 187 883 203 917
rect 271 883 287 917
rect 187 836 287 883
rect 345 917 445 933
rect 345 883 361 917
rect 429 883 445 917
rect 345 836 445 883
rect 503 917 603 933
rect 503 883 519 917
rect 587 883 603 917
rect 503 836 603 883
rect 661 917 761 933
rect 661 883 677 917
rect 745 883 761 917
rect 661 836 761 883
rect -761 389 -661 436
rect -761 355 -745 389
rect -677 355 -661 389
rect -761 339 -661 355
rect -603 389 -503 436
rect -603 355 -587 389
rect -519 355 -503 389
rect -603 339 -503 355
rect -445 389 -345 436
rect -445 355 -429 389
rect -361 355 -345 389
rect -445 339 -345 355
rect -287 389 -187 436
rect -287 355 -271 389
rect -203 355 -187 389
rect -287 339 -187 355
rect -129 389 -29 436
rect -129 355 -113 389
rect -45 355 -29 389
rect -129 339 -29 355
rect 29 389 129 436
rect 29 355 45 389
rect 113 355 129 389
rect 29 339 129 355
rect 187 389 287 436
rect 187 355 203 389
rect 271 355 287 389
rect 187 339 287 355
rect 345 389 445 436
rect 345 355 361 389
rect 429 355 445 389
rect 345 339 445 355
rect 503 389 603 436
rect 503 355 519 389
rect 587 355 603 389
rect 503 339 603 355
rect 661 389 761 436
rect 661 355 677 389
rect 745 355 761 389
rect 661 339 761 355
rect -761 281 -661 297
rect -761 247 -745 281
rect -677 247 -661 281
rect -761 200 -661 247
rect -603 281 -503 297
rect -603 247 -587 281
rect -519 247 -503 281
rect -603 200 -503 247
rect -445 281 -345 297
rect -445 247 -429 281
rect -361 247 -345 281
rect -445 200 -345 247
rect -287 281 -187 297
rect -287 247 -271 281
rect -203 247 -187 281
rect -287 200 -187 247
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect 187 281 287 297
rect 187 247 203 281
rect 271 247 287 281
rect 187 200 287 247
rect 345 281 445 297
rect 345 247 361 281
rect 429 247 445 281
rect 345 200 445 247
rect 503 281 603 297
rect 503 247 519 281
rect 587 247 603 281
rect 503 200 603 247
rect 661 281 761 297
rect 661 247 677 281
rect 745 247 761 281
rect 661 200 761 247
rect -761 -247 -661 -200
rect -761 -281 -745 -247
rect -677 -281 -661 -247
rect -761 -297 -661 -281
rect -603 -247 -503 -200
rect -603 -281 -587 -247
rect -519 -281 -503 -247
rect -603 -297 -503 -281
rect -445 -247 -345 -200
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -445 -297 -345 -281
rect -287 -247 -187 -200
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -287 -297 -187 -281
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
rect 187 -247 287 -200
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 187 -297 287 -281
rect 345 -247 445 -200
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 345 -297 445 -281
rect 503 -247 603 -200
rect 503 -281 519 -247
rect 587 -281 603 -247
rect 503 -297 603 -281
rect 661 -247 761 -200
rect 661 -281 677 -247
rect 745 -281 761 -247
rect 661 -297 761 -281
rect -761 -355 -661 -339
rect -761 -389 -745 -355
rect -677 -389 -661 -355
rect -761 -436 -661 -389
rect -603 -355 -503 -339
rect -603 -389 -587 -355
rect -519 -389 -503 -355
rect -603 -436 -503 -389
rect -445 -355 -345 -339
rect -445 -389 -429 -355
rect -361 -389 -345 -355
rect -445 -436 -345 -389
rect -287 -355 -187 -339
rect -287 -389 -271 -355
rect -203 -389 -187 -355
rect -287 -436 -187 -389
rect -129 -355 -29 -339
rect -129 -389 -113 -355
rect -45 -389 -29 -355
rect -129 -436 -29 -389
rect 29 -355 129 -339
rect 29 -389 45 -355
rect 113 -389 129 -355
rect 29 -436 129 -389
rect 187 -355 287 -339
rect 187 -389 203 -355
rect 271 -389 287 -355
rect 187 -436 287 -389
rect 345 -355 445 -339
rect 345 -389 361 -355
rect 429 -389 445 -355
rect 345 -436 445 -389
rect 503 -355 603 -339
rect 503 -389 519 -355
rect 587 -389 603 -355
rect 503 -436 603 -389
rect 661 -355 761 -339
rect 661 -389 677 -355
rect 745 -389 761 -355
rect 661 -436 761 -389
rect -761 -883 -661 -836
rect -761 -917 -745 -883
rect -677 -917 -661 -883
rect -761 -933 -661 -917
rect -603 -883 -503 -836
rect -603 -917 -587 -883
rect -519 -917 -503 -883
rect -603 -933 -503 -917
rect -445 -883 -345 -836
rect -445 -917 -429 -883
rect -361 -917 -345 -883
rect -445 -933 -345 -917
rect -287 -883 -187 -836
rect -287 -917 -271 -883
rect -203 -917 -187 -883
rect -287 -933 -187 -917
rect -129 -883 -29 -836
rect -129 -917 -113 -883
rect -45 -917 -29 -883
rect -129 -933 -29 -917
rect 29 -883 129 -836
rect 29 -917 45 -883
rect 113 -917 129 -883
rect 29 -933 129 -917
rect 187 -883 287 -836
rect 187 -917 203 -883
rect 271 -917 287 -883
rect 187 -933 287 -917
rect 345 -883 445 -836
rect 345 -917 361 -883
rect 429 -917 445 -883
rect 345 -933 445 -917
rect 503 -883 603 -836
rect 503 -917 519 -883
rect 587 -917 603 -883
rect 503 -933 603 -917
rect 661 -883 761 -836
rect 661 -917 677 -883
rect 745 -917 761 -883
rect 661 -933 761 -917
<< polycont >>
rect -745 883 -677 917
rect -587 883 -519 917
rect -429 883 -361 917
rect -271 883 -203 917
rect -113 883 -45 917
rect 45 883 113 917
rect 203 883 271 917
rect 361 883 429 917
rect 519 883 587 917
rect 677 883 745 917
rect -745 355 -677 389
rect -587 355 -519 389
rect -429 355 -361 389
rect -271 355 -203 389
rect -113 355 -45 389
rect 45 355 113 389
rect 203 355 271 389
rect 361 355 429 389
rect 519 355 587 389
rect 677 355 745 389
rect -745 247 -677 281
rect -587 247 -519 281
rect -429 247 -361 281
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect 361 247 429 281
rect 519 247 587 281
rect 677 247 745 281
rect -745 -281 -677 -247
rect -587 -281 -519 -247
rect -429 -281 -361 -247
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
rect 361 -281 429 -247
rect 519 -281 587 -247
rect 677 -281 745 -247
rect -745 -389 -677 -355
rect -587 -389 -519 -355
rect -429 -389 -361 -355
rect -271 -389 -203 -355
rect -113 -389 -45 -355
rect 45 -389 113 -355
rect 203 -389 271 -355
rect 361 -389 429 -355
rect 519 -389 587 -355
rect 677 -389 745 -355
rect -745 -917 -677 -883
rect -587 -917 -519 -883
rect -429 -917 -361 -883
rect -271 -917 -203 -883
rect -113 -917 -45 -883
rect 45 -917 113 -883
rect 203 -917 271 -883
rect 361 -917 429 -883
rect 519 -917 587 -883
rect 677 -917 745 -883
<< locali >>
rect -921 985 -825 1019
rect 825 985 921 1019
rect -921 923 -887 985
rect 887 923 921 985
rect -761 883 -745 917
rect -677 883 -661 917
rect -603 883 -587 917
rect -519 883 -503 917
rect -445 883 -429 917
rect -361 883 -345 917
rect -287 883 -271 917
rect -203 883 -187 917
rect -129 883 -113 917
rect -45 883 -29 917
rect 29 883 45 917
rect 113 883 129 917
rect 187 883 203 917
rect 271 883 287 917
rect 345 883 361 917
rect 429 883 445 917
rect 503 883 519 917
rect 587 883 603 917
rect 661 883 677 917
rect 745 883 761 917
rect -807 824 -773 840
rect -807 432 -773 448
rect -649 824 -615 840
rect -649 432 -615 448
rect -491 824 -457 840
rect -491 432 -457 448
rect -333 824 -299 840
rect -333 432 -299 448
rect -175 824 -141 840
rect -175 432 -141 448
rect -17 824 17 840
rect -17 432 17 448
rect 141 824 175 840
rect 141 432 175 448
rect 299 824 333 840
rect 299 432 333 448
rect 457 824 491 840
rect 457 432 491 448
rect 615 824 649 840
rect 615 432 649 448
rect 773 824 807 840
rect 773 432 807 448
rect -761 355 -745 389
rect -677 355 -661 389
rect -603 355 -587 389
rect -519 355 -503 389
rect -445 355 -429 389
rect -361 355 -345 389
rect -287 355 -271 389
rect -203 355 -187 389
rect -129 355 -113 389
rect -45 355 -29 389
rect 29 355 45 389
rect 113 355 129 389
rect 187 355 203 389
rect 271 355 287 389
rect 345 355 361 389
rect 429 355 445 389
rect 503 355 519 389
rect 587 355 603 389
rect 661 355 677 389
rect 745 355 761 389
rect -761 247 -745 281
rect -677 247 -661 281
rect -603 247 -587 281
rect -519 247 -503 281
rect -445 247 -429 281
rect -361 247 -345 281
rect -287 247 -271 281
rect -203 247 -187 281
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect 187 247 203 281
rect 271 247 287 281
rect 345 247 361 281
rect 429 247 445 281
rect 503 247 519 281
rect 587 247 603 281
rect 661 247 677 281
rect 745 247 761 281
rect -807 188 -773 204
rect -807 -204 -773 -188
rect -649 188 -615 204
rect -649 -204 -615 -188
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect 615 188 649 204
rect 615 -204 649 -188
rect 773 188 807 204
rect 773 -204 807 -188
rect -761 -281 -745 -247
rect -677 -281 -661 -247
rect -603 -281 -587 -247
rect -519 -281 -503 -247
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 503 -281 519 -247
rect 587 -281 603 -247
rect 661 -281 677 -247
rect 745 -281 761 -247
rect -761 -389 -745 -355
rect -677 -389 -661 -355
rect -603 -389 -587 -355
rect -519 -389 -503 -355
rect -445 -389 -429 -355
rect -361 -389 -345 -355
rect -287 -389 -271 -355
rect -203 -389 -187 -355
rect -129 -389 -113 -355
rect -45 -389 -29 -355
rect 29 -389 45 -355
rect 113 -389 129 -355
rect 187 -389 203 -355
rect 271 -389 287 -355
rect 345 -389 361 -355
rect 429 -389 445 -355
rect 503 -389 519 -355
rect 587 -389 603 -355
rect 661 -389 677 -355
rect 745 -389 761 -355
rect -807 -448 -773 -432
rect -807 -840 -773 -824
rect -649 -448 -615 -432
rect -649 -840 -615 -824
rect -491 -448 -457 -432
rect -491 -840 -457 -824
rect -333 -448 -299 -432
rect -333 -840 -299 -824
rect -175 -448 -141 -432
rect -175 -840 -141 -824
rect -17 -448 17 -432
rect -17 -840 17 -824
rect 141 -448 175 -432
rect 141 -840 175 -824
rect 299 -448 333 -432
rect 299 -840 333 -824
rect 457 -448 491 -432
rect 457 -840 491 -824
rect 615 -448 649 -432
rect 615 -840 649 -824
rect 773 -448 807 -432
rect 773 -840 807 -824
rect -761 -917 -745 -883
rect -677 -917 -661 -883
rect -603 -917 -587 -883
rect -519 -917 -503 -883
rect -445 -917 -429 -883
rect -361 -917 -345 -883
rect -287 -917 -271 -883
rect -203 -917 -187 -883
rect -129 -917 -113 -883
rect -45 -917 -29 -883
rect 29 -917 45 -883
rect 113 -917 129 -883
rect 187 -917 203 -883
rect 271 -917 287 -883
rect 345 -917 361 -883
rect 429 -917 445 -883
rect 503 -917 519 -883
rect 587 -917 603 -883
rect 661 -917 677 -883
rect 745 -917 761 -883
rect -921 -985 -887 -923
rect 887 -985 921 -923
rect -921 -1019 -825 -985
rect 825 -1019 921 -985
<< viali >>
rect -745 883 -677 917
rect -587 883 -519 917
rect -429 883 -361 917
rect -271 883 -203 917
rect -113 883 -45 917
rect 45 883 113 917
rect 203 883 271 917
rect 361 883 429 917
rect 519 883 587 917
rect 677 883 745 917
rect -807 448 -773 824
rect -649 448 -615 824
rect -491 448 -457 824
rect -333 448 -299 824
rect -175 448 -141 824
rect -17 448 17 824
rect 141 448 175 824
rect 299 448 333 824
rect 457 448 491 824
rect 615 448 649 824
rect 773 448 807 824
rect -745 355 -677 389
rect -587 355 -519 389
rect -429 355 -361 389
rect -271 355 -203 389
rect -113 355 -45 389
rect 45 355 113 389
rect 203 355 271 389
rect 361 355 429 389
rect 519 355 587 389
rect 677 355 745 389
rect -745 247 -677 281
rect -587 247 -519 281
rect -429 247 -361 281
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect 361 247 429 281
rect 519 247 587 281
rect 677 247 745 281
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect -745 -281 -677 -247
rect -587 -281 -519 -247
rect -429 -281 -361 -247
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
rect 361 -281 429 -247
rect 519 -281 587 -247
rect 677 -281 745 -247
rect -745 -389 -677 -355
rect -587 -389 -519 -355
rect -429 -389 -361 -355
rect -271 -389 -203 -355
rect -113 -389 -45 -355
rect 45 -389 113 -355
rect 203 -389 271 -355
rect 361 -389 429 -355
rect 519 -389 587 -355
rect 677 -389 745 -355
rect -807 -824 -773 -448
rect -649 -824 -615 -448
rect -491 -824 -457 -448
rect -333 -824 -299 -448
rect -175 -824 -141 -448
rect -17 -824 17 -448
rect 141 -824 175 -448
rect 299 -824 333 -448
rect 457 -824 491 -448
rect 615 -824 649 -448
rect 773 -824 807 -448
rect -745 -917 -677 -883
rect -587 -917 -519 -883
rect -429 -917 -361 -883
rect -271 -917 -203 -883
rect -113 -917 -45 -883
rect 45 -917 113 -883
rect 203 -917 271 -883
rect 361 -917 429 -883
rect 519 -917 587 -883
rect 677 -917 745 -883
<< metal1 >>
rect -757 917 -665 923
rect -757 883 -745 917
rect -677 883 -665 917
rect -757 877 -665 883
rect -599 917 -507 923
rect -599 883 -587 917
rect -519 883 -507 917
rect -599 877 -507 883
rect -441 917 -349 923
rect -441 883 -429 917
rect -361 883 -349 917
rect -441 877 -349 883
rect -283 917 -191 923
rect -283 883 -271 917
rect -203 883 -191 917
rect -283 877 -191 883
rect -125 917 -33 923
rect -125 883 -113 917
rect -45 883 -33 917
rect -125 877 -33 883
rect 33 917 125 923
rect 33 883 45 917
rect 113 883 125 917
rect 33 877 125 883
rect 191 917 283 923
rect 191 883 203 917
rect 271 883 283 917
rect 191 877 283 883
rect 349 917 441 923
rect 349 883 361 917
rect 429 883 441 917
rect 349 877 441 883
rect 507 917 599 923
rect 507 883 519 917
rect 587 883 599 917
rect 507 877 599 883
rect 665 917 757 923
rect 665 883 677 917
rect 745 883 757 917
rect 665 877 757 883
rect -813 824 -767 836
rect -813 448 -807 824
rect -773 448 -767 824
rect -813 436 -767 448
rect -655 824 -609 836
rect -655 448 -649 824
rect -615 448 -609 824
rect -655 436 -609 448
rect -497 824 -451 836
rect -497 448 -491 824
rect -457 448 -451 824
rect -497 436 -451 448
rect -339 824 -293 836
rect -339 448 -333 824
rect -299 448 -293 824
rect -339 436 -293 448
rect -181 824 -135 836
rect -181 448 -175 824
rect -141 448 -135 824
rect -181 436 -135 448
rect -23 824 23 836
rect -23 448 -17 824
rect 17 448 23 824
rect -23 436 23 448
rect 135 824 181 836
rect 135 448 141 824
rect 175 448 181 824
rect 135 436 181 448
rect 293 824 339 836
rect 293 448 299 824
rect 333 448 339 824
rect 293 436 339 448
rect 451 824 497 836
rect 451 448 457 824
rect 491 448 497 824
rect 451 436 497 448
rect 609 824 655 836
rect 609 448 615 824
rect 649 448 655 824
rect 609 436 655 448
rect 767 824 813 836
rect 767 448 773 824
rect 807 448 813 824
rect 767 436 813 448
rect -757 389 -665 395
rect -757 355 -745 389
rect -677 355 -665 389
rect -757 349 -665 355
rect -599 389 -507 395
rect -599 355 -587 389
rect -519 355 -507 389
rect -599 349 -507 355
rect -441 389 -349 395
rect -441 355 -429 389
rect -361 355 -349 389
rect -441 349 -349 355
rect -283 389 -191 395
rect -283 355 -271 389
rect -203 355 -191 389
rect -283 349 -191 355
rect -125 389 -33 395
rect -125 355 -113 389
rect -45 355 -33 389
rect -125 349 -33 355
rect 33 389 125 395
rect 33 355 45 389
rect 113 355 125 389
rect 33 349 125 355
rect 191 389 283 395
rect 191 355 203 389
rect 271 355 283 389
rect 191 349 283 355
rect 349 389 441 395
rect 349 355 361 389
rect 429 355 441 389
rect 349 349 441 355
rect 507 389 599 395
rect 507 355 519 389
rect 587 355 599 389
rect 507 349 599 355
rect 665 389 757 395
rect 665 355 677 389
rect 745 355 757 389
rect 665 349 757 355
rect -757 281 -665 287
rect -757 247 -745 281
rect -677 247 -665 281
rect -757 241 -665 247
rect -599 281 -507 287
rect -599 247 -587 281
rect -519 247 -507 281
rect -599 241 -507 247
rect -441 281 -349 287
rect -441 247 -429 281
rect -361 247 -349 281
rect -441 241 -349 247
rect -283 281 -191 287
rect -283 247 -271 281
rect -203 247 -191 281
rect -283 241 -191 247
rect -125 281 -33 287
rect -125 247 -113 281
rect -45 247 -33 281
rect -125 241 -33 247
rect 33 281 125 287
rect 33 247 45 281
rect 113 247 125 281
rect 33 241 125 247
rect 191 281 283 287
rect 191 247 203 281
rect 271 247 283 281
rect 191 241 283 247
rect 349 281 441 287
rect 349 247 361 281
rect 429 247 441 281
rect 349 241 441 247
rect 507 281 599 287
rect 507 247 519 281
rect 587 247 599 281
rect 507 241 599 247
rect 665 281 757 287
rect 665 247 677 281
rect 745 247 757 281
rect 665 241 757 247
rect -813 188 -767 200
rect -813 -188 -807 188
rect -773 -188 -767 188
rect -813 -200 -767 -188
rect -655 188 -609 200
rect -655 -188 -649 188
rect -615 -188 -609 188
rect -655 -200 -609 -188
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect 609 188 655 200
rect 609 -188 615 188
rect 649 -188 655 188
rect 609 -200 655 -188
rect 767 188 813 200
rect 767 -188 773 188
rect 807 -188 813 188
rect 767 -200 813 -188
rect -757 -247 -665 -241
rect -757 -281 -745 -247
rect -677 -281 -665 -247
rect -757 -287 -665 -281
rect -599 -247 -507 -241
rect -599 -281 -587 -247
rect -519 -281 -507 -247
rect -599 -287 -507 -281
rect -441 -247 -349 -241
rect -441 -281 -429 -247
rect -361 -281 -349 -247
rect -441 -287 -349 -281
rect -283 -247 -191 -241
rect -283 -281 -271 -247
rect -203 -281 -191 -247
rect -283 -287 -191 -281
rect -125 -247 -33 -241
rect -125 -281 -113 -247
rect -45 -281 -33 -247
rect -125 -287 -33 -281
rect 33 -247 125 -241
rect 33 -281 45 -247
rect 113 -281 125 -247
rect 33 -287 125 -281
rect 191 -247 283 -241
rect 191 -281 203 -247
rect 271 -281 283 -247
rect 191 -287 283 -281
rect 349 -247 441 -241
rect 349 -281 361 -247
rect 429 -281 441 -247
rect 349 -287 441 -281
rect 507 -247 599 -241
rect 507 -281 519 -247
rect 587 -281 599 -247
rect 507 -287 599 -281
rect 665 -247 757 -241
rect 665 -281 677 -247
rect 745 -281 757 -247
rect 665 -287 757 -281
rect -757 -355 -665 -349
rect -757 -389 -745 -355
rect -677 -389 -665 -355
rect -757 -395 -665 -389
rect -599 -355 -507 -349
rect -599 -389 -587 -355
rect -519 -389 -507 -355
rect -599 -395 -507 -389
rect -441 -355 -349 -349
rect -441 -389 -429 -355
rect -361 -389 -349 -355
rect -441 -395 -349 -389
rect -283 -355 -191 -349
rect -283 -389 -271 -355
rect -203 -389 -191 -355
rect -283 -395 -191 -389
rect -125 -355 -33 -349
rect -125 -389 -113 -355
rect -45 -389 -33 -355
rect -125 -395 -33 -389
rect 33 -355 125 -349
rect 33 -389 45 -355
rect 113 -389 125 -355
rect 33 -395 125 -389
rect 191 -355 283 -349
rect 191 -389 203 -355
rect 271 -389 283 -355
rect 191 -395 283 -389
rect 349 -355 441 -349
rect 349 -389 361 -355
rect 429 -389 441 -355
rect 349 -395 441 -389
rect 507 -355 599 -349
rect 507 -389 519 -355
rect 587 -389 599 -355
rect 507 -395 599 -389
rect 665 -355 757 -349
rect 665 -389 677 -355
rect 745 -389 757 -355
rect 665 -395 757 -389
rect -813 -448 -767 -436
rect -813 -824 -807 -448
rect -773 -824 -767 -448
rect -813 -836 -767 -824
rect -655 -448 -609 -436
rect -655 -824 -649 -448
rect -615 -824 -609 -448
rect -655 -836 -609 -824
rect -497 -448 -451 -436
rect -497 -824 -491 -448
rect -457 -824 -451 -448
rect -497 -836 -451 -824
rect -339 -448 -293 -436
rect -339 -824 -333 -448
rect -299 -824 -293 -448
rect -339 -836 -293 -824
rect -181 -448 -135 -436
rect -181 -824 -175 -448
rect -141 -824 -135 -448
rect -181 -836 -135 -824
rect -23 -448 23 -436
rect -23 -824 -17 -448
rect 17 -824 23 -448
rect -23 -836 23 -824
rect 135 -448 181 -436
rect 135 -824 141 -448
rect 175 -824 181 -448
rect 135 -836 181 -824
rect 293 -448 339 -436
rect 293 -824 299 -448
rect 333 -824 339 -448
rect 293 -836 339 -824
rect 451 -448 497 -436
rect 451 -824 457 -448
rect 491 -824 497 -448
rect 451 -836 497 -824
rect 609 -448 655 -436
rect 609 -824 615 -448
rect 649 -824 655 -448
rect 609 -836 655 -824
rect 767 -448 813 -436
rect 767 -824 773 -448
rect 807 -824 813 -448
rect 767 -836 813 -824
rect -757 -883 -665 -877
rect -757 -917 -745 -883
rect -677 -917 -665 -883
rect -757 -923 -665 -917
rect -599 -883 -507 -877
rect -599 -917 -587 -883
rect -519 -917 -507 -883
rect -599 -923 -507 -917
rect -441 -883 -349 -877
rect -441 -917 -429 -883
rect -361 -917 -349 -883
rect -441 -923 -349 -917
rect -283 -883 -191 -877
rect -283 -917 -271 -883
rect -203 -917 -191 -883
rect -283 -923 -191 -917
rect -125 -883 -33 -877
rect -125 -917 -113 -883
rect -45 -917 -33 -883
rect -125 -923 -33 -917
rect 33 -883 125 -877
rect 33 -917 45 -883
rect 113 -917 125 -883
rect 33 -923 125 -917
rect 191 -883 283 -877
rect 191 -917 203 -883
rect 271 -917 283 -883
rect 191 -923 283 -917
rect 349 -883 441 -877
rect 349 -917 361 -883
rect 429 -917 441 -883
rect 349 -923 441 -917
rect 507 -883 599 -877
rect 507 -917 519 -883
rect 587 -917 599 -883
rect 507 -923 599 -917
rect 665 -883 757 -877
rect 665 -917 677 -883
rect 745 -917 757 -883
rect 665 -923 757 -917
<< properties >>
string FIXED_BBOX -904 -1002 904 1002
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.5 m 3 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
