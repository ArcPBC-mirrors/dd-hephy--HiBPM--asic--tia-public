magic
tech sky130A
magscale 1 2
timestamp 1685108691
<< metal3 >>
rect -1686 7832 1686 7860
rect -1686 2808 1602 7832
rect 1666 2808 1686 7832
rect -1686 2780 1686 2808
rect -1686 2512 1686 2540
rect -1686 -2512 1602 2512
rect 1666 -2512 1686 2512
rect -1686 -2540 1686 -2512
rect -1686 -2808 1686 -2780
rect -1686 -7832 1602 -2808
rect 1666 -7832 1686 -2808
rect -1686 -7860 1686 -7832
<< via3 >>
rect 1602 2808 1666 7832
rect 1602 -2512 1666 2512
rect 1602 -7832 1666 -2808
<< mimcap >>
rect -1646 7780 1354 7820
rect -1646 2860 -1606 7780
rect 1314 2860 1354 7780
rect -1646 2820 1354 2860
rect -1646 2460 1354 2500
rect -1646 -2460 -1606 2460
rect 1314 -2460 1354 2460
rect -1646 -2500 1354 -2460
rect -1646 -2860 1354 -2820
rect -1646 -7780 -1606 -2860
rect 1314 -7780 1354 -2860
rect -1646 -7820 1354 -7780
<< mimcapcontact >>
rect -1606 2860 1314 7780
rect -1606 -2460 1314 2460
rect -1606 -7780 1314 -2860
<< metal4 >>
rect -198 7781 -94 7980
rect 1582 7832 1686 7980
rect -1607 7780 1315 7781
rect -1607 2860 -1606 7780
rect 1314 2860 1315 7780
rect -1607 2859 1315 2860
rect -198 2461 -94 2859
rect 1582 2808 1602 7832
rect 1666 2808 1686 7832
rect 1582 2512 1686 2808
rect -1607 2460 1315 2461
rect -1607 -2460 -1606 2460
rect 1314 -2460 1315 2460
rect -1607 -2461 1315 -2460
rect -198 -2859 -94 -2461
rect 1582 -2512 1602 2512
rect 1666 -2512 1686 2512
rect 1582 -2808 1686 -2512
rect -1607 -2860 1315 -2859
rect -1607 -7780 -1606 -2860
rect 1314 -7780 1315 -2860
rect -1607 -7781 1315 -7780
rect -198 -7980 -94 -7781
rect 1582 -7832 1602 -2808
rect 1666 -7832 1686 -2808
rect 1582 -7980 1686 -7832
<< properties >>
string FIXED_BBOX -1686 2780 1394 7860
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15 l 25 val 765.2 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
