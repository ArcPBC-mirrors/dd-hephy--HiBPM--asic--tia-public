magic
tech sky130A
timestamp 1689606798
<< metal4 >>
rect -200 2300 800 2500
rect 3800 2300 4800 2500
rect -200 -1700 800 -1500
rect 3800 -1700 4800 -1500
<< via4 >>
rect -800 2500 -600 2900
rect -1200 2300 -200 2500
rect -800 1900 -600 2300
rect 800 1900 1800 2900
rect 2800 1900 3800 2900
rect 5200 2500 5400 2900
rect 4800 2300 5800 2500
rect 5200 1900 5400 2300
rect -600 -100 400 900
rect 4200 -100 5200 900
rect -1600 -1300 -200 -1100
rect -1600 -2300 -1400 -1300
rect -400 -2300 -200 -1300
rect 800 -2100 1800 -1100
rect 2800 -2100 3800 -1100
rect 5200 -1500 5400 -1100
rect 4800 -1700 5800 -1500
rect 5200 -2100 5400 -1700
rect -1600 -2500 -200 -2300
<< metal5 >>
rect -812 2900 -588 2912
rect -812 2512 -800 2900
rect -1212 2500 -800 2512
rect -600 2512 -588 2900
rect 788 2900 1812 2912
rect -600 2500 -188 2512
rect -1212 2300 -1200 2500
rect -200 2300 -188 2500
rect -1212 2288 -800 2300
rect -812 1900 -800 2288
rect -600 2288 -188 2300
rect -600 1900 -588 2288
rect -812 1888 -588 1900
rect 788 1900 800 2900
rect 1800 1900 1812 2900
rect 788 1888 1812 1900
rect 2788 2900 3812 2912
rect 2788 1900 2800 2900
rect 3800 1900 3812 2900
rect 5188 2900 5412 2912
rect 5188 2512 5200 2900
rect 4788 2500 5200 2512
rect 5400 2512 5412 2900
rect 5400 2500 5812 2512
rect 4788 2300 4800 2500
rect 5800 2300 5812 2500
rect 4788 2288 5200 2300
rect 2788 1888 3812 1900
rect 5188 1900 5200 2288
rect 5400 2288 5812 2300
rect 5400 1900 5412 2288
rect 5188 1888 5412 1900
rect -612 900 412 912
rect -612 -100 -600 900
rect 400 -100 412 900
rect -612 -112 412 -100
rect 4188 900 5212 912
rect 4188 -100 4200 900
rect 5200 -100 5212 900
rect 4188 -112 5212 -100
rect -1612 -1100 -188 -1088
rect -1612 -2500 -1600 -1100
rect -1400 -1312 -400 -1300
rect -1400 -2288 -1388 -1312
rect -412 -2288 -400 -1312
rect -1400 -2300 -400 -2288
rect -200 -2500 -188 -1100
rect 788 -1100 1812 -1088
rect 788 -2100 800 -1100
rect 1800 -2100 1812 -1100
rect 788 -2112 1812 -2100
rect 2788 -1100 3812 -1088
rect 2788 -2100 2800 -1100
rect 3800 -2100 3812 -1100
rect 5188 -1100 5412 -1088
rect 5188 -1488 5200 -1100
rect 4788 -1500 5200 -1488
rect 5400 -1488 5412 -1100
rect 5400 -1500 5812 -1488
rect 4788 -1700 4800 -1500
rect 5800 -1700 5812 -1500
rect 4788 -1712 5200 -1700
rect 2788 -2112 3812 -2100
rect 5188 -2100 5200 -1712
rect 5400 -1712 5812 -1700
rect 5400 -2100 5412 -1712
rect 5188 -2112 5412 -2100
rect -1612 -2512 -188 -2500
<< end >>
