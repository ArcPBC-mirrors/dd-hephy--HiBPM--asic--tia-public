magic
tech sky130A
magscale 1 2
timestamp 1684830260
<< error_p >>
rect -461 272 -403 278
rect -269 272 -211 278
rect -77 272 -19 278
rect 115 272 173 278
rect 307 272 365 278
rect 499 272 557 278
rect -461 238 -449 272
rect -269 238 -257 272
rect -77 238 -65 272
rect 115 238 127 272
rect 307 238 319 272
rect 499 238 511 272
rect -461 232 -403 238
rect -269 232 -211 238
rect -77 232 -19 238
rect 115 232 173 238
rect 307 232 365 238
rect 499 232 557 238
rect -557 -238 -499 -232
rect -365 -238 -307 -232
rect -173 -238 -115 -232
rect 19 -238 77 -232
rect 211 -238 269 -232
rect 403 -238 461 -232
rect -557 -272 -545 -238
rect -365 -272 -353 -238
rect -173 -272 -161 -238
rect 19 -272 31 -238
rect 211 -272 223 -238
rect 403 -272 415 -238
rect -557 -278 -499 -272
rect -365 -278 -307 -272
rect -173 -278 -115 -272
rect 19 -278 77 -272
rect 211 -278 269 -272
rect 403 -278 461 -272
<< pwell >>
rect -743 -410 743 410
<< nmoslvt >>
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
<< ndiff >>
rect -605 188 -543 200
rect -605 -188 -593 188
rect -559 -188 -543 188
rect -605 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 605 200
rect 543 -188 559 188
rect 593 -188 605 188
rect 543 -200 605 -188
<< ndiffc >>
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
<< psubdiff >>
rect -707 340 -611 374
rect 611 340 707 374
rect -707 278 -673 340
rect 673 278 707 340
rect -707 -340 -673 -278
rect 673 -340 707 -278
rect -707 -374 -611 -340
rect 611 -374 707 -340
<< psubdiffcont >>
rect -611 340 611 374
rect -707 -278 -673 278
rect 673 -278 707 278
rect -611 -374 611 -340
<< poly >>
rect -465 272 -399 288
rect -465 238 -449 272
rect -415 238 -399 272
rect -543 200 -513 226
rect -465 222 -399 238
rect -273 272 -207 288
rect -273 238 -257 272
rect -223 238 -207 272
rect -447 200 -417 222
rect -351 200 -321 226
rect -273 222 -207 238
rect -81 272 -15 288
rect -81 238 -65 272
rect -31 238 -15 272
rect -255 200 -225 222
rect -159 200 -129 226
rect -81 222 -15 238
rect 111 272 177 288
rect 111 238 127 272
rect 161 238 177 272
rect -63 200 -33 222
rect 33 200 63 226
rect 111 222 177 238
rect 303 272 369 288
rect 303 238 319 272
rect 353 238 369 272
rect 129 200 159 222
rect 225 200 255 226
rect 303 222 369 238
rect 495 272 561 288
rect 495 238 511 272
rect 545 238 561 272
rect 321 200 351 222
rect 417 200 447 226
rect 495 222 561 238
rect 513 200 543 222
rect -543 -222 -513 -200
rect -561 -238 -495 -222
rect -447 -226 -417 -200
rect -351 -222 -321 -200
rect -561 -272 -545 -238
rect -511 -272 -495 -238
rect -561 -288 -495 -272
rect -369 -238 -303 -222
rect -255 -226 -225 -200
rect -159 -222 -129 -200
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -369 -288 -303 -272
rect -177 -238 -111 -222
rect -63 -226 -33 -200
rect 33 -222 63 -200
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect -177 -288 -111 -272
rect 15 -238 81 -222
rect 129 -226 159 -200
rect 225 -222 255 -200
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 15 -288 81 -272
rect 207 -238 273 -222
rect 321 -226 351 -200
rect 417 -222 447 -200
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 207 -288 273 -272
rect 399 -238 465 -222
rect 513 -226 543 -200
rect 399 -272 415 -238
rect 449 -272 465 -238
rect 399 -288 465 -272
<< polycont >>
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect 511 238 545 272
rect -545 -272 -511 -238
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
<< locali >>
rect -707 340 -611 374
rect 611 340 707 374
rect -707 278 -673 340
rect 673 278 707 340
rect -465 238 -449 272
rect -415 238 -399 272
rect -273 238 -257 272
rect -223 238 -207 272
rect -81 238 -65 272
rect -31 238 -15 272
rect 111 238 127 272
rect 161 238 177 272
rect 303 238 319 272
rect 353 238 369 272
rect 495 238 511 272
rect 545 238 561 272
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect -561 -272 -545 -238
rect -511 -272 -495 -238
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 399 -272 415 -238
rect 449 -272 465 -238
rect -707 -340 -673 -278
rect 673 -340 707 -278
rect -707 -374 -611 -340
rect 611 -374 707 -340
<< viali >>
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect 511 238 545 272
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect -545 -272 -511 -238
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
<< metal1 >>
rect -461 272 -403 278
rect -461 238 -449 272
rect -415 238 -403 272
rect -461 232 -403 238
rect -269 272 -211 278
rect -269 238 -257 272
rect -223 238 -211 272
rect -269 232 -211 238
rect -77 272 -19 278
rect -77 238 -65 272
rect -31 238 -19 272
rect -77 232 -19 238
rect 115 272 173 278
rect 115 238 127 272
rect 161 238 173 272
rect 115 232 173 238
rect 307 272 365 278
rect 307 238 319 272
rect 353 238 365 272
rect 307 232 365 238
rect 499 272 557 278
rect 499 238 511 272
rect 545 238 557 272
rect 499 232 557 238
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect -557 -238 -499 -232
rect -557 -272 -545 -238
rect -511 -272 -499 -238
rect -557 -278 -499 -272
rect -365 -238 -307 -232
rect -365 -272 -353 -238
rect -319 -272 -307 -238
rect -365 -278 -307 -272
rect -173 -238 -115 -232
rect -173 -272 -161 -238
rect -127 -272 -115 -238
rect -173 -278 -115 -272
rect 19 -238 77 -232
rect 19 -272 31 -238
rect 65 -272 77 -238
rect 19 -278 77 -272
rect 211 -238 269 -232
rect 211 -272 223 -238
rect 257 -272 269 -238
rect 211 -278 269 -272
rect 403 -238 461 -232
rect 403 -272 415 -238
rect 449 -272 461 -238
rect 403 -278 461 -272
<< properties >>
string FIXED_BBOX -690 -357 690 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
