magic
tech sky130A
magscale 1 2
timestamp 1685113734
<< metal1 >>
rect -3398 4370 -2564 4376
rect -3398 4268 -3102 4370
rect -2912 4268 -2564 4370
rect -3398 4260 -2564 4268
rect -1658 4370 -824 4376
rect -1658 4268 -1368 4370
rect -1178 4268 -824 4370
rect -1658 4260 -824 4268
rect 90 4372 924 4376
rect 90 4270 374 4372
rect 564 4270 924 4372
rect 90 4260 924 4270
rect -3442 3792 -2608 3800
rect -3442 3690 -3104 3792
rect -2914 3690 -2608 3792
rect -3442 3684 -2608 3690
rect -1688 3794 -854 3800
rect -1688 3692 -1366 3794
rect -1176 3692 -854 3794
rect -1688 3684 -854 3692
rect 48 3794 882 3800
rect 48 3692 374 3794
rect 564 3692 882 3794
rect 48 3684 882 3692
<< via1 >>
rect -3102 4268 -2912 4370
rect -1368 4268 -1178 4370
rect 374 4270 564 4372
rect -3104 3690 -2914 3792
rect -1366 3692 -1176 3794
rect 374 3692 564 3794
<< metal2 >>
rect -3110 4378 -2906 4388
rect -4480 3976 -3278 3986
rect -3110 3792 -2906 4102
rect -1374 4378 -1170 4388
rect -3110 3690 -3104 3792
rect -2914 3690 -2906 3792
rect -3110 3684 -2906 3690
rect -2738 3976 -1536 3986
rect -3104 3680 -2914 3684
rect -4480 3612 -3278 3622
rect -1374 3794 -1170 4102
rect 368 4376 572 4386
rect -1374 3692 -1366 3794
rect -1176 3692 -1170 3794
rect -1374 3684 -1170 3692
rect -1000 3976 202 3986
rect -1366 3682 -1176 3684
rect -2738 3612 -1536 3622
rect 368 3794 572 4100
rect 368 3692 374 3794
rect 564 3692 572 3794
rect 368 3684 572 3692
rect 740 3976 1942 3986
rect 374 3682 564 3684
rect -1000 3612 202 3622
rect 740 3612 1942 3622
<< via2 >>
rect -3110 4370 -2906 4378
rect -3110 4268 -3102 4370
rect -3102 4268 -2912 4370
rect -2912 4268 -2906 4370
rect -3110 4102 -2906 4268
rect -4480 3622 -3278 3976
rect -1374 4370 -1170 4378
rect -1374 4268 -1368 4370
rect -1368 4268 -1178 4370
rect -1178 4268 -1170 4370
rect -1374 4102 -1170 4268
rect -2738 3622 -1536 3976
rect 368 4372 572 4376
rect 368 4270 374 4372
rect 374 4270 564 4372
rect 564 4270 572 4372
rect 368 4100 572 4270
rect -1000 3622 202 3976
rect 740 3622 1942 3976
<< metal3 >>
rect -4596 4592 2044 5040
rect -3120 4378 -2896 4383
rect -3120 4102 -3110 4378
rect -2906 4102 -2896 4378
rect -3120 4097 -2896 4102
rect -1384 4378 -1160 4383
rect -1384 4102 -1374 4378
rect -1170 4102 -1160 4378
rect -1384 4097 -1160 4102
rect 358 4376 582 4381
rect 358 4100 368 4376
rect 572 4100 582 4376
rect 358 4095 582 4100
rect -4490 3976 -3268 3981
rect -4490 3622 -4480 3976
rect -3278 3622 -3268 3976
rect -4490 3617 -3268 3622
rect -2748 3976 -1526 3981
rect -2748 3622 -2738 3976
rect -1536 3622 -1526 3976
rect -2748 3617 -1526 3622
rect -1010 3976 212 3981
rect -1010 3622 -1000 3976
rect 202 3622 212 3976
rect -1010 3617 212 3622
rect 730 3976 1952 3981
rect 730 3622 740 3976
rect 1942 3622 1952 3976
rect 730 3617 1952 3622
<< via3 >>
rect -3110 4102 -2906 4378
rect -1374 4102 -1170 4378
rect 368 4100 572 4376
<< metal4 >>
rect -3111 4378 -2905 4379
rect -1375 4378 -1169 4379
rect -4422 4102 -3110 4378
rect -2906 4102 -1374 4378
rect -1170 4376 574 4378
rect -1170 4102 368 4376
rect -3111 4101 -2905 4102
rect -1375 4101 -1169 4102
rect 367 4100 368 4102
rect 572 4102 574 4376
rect 572 4100 573 4102
rect 367 4099 573 4100
use outd_diffamp_10#0  outd_diffamp_10_6
timestamp 1685113734
transform 1 0 -4680 0 1 3600
box -80 20 1668 3804
use outd_diffamp_10#0  outd_diffamp_10_7
timestamp 1685113734
transform 1 0 -2940 0 1 3600
box -80 20 1668 3804
use outd_diffamp_10#0  outd_diffamp_10_8
timestamp 1685113734
transform 1 0 540 0 1 3600
box -80 20 1668 3804
use outd_diffamp_10#0  outd_diffamp_10_9
timestamp 1685113734
transform 1 0 -1200 0 1 3600
box -80 20 1668 3804
<< end >>
