magic
tech sky130A
magscale 1 2
timestamp 1683131499
<< error_p >>
rect -941 581 -883 587
rect -749 581 -691 587
rect -557 581 -499 587
rect -365 581 -307 587
rect -173 581 -115 587
rect 19 581 77 587
rect 211 581 269 587
rect 403 581 461 587
rect 595 581 653 587
rect 787 581 845 587
rect -941 547 -929 581
rect -749 547 -737 581
rect -557 547 -545 581
rect -365 547 -353 581
rect -173 547 -161 581
rect 19 547 31 581
rect 211 547 223 581
rect 403 547 415 581
rect 595 547 607 581
rect 787 547 799 581
rect -941 541 -883 547
rect -749 541 -691 547
rect -557 541 -499 547
rect -365 541 -307 547
rect -173 541 -115 547
rect 19 541 77 547
rect 211 541 269 547
rect 403 541 461 547
rect 595 541 653 547
rect 787 541 845 547
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect -941 -547 -883 -541
rect -749 -547 -691 -541
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect 595 -547 653 -541
rect 787 -547 845 -541
rect -941 -581 -929 -547
rect -749 -581 -737 -547
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect 595 -581 607 -547
rect 787 -581 799 -547
rect -941 -587 -883 -581
rect -749 -587 -691 -581
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
rect 595 -587 653 -581
rect 787 -587 845 -581
<< pwell >>
rect -1127 -719 1127 719
<< nmos >>
rect -927 109 -897 509
rect -831 109 -801 509
rect -735 109 -705 509
rect -639 109 -609 509
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect 609 109 639 509
rect 705 109 735 509
rect 801 109 831 509
rect 897 109 927 509
rect -927 -509 -897 -109
rect -831 -509 -801 -109
rect -735 -509 -705 -109
rect -639 -509 -609 -109
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect 609 -509 639 -109
rect 705 -509 735 -109
rect 801 -509 831 -109
rect 897 -509 927 -109
<< ndiff >>
rect -989 497 -927 509
rect -989 121 -977 497
rect -943 121 -927 497
rect -989 109 -927 121
rect -897 497 -831 509
rect -897 121 -881 497
rect -847 121 -831 497
rect -897 109 -831 121
rect -801 497 -735 509
rect -801 121 -785 497
rect -751 121 -735 497
rect -801 109 -735 121
rect -705 497 -639 509
rect -705 121 -689 497
rect -655 121 -639 497
rect -705 109 -639 121
rect -609 497 -543 509
rect -609 121 -593 497
rect -559 121 -543 497
rect -609 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 609 509
rect 543 121 559 497
rect 593 121 609 497
rect 543 109 609 121
rect 639 497 705 509
rect 639 121 655 497
rect 689 121 705 497
rect 639 109 705 121
rect 735 497 801 509
rect 735 121 751 497
rect 785 121 801 497
rect 735 109 801 121
rect 831 497 897 509
rect 831 121 847 497
rect 881 121 897 497
rect 831 109 897 121
rect 927 497 989 509
rect 927 121 943 497
rect 977 121 989 497
rect 927 109 989 121
rect -989 -121 -927 -109
rect -989 -497 -977 -121
rect -943 -497 -927 -121
rect -989 -509 -927 -497
rect -897 -121 -831 -109
rect -897 -497 -881 -121
rect -847 -497 -831 -121
rect -897 -509 -831 -497
rect -801 -121 -735 -109
rect -801 -497 -785 -121
rect -751 -497 -735 -121
rect -801 -509 -735 -497
rect -705 -121 -639 -109
rect -705 -497 -689 -121
rect -655 -497 -639 -121
rect -705 -509 -639 -497
rect -609 -121 -543 -109
rect -609 -497 -593 -121
rect -559 -497 -543 -121
rect -609 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 609 -109
rect 543 -497 559 -121
rect 593 -497 609 -121
rect 543 -509 609 -497
rect 639 -121 705 -109
rect 639 -497 655 -121
rect 689 -497 705 -121
rect 639 -509 705 -497
rect 735 -121 801 -109
rect 735 -497 751 -121
rect 785 -497 801 -121
rect 735 -509 801 -497
rect 831 -121 897 -109
rect 831 -497 847 -121
rect 881 -497 897 -121
rect 831 -509 897 -497
rect 927 -121 989 -109
rect 927 -497 943 -121
rect 977 -497 989 -121
rect 927 -509 989 -497
<< ndiffc >>
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
<< psubdiff >>
rect -1091 649 -995 683
rect 995 649 1091 683
rect -1091 587 -1057 649
rect 1057 587 1091 649
rect -1091 -649 -1057 -587
rect 1057 -649 1091 -587
rect -1091 -683 -995 -649
rect 995 -683 1091 -649
<< psubdiffcont >>
rect -995 649 995 683
rect -1091 -587 -1057 587
rect 1057 -587 1091 587
rect -995 -683 995 -649
<< poly >>
rect -945 581 -879 597
rect -945 547 -929 581
rect -895 547 -879 581
rect -945 531 -879 547
rect -753 581 -687 597
rect -753 547 -737 581
rect -703 547 -687 581
rect -927 509 -897 531
rect -831 509 -801 535
rect -753 531 -687 547
rect -561 581 -495 597
rect -561 547 -545 581
rect -511 547 -495 581
rect -735 509 -705 531
rect -639 509 -609 535
rect -561 531 -495 547
rect -369 581 -303 597
rect -369 547 -353 581
rect -319 547 -303 581
rect -543 509 -513 531
rect -447 509 -417 535
rect -369 531 -303 547
rect -177 581 -111 597
rect -177 547 -161 581
rect -127 547 -111 581
rect -351 509 -321 531
rect -255 509 -225 535
rect -177 531 -111 547
rect 15 581 81 597
rect 15 547 31 581
rect 65 547 81 581
rect -159 509 -129 531
rect -63 509 -33 535
rect 15 531 81 547
rect 207 581 273 597
rect 207 547 223 581
rect 257 547 273 581
rect 33 509 63 531
rect 129 509 159 535
rect 207 531 273 547
rect 399 581 465 597
rect 399 547 415 581
rect 449 547 465 581
rect 225 509 255 531
rect 321 509 351 535
rect 399 531 465 547
rect 591 581 657 597
rect 591 547 607 581
rect 641 547 657 581
rect 417 509 447 531
rect 513 509 543 535
rect 591 531 657 547
rect 783 581 849 597
rect 783 547 799 581
rect 833 547 849 581
rect 609 509 639 531
rect 705 509 735 535
rect 783 531 849 547
rect 801 509 831 531
rect 897 509 927 535
rect -927 83 -897 109
rect -831 87 -801 109
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 897 -109 927 -87
rect -927 -531 -897 -509
rect -945 -547 -879 -531
rect -831 -535 -801 -509
rect -735 -531 -705 -509
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -945 -597 -879 -581
rect -753 -547 -687 -531
rect -639 -535 -609 -509
rect -543 -531 -513 -509
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -753 -597 -687 -581
rect -561 -547 -495 -531
rect -447 -535 -417 -509
rect -351 -531 -321 -509
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -255 -535 -225 -509
rect -159 -531 -129 -509
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -63 -535 -33 -509
rect 33 -531 63 -509
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 129 -535 159 -509
rect 225 -531 255 -509
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 321 -535 351 -509
rect 417 -531 447 -509
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 513 -535 543 -509
rect 609 -531 639 -509
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
rect 591 -547 657 -531
rect 705 -535 735 -509
rect 801 -531 831 -509
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 591 -597 657 -581
rect 783 -547 849 -531
rect 897 -535 927 -509
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 783 -597 849 -581
<< polycont >>
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
<< locali >>
rect -1091 649 -995 683
rect 995 649 1091 683
rect -1091 587 -1057 649
rect 1057 587 1091 649
rect -945 547 -929 581
rect -895 547 -879 581
rect -753 547 -737 581
rect -703 547 -687 581
rect -561 547 -545 581
rect -511 547 -495 581
rect -369 547 -353 581
rect -319 547 -303 581
rect -177 547 -161 581
rect -127 547 -111 581
rect 15 547 31 581
rect 65 547 81 581
rect 207 547 223 581
rect 257 547 273 581
rect 399 547 415 581
rect 449 547 465 581
rect 591 547 607 581
rect 641 547 657 581
rect 783 547 799 581
rect 833 547 849 581
rect -977 497 -943 513
rect -977 105 -943 121
rect -881 497 -847 513
rect -881 105 -847 121
rect -785 497 -751 513
rect -785 105 -751 121
rect -689 497 -655 513
rect -689 105 -655 121
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect 655 497 689 513
rect 655 105 689 121
rect 751 497 785 513
rect 751 105 785 121
rect 847 497 881 513
rect 847 105 881 121
rect 943 497 977 513
rect 943 105 977 121
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect -977 -121 -943 -105
rect -977 -513 -943 -497
rect -881 -121 -847 -105
rect -881 -513 -847 -497
rect -785 -121 -751 -105
rect -785 -513 -751 -497
rect -689 -121 -655 -105
rect -689 -513 -655 -497
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect 655 -121 689 -105
rect 655 -513 689 -497
rect 751 -121 785 -105
rect 751 -513 785 -497
rect 847 -121 881 -105
rect 847 -513 881 -497
rect 943 -121 977 -105
rect 943 -513 977 -497
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 783 -581 799 -547
rect 833 -581 849 -547
rect -1091 -649 -1057 -587
rect 1057 -649 1091 -587
rect -1091 -683 -995 -649
rect 995 -683 1091 -649
<< viali >>
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
<< metal1 >>
rect -941 581 -883 587
rect -941 547 -929 581
rect -895 547 -883 581
rect -941 541 -883 547
rect -749 581 -691 587
rect -749 547 -737 581
rect -703 547 -691 581
rect -749 541 -691 547
rect -557 581 -499 587
rect -557 547 -545 581
rect -511 547 -499 581
rect -557 541 -499 547
rect -365 581 -307 587
rect -365 547 -353 581
rect -319 547 -307 581
rect -365 541 -307 547
rect -173 581 -115 587
rect -173 547 -161 581
rect -127 547 -115 581
rect -173 541 -115 547
rect 19 581 77 587
rect 19 547 31 581
rect 65 547 77 581
rect 19 541 77 547
rect 211 581 269 587
rect 211 547 223 581
rect 257 547 269 581
rect 211 541 269 547
rect 403 581 461 587
rect 403 547 415 581
rect 449 547 461 581
rect 403 541 461 547
rect 595 581 653 587
rect 595 547 607 581
rect 641 547 653 581
rect 595 541 653 547
rect 787 581 845 587
rect 787 547 799 581
rect 833 547 845 581
rect 787 541 845 547
rect -983 497 -937 509
rect -983 121 -977 497
rect -943 121 -937 497
rect -983 109 -937 121
rect -887 497 -841 509
rect -887 121 -881 497
rect -847 121 -841 497
rect -887 109 -841 121
rect -791 497 -745 509
rect -791 121 -785 497
rect -751 121 -745 497
rect -791 109 -745 121
rect -695 497 -649 509
rect -695 121 -689 497
rect -655 121 -649 497
rect -695 109 -649 121
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect 649 497 695 509
rect 649 121 655 497
rect 689 121 695 497
rect 649 109 695 121
rect 745 497 791 509
rect 745 121 751 497
rect 785 121 791 497
rect 745 109 791 121
rect 841 497 887 509
rect 841 121 847 497
rect 881 121 887 497
rect 841 109 887 121
rect 937 497 983 509
rect 937 121 943 497
rect 977 121 983 497
rect 937 109 983 121
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect -983 -121 -937 -109
rect -983 -497 -977 -121
rect -943 -497 -937 -121
rect -983 -509 -937 -497
rect -887 -121 -841 -109
rect -887 -497 -881 -121
rect -847 -497 -841 -121
rect -887 -509 -841 -497
rect -791 -121 -745 -109
rect -791 -497 -785 -121
rect -751 -497 -745 -121
rect -791 -509 -745 -497
rect -695 -121 -649 -109
rect -695 -497 -689 -121
rect -655 -497 -649 -121
rect -695 -509 -649 -497
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect 649 -121 695 -109
rect 649 -497 655 -121
rect 689 -497 695 -121
rect 649 -509 695 -497
rect 745 -121 791 -109
rect 745 -497 751 -121
rect 785 -497 791 -121
rect 745 -509 791 -497
rect 841 -121 887 -109
rect 841 -497 847 -121
rect 881 -497 887 -121
rect 841 -509 887 -497
rect 937 -121 983 -109
rect 937 -497 943 -121
rect 977 -497 983 -121
rect 937 -509 983 -497
rect -941 -547 -883 -541
rect -941 -581 -929 -547
rect -895 -581 -883 -547
rect -941 -587 -883 -581
rect -749 -547 -691 -541
rect -749 -581 -737 -547
rect -703 -581 -691 -547
rect -749 -587 -691 -581
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
rect 595 -547 653 -541
rect 595 -581 607 -547
rect 641 -581 653 -547
rect 595 -587 653 -581
rect 787 -547 845 -541
rect 787 -581 799 -547
rect 833 -581 845 -547
rect 787 -587 845 -581
<< properties >>
string FIXED_BBOX -1074 -666 1074 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 2 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
