magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< pwell >>
rect 188 -1284 1428 -1240
rect 752 -4264 872 -3752
<< poly >>
rect 752 -4264 872 -3752
<< metal1 >>
rect 140 1480 1292 1560
rect 226 1268 236 1448
rect 288 1268 298 1448
rect 418 1268 428 1448
rect 480 1268 490 1448
rect 610 1268 620 1448
rect 672 1268 682 1448
rect 802 1268 812 1448
rect 864 1268 874 1448
rect 994 1268 1004 1448
rect 1056 1268 1066 1448
rect 130 1044 140 1224
rect 192 1044 202 1224
rect 322 1044 332 1224
rect 384 1044 394 1224
rect 514 1044 524 1224
rect 576 1044 586 1224
rect 706 1044 716 1224
rect 768 1044 778 1224
rect 898 1044 908 1224
rect 960 1044 970 1224
rect 1090 1044 1100 1224
rect 1152 1044 1162 1224
rect 1192 1008 1292 1480
rect 176 864 1292 1008
rect 226 652 236 832
rect 288 652 298 832
rect 418 652 428 832
rect 480 652 490 832
rect 610 652 620 832
rect 672 652 682 832
rect 802 652 812 832
rect 864 652 874 832
rect 994 652 1004 832
rect 1056 652 1066 832
rect 130 428 140 608
rect 192 428 202 608
rect 322 428 332 608
rect 384 428 394 608
rect 514 428 524 608
rect 576 428 586 608
rect 706 428 716 608
rect 768 428 778 608
rect 898 428 908 608
rect 960 428 970 608
rect 1090 428 1100 608
rect 1152 428 1162 608
rect 1192 392 1292 864
rect 276 248 1292 392
rect 226 32 236 212
rect 288 32 298 212
rect 418 32 428 212
rect 480 32 490 212
rect 610 32 620 212
rect 672 32 682 212
rect 802 32 812 212
rect 864 32 874 212
rect 994 32 1004 212
rect 1056 32 1066 212
rect 130 -192 140 -12
rect 192 -192 202 -12
rect 322 -192 332 -12
rect 384 -192 394 -12
rect 514 -192 524 -12
rect 576 -192 586 -12
rect 706 -192 716 -12
rect 768 -192 778 -12
rect 898 -192 908 -12
rect 960 -192 970 -12
rect 1090 -192 1100 -12
rect 1152 -192 1162 -12
rect 1192 -228 1292 248
rect 180 -360 1292 -228
rect 740 -608 884 -360
rect 188 -668 1428 -608
rect 130 -880 140 -700
rect 192 -880 202 -700
rect 390 -1100 400 -920
rect 452 -1100 462 -920
rect 492 -1132 612 -668
rect 646 -880 656 -700
rect 708 -880 718 -700
rect 752 -1132 872 -668
rect 906 -1100 916 -920
rect 968 -1100 978 -920
rect 1012 -1132 1132 -668
rect 1162 -880 1172 -700
rect 1224 -880 1234 -700
rect 1422 -1100 1432 -920
rect 1484 -1100 1494 -920
rect 188 -1136 1428 -1132
rect 184 -1284 1428 -1136
rect 130 -1496 140 -1316
rect 192 -1496 202 -1316
rect 390 -1716 400 -1536
rect 452 -1716 462 -1536
rect 492 -1752 612 -1284
rect 646 -1496 656 -1316
rect 708 -1496 718 -1316
rect 752 -1748 872 -1284
rect 906 -1716 916 -1536
rect 968 -1716 978 -1536
rect 740 -1752 884 -1748
rect 1012 -1752 1132 -1284
rect 1162 -1496 1172 -1316
rect 1224 -1496 1234 -1316
rect 1422 -1716 1432 -1536
rect 1484 -1716 1494 -1536
rect 188 -1756 1428 -1752
rect 188 -1904 1432 -1756
rect 130 -2116 140 -1936
rect 192 -2116 202 -1936
rect 390 -2336 400 -2156
rect 452 -2336 462 -2156
rect 492 -2368 612 -1904
rect 646 -2116 656 -1936
rect 708 -2116 718 -1936
rect 752 -2368 872 -1904
rect 906 -2336 916 -2156
rect 968 -2336 978 -2156
rect 1012 -2368 1132 -1904
rect 1162 -2116 1172 -1936
rect 1224 -2116 1234 -1936
rect 1422 -2336 1432 -2156
rect 1484 -2336 1494 -2156
rect 188 -2372 386 -2368
rect 184 -2404 386 -2372
rect 458 -2404 902 -2368
rect 974 -2404 1418 -2368
rect 184 -2520 1428 -2404
rect 130 -2732 140 -2552
rect 192 -2732 202 -2552
rect 390 -2952 400 -2772
rect 452 -2952 462 -2772
rect 492 -2988 612 -2520
rect 740 -2524 884 -2520
rect 646 -2732 656 -2552
rect 708 -2732 718 -2552
rect 752 -2988 872 -2524
rect 906 -2952 916 -2772
rect 968 -2952 978 -2772
rect 1012 -2988 1132 -2520
rect 1162 -2732 1172 -2552
rect 1224 -2732 1234 -2552
rect 1422 -2952 1432 -2772
rect 1484 -2952 1494 -2772
rect 188 -2992 1428 -2988
rect 188 -3140 1432 -2992
rect 130 -3352 140 -3172
rect 192 -3352 202 -3172
rect 390 -3572 400 -3392
rect 452 -3572 462 -3392
rect 492 -3604 612 -3140
rect 646 -3352 656 -3172
rect 708 -3352 718 -3172
rect 752 -3604 872 -3140
rect 906 -3572 916 -3392
rect 968 -3572 978 -3392
rect 1012 -3604 1132 -3140
rect 1162 -3352 1172 -3172
rect 1224 -3352 1234 -3172
rect 1422 -3572 1432 -3392
rect 1484 -3572 1494 -3392
rect 188 -3620 386 -3604
rect 458 -3620 902 -3604
rect 974 -3620 1418 -3604
rect 188 -3756 1432 -3620
rect 130 -3968 140 -3788
rect 192 -3968 202 -3788
rect 390 -4188 400 -4008
rect 452 -4188 462 -4008
rect 492 -4220 612 -3756
rect 646 -3968 656 -3788
rect 708 -3968 718 -3788
rect 752 -4220 872 -3756
rect 906 -4188 916 -4008
rect 968 -4188 978 -4008
rect 1012 -4220 1132 -3756
rect 1162 -3968 1172 -3788
rect 1224 -3968 1234 -3788
rect 1422 -4188 1432 -4008
rect 1484 -4188 1494 -4008
rect 188 -4280 1428 -4220
<< via1 >>
rect 236 1268 288 1448
rect 428 1268 480 1448
rect 620 1268 672 1448
rect 812 1268 864 1448
rect 1004 1268 1056 1448
rect 140 1044 192 1224
rect 332 1044 384 1224
rect 524 1044 576 1224
rect 716 1044 768 1224
rect 908 1044 960 1224
rect 1100 1044 1152 1224
rect 236 652 288 832
rect 428 652 480 832
rect 620 652 672 832
rect 812 652 864 832
rect 1004 652 1056 832
rect 140 428 192 608
rect 332 428 384 608
rect 524 428 576 608
rect 716 428 768 608
rect 908 428 960 608
rect 1100 428 1152 608
rect 236 32 288 212
rect 428 32 480 212
rect 620 32 672 212
rect 812 32 864 212
rect 1004 32 1056 212
rect 140 -192 192 -12
rect 332 -192 384 -12
rect 524 -192 576 -12
rect 716 -192 768 -12
rect 908 -192 960 -12
rect 1100 -192 1152 -12
rect 140 -880 192 -700
rect 400 -1100 452 -920
rect 656 -880 708 -700
rect 916 -1100 968 -920
rect 1172 -880 1224 -700
rect 1432 -1100 1484 -920
rect 140 -1496 192 -1316
rect 400 -1716 452 -1536
rect 656 -1496 708 -1316
rect 916 -1716 968 -1536
rect 1172 -1496 1224 -1316
rect 1432 -1716 1484 -1536
rect 140 -2116 192 -1936
rect 400 -2336 452 -2156
rect 656 -2116 708 -1936
rect 916 -2336 968 -2156
rect 1172 -2116 1224 -1936
rect 1432 -2336 1484 -2156
rect 140 -2732 192 -2552
rect 400 -2952 452 -2772
rect 656 -2732 708 -2552
rect 916 -2952 968 -2772
rect 1172 -2732 1224 -2552
rect 1432 -2952 1484 -2772
rect 140 -3352 192 -3172
rect 400 -3572 452 -3392
rect 656 -3352 708 -3172
rect 916 -3572 968 -3392
rect 1172 -3352 1224 -3172
rect 1432 -3572 1484 -3392
rect 140 -3968 192 -3788
rect 400 -4188 452 -4008
rect 656 -3968 708 -3788
rect 916 -4188 968 -4008
rect 1172 -3968 1224 -3788
rect 1432 -4188 1484 -4008
<< metal2 >>
rect 236 1456 1056 1460
rect 236 1448 1496 1456
rect 288 1284 428 1448
rect 236 1258 288 1268
rect 480 1284 620 1448
rect 428 1258 480 1268
rect 672 1284 812 1448
rect 620 1258 672 1268
rect 864 1284 1004 1448
rect 812 1258 864 1268
rect 1056 1284 1496 1448
rect 1004 1258 1056 1268
rect 140 1226 192 1234
rect 332 1226 384 1234
rect 524 1226 576 1234
rect 716 1226 768 1234
rect 136 1224 768 1226
rect 908 1224 960 1234
rect 1100 1224 1152 1234
rect 136 1216 140 1224
rect 192 1216 332 1224
rect 384 1216 524 1224
rect 576 1216 716 1224
rect 768 1044 908 1224
rect 960 1044 1100 1224
rect 740 1036 1152 1044
rect 740 1034 768 1036
rect 908 1034 960 1036
rect 1100 1034 1152 1036
rect 136 1022 740 1032
rect 236 840 1056 844
rect 1184 840 1496 1284
rect 236 832 1496 840
rect 288 652 428 832
rect 480 652 620 832
rect 672 652 812 832
rect 864 652 1004 832
rect 1056 652 1496 832
rect 236 642 288 652
rect 428 642 480 652
rect 620 642 672 652
rect 812 642 864 652
rect 1004 642 1056 652
rect 140 610 192 618
rect 332 610 384 618
rect 524 610 576 618
rect 716 610 768 618
rect 136 608 768 610
rect 908 608 960 618
rect 1100 608 1152 618
rect 136 600 140 608
rect 192 600 332 608
rect 384 600 524 608
rect 576 600 716 608
rect 768 428 908 608
rect 960 428 1100 608
rect 740 420 1152 428
rect 740 418 768 420
rect 908 418 960 420
rect 1100 418 1152 420
rect 136 406 740 416
rect 236 216 288 222
rect 428 216 480 222
rect 620 216 672 222
rect 812 216 864 222
rect 1004 216 1056 222
rect 1184 216 1496 652
rect 236 212 1496 216
rect 288 32 428 212
rect 480 32 620 212
rect 672 32 812 212
rect 864 32 1004 212
rect 1056 32 1496 212
rect 236 28 1496 32
rect 236 22 288 28
rect 428 22 480 28
rect 620 22 672 28
rect 812 22 864 28
rect 1004 22 1056 28
rect 140 -10 192 -2
rect 332 -10 384 -2
rect 524 -10 576 -2
rect 716 -10 768 -2
rect 132 -12 768 -10
rect 908 -12 960 -2
rect 1100 -12 1152 -2
rect 132 -20 140 -12
rect 192 -20 332 -12
rect 384 -20 524 -12
rect 576 -20 716 -12
rect 768 -192 908 -12
rect 960 -192 1100 -12
rect 736 -200 1152 -192
rect 736 -202 768 -200
rect 908 -202 960 -200
rect 1100 -202 1152 -200
rect 132 -214 736 -204
rect 140 -688 740 -678
rect 740 -700 1224 -688
rect 740 -872 1172 -700
rect 192 -880 656 -872
rect 708 -880 1172 -872
rect 140 -882 740 -880
rect 140 -890 192 -882
rect 656 -890 708 -882
rect 1172 -890 1224 -880
rect 400 -920 452 -910
rect 916 -918 968 -910
rect 1432 -918 1484 -910
rect 884 -920 1484 -918
rect 452 -928 916 -920
rect 968 -928 1432 -920
rect 452 -1100 884 -928
rect 400 -1112 884 -1100
rect 884 -1122 1484 -1112
rect 140 -1304 740 -1294
rect 740 -1316 1224 -1304
rect 740 -1488 1172 -1316
rect 192 -1496 656 -1488
rect 708 -1496 1172 -1488
rect 140 -1498 740 -1496
rect 140 -1506 192 -1498
rect 656 -1506 708 -1498
rect 1172 -1506 1224 -1496
rect 400 -1536 452 -1526
rect 916 -1534 968 -1526
rect 1432 -1534 1484 -1526
rect 884 -1536 1484 -1534
rect 452 -1544 916 -1536
rect 968 -1544 1432 -1536
rect 452 -1716 884 -1544
rect 400 -1728 884 -1716
rect 884 -1738 1484 -1728
rect 140 -1924 740 -1914
rect 740 -1936 1224 -1924
rect 740 -2108 1172 -1936
rect 192 -2116 656 -2108
rect 708 -2116 1172 -2108
rect 140 -2118 740 -2116
rect 140 -2126 192 -2118
rect 656 -2126 708 -2118
rect 1172 -2126 1224 -2116
rect 400 -2156 452 -2146
rect 916 -2154 968 -2146
rect 1432 -2154 1484 -2146
rect 884 -2156 1484 -2154
rect 452 -2164 916 -2156
rect 968 -2164 1432 -2156
rect 452 -2336 884 -2164
rect 400 -2348 884 -2336
rect 884 -2358 1484 -2348
rect 140 -2540 740 -2530
rect 740 -2552 1224 -2540
rect 740 -2724 1172 -2552
rect 192 -2732 656 -2724
rect 708 -2732 1172 -2724
rect 140 -2734 740 -2732
rect 140 -2742 192 -2734
rect 656 -2742 708 -2734
rect 1172 -2742 1224 -2732
rect 400 -2772 452 -2762
rect 916 -2770 968 -2762
rect 1432 -2770 1484 -2762
rect 884 -2772 1484 -2770
rect 452 -2780 916 -2772
rect 968 -2780 1432 -2772
rect 452 -2952 884 -2780
rect 400 -2964 884 -2952
rect 884 -2974 1484 -2964
rect 140 -3160 740 -3150
rect 740 -3172 1224 -3160
rect 740 -3344 1172 -3172
rect 192 -3352 656 -3344
rect 708 -3352 1172 -3344
rect 140 -3354 740 -3352
rect 140 -3362 192 -3354
rect 656 -3362 708 -3354
rect 1172 -3362 1224 -3352
rect 400 -3392 452 -3382
rect 916 -3390 968 -3382
rect 1432 -3390 1484 -3382
rect 884 -3392 1484 -3390
rect 452 -3400 916 -3392
rect 968 -3400 1432 -3392
rect 452 -3572 884 -3400
rect 400 -3584 884 -3572
rect 884 -3594 1484 -3584
rect 140 -3776 740 -3766
rect 740 -3788 1224 -3776
rect 740 -3960 1172 -3788
rect 192 -3968 656 -3960
rect 708 -3968 1172 -3960
rect 140 -3970 740 -3968
rect 140 -3978 192 -3970
rect 656 -3978 708 -3970
rect 1172 -3978 1224 -3968
rect 400 -4008 452 -3998
rect 916 -4006 968 -3998
rect 1432 -4006 1484 -3998
rect 884 -4008 1484 -4006
rect 452 -4016 916 -4008
rect 968 -4016 1432 -4008
rect 452 -4188 884 -4016
rect 400 -4200 884 -4188
rect 884 -4210 1484 -4200
<< via2 >>
rect 136 1044 140 1216
rect 140 1044 192 1216
rect 192 1044 332 1216
rect 332 1044 384 1216
rect 384 1044 524 1216
rect 524 1044 576 1216
rect 576 1044 716 1216
rect 716 1044 740 1216
rect 136 1032 740 1044
rect 136 428 140 600
rect 140 428 192 600
rect 192 428 332 600
rect 332 428 384 600
rect 384 428 524 600
rect 524 428 576 600
rect 576 428 716 600
rect 716 428 740 600
rect 136 416 740 428
rect 132 -192 140 -20
rect 140 -192 192 -20
rect 192 -192 332 -20
rect 332 -192 384 -20
rect 384 -192 524 -20
rect 524 -192 576 -20
rect 576 -192 716 -20
rect 716 -192 736 -20
rect 132 -204 736 -192
rect 140 -700 740 -688
rect 140 -872 192 -700
rect 192 -872 656 -700
rect 656 -872 708 -700
rect 708 -872 740 -700
rect 884 -1100 916 -928
rect 916 -1100 968 -928
rect 968 -1100 1432 -928
rect 1432 -1100 1484 -928
rect 884 -1112 1484 -1100
rect 140 -1316 740 -1304
rect 140 -1488 192 -1316
rect 192 -1488 656 -1316
rect 656 -1488 708 -1316
rect 708 -1488 740 -1316
rect 884 -1716 916 -1544
rect 916 -1716 968 -1544
rect 968 -1716 1432 -1544
rect 1432 -1716 1484 -1544
rect 884 -1728 1484 -1716
rect 140 -1936 740 -1924
rect 140 -2108 192 -1936
rect 192 -2108 656 -1936
rect 656 -2108 708 -1936
rect 708 -2108 740 -1936
rect 884 -2336 916 -2164
rect 916 -2336 968 -2164
rect 968 -2336 1432 -2164
rect 1432 -2336 1484 -2164
rect 884 -2348 1484 -2336
rect 140 -2552 740 -2540
rect 140 -2724 192 -2552
rect 192 -2724 656 -2552
rect 656 -2724 708 -2552
rect 708 -2724 740 -2552
rect 884 -2952 916 -2780
rect 916 -2952 968 -2780
rect 968 -2952 1432 -2780
rect 1432 -2952 1484 -2780
rect 884 -2964 1484 -2952
rect 140 -3172 740 -3160
rect 140 -3344 192 -3172
rect 192 -3344 656 -3172
rect 656 -3344 708 -3172
rect 708 -3344 740 -3172
rect 884 -3572 916 -3400
rect 916 -3572 968 -3400
rect 968 -3572 1432 -3400
rect 1432 -3572 1484 -3400
rect 884 -3584 1484 -3572
rect 140 -3788 740 -3776
rect 140 -3960 192 -3788
rect 192 -3960 656 -3788
rect 656 -3960 708 -3788
rect 708 -3960 740 -3788
rect 884 -4188 916 -4016
rect 916 -4188 968 -4016
rect 968 -4188 1432 -4016
rect 1432 -4188 1484 -4016
rect 884 -4200 1484 -4188
<< metal3 >>
rect 136 1221 740 1224
rect 126 1216 750 1221
rect 126 1032 136 1216
rect 740 1032 750 1216
rect 126 1027 750 1032
rect 136 605 740 1027
rect 126 600 750 605
rect 126 416 136 600
rect 740 416 750 600
rect 126 411 750 416
rect 136 -15 740 411
rect 122 -20 746 -15
rect 122 -204 132 -20
rect 736 -204 746 -20
rect 122 -209 746 -204
rect 136 -683 740 -209
rect 130 -688 750 -683
rect 130 -872 140 -688
rect 740 -872 750 -688
rect 130 -877 750 -872
rect 136 -1299 740 -877
rect 874 -928 1494 -923
rect 874 -1112 884 -928
rect 1484 -1112 1494 -928
rect 874 -1117 1494 -1112
rect 130 -1304 750 -1299
rect 130 -1488 140 -1304
rect 740 -1488 750 -1304
rect 130 -1493 750 -1488
rect 136 -1919 740 -1493
rect 884 -1539 1484 -1117
rect 874 -1544 1494 -1539
rect 874 -1728 884 -1544
rect 1484 -1728 1494 -1544
rect 874 -1733 1494 -1728
rect 130 -1924 750 -1919
rect 130 -2108 140 -1924
rect 740 -2108 750 -1924
rect 130 -2113 750 -2108
rect 136 -2535 740 -2113
rect 884 -2159 1484 -1733
rect 874 -2164 1494 -2159
rect 874 -2348 884 -2164
rect 1484 -2348 1494 -2164
rect 874 -2353 1494 -2348
rect 130 -2540 750 -2535
rect 130 -2724 140 -2540
rect 740 -2724 750 -2540
rect 130 -2729 750 -2724
rect 136 -3155 740 -2729
rect 884 -2775 1484 -2353
rect 874 -2780 1494 -2775
rect 874 -2964 884 -2780
rect 1484 -2964 1494 -2780
rect 874 -2969 1494 -2964
rect 130 -3160 750 -3155
rect 130 -3344 140 -3160
rect 740 -3344 750 -3160
rect 130 -3349 750 -3344
rect 136 -3771 740 -3349
rect 884 -3395 1484 -2969
rect 874 -3400 1494 -3395
rect 874 -3584 884 -3400
rect 1484 -3584 1494 -3400
rect 874 -3589 1494 -3584
rect 130 -3776 750 -3771
rect 130 -3960 140 -3776
rect 740 -3960 750 -3776
rect 130 -3965 750 -3960
rect 136 -3984 740 -3965
rect 884 -4011 1484 -3589
rect 874 -4016 1494 -4011
rect 874 -4200 884 -4016
rect 1484 -4200 1494 -4016
rect 874 -4205 1494 -4200
use sky130_fd_pr__nfet_01v8_lvt_R2KHEY  sky130_fd_pr__nfet_01v8_lvt_R2KHEY_1
timestamp 1686659968
transform 1 0 647 0 1 628
box -647 -1028 647 1028
use sky130_fd_pr__nfet_01v8_lvt_YSJU6R  sky130_fd_pr__nfet_01v8_lvt_YSJU6R_0
timestamp 1686659968
transform 1 0 812 0 1 -2445
box -812 -1955 812 1955
<< end >>
