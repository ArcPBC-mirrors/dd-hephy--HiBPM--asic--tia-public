magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< metal3 >>
rect -3186 1012 3186 1040
rect -3186 -1012 3102 1012
rect 3166 -1012 3186 1012
rect -3186 -1040 3186 -1012
<< via3 >>
rect 3102 -1012 3166 1012
<< mimcap >>
rect -3146 960 2854 1000
rect -3146 -960 -3106 960
rect 2814 -960 2854 960
rect -3146 -1000 2854 -960
<< mimcapcontact >>
rect -3106 -960 2814 960
<< metal4 >>
rect 3086 1012 3182 1028
rect -3107 960 2815 961
rect -3107 -960 -3106 960
rect 2814 -960 2815 960
rect -3107 -961 2815 -960
rect 3086 -1012 3102 1012
rect 3166 -1012 3182 1012
rect 3086 -1028 3182 -1012
<< properties >>
string FIXED_BBOX -3186 -1040 2894 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 10 val 615.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
