magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< dnwell >>
rect 1480 -2240 4180 660
<< nwell >>
rect 1400 454 4260 740
rect 1400 -2034 1686 454
rect 3974 -2034 4260 454
rect 1400 -2320 4260 -2034
<< nsubdiff >>
rect 1437 683 4223 703
rect 1437 649 1517 683
rect 4143 649 4223 683
rect 1437 629 4223 649
rect 1437 623 1511 629
rect 1437 -2203 1457 623
rect 1491 -2203 1511 623
rect 1437 -2209 1511 -2203
rect 4149 623 4223 629
rect 4149 -2203 4169 623
rect 4203 -2203 4223 623
rect 4149 -2209 4223 -2203
rect 1437 -2229 4223 -2209
rect 1437 -2263 1517 -2229
rect 4143 -2263 4223 -2229
rect 1437 -2283 4223 -2263
<< nsubdiffcont >>
rect 1517 649 4143 683
rect 1457 -2203 1491 623
rect 4169 -2203 4203 623
rect 1517 -2263 4143 -2229
<< locali >>
rect 1457 649 1517 683
rect 4143 649 4203 683
rect 1457 623 1491 649
rect 4169 623 4203 649
rect 1688 404 1832 456
rect 2124 404 2700 456
rect 2992 404 3636 456
rect 3928 404 3976 456
rect 1688 376 3976 404
rect 1688 204 1764 376
rect 1688 -144 1700 204
rect 1756 -144 1764 204
rect 1688 -336 1764 -144
rect 3888 172 3976 376
rect 3888 -84 3900 172
rect 3960 -84 3976 172
rect 3888 -336 3976 -84
rect 1688 -348 3976 -336
rect 1688 -352 3636 -348
rect 1688 -412 1832 -352
rect 2124 -412 2700 -352
rect 3020 -408 3636 -352
rect 3928 -408 3976 -348
rect 3020 -412 3976 -408
rect 1688 -444 3976 -412
rect 1688 -656 1764 -444
rect 1688 -912 1700 -656
rect 1760 -912 1764 -656
rect 1688 -1148 1764 -912
rect 3888 -676 3976 -444
rect 3888 -932 3900 -676
rect 3960 -932 3976 -676
rect 3888 -1148 3976 -932
rect 1688 -1172 3976 -1148
rect 1688 -1232 1832 -1172
rect 2124 -1232 2700 -1172
rect 2992 -1232 3636 -1172
rect 3928 -1232 3976 -1172
rect 1688 -1248 3976 -1232
rect 1688 -1496 1764 -1248
rect 1688 -1752 1696 -1496
rect 1756 -1752 1764 -1496
rect 1688 -1952 1764 -1752
rect 3888 -1488 3976 -1248
rect 3888 -1744 3900 -1488
rect 3960 -1744 3976 -1488
rect 3888 -1952 3976 -1744
rect 1688 -1984 3976 -1952
rect 1688 -2032 1832 -1984
rect 2124 -2032 2700 -1984
rect 2992 -1988 3976 -1984
rect 2992 -2032 3636 -1988
rect 3928 -2032 3976 -1988
rect 1457 -2229 1491 -2203
rect 4169 -2229 4203 -2203
rect 1457 -2263 1517 -2229
rect 4143 -2263 4203 -2229
<< viali >>
rect 1832 404 2124 464
rect 2700 404 2992 464
rect 3636 404 3928 464
rect 1700 -144 1756 204
rect 3900 -84 3960 172
rect 1832 -412 2124 -352
rect 2700 -412 3020 -352
rect 3636 -408 3928 -348
rect 1700 -912 1760 -656
rect 3900 -932 3960 -676
rect 1832 -1232 2124 -1172
rect 2700 -1232 2992 -1172
rect 3636 -1232 3928 -1172
rect 1696 -1752 1756 -1496
rect 3900 -1744 3960 -1488
rect 1832 -2044 2124 -1984
rect 2700 -2044 2992 -1984
rect 3636 -2048 3928 -1988
<< metal1 >>
rect 1820 464 2136 470
rect 1820 404 1832 464
rect 2124 404 2136 464
rect 1820 398 2136 404
rect 2688 464 3004 470
rect 2688 404 2700 464
rect 2992 404 3004 464
rect 2688 398 3004 404
rect 3624 464 3940 470
rect 3624 404 3636 464
rect 3928 404 3940 464
rect 3624 398 3940 404
rect 1528 260 3772 368
rect 1694 204 1762 216
rect 1694 -144 1700 204
rect 1756 -144 1762 204
rect 1926 52 1936 232
rect 1988 52 1998 232
rect 2118 52 2128 232
rect 2180 52 2190 232
rect 2310 52 2320 232
rect 2372 52 2382 232
rect 2502 52 2512 232
rect 2564 52 2574 232
rect 2694 52 2704 232
rect 2756 52 2766 232
rect 2886 52 2896 232
rect 2948 52 2958 232
rect 3078 52 3088 232
rect 3140 52 3150 232
rect 3270 52 3280 232
rect 3332 52 3342 232
rect 3462 52 3472 232
rect 3524 52 3534 232
rect 3654 52 3664 232
rect 3716 52 3726 232
rect 3894 172 3966 184
rect 1694 -156 1762 -144
rect 1830 -172 1840 8
rect 1892 -172 1902 8
rect 2022 -172 2032 8
rect 2084 -172 2094 8
rect 2214 -172 2224 8
rect 2276 -172 2286 8
rect 2406 -172 2416 8
rect 2468 -172 2478 8
rect 2598 -172 2608 8
rect 2660 -172 2670 8
rect 2790 -172 2800 8
rect 2852 -172 2862 8
rect 2982 -172 2992 8
rect 3044 -172 3054 8
rect 3174 -172 3184 8
rect 3236 -172 3246 8
rect 3366 -172 3376 8
rect 3428 -172 3438 8
rect 3558 -172 3568 8
rect 3620 -172 3630 8
rect 3750 -172 3760 8
rect 3812 -172 3822 8
rect 3894 -84 3900 172
rect 3960 -84 3966 172
rect 3894 -96 3966 -84
rect 1528 -308 3676 -200
rect 1820 -352 2136 -346
rect 1820 -412 1832 -352
rect 2124 -412 2136 -352
rect 1820 -418 2136 -412
rect 2688 -352 3032 -346
rect 2688 -412 2700 -352
rect 3020 -412 3032 -352
rect 2688 -418 3032 -412
rect 3624 -348 3940 -342
rect 3624 -408 3636 -348
rect 3928 -408 3940 -348
rect 3624 -414 3940 -408
rect 1528 -560 3772 -456
rect 1694 -656 1766 -644
rect 1694 -912 1700 -656
rect 1760 -912 1766 -656
rect 1926 -768 1936 -588
rect 1988 -768 1998 -588
rect 2118 -768 2128 -588
rect 2180 -768 2190 -588
rect 2310 -768 2320 -588
rect 2372 -768 2382 -588
rect 2502 -768 2512 -588
rect 2564 -768 2574 -588
rect 2694 -768 2704 -588
rect 2756 -768 2766 -588
rect 2886 -768 2896 -588
rect 2948 -768 2958 -588
rect 3078 -768 3088 -588
rect 3140 -768 3150 -588
rect 3270 -768 3280 -588
rect 3332 -768 3342 -588
rect 3462 -768 3472 -588
rect 3524 -768 3534 -588
rect 3654 -768 3664 -588
rect 3716 -768 3726 -588
rect 3894 -676 3966 -664
rect 1694 -924 1766 -912
rect 1830 -992 1840 -812
rect 1892 -992 1902 -812
rect 2022 -992 2032 -812
rect 2084 -992 2094 -812
rect 2214 -992 2224 -812
rect 2276 -992 2286 -812
rect 2406 -992 2416 -812
rect 2468 -992 2478 -812
rect 2598 -992 2608 -812
rect 2660 -992 2670 -812
rect 2790 -992 2800 -812
rect 2852 -992 2862 -812
rect 2982 -992 2992 -812
rect 3044 -992 3054 -812
rect 3174 -992 3184 -812
rect 3236 -992 3246 -812
rect 3366 -992 3376 -812
rect 3428 -992 3438 -812
rect 3558 -992 3568 -812
rect 3620 -992 3630 -812
rect 3750 -992 3760 -812
rect 3812 -992 3822 -812
rect 3894 -932 3900 -676
rect 3960 -932 3966 -676
rect 3894 -944 3966 -932
rect 1528 -1128 3676 -1020
rect 1820 -1172 2136 -1166
rect 1820 -1232 1832 -1172
rect 2124 -1232 2136 -1172
rect 1820 -1238 2136 -1232
rect 2688 -1172 3004 -1166
rect 2688 -1232 2700 -1172
rect 2992 -1232 3004 -1172
rect 2688 -1238 3004 -1232
rect 3624 -1172 3940 -1166
rect 3624 -1232 3636 -1172
rect 3928 -1232 3940 -1172
rect 3624 -1238 3940 -1232
rect 1528 -1380 3772 -1272
rect 1690 -1496 1762 -1484
rect 1690 -1752 1696 -1496
rect 1756 -1752 1762 -1496
rect 1926 -1588 1936 -1408
rect 1988 -1588 1998 -1408
rect 2118 -1588 2128 -1408
rect 2180 -1588 2190 -1408
rect 2310 -1588 2320 -1408
rect 2372 -1588 2382 -1408
rect 2502 -1588 2512 -1408
rect 2564 -1588 2574 -1408
rect 2694 -1588 2704 -1408
rect 2756 -1588 2766 -1408
rect 2886 -1588 2896 -1408
rect 2948 -1588 2958 -1408
rect 3078 -1588 3088 -1408
rect 3140 -1588 3150 -1408
rect 3270 -1588 3280 -1408
rect 3332 -1588 3342 -1408
rect 3462 -1588 3472 -1408
rect 3524 -1588 3534 -1408
rect 3654 -1588 3664 -1408
rect 3716 -1588 3726 -1408
rect 3894 -1488 3966 -1476
rect 1690 -1764 1762 -1752
rect 1830 -1812 1840 -1632
rect 1892 -1812 1902 -1632
rect 2022 -1812 2032 -1632
rect 2084 -1812 2094 -1632
rect 2214 -1812 2224 -1632
rect 2276 -1812 2286 -1632
rect 2406 -1812 2416 -1632
rect 2468 -1812 2478 -1632
rect 2598 -1812 2608 -1632
rect 2660 -1812 2670 -1632
rect 2790 -1812 2800 -1632
rect 2852 -1812 2862 -1632
rect 2982 -1812 2992 -1632
rect 3044 -1812 3054 -1632
rect 3174 -1812 3184 -1632
rect 3236 -1812 3246 -1632
rect 3366 -1812 3376 -1632
rect 3428 -1812 3438 -1632
rect 3558 -1812 3568 -1632
rect 3620 -1812 3630 -1632
rect 3750 -1812 3760 -1632
rect 3812 -1812 3822 -1632
rect 3894 -1744 3900 -1488
rect 3960 -1744 3966 -1488
rect 3894 -1756 3966 -1744
rect 1528 -1948 3676 -1840
rect 1820 -1984 2136 -1978
rect 1820 -2044 1832 -1984
rect 2124 -2044 2136 -1984
rect 1820 -2050 2136 -2044
rect 2688 -1984 3004 -1978
rect 2688 -2044 2700 -1984
rect 2992 -2044 3004 -1984
rect 2688 -2050 3004 -2044
rect 3624 -1988 3940 -1982
rect 3624 -2048 3636 -1988
rect 3928 -2048 3940 -1988
rect 3624 -2054 3940 -2048
<< via1 >>
rect 1936 52 1988 232
rect 2128 52 2180 232
rect 2320 52 2372 232
rect 2512 52 2564 232
rect 2704 52 2756 232
rect 2896 52 2948 232
rect 3088 52 3140 232
rect 3280 52 3332 232
rect 3472 52 3524 232
rect 3664 52 3716 232
rect 1840 -172 1892 8
rect 2032 -172 2084 8
rect 2224 -172 2276 8
rect 2416 -172 2468 8
rect 2608 -172 2660 8
rect 2800 -172 2852 8
rect 2992 -172 3044 8
rect 3184 -172 3236 8
rect 3376 -172 3428 8
rect 3568 -172 3620 8
rect 3760 -172 3812 8
rect 1936 -768 1988 -588
rect 2128 -768 2180 -588
rect 2320 -768 2372 -588
rect 2512 -768 2564 -588
rect 2704 -768 2756 -588
rect 2896 -768 2948 -588
rect 3088 -768 3140 -588
rect 3280 -768 3332 -588
rect 3472 -768 3524 -588
rect 3664 -768 3716 -588
rect 1840 -992 1892 -812
rect 2032 -992 2084 -812
rect 2224 -992 2276 -812
rect 2416 -992 2468 -812
rect 2608 -992 2660 -812
rect 2800 -992 2852 -812
rect 2992 -992 3044 -812
rect 3184 -992 3236 -812
rect 3376 -992 3428 -812
rect 3568 -992 3620 -812
rect 3760 -992 3812 -812
rect 1936 -1588 1988 -1408
rect 2128 -1588 2180 -1408
rect 2320 -1588 2372 -1408
rect 2512 -1588 2564 -1408
rect 2704 -1588 2756 -1408
rect 2896 -1588 2948 -1408
rect 3088 -1588 3140 -1408
rect 3280 -1588 3332 -1408
rect 3472 -1588 3524 -1408
rect 3664 -1588 3716 -1408
rect 1840 -1812 1892 -1632
rect 2032 -1812 2084 -1632
rect 2224 -1812 2276 -1632
rect 2416 -1812 2468 -1632
rect 2608 -1812 2660 -1632
rect 2800 -1812 2852 -1632
rect 2992 -1812 3044 -1632
rect 3184 -1812 3236 -1632
rect 3376 -1812 3428 -1632
rect 3568 -1812 3620 -1632
rect 3760 -1812 3812 -1632
<< metal2 >>
rect 1936 232 1988 242
rect 1936 42 1988 52
rect 2128 232 2180 242
rect 2128 42 2180 52
rect 2320 232 2372 242
rect 2320 42 2372 52
rect 2512 232 2564 242
rect 2512 42 2564 52
rect 2704 232 2756 242
rect 2704 42 2756 52
rect 2896 232 2948 242
rect 2896 42 2948 52
rect 3088 232 3140 242
rect 3088 42 3140 52
rect 3280 232 3332 242
rect 3280 42 3332 52
rect 3472 232 3524 242
rect 3472 42 3524 52
rect 3664 232 3716 242
rect 3664 42 3716 52
rect 1840 8 1892 18
rect 1840 -182 1892 -172
rect 2032 8 2084 18
rect 2032 -182 2084 -172
rect 2224 8 2276 18
rect 2224 -182 2276 -172
rect 2416 8 2468 18
rect 2416 -182 2468 -172
rect 2608 8 2660 18
rect 2608 -182 2660 -172
rect 2800 8 2852 18
rect 2800 -182 2852 -172
rect 2992 8 3044 18
rect 2992 -182 3044 -172
rect 3184 8 3236 18
rect 3184 -182 3236 -172
rect 3376 8 3428 18
rect 3376 -182 3428 -172
rect 3568 8 3620 18
rect 3568 -182 3620 -172
rect 3760 8 3812 18
rect 3760 -182 3812 -172
rect 1936 -588 1988 -578
rect 1936 -778 1988 -768
rect 2128 -588 2180 -578
rect 2128 -778 2180 -768
rect 2320 -588 2372 -578
rect 2320 -778 2372 -768
rect 2512 -588 2564 -578
rect 2512 -778 2564 -768
rect 2704 -588 2756 -578
rect 2704 -778 2756 -768
rect 2896 -588 2948 -578
rect 2896 -778 2948 -768
rect 3088 -588 3140 -578
rect 3088 -778 3140 -768
rect 3280 -588 3332 -578
rect 3280 -778 3332 -768
rect 3472 -588 3524 -578
rect 3472 -778 3524 -768
rect 3664 -588 3716 -578
rect 3664 -778 3716 -768
rect 1840 -812 1892 -802
rect 1840 -1002 1892 -992
rect 2032 -812 2084 -802
rect 2032 -1002 2084 -992
rect 2224 -812 2276 -802
rect 2224 -1002 2276 -992
rect 2416 -812 2468 -802
rect 2416 -1002 2468 -992
rect 2608 -812 2660 -802
rect 2608 -1002 2660 -992
rect 2800 -812 2852 -802
rect 2800 -1002 2852 -992
rect 2992 -812 3044 -802
rect 2992 -1002 3044 -992
rect 3184 -812 3236 -802
rect 3184 -1002 3236 -992
rect 3376 -812 3428 -802
rect 3376 -1002 3428 -992
rect 3568 -812 3620 -802
rect 3568 -1002 3620 -992
rect 3760 -812 3812 -802
rect 3760 -1002 3812 -992
rect 1936 -1408 1988 -1398
rect 1936 -1598 1988 -1588
rect 2128 -1408 2180 -1398
rect 2128 -1598 2180 -1588
rect 2320 -1408 2372 -1398
rect 2320 -1598 2372 -1588
rect 2512 -1408 2564 -1398
rect 2512 -1598 2564 -1588
rect 2704 -1408 2756 -1398
rect 2704 -1598 2756 -1588
rect 2896 -1408 2948 -1398
rect 2896 -1598 2948 -1588
rect 3088 -1408 3140 -1398
rect 3088 -1598 3140 -1588
rect 3280 -1408 3332 -1398
rect 3280 -1598 3332 -1588
rect 3472 -1408 3524 -1398
rect 3472 -1598 3524 -1588
rect 3664 -1408 3716 -1398
rect 3664 -1598 3716 -1588
rect 1840 -1632 1892 -1622
rect 1840 -1822 1892 -1812
rect 2032 -1632 2084 -1622
rect 2032 -1822 2084 -1812
rect 2224 -1632 2276 -1622
rect 2224 -1822 2276 -1812
rect 2416 -1632 2468 -1622
rect 2416 -1822 2468 -1812
rect 2608 -1632 2660 -1622
rect 2608 -1822 2660 -1812
rect 2800 -1632 2852 -1622
rect 2800 -1822 2852 -1812
rect 2992 -1632 3044 -1622
rect 2992 -1822 3044 -1812
rect 3184 -1632 3236 -1622
rect 3184 -1822 3236 -1812
rect 3376 -1632 3428 -1622
rect 3376 -1822 3428 -1812
rect 3568 -1632 3620 -1622
rect 3568 -1822 3620 -1812
rect 3760 -1632 3812 -1622
rect 3760 -1822 3812 -1812
use sky130_fd_pr__nfet_01v8_lvt_SDPJLJ  sky130_fd_pr__nfet_01v8_lvt_SDPJLJ_0
timestamp 1686659968
transform 1 0 2827 0 1 -790
box -1127 -410 1127 410
use sky130_fd_pr__nfet_01v8_lvt_SDPJLJ  sky130_fd_pr__nfet_01v8_lvt_SDPJLJ_1
timestamp 1686659968
transform 1 0 2827 0 1 -1610
box -1127 -410 1127 410
use sky130_fd_pr__nfet_01v8_lvt_SDPJLJ  sky130_fd_pr__nfet_01v8_lvt_SDPJLJ_2
timestamp 1686659968
transform 1 0 2827 0 1 30
box -1127 -410 1127 410
<< end >>
