magic
tech sky130A
magscale 1 2
timestamp 1683557511
<< nwell >>
rect -3673 127 -2407 709
rect -2153 127 -887 709
rect -633 127 633 709
rect 887 127 2153 709
rect 2407 127 3673 709
rect -3673 -709 -2407 -127
rect -2153 -709 -887 -127
rect -633 -709 633 -127
rect 887 -709 2153 -127
rect 2407 -709 3673 -127
<< pwell >>
rect -3783 709 3783 819
rect -3783 127 -3673 709
rect -2407 127 -2153 709
rect -887 127 -633 709
rect 633 127 887 709
rect 2153 127 2407 709
rect 3673 127 3783 709
rect -3783 -127 3783 127
rect -3783 -709 -3673 -127
rect -2407 -709 -2153 -127
rect -887 -709 -633 -127
rect 633 -709 887 -127
rect 2153 -709 2407 -127
rect 3673 -709 3783 -127
rect -3783 -819 3783 -709
<< varactor >>
rect -3540 218 -2540 618
rect -2020 218 -1020 618
rect -500 218 500 618
rect 1020 218 2020 618
rect 2540 218 3540 618
rect -3540 -618 -2540 -218
rect -2020 -618 -1020 -218
rect -500 -618 500 -218
rect 1020 -618 2020 -218
rect 2540 -618 3540 -218
<< psubdiff >>
rect -3747 749 -3651 783
rect 3651 749 3747 783
rect -3747 687 -3713 749
rect 3713 687 3747 749
rect -3747 -749 -3713 -687
rect 3713 -749 3747 -687
rect -3747 -783 -3651 -749
rect 3651 -783 3747 -749
<< nsubdiff >>
rect -3637 594 -3540 618
rect -3637 242 -3625 594
rect -3591 242 -3540 594
rect -3637 218 -3540 242
rect -2540 594 -2443 618
rect -2540 242 -2489 594
rect -2455 242 -2443 594
rect -2540 218 -2443 242
rect -2117 594 -2020 618
rect -2117 242 -2105 594
rect -2071 242 -2020 594
rect -2117 218 -2020 242
rect -1020 594 -923 618
rect -1020 242 -969 594
rect -935 242 -923 594
rect -1020 218 -923 242
rect -597 594 -500 618
rect -597 242 -585 594
rect -551 242 -500 594
rect -597 218 -500 242
rect 500 594 597 618
rect 500 242 551 594
rect 585 242 597 594
rect 500 218 597 242
rect 923 594 1020 618
rect 923 242 935 594
rect 969 242 1020 594
rect 923 218 1020 242
rect 2020 594 2117 618
rect 2020 242 2071 594
rect 2105 242 2117 594
rect 2020 218 2117 242
rect 2443 594 2540 618
rect 2443 242 2455 594
rect 2489 242 2540 594
rect 2443 218 2540 242
rect 3540 594 3637 618
rect 3540 242 3591 594
rect 3625 242 3637 594
rect 3540 218 3637 242
rect -3637 -242 -3540 -218
rect -3637 -594 -3625 -242
rect -3591 -594 -3540 -242
rect -3637 -618 -3540 -594
rect -2540 -242 -2443 -218
rect -2540 -594 -2489 -242
rect -2455 -594 -2443 -242
rect -2540 -618 -2443 -594
rect -2117 -242 -2020 -218
rect -2117 -594 -2105 -242
rect -2071 -594 -2020 -242
rect -2117 -618 -2020 -594
rect -1020 -242 -923 -218
rect -1020 -594 -969 -242
rect -935 -594 -923 -242
rect -1020 -618 -923 -594
rect -597 -242 -500 -218
rect -597 -594 -585 -242
rect -551 -594 -500 -242
rect -597 -618 -500 -594
rect 500 -242 597 -218
rect 500 -594 551 -242
rect 585 -594 597 -242
rect 500 -618 597 -594
rect 923 -242 1020 -218
rect 923 -594 935 -242
rect 969 -594 1020 -242
rect 923 -618 1020 -594
rect 2020 -242 2117 -218
rect 2020 -594 2071 -242
rect 2105 -594 2117 -242
rect 2020 -618 2117 -594
rect 2443 -242 2540 -218
rect 2443 -594 2455 -242
rect 2489 -594 2540 -242
rect 2443 -618 2540 -594
rect 3540 -242 3637 -218
rect 3540 -594 3591 -242
rect 3625 -594 3637 -242
rect 3540 -618 3637 -594
<< psubdiffcont >>
rect -3651 749 3651 783
rect -3747 -687 -3713 687
rect 3713 -687 3747 687
rect -3651 -783 3651 -749
<< nsubdiffcont >>
rect -3625 242 -3591 594
rect -2489 242 -2455 594
rect -2105 242 -2071 594
rect -969 242 -935 594
rect -585 242 -551 594
rect 551 242 585 594
rect 935 242 969 594
rect 2071 242 2105 594
rect 2455 242 2489 594
rect 3591 242 3625 594
rect -3625 -594 -3591 -242
rect -2489 -594 -2455 -242
rect -2105 -594 -2071 -242
rect -969 -594 -935 -242
rect -585 -594 -551 -242
rect 551 -594 585 -242
rect 935 -594 969 -242
rect 2071 -594 2105 -242
rect 2455 -594 2489 -242
rect 3591 -594 3625 -242
<< poly >>
rect -3540 690 -2540 706
rect -3540 656 -3524 690
rect -2556 656 -2540 690
rect -3540 618 -2540 656
rect -2020 690 -1020 706
rect -2020 656 -2004 690
rect -1036 656 -1020 690
rect -2020 618 -1020 656
rect -500 690 500 706
rect -500 656 -484 690
rect 484 656 500 690
rect -500 618 500 656
rect 1020 690 2020 706
rect 1020 656 1036 690
rect 2004 656 2020 690
rect 1020 618 2020 656
rect 2540 690 3540 706
rect 2540 656 2556 690
rect 3524 656 3540 690
rect 2540 618 3540 656
rect -3540 180 -2540 218
rect -3540 146 -3524 180
rect -2556 146 -2540 180
rect -3540 130 -2540 146
rect -2020 180 -1020 218
rect -2020 146 -2004 180
rect -1036 146 -1020 180
rect -2020 130 -1020 146
rect -500 180 500 218
rect -500 146 -484 180
rect 484 146 500 180
rect -500 130 500 146
rect 1020 180 2020 218
rect 1020 146 1036 180
rect 2004 146 2020 180
rect 1020 130 2020 146
rect 2540 180 3540 218
rect 2540 146 2556 180
rect 3524 146 3540 180
rect 2540 130 3540 146
rect -3540 -146 -2540 -130
rect -3540 -180 -3524 -146
rect -2556 -180 -2540 -146
rect -3540 -218 -2540 -180
rect -2020 -146 -1020 -130
rect -2020 -180 -2004 -146
rect -1036 -180 -1020 -146
rect -2020 -218 -1020 -180
rect -500 -146 500 -130
rect -500 -180 -484 -146
rect 484 -180 500 -146
rect -500 -218 500 -180
rect 1020 -146 2020 -130
rect 1020 -180 1036 -146
rect 2004 -180 2020 -146
rect 1020 -218 2020 -180
rect 2540 -146 3540 -130
rect 2540 -180 2556 -146
rect 3524 -180 3540 -146
rect 2540 -218 3540 -180
rect -3540 -656 -2540 -618
rect -3540 -690 -3524 -656
rect -2556 -690 -2540 -656
rect -3540 -706 -2540 -690
rect -2020 -656 -1020 -618
rect -2020 -690 -2004 -656
rect -1036 -690 -1020 -656
rect -2020 -706 -1020 -690
rect -500 -656 500 -618
rect -500 -690 -484 -656
rect 484 -690 500 -656
rect -500 -706 500 -690
rect 1020 -656 2020 -618
rect 1020 -690 1036 -656
rect 2004 -690 2020 -656
rect 1020 -706 2020 -690
rect 2540 -656 3540 -618
rect 2540 -690 2556 -656
rect 3524 -690 3540 -656
rect 2540 -706 3540 -690
<< polycont >>
rect -3524 656 -2556 690
rect -2004 656 -1036 690
rect -484 656 484 690
rect 1036 656 2004 690
rect 2556 656 3524 690
rect -3524 146 -2556 180
rect -2004 146 -1036 180
rect -484 146 484 180
rect 1036 146 2004 180
rect 2556 146 3524 180
rect -3524 -180 -2556 -146
rect -2004 -180 -1036 -146
rect -484 -180 484 -146
rect 1036 -180 2004 -146
rect 2556 -180 3524 -146
rect -3524 -690 -2556 -656
rect -2004 -690 -1036 -656
rect -484 -690 484 -656
rect 1036 -690 2004 -656
rect 2556 -690 3524 -656
<< locali >>
rect -3747 749 -3651 783
rect 3651 749 3747 783
rect -3747 687 -3713 749
rect -3540 656 -3524 690
rect -2556 656 -2540 690
rect -2020 656 -2004 690
rect -1036 656 -1020 690
rect -500 656 -484 690
rect 484 656 500 690
rect 1020 656 1036 690
rect 2004 656 2020 690
rect 2540 656 2556 690
rect 3524 656 3540 690
rect 3713 687 3747 749
rect -3625 594 -3591 610
rect -3625 226 -3591 242
rect -2489 594 -2455 610
rect -2489 226 -2455 242
rect -2105 594 -2071 610
rect -2105 226 -2071 242
rect -969 594 -935 610
rect -969 226 -935 242
rect -585 594 -551 610
rect -585 226 -551 242
rect 551 594 585 610
rect 551 226 585 242
rect 935 594 969 610
rect 935 226 969 242
rect 2071 594 2105 610
rect 2071 226 2105 242
rect 2455 594 2489 610
rect 2455 226 2489 242
rect 3591 594 3625 610
rect 3591 226 3625 242
rect -3540 146 -3524 180
rect -2556 146 -2540 180
rect -2020 146 -2004 180
rect -1036 146 -1020 180
rect -500 146 -484 180
rect 484 146 500 180
rect 1020 146 1036 180
rect 2004 146 2020 180
rect 2540 146 2556 180
rect 3524 146 3540 180
rect -3540 -180 -3524 -146
rect -2556 -180 -2540 -146
rect -2020 -180 -2004 -146
rect -1036 -180 -1020 -146
rect -500 -180 -484 -146
rect 484 -180 500 -146
rect 1020 -180 1036 -146
rect 2004 -180 2020 -146
rect 2540 -180 2556 -146
rect 3524 -180 3540 -146
rect -3625 -242 -3591 -226
rect -3625 -610 -3591 -594
rect -2489 -242 -2455 -226
rect -2489 -610 -2455 -594
rect -2105 -242 -2071 -226
rect -2105 -610 -2071 -594
rect -969 -242 -935 -226
rect -969 -610 -935 -594
rect -585 -242 -551 -226
rect -585 -610 -551 -594
rect 551 -242 585 -226
rect 551 -610 585 -594
rect 935 -242 969 -226
rect 935 -610 969 -594
rect 2071 -242 2105 -226
rect 2071 -610 2105 -594
rect 2455 -242 2489 -226
rect 2455 -610 2489 -594
rect 3591 -242 3625 -226
rect 3591 -610 3625 -594
rect -3747 -749 -3713 -687
rect -3540 -690 -3524 -656
rect -2556 -690 -2540 -656
rect -2020 -690 -2004 -656
rect -1036 -690 -1020 -656
rect -500 -690 -484 -656
rect 484 -690 500 -656
rect 1020 -690 1036 -656
rect 2004 -690 2020 -656
rect 2540 -690 2556 -656
rect 3524 -690 3540 -656
rect 3713 -749 3747 -687
rect -3747 -783 -3651 -749
rect 3651 -783 3747 -749
<< viali >>
rect -3524 656 -2556 690
rect -2004 656 -1036 690
rect -484 656 484 690
rect 1036 656 2004 690
rect 2556 656 3524 690
rect -3625 242 -3591 594
rect -2489 242 -2455 594
rect -2105 242 -2071 594
rect -969 242 -935 594
rect -585 242 -551 594
rect 551 242 585 594
rect 935 242 969 594
rect 2071 242 2105 594
rect 2455 242 2489 594
rect 3591 242 3625 594
rect -3524 146 -2556 180
rect -2004 146 -1036 180
rect -484 146 484 180
rect 1036 146 2004 180
rect 2556 146 3524 180
rect -3524 -180 -2556 -146
rect -2004 -180 -1036 -146
rect -484 -180 484 -146
rect 1036 -180 2004 -146
rect 2556 -180 3524 -146
rect -3625 -594 -3591 -242
rect -2489 -594 -2455 -242
rect -2105 -594 -2071 -242
rect -969 -594 -935 -242
rect -585 -594 -551 -242
rect 551 -594 585 -242
rect 935 -594 969 -242
rect 2071 -594 2105 -242
rect 2455 -594 2489 -242
rect 3591 -594 3625 -242
rect -3524 -690 -2556 -656
rect -2004 -690 -1036 -656
rect -484 -690 484 -656
rect 1036 -690 2004 -656
rect 2556 -690 3524 -656
<< metal1 >>
rect -3536 690 -2544 696
rect -3536 656 -3524 690
rect -2556 656 -2544 690
rect -3536 650 -2544 656
rect -2016 690 -1024 696
rect -2016 656 -2004 690
rect -1036 656 -1024 690
rect -2016 650 -1024 656
rect -496 690 496 696
rect -496 656 -484 690
rect 484 656 496 690
rect -496 650 496 656
rect 1024 690 2016 696
rect 1024 656 1036 690
rect 2004 656 2016 690
rect 1024 650 2016 656
rect 2544 690 3536 696
rect 2544 656 2556 690
rect 3524 656 3536 690
rect 2544 650 3536 656
rect -3631 594 -3585 606
rect -2495 594 -2449 606
rect -3631 242 -3625 594
rect -3591 242 -2489 594
rect -2455 242 -2449 594
rect -3631 230 -3585 242
rect -2495 230 -2449 242
rect -2111 594 -2065 606
rect -975 594 -929 606
rect -2111 242 -2105 594
rect -2071 242 -969 594
rect -935 242 -929 594
rect -2111 230 -2065 242
rect -975 230 -929 242
rect -591 594 -545 606
rect 545 594 591 606
rect -591 242 -585 594
rect -551 242 551 594
rect 585 242 591 594
rect -591 230 -545 242
rect 545 230 591 242
rect 929 594 975 606
rect 2065 594 2111 606
rect 929 242 935 594
rect 969 242 2071 594
rect 2105 242 2111 594
rect 929 230 975 242
rect 2065 230 2111 242
rect 2449 594 2495 606
rect 3585 594 3631 606
rect 2449 242 2455 594
rect 2489 242 3591 594
rect 3625 242 3631 594
rect 2449 230 2495 242
rect 3585 230 3631 242
rect -3536 180 -2544 186
rect -3536 146 -3524 180
rect -2556 146 -2544 180
rect -3536 140 -2544 146
rect -2016 180 -1024 186
rect -2016 146 -2004 180
rect -1036 146 -1024 180
rect -2016 140 -1024 146
rect -496 180 496 186
rect -496 146 -484 180
rect 484 146 496 180
rect -496 140 496 146
rect 1024 180 2016 186
rect 1024 146 1036 180
rect 2004 146 2016 180
rect 1024 140 2016 146
rect 2544 180 3536 186
rect 2544 146 2556 180
rect 3524 146 3536 180
rect 2544 140 3536 146
rect -3536 -146 -2544 -140
rect -3536 -180 -3524 -146
rect -2556 -180 -2544 -146
rect -3536 -186 -2544 -180
rect -2016 -146 -1024 -140
rect -2016 -180 -2004 -146
rect -1036 -180 -1024 -146
rect -2016 -186 -1024 -180
rect -496 -146 496 -140
rect -496 -180 -484 -146
rect 484 -180 496 -146
rect -496 -186 496 -180
rect 1024 -146 2016 -140
rect 1024 -180 1036 -146
rect 2004 -180 2016 -146
rect 1024 -186 2016 -180
rect 2544 -146 3536 -140
rect 2544 -180 2556 -146
rect 3524 -180 3536 -146
rect 2544 -186 3536 -180
rect -3631 -242 -3585 -230
rect -2495 -242 -2449 -230
rect -3631 -594 -3625 -242
rect -3591 -594 -2489 -242
rect -2455 -594 -2449 -242
rect -3631 -606 -3585 -594
rect -2495 -606 -2449 -594
rect -2111 -242 -2065 -230
rect -975 -242 -929 -230
rect -2111 -594 -2105 -242
rect -2071 -594 -969 -242
rect -935 -594 -929 -242
rect -2111 -606 -2065 -594
rect -975 -606 -929 -594
rect -591 -242 -545 -230
rect 545 -242 591 -230
rect -591 -594 -585 -242
rect -551 -594 551 -242
rect 585 -594 591 -242
rect -591 -606 -545 -594
rect 545 -606 591 -594
rect 929 -242 975 -230
rect 2065 -242 2111 -230
rect 929 -594 935 -242
rect 969 -594 2071 -242
rect 2105 -594 2111 -242
rect 929 -606 975 -594
rect 2065 -606 2111 -594
rect 2449 -242 2495 -230
rect 3585 -242 3631 -230
rect 2449 -594 2455 -242
rect 2489 -594 3591 -242
rect 3625 -594 3631 -242
rect 2449 -606 2495 -594
rect 3585 -606 3631 -594
rect -3536 -656 -2544 -650
rect -3536 -690 -3524 -656
rect -2556 -690 -2544 -656
rect -3536 -696 -2544 -690
rect -2016 -656 -1024 -650
rect -2016 -690 -2004 -656
rect -1036 -690 -1024 -656
rect -2016 -696 -1024 -690
rect -496 -656 496 -650
rect -496 -690 -484 -656
rect 484 -690 496 -656
rect -496 -696 496 -690
rect 1024 -656 2016 -650
rect 1024 -690 1036 -656
rect 2004 -690 2016 -656
rect 1024 -696 2016 -690
rect 2544 -656 3536 -650
rect 2544 -690 2556 -656
rect 3524 -690 3536 -656
rect 2544 -696 3536 -690
<< properties >>
string FIXED_BBOX -3730 -766 3730 766
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 5 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
