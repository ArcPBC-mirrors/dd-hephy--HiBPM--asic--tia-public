magic
tech sky130A
magscale 1 2
timestamp 1684500887
<< metal1 >>
rect 18270 24600 18280 25120
rect 18640 24600 18650 25120
rect 19030 25040 19040 25260
rect 19240 25040 19250 25260
rect 8964 21556 18208 21688
rect 8964 21460 18224 21556
rect 10320 21220 11900 21300
rect 10320 20860 10380 21220
rect 10840 20860 11900 21220
rect 10320 20780 11900 20860
rect 9400 17280 9600 17720
rect 9400 16980 10160 17280
rect -3192 4532 -3008 4568
rect -3192 4420 -3172 4532
rect -3028 4420 -3008 4532
rect -3192 4200 -3008 4420
rect 9840 4200 10160 16980
rect 10800 7928 11300 17712
rect 11480 11940 11900 20780
rect 11480 11500 24900 11940
rect 10790 7472 10800 7928
rect 11300 7472 11310 7928
rect 11480 4920 11900 11500
rect 11400 4860 11900 4920
rect 11400 4580 11480 4860
rect 11820 4580 11900 4860
rect 24520 4700 24900 11500
rect 11400 4520 11900 4580
rect 11480 4500 11900 4520
rect 24510 4360 24520 4700
rect 24900 4360 24910 4700
rect -3192 4048 80 4200
rect -3224 3780 80 4048
rect 7040 3780 14220 4200
rect 24520 3420 24900 4360
<< via1 >>
rect 18280 24600 18640 25120
rect 19040 25040 19240 25260
rect 10380 20860 10840 21220
rect -3172 4420 -3028 4532
rect 10800 7472 11300 7928
rect 11480 4580 11820 4860
rect 24520 4360 24900 4700
<< metal2 >>
rect 18940 25260 19360 25280
rect 18280 25120 18640 25130
rect 18280 24590 18640 24600
rect 18940 25040 19040 25260
rect 19240 25040 19360 25260
rect 18940 24420 19360 25040
rect 17480 24040 19360 24420
rect 17480 23300 17840 24040
rect 15900 22940 17840 23300
rect 15900 22180 16300 22940
rect 15900 21730 16300 21740
rect 24560 21500 24880 21510
rect 10380 21220 10840 21230
rect 24880 21140 25620 21500
rect 24560 21130 24880 21140
rect 10380 20850 10840 20860
rect 15580 18860 15980 18870
rect 15580 18410 15980 18420
rect 15620 11760 15980 18410
rect 1980 11400 15980 11760
rect 16220 18860 16620 18870
rect 1980 9800 2300 11400
rect -10000 8800 -8800 9400
rect -3300 9120 2320 9800
rect 16220 9120 16620 18420
rect 21460 9780 21490 10040
rect -9200 8200 -8860 8800
rect 10800 7928 11300 7938
rect 10580 7472 10800 7600
rect 11300 7472 12028 7580
rect -3090 6270 -2352 6910
rect 10580 6140 12028 7472
rect 11130 6130 12028 6140
rect 11480 4860 11820 4870
rect 11480 4570 11820 4580
rect 24520 4700 24900 4710
rect -3172 4532 -3028 4542
rect -3172 4410 -3028 4420
rect 24520 4350 24900 4360
<< via2 >>
rect 18280 24600 18640 25120
rect 15900 21740 16300 22180
rect 10380 20860 10840 21220
rect 24560 21140 24880 21500
rect 15580 18420 15980 18860
rect 16220 18420 16620 18860
rect 11480 4580 11820 4860
rect -3172 4420 -3028 4532
rect 24520 4360 24900 4700
<< metal3 >>
rect 6460 27440 28460 29380
rect 18220 25120 18680 27440
rect 18220 24600 18280 25120
rect 18640 24600 18680 25120
rect 18220 24560 18680 24600
rect 15890 22180 16310 22185
rect 15890 21740 15900 22180
rect 16300 21740 16310 22180
rect 15890 21735 16310 21740
rect 24550 21500 24890 21505
rect 10370 21220 10850 21225
rect 10370 20860 10380 21220
rect 10840 20860 10850 21220
rect 23980 21140 24560 21500
rect 24880 21140 24890 21500
rect 24550 21135 24890 21140
rect 10370 20855 10850 20860
rect 15570 18860 15990 18865
rect 15570 18420 15580 18860
rect 15980 18420 15990 18860
rect 15570 18415 15990 18420
rect 16210 18860 16630 18865
rect 16210 18420 16220 18860
rect 16620 18420 16630 18860
rect 16210 18415 16630 18420
rect 18290 17720 18300 18180
rect 18900 17720 18910 18180
rect 26380 14740 28460 27440
rect -10460 10740 28460 14740
rect -1860 9960 -540 10740
rect 12540 10000 13920 10740
rect 24540 10720 28460 10740
rect 5110 8740 5120 9180
rect 6060 8740 6070 9180
rect 10200 4860 11860 4900
rect 10200 4580 11480 4860
rect 11820 4580 11860 4860
rect -3182 4532 -3018 4537
rect -3182 4420 -3172 4532
rect -3028 4420 -3018 4532
rect -3182 4415 -3018 4420
rect 10200 4520 11860 4580
rect 24510 4700 24910 4705
rect 10200 4060 10520 4520
rect 24510 4360 24520 4700
rect 24900 4360 24910 4700
rect 24510 4355 24910 4360
rect 24520 3440 24900 4355
<< via3 >>
rect 15900 21740 16300 22180
rect 15580 18420 15980 18860
rect 16220 18420 16620 18860
rect 18300 17720 18900 18180
rect 5120 8740 6060 9180
rect -3172 4420 -3028 4532
<< metal4 >>
rect 15899 22180 16301 22181
rect 15899 21740 15900 22180
rect 16300 21740 16301 22180
rect 15899 21739 16301 21740
rect 15900 20520 16300 21739
rect 15580 18861 15980 20000
rect 16220 18861 16620 20000
rect 15579 18860 15981 18861
rect 15579 18420 15580 18860
rect 15980 18420 15981 18860
rect 15579 18419 15981 18420
rect 16219 18860 16621 18861
rect 16219 18420 16220 18860
rect 16620 18420 16621 18860
rect 16219 18419 16621 18420
rect 18299 18180 18901 18181
rect 18299 17720 18300 18180
rect 18900 17720 18901 18180
rect 18299 17719 18901 17720
rect 18300 17480 18900 17719
rect 19992 17480 21096 18848
rect 6660 15540 28600 17480
rect 5120 9181 10640 9460
rect 5119 9180 10640 9181
rect 5119 8740 5120 9180
rect 6060 8740 10640 9180
rect 5119 8739 6061 8740
rect -3192 4532 -3008 4568
rect -3192 4420 -3172 4532
rect -3028 4420 -3008 4532
rect -3192 4368 -3008 4420
rect -3884 4272 -3008 4368
rect -8520 280 -8340 540
rect -9320 -80 -7620 280
rect 26000 -80 28600 15540
rect -10640 -4080 28600 -80
use curr_filter  curr_filter_0
timestamp 1684252655
transform 1 0 -11340 0 1 148
box 1140 -148 7552 8540
use tia_bias  tia_bias_1
timestamp 1684252655
transform 1 0 6460 0 1 23756
box -120 -6836 10684 4104
use tia_core  tia_core_0
timestamp 1684500887
transform 1 0 17076 0 1 8228
box -6076 -9628 7964 3244
use tia_core  tia_core_1
timestamp 1684500887
transform 1 0 2676 0 1 8228
box -6076 -9628 7964 3244
use tia_outfilter  tia_outfilter_0
timestamp 1684252655
transform 1 0 18220 0 1 21076
box -160 -3030 6012 6060
<< labels >>
rlabel metal3 -10000 12200 -8800 13600 1 VP
port 1 n
rlabel metal2 -10000 8800 -9600 9400 1 I_Bias1
port 6 n
rlabel metal4 -10400 -2800 -9600 -1400 1 VN
port 7 n
rlabel metal2 10600 6400 11200 7400 1 Input_ref
port 4 n
rlabel metal2 -3020 6340 -2520 6830 1 Input
port 5 n
rlabel metal1 9884 5220 10104 5448 1 VM9G
rlabel metal2 -3220 9220 -2700 9740 1 Out_2
port 8 n
rlabel metal4 15940 20560 16260 21000 1 Filter_in
port 10 n
rlabel metal2 24960 21180 25560 21460 1 Filter_out
port 12 n
rlabel metal4 16260 19520 16580 19960 1 Out_ref
port 13 n
<< end >>
