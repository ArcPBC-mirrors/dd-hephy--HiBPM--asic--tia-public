magic
tech sky130A
magscale 1 2
timestamp 1683564698
<< error_p >>
rect -3570 2345 -2510 2372
rect -2050 2345 -990 2372
rect -530 2345 530 2372
rect 990 2345 2050 2372
rect 2510 2345 3570 2372
rect -3570 1336 -2510 1363
rect -2050 1336 -990 1363
rect -530 1336 530 1363
rect 990 1336 2050 1363
rect 2510 1336 3570 1363
rect -3570 1109 -2510 1136
rect -2050 1109 -990 1136
rect -530 1109 530 1136
rect 990 1109 2050 1136
rect 2510 1109 3570 1136
rect -3570 100 -2510 127
rect -2050 100 -990 127
rect -530 100 530 127
rect 990 100 2050 127
rect 2510 100 3570 127
rect -3570 -127 -2510 -100
rect -2050 -127 -990 -100
rect -530 -127 530 -100
rect 990 -127 2050 -100
rect 2510 -127 3570 -100
rect -3570 -1136 -2510 -1109
rect -2050 -1136 -990 -1109
rect -530 -1136 530 -1109
rect 990 -1136 2050 -1109
rect 2510 -1136 3570 -1109
rect -3570 -1363 -2510 -1336
rect -2050 -1363 -990 -1336
rect -530 -1363 530 -1336
rect 990 -1363 2050 -1336
rect 2510 -1363 3570 -1336
rect -3570 -2372 -2510 -2345
rect -2050 -2372 -990 -2345
rect -530 -2372 530 -2345
rect 990 -2372 2050 -2345
rect 2510 -2372 3570 -2345
<< nwell >>
rect -3673 1363 -2407 2345
rect -2153 1363 -887 2345
rect -633 1363 633 2345
rect 887 1363 2153 2345
rect 2407 1363 3673 2345
rect -3673 127 -2407 1109
rect -2153 127 -887 1109
rect -633 127 633 1109
rect 887 127 2153 1109
rect 2407 127 3673 1109
rect -3673 -1109 -2407 -127
rect -2153 -1109 -887 -127
rect -633 -1109 633 -127
rect 887 -1109 2153 -127
rect 2407 -1109 3673 -127
rect -3673 -2345 -2407 -1363
rect -2153 -2345 -887 -1363
rect -633 -2345 633 -1363
rect 887 -2345 2153 -1363
rect 2407 -2345 3673 -1363
<< pwell >>
rect -3783 2345 3783 2455
rect -3783 1363 -3673 2345
rect -2407 1363 -2153 2345
rect -887 1363 -633 2345
rect 633 1363 887 2345
rect 2153 1363 2407 2345
rect 3673 1363 3783 2345
rect -3783 1109 3783 1363
rect -3783 127 -3673 1109
rect -2407 127 -2153 1109
rect -887 127 -633 1109
rect 633 127 887 1109
rect 2153 127 2407 1109
rect 3673 127 3783 1109
rect -3783 -127 3783 127
rect -3783 -1109 -3673 -127
rect -2407 -1109 -2153 -127
rect -887 -1109 -633 -127
rect 633 -1109 887 -127
rect 2153 -1109 2407 -127
rect 3673 -1109 3783 -127
rect -3783 -1363 3783 -1109
rect -3783 -2345 -3673 -1363
rect -2407 -2345 -2153 -1363
rect -887 -2345 -633 -1363
rect 633 -2345 887 -1363
rect 2153 -2345 2407 -1363
rect 3673 -2345 3783 -1363
rect -3783 -2455 3783 -2345
<< varactor >>
rect -3540 1454 -2540 2254
rect -2020 1454 -1020 2254
rect -500 1454 500 2254
rect 1020 1454 2020 2254
rect 2540 1454 3540 2254
rect -3540 218 -2540 1018
rect -2020 218 -1020 1018
rect -500 218 500 1018
rect 1020 218 2020 1018
rect 2540 218 3540 1018
rect -3540 -1018 -2540 -218
rect -2020 -1018 -1020 -218
rect -500 -1018 500 -218
rect 1020 -1018 2020 -218
rect 2540 -1018 3540 -218
rect -3540 -2254 -2540 -1454
rect -2020 -2254 -1020 -1454
rect -500 -2254 500 -1454
rect 1020 -2254 2020 -1454
rect 2540 -2254 3540 -1454
<< psubdiff >>
rect -3747 2385 -3651 2419
rect 3651 2385 3747 2419
rect -3747 2323 -3713 2385
rect 3713 2323 3747 2385
rect -3747 -2385 -3713 -2323
rect 3713 -2385 3747 -2323
rect -3747 -2419 -3651 -2385
rect 3651 -2419 3747 -2385
<< nsubdiff >>
rect -3637 2230 -3540 2254
rect -3637 1478 -3625 2230
rect -3591 1478 -3540 2230
rect -3637 1454 -3540 1478
rect -2540 2230 -2443 2254
rect -2540 1478 -2489 2230
rect -2455 1478 -2443 2230
rect -2540 1454 -2443 1478
rect -2117 2230 -2020 2254
rect -2117 1478 -2105 2230
rect -2071 1478 -2020 2230
rect -2117 1454 -2020 1478
rect -1020 2230 -923 2254
rect -1020 1478 -969 2230
rect -935 1478 -923 2230
rect -1020 1454 -923 1478
rect -597 2230 -500 2254
rect -597 1478 -585 2230
rect -551 1478 -500 2230
rect -597 1454 -500 1478
rect 500 2230 597 2254
rect 500 1478 551 2230
rect 585 1478 597 2230
rect 500 1454 597 1478
rect 923 2230 1020 2254
rect 923 1478 935 2230
rect 969 1478 1020 2230
rect 923 1454 1020 1478
rect 2020 2230 2117 2254
rect 2020 1478 2071 2230
rect 2105 1478 2117 2230
rect 2020 1454 2117 1478
rect 2443 2230 2540 2254
rect 2443 1478 2455 2230
rect 2489 1478 2540 2230
rect 2443 1454 2540 1478
rect 3540 2230 3637 2254
rect 3540 1478 3591 2230
rect 3625 1478 3637 2230
rect 3540 1454 3637 1478
rect -3637 994 -3540 1018
rect -3637 242 -3625 994
rect -3591 242 -3540 994
rect -3637 218 -3540 242
rect -2540 994 -2443 1018
rect -2540 242 -2489 994
rect -2455 242 -2443 994
rect -2540 218 -2443 242
rect -2117 994 -2020 1018
rect -2117 242 -2105 994
rect -2071 242 -2020 994
rect -2117 218 -2020 242
rect -1020 994 -923 1018
rect -1020 242 -969 994
rect -935 242 -923 994
rect -1020 218 -923 242
rect -597 994 -500 1018
rect -597 242 -585 994
rect -551 242 -500 994
rect -597 218 -500 242
rect 500 994 597 1018
rect 500 242 551 994
rect 585 242 597 994
rect 500 218 597 242
rect 923 994 1020 1018
rect 923 242 935 994
rect 969 242 1020 994
rect 923 218 1020 242
rect 2020 994 2117 1018
rect 2020 242 2071 994
rect 2105 242 2117 994
rect 2020 218 2117 242
rect 2443 994 2540 1018
rect 2443 242 2455 994
rect 2489 242 2540 994
rect 2443 218 2540 242
rect 3540 994 3637 1018
rect 3540 242 3591 994
rect 3625 242 3637 994
rect 3540 218 3637 242
rect -3637 -242 -3540 -218
rect -3637 -994 -3625 -242
rect -3591 -994 -3540 -242
rect -3637 -1018 -3540 -994
rect -2540 -242 -2443 -218
rect -2540 -994 -2489 -242
rect -2455 -994 -2443 -242
rect -2540 -1018 -2443 -994
rect -2117 -242 -2020 -218
rect -2117 -994 -2105 -242
rect -2071 -994 -2020 -242
rect -2117 -1018 -2020 -994
rect -1020 -242 -923 -218
rect -1020 -994 -969 -242
rect -935 -994 -923 -242
rect -1020 -1018 -923 -994
rect -597 -242 -500 -218
rect -597 -994 -585 -242
rect -551 -994 -500 -242
rect -597 -1018 -500 -994
rect 500 -242 597 -218
rect 500 -994 551 -242
rect 585 -994 597 -242
rect 500 -1018 597 -994
rect 923 -242 1020 -218
rect 923 -994 935 -242
rect 969 -994 1020 -242
rect 923 -1018 1020 -994
rect 2020 -242 2117 -218
rect 2020 -994 2071 -242
rect 2105 -994 2117 -242
rect 2020 -1018 2117 -994
rect 2443 -242 2540 -218
rect 2443 -994 2455 -242
rect 2489 -994 2540 -242
rect 2443 -1018 2540 -994
rect 3540 -242 3637 -218
rect 3540 -994 3591 -242
rect 3625 -994 3637 -242
rect 3540 -1018 3637 -994
rect -3637 -1478 -3540 -1454
rect -3637 -2230 -3625 -1478
rect -3591 -2230 -3540 -1478
rect -3637 -2254 -3540 -2230
rect -2540 -1478 -2443 -1454
rect -2540 -2230 -2489 -1478
rect -2455 -2230 -2443 -1478
rect -2540 -2254 -2443 -2230
rect -2117 -1478 -2020 -1454
rect -2117 -2230 -2105 -1478
rect -2071 -2230 -2020 -1478
rect -2117 -2254 -2020 -2230
rect -1020 -1478 -923 -1454
rect -1020 -2230 -969 -1478
rect -935 -2230 -923 -1478
rect -1020 -2254 -923 -2230
rect -597 -1478 -500 -1454
rect -597 -2230 -585 -1478
rect -551 -2230 -500 -1478
rect -597 -2254 -500 -2230
rect 500 -1478 597 -1454
rect 500 -2230 551 -1478
rect 585 -2230 597 -1478
rect 500 -2254 597 -2230
rect 923 -1478 1020 -1454
rect 923 -2230 935 -1478
rect 969 -2230 1020 -1478
rect 923 -2254 1020 -2230
rect 2020 -1478 2117 -1454
rect 2020 -2230 2071 -1478
rect 2105 -2230 2117 -1478
rect 2020 -2254 2117 -2230
rect 2443 -1478 2540 -1454
rect 2443 -2230 2455 -1478
rect 2489 -2230 2540 -1478
rect 2443 -2254 2540 -2230
rect 3540 -1478 3637 -1454
rect 3540 -2230 3591 -1478
rect 3625 -2230 3637 -1478
rect 3540 -2254 3637 -2230
<< psubdiffcont >>
rect -3651 2385 3651 2419
rect -3747 -2323 -3713 2323
rect 3713 -2323 3747 2323
rect -3651 -2419 3651 -2385
<< nsubdiffcont >>
rect -3625 1478 -3591 2230
rect -2489 1478 -2455 2230
rect -2105 1478 -2071 2230
rect -969 1478 -935 2230
rect -585 1478 -551 2230
rect 551 1478 585 2230
rect 935 1478 969 2230
rect 2071 1478 2105 2230
rect 2455 1478 2489 2230
rect 3591 1478 3625 2230
rect -3625 242 -3591 994
rect -2489 242 -2455 994
rect -2105 242 -2071 994
rect -969 242 -935 994
rect -585 242 -551 994
rect 551 242 585 994
rect 935 242 969 994
rect 2071 242 2105 994
rect 2455 242 2489 994
rect 3591 242 3625 994
rect -3625 -994 -3591 -242
rect -2489 -994 -2455 -242
rect -2105 -994 -2071 -242
rect -969 -994 -935 -242
rect -585 -994 -551 -242
rect 551 -994 585 -242
rect 935 -994 969 -242
rect 2071 -994 2105 -242
rect 2455 -994 2489 -242
rect 3591 -994 3625 -242
rect -3625 -2230 -3591 -1478
rect -2489 -2230 -2455 -1478
rect -2105 -2230 -2071 -1478
rect -969 -2230 -935 -1478
rect -585 -2230 -551 -1478
rect 551 -2230 585 -1478
rect 935 -2230 969 -1478
rect 2071 -2230 2105 -1478
rect 2455 -2230 2489 -1478
rect 3591 -2230 3625 -1478
<< poly >>
rect -3540 2326 -2540 2342
rect -3540 2292 -3524 2326
rect -2556 2292 -2540 2326
rect -3540 2254 -2540 2292
rect -2020 2326 -1020 2342
rect -2020 2292 -2004 2326
rect -1036 2292 -1020 2326
rect -2020 2254 -1020 2292
rect -500 2326 500 2342
rect -500 2292 -484 2326
rect 484 2292 500 2326
rect -500 2254 500 2292
rect 1020 2326 2020 2342
rect 1020 2292 1036 2326
rect 2004 2292 2020 2326
rect 1020 2254 2020 2292
rect 2540 2326 3540 2342
rect 2540 2292 2556 2326
rect 3524 2292 3540 2326
rect 2540 2254 3540 2292
rect -3540 1416 -2540 1454
rect -3540 1382 -3524 1416
rect -2556 1382 -2540 1416
rect -3540 1366 -2540 1382
rect -2020 1416 -1020 1454
rect -2020 1382 -2004 1416
rect -1036 1382 -1020 1416
rect -2020 1366 -1020 1382
rect -500 1416 500 1454
rect -500 1382 -484 1416
rect 484 1382 500 1416
rect -500 1366 500 1382
rect 1020 1416 2020 1454
rect 1020 1382 1036 1416
rect 2004 1382 2020 1416
rect 1020 1366 2020 1382
rect 2540 1416 3540 1454
rect 2540 1382 2556 1416
rect 3524 1382 3540 1416
rect 2540 1366 3540 1382
rect -3540 1090 -2540 1106
rect -3540 1056 -3524 1090
rect -2556 1056 -2540 1090
rect -3540 1018 -2540 1056
rect -2020 1090 -1020 1106
rect -2020 1056 -2004 1090
rect -1036 1056 -1020 1090
rect -2020 1018 -1020 1056
rect -500 1090 500 1106
rect -500 1056 -484 1090
rect 484 1056 500 1090
rect -500 1018 500 1056
rect 1020 1090 2020 1106
rect 1020 1056 1036 1090
rect 2004 1056 2020 1090
rect 1020 1018 2020 1056
rect 2540 1090 3540 1106
rect 2540 1056 2556 1090
rect 3524 1056 3540 1090
rect 2540 1018 3540 1056
rect -3540 180 -2540 218
rect -3540 146 -3524 180
rect -2556 146 -2540 180
rect -3540 130 -2540 146
rect -2020 180 -1020 218
rect -2020 146 -2004 180
rect -1036 146 -1020 180
rect -2020 130 -1020 146
rect -500 180 500 218
rect -500 146 -484 180
rect 484 146 500 180
rect -500 130 500 146
rect 1020 180 2020 218
rect 1020 146 1036 180
rect 2004 146 2020 180
rect 1020 130 2020 146
rect 2540 180 3540 218
rect 2540 146 2556 180
rect 3524 146 3540 180
rect 2540 130 3540 146
rect -3540 -146 -2540 -130
rect -3540 -180 -3524 -146
rect -2556 -180 -2540 -146
rect -3540 -218 -2540 -180
rect -2020 -146 -1020 -130
rect -2020 -180 -2004 -146
rect -1036 -180 -1020 -146
rect -2020 -218 -1020 -180
rect -500 -146 500 -130
rect -500 -180 -484 -146
rect 484 -180 500 -146
rect -500 -218 500 -180
rect 1020 -146 2020 -130
rect 1020 -180 1036 -146
rect 2004 -180 2020 -146
rect 1020 -218 2020 -180
rect 2540 -146 3540 -130
rect 2540 -180 2556 -146
rect 3524 -180 3540 -146
rect 2540 -218 3540 -180
rect -3540 -1056 -2540 -1018
rect -3540 -1090 -3524 -1056
rect -2556 -1090 -2540 -1056
rect -3540 -1106 -2540 -1090
rect -2020 -1056 -1020 -1018
rect -2020 -1090 -2004 -1056
rect -1036 -1090 -1020 -1056
rect -2020 -1106 -1020 -1090
rect -500 -1056 500 -1018
rect -500 -1090 -484 -1056
rect 484 -1090 500 -1056
rect -500 -1106 500 -1090
rect 1020 -1056 2020 -1018
rect 1020 -1090 1036 -1056
rect 2004 -1090 2020 -1056
rect 1020 -1106 2020 -1090
rect 2540 -1056 3540 -1018
rect 2540 -1090 2556 -1056
rect 3524 -1090 3540 -1056
rect 2540 -1106 3540 -1090
rect -3540 -1382 -2540 -1366
rect -3540 -1416 -3524 -1382
rect -2556 -1416 -2540 -1382
rect -3540 -1454 -2540 -1416
rect -2020 -1382 -1020 -1366
rect -2020 -1416 -2004 -1382
rect -1036 -1416 -1020 -1382
rect -2020 -1454 -1020 -1416
rect -500 -1382 500 -1366
rect -500 -1416 -484 -1382
rect 484 -1416 500 -1382
rect -500 -1454 500 -1416
rect 1020 -1382 2020 -1366
rect 1020 -1416 1036 -1382
rect 2004 -1416 2020 -1382
rect 1020 -1454 2020 -1416
rect 2540 -1382 3540 -1366
rect 2540 -1416 2556 -1382
rect 3524 -1416 3540 -1382
rect 2540 -1454 3540 -1416
rect -3540 -2292 -2540 -2254
rect -3540 -2326 -3524 -2292
rect -2556 -2326 -2540 -2292
rect -3540 -2342 -2540 -2326
rect -2020 -2292 -1020 -2254
rect -2020 -2326 -2004 -2292
rect -1036 -2326 -1020 -2292
rect -2020 -2342 -1020 -2326
rect -500 -2292 500 -2254
rect -500 -2326 -484 -2292
rect 484 -2326 500 -2292
rect -500 -2342 500 -2326
rect 1020 -2292 2020 -2254
rect 1020 -2326 1036 -2292
rect 2004 -2326 2020 -2292
rect 1020 -2342 2020 -2326
rect 2540 -2292 3540 -2254
rect 2540 -2326 2556 -2292
rect 3524 -2326 3540 -2292
rect 2540 -2342 3540 -2326
<< polycont >>
rect -3524 2292 -2556 2326
rect -2004 2292 -1036 2326
rect -484 2292 484 2326
rect 1036 2292 2004 2326
rect 2556 2292 3524 2326
rect -3524 1382 -2556 1416
rect -2004 1382 -1036 1416
rect -484 1382 484 1416
rect 1036 1382 2004 1416
rect 2556 1382 3524 1416
rect -3524 1056 -2556 1090
rect -2004 1056 -1036 1090
rect -484 1056 484 1090
rect 1036 1056 2004 1090
rect 2556 1056 3524 1090
rect -3524 146 -2556 180
rect -2004 146 -1036 180
rect -484 146 484 180
rect 1036 146 2004 180
rect 2556 146 3524 180
rect -3524 -180 -2556 -146
rect -2004 -180 -1036 -146
rect -484 -180 484 -146
rect 1036 -180 2004 -146
rect 2556 -180 3524 -146
rect -3524 -1090 -2556 -1056
rect -2004 -1090 -1036 -1056
rect -484 -1090 484 -1056
rect 1036 -1090 2004 -1056
rect 2556 -1090 3524 -1056
rect -3524 -1416 -2556 -1382
rect -2004 -1416 -1036 -1382
rect -484 -1416 484 -1382
rect 1036 -1416 2004 -1382
rect 2556 -1416 3524 -1382
rect -3524 -2326 -2556 -2292
rect -2004 -2326 -1036 -2292
rect -484 -2326 484 -2292
rect 1036 -2326 2004 -2292
rect 2556 -2326 3524 -2292
<< locali >>
rect -3747 2385 -3651 2419
rect 3651 2385 3747 2419
rect -3747 2323 -3713 2385
rect -3540 2292 -3524 2326
rect -2556 2292 -2540 2326
rect -2020 2292 -2004 2326
rect -1036 2292 -1020 2326
rect -500 2292 -484 2326
rect 484 2292 500 2326
rect 1020 2292 1036 2326
rect 2004 2292 2020 2326
rect 2540 2292 2556 2326
rect 3524 2292 3540 2326
rect 3713 2323 3747 2385
rect -3625 2230 -3591 2246
rect -3625 1462 -3591 1478
rect -2489 2230 -2455 2246
rect -2489 1462 -2455 1478
rect -2105 2230 -2071 2246
rect -2105 1462 -2071 1478
rect -969 2230 -935 2246
rect -969 1462 -935 1478
rect -585 2230 -551 2246
rect -585 1462 -551 1478
rect 551 2230 585 2246
rect 551 1462 585 1478
rect 935 2230 969 2246
rect 935 1462 969 1478
rect 2071 2230 2105 2246
rect 2071 1462 2105 1478
rect 2455 2230 2489 2246
rect 2455 1462 2489 1478
rect 3591 2230 3625 2246
rect 3591 1462 3625 1478
rect -3540 1382 -3524 1416
rect -2556 1382 -2540 1416
rect -2020 1382 -2004 1416
rect -1036 1382 -1020 1416
rect -500 1382 -484 1416
rect 484 1382 500 1416
rect 1020 1382 1036 1416
rect 2004 1382 2020 1416
rect 2540 1382 2556 1416
rect 3524 1382 3540 1416
rect -3540 1056 -3524 1090
rect -2556 1056 -2540 1090
rect -2020 1056 -2004 1090
rect -1036 1056 -1020 1090
rect -500 1056 -484 1090
rect 484 1056 500 1090
rect 1020 1056 1036 1090
rect 2004 1056 2020 1090
rect 2540 1056 2556 1090
rect 3524 1056 3540 1090
rect -3625 994 -3591 1010
rect -3625 226 -3591 242
rect -2489 994 -2455 1010
rect -2489 226 -2455 242
rect -2105 994 -2071 1010
rect -2105 226 -2071 242
rect -969 994 -935 1010
rect -969 226 -935 242
rect -585 994 -551 1010
rect -585 226 -551 242
rect 551 994 585 1010
rect 551 226 585 242
rect 935 994 969 1010
rect 935 226 969 242
rect 2071 994 2105 1010
rect 2071 226 2105 242
rect 2455 994 2489 1010
rect 2455 226 2489 242
rect 3591 994 3625 1010
rect 3591 226 3625 242
rect -3540 146 -3524 180
rect -2556 146 -2540 180
rect -2020 146 -2004 180
rect -1036 146 -1020 180
rect -500 146 -484 180
rect 484 146 500 180
rect 1020 146 1036 180
rect 2004 146 2020 180
rect 2540 146 2556 180
rect 3524 146 3540 180
rect -3540 -180 -3524 -146
rect -2556 -180 -2540 -146
rect -2020 -180 -2004 -146
rect -1036 -180 -1020 -146
rect -500 -180 -484 -146
rect 484 -180 500 -146
rect 1020 -180 1036 -146
rect 2004 -180 2020 -146
rect 2540 -180 2556 -146
rect 3524 -180 3540 -146
rect -3625 -242 -3591 -226
rect -3625 -1010 -3591 -994
rect -2489 -242 -2455 -226
rect -2489 -1010 -2455 -994
rect -2105 -242 -2071 -226
rect -2105 -1010 -2071 -994
rect -969 -242 -935 -226
rect -969 -1010 -935 -994
rect -585 -242 -551 -226
rect -585 -1010 -551 -994
rect 551 -242 585 -226
rect 551 -1010 585 -994
rect 935 -242 969 -226
rect 935 -1010 969 -994
rect 2071 -242 2105 -226
rect 2071 -1010 2105 -994
rect 2455 -242 2489 -226
rect 2455 -1010 2489 -994
rect 3591 -242 3625 -226
rect 3591 -1010 3625 -994
rect -3540 -1090 -3524 -1056
rect -2556 -1090 -2540 -1056
rect -2020 -1090 -2004 -1056
rect -1036 -1090 -1020 -1056
rect -500 -1090 -484 -1056
rect 484 -1090 500 -1056
rect 1020 -1090 1036 -1056
rect 2004 -1090 2020 -1056
rect 2540 -1090 2556 -1056
rect 3524 -1090 3540 -1056
rect -3540 -1416 -3524 -1382
rect -2556 -1416 -2540 -1382
rect -2020 -1416 -2004 -1382
rect -1036 -1416 -1020 -1382
rect -500 -1416 -484 -1382
rect 484 -1416 500 -1382
rect 1020 -1416 1036 -1382
rect 2004 -1416 2020 -1382
rect 2540 -1416 2556 -1382
rect 3524 -1416 3540 -1382
rect -3625 -1478 -3591 -1462
rect -3625 -2246 -3591 -2230
rect -2489 -1478 -2455 -1462
rect -2489 -2246 -2455 -2230
rect -2105 -1478 -2071 -1462
rect -2105 -2246 -2071 -2230
rect -969 -1478 -935 -1462
rect -969 -2246 -935 -2230
rect -585 -1478 -551 -1462
rect -585 -2246 -551 -2230
rect 551 -1478 585 -1462
rect 551 -2246 585 -2230
rect 935 -1478 969 -1462
rect 935 -2246 969 -2230
rect 2071 -1478 2105 -1462
rect 2071 -2246 2105 -2230
rect 2455 -1478 2489 -1462
rect 2455 -2246 2489 -2230
rect 3591 -1478 3625 -1462
rect 3591 -2246 3625 -2230
rect -3747 -2385 -3713 -2323
rect -3540 -2326 -3524 -2292
rect -2556 -2326 -2540 -2292
rect -2020 -2326 -2004 -2292
rect -1036 -2326 -1020 -2292
rect -500 -2326 -484 -2292
rect 484 -2326 500 -2292
rect 1020 -2326 1036 -2292
rect 2004 -2326 2020 -2292
rect 2540 -2326 2556 -2292
rect 3524 -2326 3540 -2292
rect 3713 -2385 3747 -2323
rect -3747 -2419 -3651 -2385
rect 3651 -2419 3747 -2385
<< viali >>
rect -3524 2292 -2556 2326
rect -2004 2292 -1036 2326
rect -484 2292 484 2326
rect 1036 2292 2004 2326
rect 2556 2292 3524 2326
rect -3625 1478 -3591 2230
rect -2489 1478 -2455 2230
rect -2105 1478 -2071 2230
rect -969 1478 -935 2230
rect -585 1478 -551 2230
rect 551 1478 585 2230
rect 935 1478 969 2230
rect 2071 1478 2105 2230
rect 2455 1478 2489 2230
rect 3591 1478 3625 2230
rect -3524 1382 -2556 1416
rect -2004 1382 -1036 1416
rect -484 1382 484 1416
rect 1036 1382 2004 1416
rect 2556 1382 3524 1416
rect -3524 1056 -2556 1090
rect -2004 1056 -1036 1090
rect -484 1056 484 1090
rect 1036 1056 2004 1090
rect 2556 1056 3524 1090
rect -3625 242 -3591 994
rect -2489 242 -2455 994
rect -2105 242 -2071 994
rect -969 242 -935 994
rect -585 242 -551 994
rect 551 242 585 994
rect 935 242 969 994
rect 2071 242 2105 994
rect 2455 242 2489 994
rect 3591 242 3625 994
rect -3524 146 -2556 180
rect -2004 146 -1036 180
rect -484 146 484 180
rect 1036 146 2004 180
rect 2556 146 3524 180
rect -3524 -180 -2556 -146
rect -2004 -180 -1036 -146
rect -484 -180 484 -146
rect 1036 -180 2004 -146
rect 2556 -180 3524 -146
rect -3625 -994 -3591 -242
rect -2489 -994 -2455 -242
rect -2105 -994 -2071 -242
rect -969 -994 -935 -242
rect -585 -994 -551 -242
rect 551 -994 585 -242
rect 935 -994 969 -242
rect 2071 -994 2105 -242
rect 2455 -994 2489 -242
rect 3591 -994 3625 -242
rect -3524 -1090 -2556 -1056
rect -2004 -1090 -1036 -1056
rect -484 -1090 484 -1056
rect 1036 -1090 2004 -1056
rect 2556 -1090 3524 -1056
rect -3524 -1416 -2556 -1382
rect -2004 -1416 -1036 -1382
rect -484 -1416 484 -1382
rect 1036 -1416 2004 -1382
rect 2556 -1416 3524 -1382
rect -3625 -2230 -3591 -1478
rect -2489 -2230 -2455 -1478
rect -2105 -2230 -2071 -1478
rect -969 -2230 -935 -1478
rect -585 -2230 -551 -1478
rect 551 -2230 585 -1478
rect 935 -2230 969 -1478
rect 2071 -2230 2105 -1478
rect 2455 -2230 2489 -1478
rect 3591 -2230 3625 -1478
rect -3524 -2326 -2556 -2292
rect -2004 -2326 -1036 -2292
rect -484 -2326 484 -2292
rect 1036 -2326 2004 -2292
rect 2556 -2326 3524 -2292
<< metal1 >>
rect -3536 2326 -2544 2332
rect -3536 2292 -3524 2326
rect -2556 2292 -2544 2326
rect -3536 2286 -2544 2292
rect -2016 2326 -1024 2332
rect -2016 2292 -2004 2326
rect -1036 2292 -1024 2326
rect -2016 2286 -1024 2292
rect -496 2326 496 2332
rect -496 2292 -484 2326
rect 484 2292 496 2326
rect -496 2286 496 2292
rect 1024 2326 2016 2332
rect 1024 2292 1036 2326
rect 2004 2292 2016 2326
rect 1024 2286 2016 2292
rect 2544 2326 3536 2332
rect 2544 2292 2556 2326
rect 3524 2292 3536 2326
rect 2544 2286 3536 2292
rect -3631 2230 -3585 2242
rect -2495 2230 -2449 2242
rect -3631 1478 -3625 2230
rect -3591 1478 -2489 2230
rect -2455 1478 -2449 2230
rect -3631 1466 -3585 1478
rect -2495 1466 -2449 1478
rect -2111 2230 -2065 2242
rect -975 2230 -929 2242
rect -2111 1478 -2105 2230
rect -2071 1478 -969 2230
rect -935 1478 -929 2230
rect -2111 1466 -2065 1478
rect -975 1466 -929 1478
rect -591 2230 -545 2242
rect 545 2230 591 2242
rect -591 1478 -585 2230
rect -551 1478 551 2230
rect 585 1478 591 2230
rect -591 1466 -545 1478
rect 545 1466 591 1478
rect 929 2230 975 2242
rect 2065 2230 2111 2242
rect 929 1478 935 2230
rect 969 1478 2071 2230
rect 2105 1478 2111 2230
rect 929 1466 975 1478
rect 2065 1466 2111 1478
rect 2449 2230 2495 2242
rect 3585 2230 3631 2242
rect 2449 1478 2455 2230
rect 2489 1478 3591 2230
rect 3625 1478 3631 2230
rect 2449 1466 2495 1478
rect 3585 1466 3631 1478
rect -3536 1416 -2544 1422
rect -3536 1382 -3524 1416
rect -2556 1382 -2544 1416
rect -3536 1376 -2544 1382
rect -2016 1416 -1024 1422
rect -2016 1382 -2004 1416
rect -1036 1382 -1024 1416
rect -2016 1376 -1024 1382
rect -496 1416 496 1422
rect -496 1382 -484 1416
rect 484 1382 496 1416
rect -496 1376 496 1382
rect 1024 1416 2016 1422
rect 1024 1382 1036 1416
rect 2004 1382 2016 1416
rect 1024 1376 2016 1382
rect 2544 1416 3536 1422
rect 2544 1382 2556 1416
rect 3524 1382 3536 1416
rect 2544 1376 3536 1382
rect -3536 1090 -2544 1096
rect -3536 1056 -3524 1090
rect -2556 1056 -2544 1090
rect -3536 1050 -2544 1056
rect -2016 1090 -1024 1096
rect -2016 1056 -2004 1090
rect -1036 1056 -1024 1090
rect -2016 1050 -1024 1056
rect -496 1090 496 1096
rect -496 1056 -484 1090
rect 484 1056 496 1090
rect -496 1050 496 1056
rect 1024 1090 2016 1096
rect 1024 1056 1036 1090
rect 2004 1056 2016 1090
rect 1024 1050 2016 1056
rect 2544 1090 3536 1096
rect 2544 1056 2556 1090
rect 3524 1056 3536 1090
rect 2544 1050 3536 1056
rect -3631 994 -3585 1006
rect -2495 994 -2449 1006
rect -3631 242 -3625 994
rect -3591 242 -2489 994
rect -2455 242 -2449 994
rect -3631 230 -3585 242
rect -2495 230 -2449 242
rect -2111 994 -2065 1006
rect -975 994 -929 1006
rect -2111 242 -2105 994
rect -2071 242 -969 994
rect -935 242 -929 994
rect -2111 230 -2065 242
rect -975 230 -929 242
rect -591 994 -545 1006
rect 545 994 591 1006
rect -591 242 -585 994
rect -551 242 551 994
rect 585 242 591 994
rect -591 230 -545 242
rect 545 230 591 242
rect 929 994 975 1006
rect 2065 994 2111 1006
rect 929 242 935 994
rect 969 242 2071 994
rect 2105 242 2111 994
rect 929 230 975 242
rect 2065 230 2111 242
rect 2449 994 2495 1006
rect 3585 994 3631 1006
rect 2449 242 2455 994
rect 2489 242 3591 994
rect 3625 242 3631 994
rect 2449 230 2495 242
rect 3585 230 3631 242
rect -3536 180 -2544 186
rect -3536 146 -3524 180
rect -2556 146 -2544 180
rect -3536 140 -2544 146
rect -2016 180 -1024 186
rect -2016 146 -2004 180
rect -1036 146 -1024 180
rect -2016 140 -1024 146
rect -496 180 496 186
rect -496 146 -484 180
rect 484 146 496 180
rect -496 140 496 146
rect 1024 180 2016 186
rect 1024 146 1036 180
rect 2004 146 2016 180
rect 1024 140 2016 146
rect 2544 180 3536 186
rect 2544 146 2556 180
rect 3524 146 3536 180
rect 2544 140 3536 146
rect -3536 -146 -2544 -140
rect -3536 -180 -3524 -146
rect -2556 -180 -2544 -146
rect -3536 -186 -2544 -180
rect -2016 -146 -1024 -140
rect -2016 -180 -2004 -146
rect -1036 -180 -1024 -146
rect -2016 -186 -1024 -180
rect -496 -146 496 -140
rect -496 -180 -484 -146
rect 484 -180 496 -146
rect -496 -186 496 -180
rect 1024 -146 2016 -140
rect 1024 -180 1036 -146
rect 2004 -180 2016 -146
rect 1024 -186 2016 -180
rect 2544 -146 3536 -140
rect 2544 -180 2556 -146
rect 3524 -180 3536 -146
rect 2544 -186 3536 -180
rect -3631 -242 -3585 -230
rect -2495 -242 -2449 -230
rect -3631 -994 -3625 -242
rect -3591 -994 -2489 -242
rect -2455 -994 -2449 -242
rect -3631 -1006 -3585 -994
rect -2495 -1006 -2449 -994
rect -2111 -242 -2065 -230
rect -975 -242 -929 -230
rect -2111 -994 -2105 -242
rect -2071 -994 -969 -242
rect -935 -994 -929 -242
rect -2111 -1006 -2065 -994
rect -975 -1006 -929 -994
rect -591 -242 -545 -230
rect 545 -242 591 -230
rect -591 -994 -585 -242
rect -551 -994 551 -242
rect 585 -994 591 -242
rect -591 -1006 -545 -994
rect 545 -1006 591 -994
rect 929 -242 975 -230
rect 2065 -242 2111 -230
rect 929 -994 935 -242
rect 969 -994 2071 -242
rect 2105 -994 2111 -242
rect 929 -1006 975 -994
rect 2065 -1006 2111 -994
rect 2449 -242 2495 -230
rect 3585 -242 3631 -230
rect 2449 -994 2455 -242
rect 2489 -994 3591 -242
rect 3625 -994 3631 -242
rect 2449 -1006 2495 -994
rect 3585 -1006 3631 -994
rect -3536 -1056 -2544 -1050
rect -3536 -1090 -3524 -1056
rect -2556 -1090 -2544 -1056
rect -3536 -1096 -2544 -1090
rect -2016 -1056 -1024 -1050
rect -2016 -1090 -2004 -1056
rect -1036 -1090 -1024 -1056
rect -2016 -1096 -1024 -1090
rect -496 -1056 496 -1050
rect -496 -1090 -484 -1056
rect 484 -1090 496 -1056
rect -496 -1096 496 -1090
rect 1024 -1056 2016 -1050
rect 1024 -1090 1036 -1056
rect 2004 -1090 2016 -1056
rect 1024 -1096 2016 -1090
rect 2544 -1056 3536 -1050
rect 2544 -1090 2556 -1056
rect 3524 -1090 3536 -1056
rect 2544 -1096 3536 -1090
rect -3536 -1382 -2544 -1376
rect -3536 -1416 -3524 -1382
rect -2556 -1416 -2544 -1382
rect -3536 -1422 -2544 -1416
rect -2016 -1382 -1024 -1376
rect -2016 -1416 -2004 -1382
rect -1036 -1416 -1024 -1382
rect -2016 -1422 -1024 -1416
rect -496 -1382 496 -1376
rect -496 -1416 -484 -1382
rect 484 -1416 496 -1382
rect -496 -1422 496 -1416
rect 1024 -1382 2016 -1376
rect 1024 -1416 1036 -1382
rect 2004 -1416 2016 -1382
rect 1024 -1422 2016 -1416
rect 2544 -1382 3536 -1376
rect 2544 -1416 2556 -1382
rect 3524 -1416 3536 -1382
rect 2544 -1422 3536 -1416
rect -3631 -1478 -3585 -1466
rect -2495 -1478 -2449 -1466
rect -3631 -2230 -3625 -1478
rect -3591 -2230 -2489 -1478
rect -2455 -2230 -2449 -1478
rect -3631 -2242 -3585 -2230
rect -2495 -2242 -2449 -2230
rect -2111 -1478 -2065 -1466
rect -975 -1478 -929 -1466
rect -2111 -2230 -2105 -1478
rect -2071 -2230 -969 -1478
rect -935 -2230 -929 -1478
rect -2111 -2242 -2065 -2230
rect -975 -2242 -929 -2230
rect -591 -1478 -545 -1466
rect 545 -1478 591 -1466
rect -591 -2230 -585 -1478
rect -551 -2230 551 -1478
rect 585 -2230 591 -1478
rect -591 -2242 -545 -2230
rect 545 -2242 591 -2230
rect 929 -1478 975 -1466
rect 2065 -1478 2111 -1466
rect 929 -2230 935 -1478
rect 969 -2230 2071 -1478
rect 2105 -2230 2111 -1478
rect 929 -2242 975 -2230
rect 2065 -2242 2111 -2230
rect 2449 -1478 2495 -1466
rect 3585 -1478 3631 -1466
rect 2449 -2230 2455 -1478
rect 2489 -2230 3591 -1478
rect 3625 -2230 3631 -1478
rect 2449 -2242 2495 -2230
rect 3585 -2242 3631 -2230
rect -3536 -2292 -2544 -2286
rect -3536 -2326 -3524 -2292
rect -2556 -2326 -2544 -2292
rect -3536 -2332 -2544 -2326
rect -2016 -2292 -1024 -2286
rect -2016 -2326 -2004 -2292
rect -1036 -2326 -1024 -2292
rect -2016 -2332 -1024 -2326
rect -496 -2292 496 -2286
rect -496 -2326 -484 -2292
rect 484 -2326 496 -2292
rect -496 -2332 496 -2326
rect 1024 -2292 2016 -2286
rect 1024 -2326 1036 -2292
rect 2004 -2326 2016 -2292
rect 1024 -2332 2016 -2326
rect 2544 -2292 3536 -2286
rect 2544 -2326 2556 -2292
rect 3524 -2326 3536 -2292
rect 2544 -2332 3536 -2326
<< properties >>
string FIXED_BBOX -3730 -2402 3730 2402
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 4 l 5 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
