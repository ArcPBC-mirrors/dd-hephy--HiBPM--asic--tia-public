magic
tech sky130A
magscale 1 2
timestamp 1685113734
<< locali >>
rect 260 6680 3320 6780
rect 40 4420 860 4520
rect 1100 4420 1900 4520
rect 2140 4420 2880 4540
rect 3180 4420 4100 4540
rect 1000 2280 1080 3020
rect 100 2180 820 2280
rect 1140 2200 1860 2300
rect 2040 2280 2120 3020
rect 2140 2200 2860 2300
rect 40 0 3080 60
rect 40 -40 840 0
rect 1140 -40 3080 0
<< viali >>
rect 840 -120 1140 0
<< metal1 >>
rect -84 5944 3940 6060
rect -84 3820 72 5944
rect -84 3704 2920 3820
rect -84 1580 72 3704
rect -84 1464 2940 1580
rect 828 0 1152 6
rect 828 -120 840 0
rect 1140 -120 1152 0
rect 828 -126 1152 -120
<< via1 >>
rect 840 -120 1140 0
<< metal2 >>
rect 780 9260 1180 9270
rect 780 9030 1180 9040
rect 1800 9260 2200 9270
rect 1800 9030 2200 9040
rect 2840 9260 3240 9270
rect 2840 9030 3240 9040
rect 220 8940 660 8950
rect 220 8690 660 8700
rect 1300 8920 1700 8930
rect 1300 8690 1700 8700
rect 2340 8920 2740 8930
rect 2340 8690 2740 8700
rect 780 8640 1180 8650
rect 780 8410 1180 8420
rect 1800 8640 2200 8650
rect 1800 8410 2200 8420
rect 2840 8640 3240 8650
rect 2840 8410 3240 8420
rect 220 8320 660 8330
rect 220 8090 660 8100
rect 1300 8320 1700 8330
rect 1300 8090 1700 8100
rect 2340 8320 2740 8330
rect 2340 8090 2740 8100
rect 780 8020 1180 8030
rect 780 7790 1180 7800
rect 1800 8020 2200 8030
rect 1800 7790 2200 7800
rect 2840 8020 3240 8030
rect 2840 7790 3240 7800
rect 220 7700 660 7710
rect 220 7470 660 7480
rect 1300 7700 1700 7710
rect 1300 7470 1700 7480
rect 2340 7700 2740 7710
rect 2340 7470 2740 7480
rect 780 7400 1180 7410
rect 780 7170 1180 7180
rect 1800 7400 2200 7410
rect 1800 7170 2200 7180
rect 2840 7400 3240 7410
rect 2840 7170 3240 7180
rect 220 7080 660 7090
rect 220 6850 660 6860
rect 1300 7080 1700 7090
rect 1300 6850 1700 6860
rect 2340 7080 2740 7090
rect 2340 6850 2740 6860
rect 244 6270 664 6280
rect 244 5726 664 5736
rect 1284 6270 1704 6280
rect 1284 5726 1704 5736
rect 2324 6270 2744 6280
rect 2324 5726 2744 5736
rect 3364 6270 3784 6280
rect 3364 5726 3784 5736
rect -84 3288 72 5528
rect 220 5384 3940 5528
rect 780 4840 1200 4850
rect 140 4500 780 4740
rect 1180 4740 1200 4840
rect 1820 4840 2240 4850
rect 1180 4520 1820 4740
rect 2840 4840 3260 4850
rect 2240 4520 2840 4740
rect 3820 4800 4220 4810
rect 3260 4560 3820 4740
rect 3260 4520 4220 4560
rect 1180 4500 4220 4520
rect 140 4440 4220 4500
rect 248 4030 668 4040
rect 248 3486 668 3496
rect 1292 4030 1712 4040
rect 1292 3486 1712 3496
rect 2328 4030 2748 4040
rect 2328 3486 2748 3496
rect -84 3144 2920 3288
rect -84 1048 72 3144
rect 760 2600 1180 2610
rect 760 2270 1180 2280
rect 1820 2600 2240 2610
rect 1820 2270 2240 2280
rect 2840 2600 3260 2610
rect 2840 2270 3260 2280
rect 248 1784 648 1794
rect 248 1250 648 1260
rect 1288 1784 1688 1794
rect 1288 1250 1688 1260
rect 2328 1784 2728 1794
rect 2328 1250 2728 1260
rect -84 904 2940 1048
rect 760 360 1200 370
rect 120 340 760 350
rect 1800 350 2240 370
rect 1200 340 3260 350
rect 120 70 1820 80
rect 2220 70 2840 80
rect 1820 10 2220 20
rect 2840 10 3260 20
rect 840 0 1140 10
rect 840 -130 1140 -120
<< via2 >>
rect 780 9040 1180 9260
rect 1800 9040 2200 9260
rect 2840 9040 3240 9260
rect 220 8700 660 8940
rect 1300 8700 1700 8920
rect 2340 8700 2740 8920
rect 780 8420 1180 8640
rect 1800 8420 2200 8640
rect 2840 8420 3240 8640
rect 220 8100 660 8320
rect 1300 8100 1700 8320
rect 2340 8100 2740 8320
rect 780 7800 1180 8020
rect 1800 7800 2200 8020
rect 2840 7800 3240 8020
rect 220 7480 660 7700
rect 1300 7480 1700 7700
rect 2340 7480 2740 7700
rect 780 7180 1180 7400
rect 1800 7180 2200 7400
rect 2840 7180 3240 7400
rect 220 6860 660 7080
rect 1300 6860 1700 7080
rect 2340 6860 2740 7080
rect 244 5736 664 6270
rect 1284 5736 1704 6270
rect 2324 5736 2744 6270
rect 3364 5736 3784 6270
rect 780 4500 1180 4840
rect 1820 4520 2240 4840
rect 2840 4520 3260 4840
rect 3820 4560 4220 4800
rect 248 3496 668 4030
rect 1292 3496 1712 4030
rect 2328 3496 2748 4030
rect 760 2280 1180 2600
rect 1820 2280 2240 2600
rect 2840 2280 3260 2600
rect 248 1260 648 1784
rect 1288 1260 1688 1784
rect 2328 1260 2728 1784
rect 760 340 1200 360
rect 120 80 3260 340
rect 1820 20 2220 80
rect 2840 20 3260 80
rect 840 -120 1140 0
<< metal3 >>
rect 200 9400 3380 10600
rect 760 9260 1200 9400
rect 760 9040 780 9260
rect 1180 9040 1200 9260
rect 240 8945 680 8960
rect 210 8940 680 8945
rect 210 8700 220 8940
rect 660 8700 680 8940
rect 210 8695 680 8700
rect 240 8325 680 8695
rect 210 8320 680 8325
rect 210 8100 220 8320
rect 660 8100 680 8320
rect 210 8095 680 8100
rect 240 7705 680 8095
rect 210 7700 680 7705
rect 210 7480 220 7700
rect 660 7480 680 7700
rect 210 7475 680 7480
rect 240 7085 680 7475
rect 760 8640 1200 9040
rect 1780 9260 2220 9400
rect 1780 9040 1800 9260
rect 2200 9040 2220 9260
rect 760 8420 780 8640
rect 1180 8420 1200 8640
rect 760 8020 1200 8420
rect 760 7800 780 8020
rect 1180 7800 1200 8020
rect 760 7400 1200 7800
rect 760 7180 780 7400
rect 1180 7180 1200 7400
rect 760 7160 1200 7180
rect 1280 8920 1720 8960
rect 1280 8700 1300 8920
rect 1700 8700 1720 8920
rect 1280 8320 1720 8700
rect 1280 8100 1300 8320
rect 1700 8100 1720 8320
rect 1280 7700 1720 8100
rect 1280 7480 1300 7700
rect 1700 7480 1720 7700
rect 210 7080 680 7085
rect 210 6860 220 7080
rect 660 7040 680 7080
rect 1280 7080 1720 7480
rect 1780 8640 2220 9040
rect 2820 9260 3260 9400
rect 2820 9040 2840 9260
rect 3240 9040 3260 9260
rect 1780 8420 1800 8640
rect 2200 8420 2220 8640
rect 1780 8020 2220 8420
rect 1780 7800 1800 8020
rect 2200 7800 2220 8020
rect 1780 7400 2220 7800
rect 1780 7180 1800 7400
rect 2200 7180 2220 7400
rect 1780 7160 2220 7180
rect 2320 8920 2760 8960
rect 2320 8700 2340 8920
rect 2740 8700 2760 8920
rect 2320 8320 2760 8700
rect 2320 8100 2340 8320
rect 2740 8100 2760 8320
rect 2320 7700 2760 8100
rect 2320 7480 2340 7700
rect 2740 7480 2760 7700
rect 1280 7056 1300 7080
rect 1276 7040 1300 7056
rect 660 6860 1300 7040
rect 1700 7040 1720 7080
rect 2320 7080 2760 7480
rect 2820 8640 3260 9040
rect 2820 8420 2840 8640
rect 3240 8420 3260 8640
rect 2820 8020 3260 8420
rect 2820 7800 2840 8020
rect 3240 7800 3260 8020
rect 2820 7400 3260 7800
rect 2820 7180 2840 7400
rect 3240 7180 3260 7400
rect 2820 7160 3260 7180
rect 2320 7056 2340 7080
rect 2312 7040 2340 7056
rect 1700 6860 2340 7040
rect 2740 7040 2760 7080
rect 2740 6860 3800 7040
rect 210 6855 3800 6860
rect 232 6680 3800 6855
rect 232 6440 3804 6680
rect 232 6270 676 6440
rect 1276 6275 1720 6440
rect 232 5736 244 6270
rect 664 5736 676 6270
rect 232 4035 676 5736
rect 1274 6270 1720 6275
rect 1274 5736 1284 6270
rect 1704 5736 1720 6270
rect 1274 5731 1720 5736
rect 760 4840 1200 4860
rect 760 4500 780 4840
rect 1180 4500 1200 4840
rect 232 4030 678 4035
rect 232 3496 248 4030
rect 668 3496 678 4030
rect 760 3600 1200 4500
rect 232 3491 678 3496
rect 232 1784 676 3491
rect 232 1260 248 1784
rect 648 1260 676 1784
rect 232 1240 676 1260
rect 740 2600 1200 3600
rect 740 2280 760 2600
rect 1180 2280 1200 2600
rect 740 1020 1200 2280
rect 1276 4035 1720 5731
rect 2312 6270 2756 6440
rect 3360 6275 3804 6440
rect 2312 5736 2324 6270
rect 2744 5736 2756 6270
rect 1800 4845 2240 4860
rect 1800 4840 2250 4845
rect 1800 4520 1820 4840
rect 2240 4520 2250 4840
rect 1800 4515 2250 4520
rect 1276 4030 1722 4035
rect 1276 3496 1292 4030
rect 1712 3496 1722 4030
rect 1276 3491 1722 3496
rect 1276 1784 1720 3491
rect 1800 3060 2240 4515
rect 1780 2780 2240 3060
rect 1276 1260 1288 1784
rect 1688 1260 1720 1784
rect 1276 1240 1720 1260
rect 1800 2605 2240 2780
rect 2312 4035 2756 5736
rect 3354 6270 3804 6275
rect 3354 5736 3364 6270
rect 3784 5736 3804 6270
rect 3354 5731 3804 5736
rect 3360 5700 3804 5731
rect 2820 4840 3280 4860
rect 2820 4520 2840 4840
rect 3260 4520 3280 4840
rect 3880 4805 4260 4840
rect 3810 4800 4260 4805
rect 3810 4560 3820 4800
rect 4220 4560 4260 4800
rect 3810 4555 4260 4560
rect 2312 4030 2758 4035
rect 2312 3496 2328 4030
rect 2748 3496 2758 4030
rect 2312 3491 2758 3496
rect 1800 2600 2250 2605
rect 1800 2280 1820 2600
rect 2240 2280 2250 2600
rect 1800 2275 2250 2280
rect 1800 1020 2240 2275
rect 2312 1784 2756 3491
rect 2312 1260 2328 1784
rect 2728 1260 2756 1784
rect 2312 1240 2756 1260
rect 2820 2600 3280 4520
rect 2820 2280 2840 2600
rect 3260 2280 3280 2600
rect 2820 1020 3280 2280
rect 3880 1020 4260 4555
rect 120 360 4260 1020
rect 120 345 760 360
rect 110 340 760 345
rect 1200 340 4260 360
rect 110 80 120 340
rect 110 75 1820 80
rect 120 20 1820 75
rect 2220 20 2840 80
rect 3260 20 4260 340
rect 120 0 4260 20
rect 120 -120 840 0
rect 1140 -120 4260 0
rect 120 -200 4260 -120
use outd_follower  outd_follower_0
timestamp 1685113734
transform 1 0 100 0 1 6740
box -100 -6740 4062 2654
<< end >>
