magic
tech sky130A
magscale 1 2
timestamp 1683553776
<< error_p >>
rect -221 1235 -163 1241
rect -29 1235 29 1241
rect 163 1235 221 1241
rect -221 1201 -209 1235
rect -29 1201 -17 1235
rect 163 1201 175 1235
rect -221 1195 -163 1201
rect -29 1195 29 1201
rect 163 1195 221 1201
rect -125 707 -67 713
rect 67 707 125 713
rect -125 673 -113 707
rect 67 673 79 707
rect -125 667 -67 673
rect 67 667 125 673
rect -125 599 -67 605
rect 67 599 125 605
rect -125 565 -113 599
rect 67 565 79 599
rect -125 559 -67 565
rect 67 559 125 565
rect -221 71 -163 77
rect -29 71 29 77
rect 163 71 221 77
rect -221 37 -209 71
rect -29 37 -17 71
rect 163 37 175 71
rect -221 31 -163 37
rect -29 31 29 37
rect 163 31 221 37
rect -221 -37 -163 -31
rect -29 -37 29 -31
rect 163 -37 221 -31
rect -221 -71 -209 -37
rect -29 -71 -17 -37
rect 163 -71 175 -37
rect -221 -77 -163 -71
rect -29 -77 29 -71
rect 163 -77 221 -71
rect -125 -565 -67 -559
rect 67 -565 125 -559
rect -125 -599 -113 -565
rect 67 -599 79 -565
rect -125 -605 -67 -599
rect 67 -605 125 -599
rect -125 -673 -67 -667
rect 67 -673 125 -667
rect -125 -707 -113 -673
rect 67 -707 79 -673
rect -125 -713 -67 -707
rect 67 -713 125 -707
rect -221 -1201 -163 -1195
rect -29 -1201 29 -1195
rect 163 -1201 221 -1195
rect -221 -1235 -209 -1201
rect -29 -1235 -17 -1201
rect 163 -1235 175 -1201
rect -221 -1241 -163 -1235
rect -29 -1241 29 -1235
rect 163 -1241 221 -1235
<< nwell >>
rect -407 -1373 407 1373
<< pmos >>
rect -207 754 -177 1154
rect -111 754 -81 1154
rect -15 754 15 1154
rect 81 754 111 1154
rect 177 754 207 1154
rect -207 118 -177 518
rect -111 118 -81 518
rect -15 118 15 518
rect 81 118 111 518
rect 177 118 207 518
rect -207 -518 -177 -118
rect -111 -518 -81 -118
rect -15 -518 15 -118
rect 81 -518 111 -118
rect 177 -518 207 -118
rect -207 -1154 -177 -754
rect -111 -1154 -81 -754
rect -15 -1154 15 -754
rect 81 -1154 111 -754
rect 177 -1154 207 -754
<< pdiff >>
rect -269 1142 -207 1154
rect -269 766 -257 1142
rect -223 766 -207 1142
rect -269 754 -207 766
rect -177 1142 -111 1154
rect -177 766 -161 1142
rect -127 766 -111 1142
rect -177 754 -111 766
rect -81 1142 -15 1154
rect -81 766 -65 1142
rect -31 766 -15 1142
rect -81 754 -15 766
rect 15 1142 81 1154
rect 15 766 31 1142
rect 65 766 81 1142
rect 15 754 81 766
rect 111 1142 177 1154
rect 111 766 127 1142
rect 161 766 177 1142
rect 111 754 177 766
rect 207 1142 269 1154
rect 207 766 223 1142
rect 257 766 269 1142
rect 207 754 269 766
rect -269 506 -207 518
rect -269 130 -257 506
rect -223 130 -207 506
rect -269 118 -207 130
rect -177 506 -111 518
rect -177 130 -161 506
rect -127 130 -111 506
rect -177 118 -111 130
rect -81 506 -15 518
rect -81 130 -65 506
rect -31 130 -15 506
rect -81 118 -15 130
rect 15 506 81 518
rect 15 130 31 506
rect 65 130 81 506
rect 15 118 81 130
rect 111 506 177 518
rect 111 130 127 506
rect 161 130 177 506
rect 111 118 177 130
rect 207 506 269 518
rect 207 130 223 506
rect 257 130 269 506
rect 207 118 269 130
rect -269 -130 -207 -118
rect -269 -506 -257 -130
rect -223 -506 -207 -130
rect -269 -518 -207 -506
rect -177 -130 -111 -118
rect -177 -506 -161 -130
rect -127 -506 -111 -130
rect -177 -518 -111 -506
rect -81 -130 -15 -118
rect -81 -506 -65 -130
rect -31 -506 -15 -130
rect -81 -518 -15 -506
rect 15 -130 81 -118
rect 15 -506 31 -130
rect 65 -506 81 -130
rect 15 -518 81 -506
rect 111 -130 177 -118
rect 111 -506 127 -130
rect 161 -506 177 -130
rect 111 -518 177 -506
rect 207 -130 269 -118
rect 207 -506 223 -130
rect 257 -506 269 -130
rect 207 -518 269 -506
rect -269 -766 -207 -754
rect -269 -1142 -257 -766
rect -223 -1142 -207 -766
rect -269 -1154 -207 -1142
rect -177 -766 -111 -754
rect -177 -1142 -161 -766
rect -127 -1142 -111 -766
rect -177 -1154 -111 -1142
rect -81 -766 -15 -754
rect -81 -1142 -65 -766
rect -31 -1142 -15 -766
rect -81 -1154 -15 -1142
rect 15 -766 81 -754
rect 15 -1142 31 -766
rect 65 -1142 81 -766
rect 15 -1154 81 -1142
rect 111 -766 177 -754
rect 111 -1142 127 -766
rect 161 -1142 177 -766
rect 111 -1154 177 -1142
rect 207 -766 269 -754
rect 207 -1142 223 -766
rect 257 -1142 269 -766
rect 207 -1154 269 -1142
<< pdiffc >>
rect -257 766 -223 1142
rect -161 766 -127 1142
rect -65 766 -31 1142
rect 31 766 65 1142
rect 127 766 161 1142
rect 223 766 257 1142
rect -257 130 -223 506
rect -161 130 -127 506
rect -65 130 -31 506
rect 31 130 65 506
rect 127 130 161 506
rect 223 130 257 506
rect -257 -506 -223 -130
rect -161 -506 -127 -130
rect -65 -506 -31 -130
rect 31 -506 65 -130
rect 127 -506 161 -130
rect 223 -506 257 -130
rect -257 -1142 -223 -766
rect -161 -1142 -127 -766
rect -65 -1142 -31 -766
rect 31 -1142 65 -766
rect 127 -1142 161 -766
rect 223 -1142 257 -766
<< nsubdiff >>
rect -371 1303 -275 1337
rect 275 1303 371 1337
rect -371 1241 -337 1303
rect 337 1241 371 1303
rect -371 -1303 -337 -1241
rect 337 -1303 371 -1241
rect -371 -1337 -275 -1303
rect 275 -1337 371 -1303
<< nsubdiffcont >>
rect -275 1303 275 1337
rect -371 -1241 -337 1241
rect 337 -1241 371 1241
rect -275 -1337 275 -1303
<< poly >>
rect -225 1235 -159 1251
rect -225 1201 -209 1235
rect -175 1201 -159 1235
rect -225 1185 -159 1201
rect -33 1235 33 1251
rect -33 1201 -17 1235
rect 17 1201 33 1235
rect -33 1185 33 1201
rect 159 1235 225 1251
rect 159 1201 175 1235
rect 209 1201 225 1235
rect 159 1185 225 1201
rect -207 1154 -177 1185
rect -111 1154 -81 1180
rect -15 1154 15 1185
rect 81 1154 111 1180
rect 177 1154 207 1185
rect -207 728 -177 754
rect -111 723 -81 754
rect -15 728 15 754
rect 81 723 111 754
rect 177 728 207 754
rect -129 707 -63 723
rect -129 673 -113 707
rect -79 673 -63 707
rect -129 657 -63 673
rect 63 707 129 723
rect 63 673 79 707
rect 113 673 129 707
rect 63 657 129 673
rect -129 599 -63 615
rect -129 565 -113 599
rect -79 565 -63 599
rect -129 549 -63 565
rect 63 599 129 615
rect 63 565 79 599
rect 113 565 129 599
rect 63 549 129 565
rect -207 518 -177 544
rect -111 518 -81 549
rect -15 518 15 544
rect 81 518 111 549
rect 177 518 207 544
rect -207 87 -177 118
rect -111 92 -81 118
rect -15 87 15 118
rect 81 92 111 118
rect 177 87 207 118
rect -225 71 -159 87
rect -225 37 -209 71
rect -175 37 -159 71
rect -225 21 -159 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 159 71 225 87
rect 159 37 175 71
rect 209 37 225 71
rect 159 21 225 37
rect -225 -37 -159 -21
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -225 -87 -159 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 159 -37 225 -21
rect 159 -71 175 -37
rect 209 -71 225 -37
rect 159 -87 225 -71
rect -207 -118 -177 -87
rect -111 -118 -81 -92
rect -15 -118 15 -87
rect 81 -118 111 -92
rect 177 -118 207 -87
rect -207 -544 -177 -518
rect -111 -549 -81 -518
rect -15 -544 15 -518
rect 81 -549 111 -518
rect 177 -544 207 -518
rect -129 -565 -63 -549
rect -129 -599 -113 -565
rect -79 -599 -63 -565
rect -129 -615 -63 -599
rect 63 -565 129 -549
rect 63 -599 79 -565
rect 113 -599 129 -565
rect 63 -615 129 -599
rect -129 -673 -63 -657
rect -129 -707 -113 -673
rect -79 -707 -63 -673
rect -129 -723 -63 -707
rect 63 -673 129 -657
rect 63 -707 79 -673
rect 113 -707 129 -673
rect 63 -723 129 -707
rect -207 -754 -177 -728
rect -111 -754 -81 -723
rect -15 -754 15 -728
rect 81 -754 111 -723
rect 177 -754 207 -728
rect -207 -1185 -177 -1154
rect -111 -1180 -81 -1154
rect -15 -1185 15 -1154
rect 81 -1180 111 -1154
rect 177 -1185 207 -1154
rect -225 -1201 -159 -1185
rect -225 -1235 -209 -1201
rect -175 -1235 -159 -1201
rect -225 -1251 -159 -1235
rect -33 -1201 33 -1185
rect -33 -1235 -17 -1201
rect 17 -1235 33 -1201
rect -33 -1251 33 -1235
rect 159 -1201 225 -1185
rect 159 -1235 175 -1201
rect 209 -1235 225 -1201
rect 159 -1251 225 -1235
<< polycont >>
rect -209 1201 -175 1235
rect -17 1201 17 1235
rect 175 1201 209 1235
rect -113 673 -79 707
rect 79 673 113 707
rect -113 565 -79 599
rect 79 565 113 599
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect -113 -599 -79 -565
rect 79 -599 113 -565
rect -113 -707 -79 -673
rect 79 -707 113 -673
rect -209 -1235 -175 -1201
rect -17 -1235 17 -1201
rect 175 -1235 209 -1201
<< locali >>
rect -371 1303 -275 1337
rect 275 1303 371 1337
rect -371 1241 -337 1303
rect 337 1241 371 1303
rect -225 1201 -209 1235
rect -175 1201 -159 1235
rect -33 1201 -17 1235
rect 17 1201 33 1235
rect 159 1201 175 1235
rect 209 1201 225 1235
rect -257 1142 -223 1158
rect -257 750 -223 766
rect -161 1142 -127 1158
rect -161 750 -127 766
rect -65 1142 -31 1158
rect -65 750 -31 766
rect 31 1142 65 1158
rect 31 750 65 766
rect 127 1142 161 1158
rect 127 750 161 766
rect 223 1142 257 1158
rect 223 750 257 766
rect -129 673 -113 707
rect -79 673 -63 707
rect 63 673 79 707
rect 113 673 129 707
rect -129 565 -113 599
rect -79 565 -63 599
rect 63 565 79 599
rect 113 565 129 599
rect -257 506 -223 522
rect -257 114 -223 130
rect -161 506 -127 522
rect -161 114 -127 130
rect -65 506 -31 522
rect -65 114 -31 130
rect 31 506 65 522
rect 31 114 65 130
rect 127 506 161 522
rect 127 114 161 130
rect 223 506 257 522
rect 223 114 257 130
rect -225 37 -209 71
rect -175 37 -159 71
rect -33 37 -17 71
rect 17 37 33 71
rect 159 37 175 71
rect 209 37 225 71
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 159 -71 175 -37
rect 209 -71 225 -37
rect -257 -130 -223 -114
rect -257 -522 -223 -506
rect -161 -130 -127 -114
rect -161 -522 -127 -506
rect -65 -130 -31 -114
rect -65 -522 -31 -506
rect 31 -130 65 -114
rect 31 -522 65 -506
rect 127 -130 161 -114
rect 127 -522 161 -506
rect 223 -130 257 -114
rect 223 -522 257 -506
rect -129 -599 -113 -565
rect -79 -599 -63 -565
rect 63 -599 79 -565
rect 113 -599 129 -565
rect -129 -707 -113 -673
rect -79 -707 -63 -673
rect 63 -707 79 -673
rect 113 -707 129 -673
rect -257 -766 -223 -750
rect -257 -1158 -223 -1142
rect -161 -766 -127 -750
rect -161 -1158 -127 -1142
rect -65 -766 -31 -750
rect -65 -1158 -31 -1142
rect 31 -766 65 -750
rect 31 -1158 65 -1142
rect 127 -766 161 -750
rect 127 -1158 161 -1142
rect 223 -766 257 -750
rect 223 -1158 257 -1142
rect -225 -1235 -209 -1201
rect -175 -1235 -159 -1201
rect -33 -1235 -17 -1201
rect 17 -1235 33 -1201
rect 159 -1235 175 -1201
rect 209 -1235 225 -1201
rect -371 -1303 -337 -1241
rect 337 -1303 371 -1241
rect -371 -1337 -275 -1303
rect 275 -1337 371 -1303
<< viali >>
rect -209 1201 -175 1235
rect -17 1201 17 1235
rect 175 1201 209 1235
rect -257 766 -223 1142
rect -161 766 -127 1142
rect -65 766 -31 1142
rect 31 766 65 1142
rect 127 766 161 1142
rect 223 766 257 1142
rect -113 673 -79 707
rect 79 673 113 707
rect -113 565 -79 599
rect 79 565 113 599
rect -257 130 -223 506
rect -161 130 -127 506
rect -65 130 -31 506
rect 31 130 65 506
rect 127 130 161 506
rect 223 130 257 506
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect -257 -506 -223 -130
rect -161 -506 -127 -130
rect -65 -506 -31 -130
rect 31 -506 65 -130
rect 127 -506 161 -130
rect 223 -506 257 -130
rect -113 -599 -79 -565
rect 79 -599 113 -565
rect -113 -707 -79 -673
rect 79 -707 113 -673
rect -257 -1142 -223 -766
rect -161 -1142 -127 -766
rect -65 -1142 -31 -766
rect 31 -1142 65 -766
rect 127 -1142 161 -766
rect 223 -1142 257 -766
rect -209 -1235 -175 -1201
rect -17 -1235 17 -1201
rect 175 -1235 209 -1201
<< metal1 >>
rect -221 1235 -163 1241
rect -221 1201 -209 1235
rect -175 1201 -163 1235
rect -221 1195 -163 1201
rect -29 1235 29 1241
rect -29 1201 -17 1235
rect 17 1201 29 1235
rect -29 1195 29 1201
rect 163 1235 221 1241
rect 163 1201 175 1235
rect 209 1201 221 1235
rect 163 1195 221 1201
rect -263 1142 -217 1154
rect -263 766 -257 1142
rect -223 766 -217 1142
rect -263 754 -217 766
rect -167 1142 -121 1154
rect -167 766 -161 1142
rect -127 766 -121 1142
rect -167 754 -121 766
rect -71 1142 -25 1154
rect -71 766 -65 1142
rect -31 766 -25 1142
rect -71 754 -25 766
rect 25 1142 71 1154
rect 25 766 31 1142
rect 65 766 71 1142
rect 25 754 71 766
rect 121 1142 167 1154
rect 121 766 127 1142
rect 161 766 167 1142
rect 121 754 167 766
rect 217 1142 263 1154
rect 217 766 223 1142
rect 257 766 263 1142
rect 217 754 263 766
rect -125 707 -67 713
rect -125 673 -113 707
rect -79 673 -67 707
rect -125 667 -67 673
rect 67 707 125 713
rect 67 673 79 707
rect 113 673 125 707
rect 67 667 125 673
rect -125 599 -67 605
rect -125 565 -113 599
rect -79 565 -67 599
rect -125 559 -67 565
rect 67 599 125 605
rect 67 565 79 599
rect 113 565 125 599
rect 67 559 125 565
rect -263 506 -217 518
rect -263 130 -257 506
rect -223 130 -217 506
rect -263 118 -217 130
rect -167 506 -121 518
rect -167 130 -161 506
rect -127 130 -121 506
rect -167 118 -121 130
rect -71 506 -25 518
rect -71 130 -65 506
rect -31 130 -25 506
rect -71 118 -25 130
rect 25 506 71 518
rect 25 130 31 506
rect 65 130 71 506
rect 25 118 71 130
rect 121 506 167 518
rect 121 130 127 506
rect 161 130 167 506
rect 121 118 167 130
rect 217 506 263 518
rect 217 130 223 506
rect 257 130 263 506
rect 217 118 263 130
rect -221 71 -163 77
rect -221 37 -209 71
rect -175 37 -163 71
rect -221 31 -163 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 163 71 221 77
rect 163 37 175 71
rect 209 37 221 71
rect 163 31 221 37
rect -221 -37 -163 -31
rect -221 -71 -209 -37
rect -175 -71 -163 -37
rect -221 -77 -163 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 163 -37 221 -31
rect 163 -71 175 -37
rect 209 -71 221 -37
rect 163 -77 221 -71
rect -263 -130 -217 -118
rect -263 -506 -257 -130
rect -223 -506 -217 -130
rect -263 -518 -217 -506
rect -167 -130 -121 -118
rect -167 -506 -161 -130
rect -127 -506 -121 -130
rect -167 -518 -121 -506
rect -71 -130 -25 -118
rect -71 -506 -65 -130
rect -31 -506 -25 -130
rect -71 -518 -25 -506
rect 25 -130 71 -118
rect 25 -506 31 -130
rect 65 -506 71 -130
rect 25 -518 71 -506
rect 121 -130 167 -118
rect 121 -506 127 -130
rect 161 -506 167 -130
rect 121 -518 167 -506
rect 217 -130 263 -118
rect 217 -506 223 -130
rect 257 -506 263 -130
rect 217 -518 263 -506
rect -125 -565 -67 -559
rect -125 -599 -113 -565
rect -79 -599 -67 -565
rect -125 -605 -67 -599
rect 67 -565 125 -559
rect 67 -599 79 -565
rect 113 -599 125 -565
rect 67 -605 125 -599
rect -125 -673 -67 -667
rect -125 -707 -113 -673
rect -79 -707 -67 -673
rect -125 -713 -67 -707
rect 67 -673 125 -667
rect 67 -707 79 -673
rect 113 -707 125 -673
rect 67 -713 125 -707
rect -263 -766 -217 -754
rect -263 -1142 -257 -766
rect -223 -1142 -217 -766
rect -263 -1154 -217 -1142
rect -167 -766 -121 -754
rect -167 -1142 -161 -766
rect -127 -1142 -121 -766
rect -167 -1154 -121 -1142
rect -71 -766 -25 -754
rect -71 -1142 -65 -766
rect -31 -1142 -25 -766
rect -71 -1154 -25 -1142
rect 25 -766 71 -754
rect 25 -1142 31 -766
rect 65 -1142 71 -766
rect 25 -1154 71 -1142
rect 121 -766 167 -754
rect 121 -1142 127 -766
rect 161 -1142 167 -766
rect 121 -1154 167 -1142
rect 217 -766 263 -754
rect 217 -1142 223 -766
rect 257 -1142 263 -766
rect 217 -1154 263 -1142
rect -221 -1201 -163 -1195
rect -221 -1235 -209 -1201
rect -175 -1235 -163 -1201
rect -221 -1241 -163 -1235
rect -29 -1201 29 -1195
rect -29 -1235 -17 -1201
rect 17 -1235 29 -1201
rect -29 -1241 29 -1235
rect 163 -1201 221 -1195
rect 163 -1235 175 -1201
rect 209 -1235 221 -1201
rect 163 -1241 221 -1235
<< properties >>
string FIXED_BBOX -354 -1320 354 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
