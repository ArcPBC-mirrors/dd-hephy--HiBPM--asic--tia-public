magic
tech sky130A
magscale 1 2
timestamp 1687287864
<< error_s >>
rect 47740 77378 47744 77394
rect 68740 77378 68744 77394
rect 89740 77378 89744 77394
rect 110740 77378 110744 77394
rect 47744 77158 47747 77378
rect 68744 77158 68747 77378
rect 89744 77158 89747 77378
rect 110744 77158 110747 77378
rect 34987 77109 35215 77125
rect 55987 77109 56215 77125
rect 76987 77109 77215 77125
rect 97987 77109 98215 77125
rect 34984 77098 34987 77109
rect 55984 77098 55987 77109
rect 76984 77098 76987 77109
rect 97984 77098 97987 77109
rect 48004 64642 48016 64662
rect 69004 64642 69016 64662
rect 90004 64642 90016 64662
rect 111004 64642 111016 64662
rect 47780 64635 48004 64642
rect 68780 64635 69004 64642
rect 89780 64635 90004 64642
rect 110780 64635 111004 64642
rect 35253 64382 35256 64390
rect 56253 64382 56256 64390
rect 77253 64382 77256 64602
rect 98253 64382 98256 64390
rect 35256 64366 35260 64382
rect 56256 64366 56260 64382
rect 77256 64366 77260 64382
rect 98256 64366 98260 64382
rect 30178 52413 30180 52497
rect 30262 52372 30264 52413
rect 115820 52372 115822 52497
rect 13138 42004 13158 42016
rect 145298 42013 145309 42016
rect 13158 41780 13165 42004
rect 145309 41785 145325 42013
rect 422 41744 642 41747
rect 132582 41744 132802 41747
rect 406 41740 422 41744
rect 132566 41740 132582 41744
rect 13418 29256 13434 29260
rect 145578 29256 145594 29260
rect 13198 29253 13418 29256
rect 145358 29253 145578 29256
rect 675 28987 691 29215
rect 132835 28996 132842 29220
rect 691 28984 702 28987
rect 132842 28984 132862 28996
rect 13138 21004 13158 21016
rect 145298 21013 145309 21016
rect 13158 20780 13165 21004
rect 145309 20785 145325 21013
rect 422 20744 642 20747
rect 132582 20744 132802 20747
rect 406 20740 422 20744
rect 132566 20740 132582 20744
rect 13418 8256 13434 8260
rect 145578 8256 145594 8260
rect 13198 8253 13418 8256
rect 145358 8253 145578 8256
rect 675 7987 691 8215
rect 132835 7996 132842 8220
rect 691 7984 702 7987
rect 132842 7984 132862 7996
rect 1583 0 2483 315
rect 13138 4 13158 16
rect 145298 13 145309 16
rect 13158 -220 13165 4
rect 145309 -215 145325 13
rect 422 -256 642 -253
rect 132582 -256 132802 -253
rect 406 -489 422 -256
rect 13252 -310 13472 -307
rect 13472 -543 13488 -310
rect 132566 -489 132582 -256
rect 145537 -310 145632 -307
rect 145632 -543 145648 -310
rect 102 -576 322 -573
rect 86 -809 102 -576
rect 132256 -582 132482 -573
rect 13572 -640 13802 -627
rect 13802 -863 13808 -640
rect 132246 -809 132256 -582
rect 145732 -630 145952 -627
rect 145952 -747 145968 -630
rect -218 -896 2 -893
rect 131942 -896 132162 -893
rect -234 -1026 -218 -896
rect 13892 -950 14112 -947
rect 14112 -1183 14128 -950
rect 131926 -1129 131942 -896
rect 146069 -950 146272 -947
rect 146272 -1016 146288 -950
rect -580 -1258 -360 -1255
rect 131580 -1258 131800 -1255
rect -596 -1282 -580 -1258
rect 14200 -1282 14436 -1269
rect 131564 -1282 131580 -1258
rect 146360 -1282 146596 -1269
rect 3275 -1477 3309 -1443
rect 6297 -1477 6331 -1443
rect 139669 -1477 139703 -1443
rect 142691 -1477 142725 -1443
rect 3275 -1515 3347 -1479
rect 6259 -1515 6331 -1479
rect 139669 -1515 139741 -1479
rect 142653 -1515 142725 -1479
rect 3275 -11521 3347 -11485
rect 6259 -11521 6331 -11485
rect 139669 -11521 139741 -11485
rect 142653 -11521 142725 -11485
rect 3275 -11557 3309 -11523
rect 6297 -11557 6331 -11523
rect 139669 -11557 139703 -11523
rect 142691 -11557 142725 -11523
rect -596 -11731 -360 -11718
rect 14420 -11742 14436 -11718
rect 131564 -11731 131800 -11718
rect 146580 -11742 146596 -11718
rect 14200 -11745 14420 -11742
rect 146360 -11745 146580 -11742
rect -288 -12050 -272 -11984
rect -272 -12053 -69 -12050
rect 14058 -12104 14074 -11871
rect 131872 -12050 131888 -11817
rect 131888 -12053 132108 -12050
rect 146218 -12104 146234 -11974
rect 13838 -12107 14058 -12104
rect 145998 -12107 146218 -12104
rect 32 -12370 48 -12253
rect 48 -12373 268 -12370
rect 13744 -12418 13754 -12191
rect 132192 -12360 132198 -12137
rect 132198 -12373 132428 -12360
rect 13518 -12427 13744 -12418
rect 145898 -12424 145914 -12191
rect 145678 -12427 145898 -12424
rect 352 -12690 368 -12457
rect 368 -12693 463 -12690
rect 13418 -12744 13434 -12511
rect 132512 -12690 132528 -12457
rect 132528 -12693 132748 -12690
rect 145578 -12744 145594 -12511
rect 13198 -12747 13418 -12744
rect 145358 -12747 145578 -12744
rect 675 -13013 691 -12785
rect 132835 -13004 132842 -12780
rect 691 -13016 702 -13013
rect 132842 -13016 132862 -13004
rect 13138 -20996 13158 -20984
rect 145298 -20987 145309 -20984
rect 13158 -21220 13165 -20996
rect 145309 -21215 145325 -20987
rect 422 -21256 642 -21253
rect 132582 -21256 132802 -21253
rect 406 -21489 422 -21256
rect 13252 -21310 13472 -21307
rect 13472 -21543 13488 -21310
rect 132566 -21489 132582 -21256
rect 145537 -21310 145632 -21307
rect 145632 -21543 145648 -21310
rect 102 -21576 322 -21573
rect 86 -21809 102 -21576
rect 132256 -21582 132482 -21573
rect 13572 -21640 13802 -21627
rect 13802 -21863 13808 -21640
rect 132246 -21809 132256 -21582
rect 145732 -21630 145952 -21627
rect 145952 -21747 145968 -21630
rect -218 -21896 2 -21893
rect 131942 -21896 132162 -21893
rect -234 -22026 -218 -21896
rect 13892 -21950 14112 -21947
rect 14112 -22183 14128 -21950
rect 131926 -22129 131942 -21896
rect 146069 -21950 146272 -21947
rect 146272 -22183 146288 -21950
rect -580 -22258 -360 -22255
rect 131580 -22258 131800 -22255
rect -596 -22282 -580 -22258
rect 14200 -22282 14436 -22269
rect 131564 -22282 131580 -22258
rect 146360 -22282 146596 -22269
rect 3275 -22477 3309 -22443
rect 6297 -22477 6331 -22443
rect 3275 -22515 3347 -22479
rect 6259 -22515 6331 -22479
rect 3275 -32521 3347 -32485
rect 6259 -32521 6331 -32485
rect 3275 -32557 3309 -32523
rect 6297 -32557 6331 -32523
rect -596 -32731 -360 -32718
rect 14420 -32742 14436 -32718
rect 131564 -32731 131800 -32718
rect 146580 -32742 146596 -32718
rect 14200 -32745 14420 -32742
rect 146360 -32745 146580 -32742
rect -288 -33050 -272 -32984
rect -272 -33053 -69 -33050
rect 14058 -33104 14074 -32871
rect 131872 -33050 131888 -32817
rect 131888 -33053 132108 -33050
rect 146218 -33104 146234 -32871
rect 13838 -33107 14058 -33104
rect 145998 -33107 146218 -33104
rect 32 -33370 48 -33253
rect 48 -33373 268 -33370
rect 13744 -33418 13754 -33191
rect 132192 -33360 132198 -33137
rect 132198 -33373 132428 -33360
rect 13518 -33427 13744 -33418
rect 145898 -33424 145914 -33191
rect 145678 -33427 145898 -33424
rect 352 -33690 368 -33457
rect 368 -33693 463 -33690
rect 13418 -33744 13434 -33511
rect 132512 -33690 132528 -33457
rect 132528 -33693 132748 -33690
rect 145578 -33744 145594 -33511
rect 13198 -33747 13418 -33744
rect 145358 -33747 145578 -33744
rect 675 -34013 691 -33785
rect 132835 -34004 132842 -33780
rect 691 -34016 702 -34013
rect 132842 -34016 132862 -34004
rect 13138 -41996 13158 -41984
rect 145298 -41987 145309 -41984
rect 13158 -42220 13165 -41996
rect 145309 -42215 145325 -41987
rect 422 -42256 642 -42253
rect 132582 -42256 132802 -42253
rect 406 -42489 422 -42256
rect 13252 -42310 13472 -42307
rect 13472 -42543 13488 -42310
rect 132566 -42489 132582 -42256
rect 145537 -42310 145632 -42307
rect 145632 -42543 145648 -42310
rect 102 -42576 322 -42573
rect 86 -42809 102 -42576
rect 132256 -42582 132482 -42573
rect 13572 -42640 13802 -42627
rect 13802 -42863 13808 -42640
rect 132246 -42809 132256 -42582
rect 145732 -42630 145952 -42627
rect 145952 -42747 145968 -42630
rect -218 -42896 2 -42893
rect 131942 -42896 132162 -42893
rect -234 -43129 -218 -42896
rect 13892 -42950 14112 -42947
rect 14112 -43183 14128 -42950
rect 131926 -43129 131942 -42896
rect 146069 -42950 146272 -42947
rect 146272 -43016 146288 -42950
rect -580 -43258 -360 -43255
rect 131580 -43258 131800 -43255
rect -596 -43282 -580 -43258
rect 14200 -43282 14436 -43269
rect 131564 -43282 131580 -43258
rect 146360 -43282 146596 -43269
rect 139669 -43477 139703 -43443
rect 142691 -43477 142725 -43443
rect 139669 -43515 139741 -43479
rect 142653 -43515 142725 -43479
rect 139669 -53521 139741 -53485
rect 142653 -53521 142725 -53485
rect 139669 -53557 139703 -53523
rect 142691 -53557 142725 -53523
rect -596 -53731 -360 -53718
rect 14420 -53742 14436 -53718
rect 131564 -53731 131800 -53718
rect 146580 -53742 146596 -53718
rect 14200 -53745 14420 -53742
rect 146360 -53745 146580 -53742
rect -288 -54050 -272 -53817
rect -272 -54053 -69 -54050
rect 14058 -54104 14074 -53871
rect 131872 -54050 131888 -53817
rect 131888 -54053 132108 -54050
rect 146218 -54104 146234 -53974
rect 13838 -54107 14058 -54104
rect 145998 -54107 146218 -54104
rect 32 -54370 48 -54253
rect 48 -54373 268 -54370
rect 13744 -54418 13754 -54191
rect 132192 -54360 132198 -54137
rect 132198 -54373 132428 -54360
rect 13518 -54427 13744 -54418
rect 145898 -54424 145914 -54191
rect 145678 -54427 145898 -54424
rect 352 -54690 368 -54457
rect 368 -54693 463 -54690
rect 13418 -54744 13434 -54511
rect 132512 -54690 132528 -54457
rect 132528 -54693 132748 -54690
rect 145578 -54744 145594 -54511
rect 13198 -54747 13418 -54744
rect 145358 -54747 145578 -54744
rect 675 -55013 691 -54785
rect 132835 -55004 132842 -54780
rect 691 -55016 702 -55013
rect 132842 -55016 132862 -55004
rect 47740 -77382 47744 -77366
rect 68740 -77382 68744 -77366
rect 89540 -77382 89744 -77366
rect 110740 -77382 110744 -77366
rect 47744 -77390 47747 -77382
rect 68744 -77390 68747 -77382
rect 89744 -77602 89747 -77382
rect 110744 -77390 110747 -77382
rect 34996 -77642 35220 -77635
rect 55996 -77642 56220 -77635
rect 76996 -77642 77220 -77635
rect 97996 -77642 98220 -77635
rect 34984 -77662 34996 -77642
rect 55984 -77662 55996 -77642
rect 76984 -77662 76996 -77642
rect 97984 -77662 97996 -77642
rect 48013 -90109 48016 -90098
rect 69013 -90109 69016 -90098
rect 90013 -90109 90016 -90098
rect 111013 -90109 111016 -90098
rect 47785 -90125 48013 -90109
rect 68785 -90125 69013 -90109
rect 89785 -90125 90013 -90109
rect 110785 -90125 111013 -90109
rect 35253 -90378 35256 -90158
rect 56253 -90378 56256 -90337
rect 77253 -90378 77256 -90158
rect 35256 -90394 35260 -90378
rect 56256 -90380 56258 -90378
rect 56258 -90394 56260 -90380
rect 77256 -90394 77260 -90378
rect 89690 -90432 89693 -90337
rect 98253 -90378 98256 -90158
rect 98256 -90394 98260 -90378
rect 89540 -90448 89690 -90432
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_0 ~/code/hibpm-sky130a-tapeout/mag/frame/io_pdk
timestamp 1683767628
transform 0 -1 34000 1 0 -35000
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_1
timestamp 1683767628
transform -1 0 112000 0 -1 -56800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_2
timestamp 1683767628
transform 0 -1 34000 1 0 -14000
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_3
timestamp 1683767628
transform -1 0 70000 0 -1 -56800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_5
timestamp 1683767628
transform 0 1 112000 -1 0 43000
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_6
timestamp 1683767628
transform 1 0 55000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_7
timestamp 1683767628
transform 1 0 97000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_8
timestamp 1683767628
transform 0 1 112000 -1 0 -41000
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_9
timestamp 1683767628
transform 1 0 34000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_10
timestamp 1683767628
transform -1 0 49000 0 -1 -56800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_13
timestamp 1683767628
transform 0 -1 34000 1 0 7000
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_14
timestamp 1683767628
transform 0 1 112000 -1 0 1000
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_0 ~/code/hibpm-sky130a-tapeout/mag/frame/io_pdk
timestamp 1683767628
transform 0 -1 33593 1 0 -37000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_1
timestamp 1683767628
transform 0 -1 33593 1 0 26000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_2
timestamp 1683767628
transform 0 -1 33593 1 0 -16000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_3
timestamp 1683767628
transform 0 -1 33593 1 0 5000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_4
timestamp 1683767628
transform 1 0 74000 0 1 44207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_5
timestamp 1683767628
transform -1 0 76000 0 -1 -57207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_6
timestamp 1683767628
transform 0 1 112407 -1 0 -35000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_7
timestamp 1683767628
transform 1 0 95000 0 1 44207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_8
timestamp 1683767628
transform 0 1 112407 -1 0 7000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_9
timestamp 1683767628
transform 1 0 53000 0 1 44207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_10
timestamp 1683767628
transform -1 0 55000 0 -1 -57207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_11
timestamp 1683767628
transform -1 0 97000 0 -1 -57207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_12
timestamp 1683767628
transform 0 1 112407 -1 0 -14000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_13
timestamp 1683767628
transform 0 1 112407 -1 0 24000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_0 ~/code/hibpm-sky130a-tapeout/mag/frame/io_pdk
timestamp 1683767628
transform 0 -1 33593 1 0 -41000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_1
timestamp 1683767628
transform 0 -1 33593 1 0 -20000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_2
timestamp 1683767628
transform 0 -1 33593 1 0 22000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_3
timestamp 1683767628
transform 0 -1 33593 1 0 1000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_4
timestamp 1683767628
transform 1 0 70000 0 1 44207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_5
timestamp 1683767628
transform -1 0 74000 0 -1 -57207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_6
timestamp 1683767628
transform 0 1 112407 -1 0 -37000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_7
timestamp 1683767628
transform 1 0 91000 0 1 44207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_8
timestamp 1683767628
transform 0 1 112407 -1 0 5000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_9
timestamp 1683767628
transform 1 0 49000 0 1 44207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_10
timestamp 1683767628
transform -1 0 53000 0 -1 -57207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_11
timestamp 1683767628
transform -1 0 94800 0 -1 -57207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_13
timestamp 1683767628
transform 0 1 112407 -1 0 28000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_14
timestamp 1683767628
transform -1 0 95000 0 -1 -57207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_15
timestamp 1683767628
transform 0 1 112407 -1 0 -16000
box 0 0 4000 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_0 ~/code/hibpm-sky130a-tapeout/mag/frame/io_pdk
timestamp 1683767628
transform 1 0 112000 0 1 43000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_1
timestamp 1683767628
transform 1 0 112000 0 -1 -56000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_3
timestamp 1683767628
transform -1 0 34000 0 -1 -56000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_4
timestamp 1683767628
transform -1 0 34000 0 1 43000
box 0 0 40000 40800
use sky130_ef_io__vddio_lvc_clamped_pad  sky130_ef_io__vddio_lvc_clamped_pad_0 ~/code/hibpm-sky130a-tapeout/mag/frame/io_pdk
timestamp 1683767628
transform 0 -1 33593 1 0 28000
box 0 -7 15000 39593
use sky130_ef_io__vssio_lvc_clamped_pad  sky130_ef_io__vssio_lvc_clamped_pad_0 ~/code/hibpm-sky130a-tapeout/mag/frame/io_pdk
timestamp 1683767628
transform 0 -1 33593 1 0 -56000
box 0 -7 15000 39593
use sky130_ef_io__vssio_lvc_clamped_pad  sky130_ef_io__vssio_lvc_clamped_pad_1
timestamp 1683767628
transform -1 0 91000 0 -1 -57207
box 0 -7 15000 39593
use sky130_ef_io__vssio_lvc_clamped_pad  sky130_ef_io__vssio_lvc_clamped_pad_2
timestamp 1683767628
transform 0 1 112407 -1 0 -20000
box 0 -7 15000 39593
use sky130_ef_io__vssio_lvc_clamped_pad  sky130_ef_io__vssio_lvc_clamped_pad_3
timestamp 1683767628
transform 0 1 112407 -1 0 22000
box 0 -7 15000 39593
use sky130_ef_io__vssio_lvc_clamped_pad  sky130_ef_io__vssio_lvc_clamped_pad_4
timestamp 1683767628
transform 1 0 76000 0 1 44207
box 0 -7 15000 39593
<< end >>
