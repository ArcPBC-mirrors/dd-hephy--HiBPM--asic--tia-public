magic
tech sky130A
magscale 1 2
timestamp 1683736741
<< pwell >>
rect -425 -1028 425 1028
<< nmoslvt >>
rect -229 418 -29 818
rect 29 418 229 818
rect -229 -200 -29 200
rect 29 -200 229 200
rect -229 -818 -29 -418
rect 29 -818 229 -418
<< ndiff >>
rect -287 806 -229 818
rect -287 430 -275 806
rect -241 430 -229 806
rect -287 418 -229 430
rect -29 806 29 818
rect -29 430 -17 806
rect 17 430 29 806
rect -29 418 29 430
rect 229 806 287 818
rect 229 430 241 806
rect 275 430 287 806
rect 229 418 287 430
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect -287 -430 -229 -418
rect -287 -806 -275 -430
rect -241 -806 -229 -430
rect -287 -818 -229 -806
rect -29 -430 29 -418
rect -29 -806 -17 -430
rect 17 -806 29 -430
rect -29 -818 29 -806
rect 229 -430 287 -418
rect 229 -806 241 -430
rect 275 -806 287 -430
rect 229 -818 287 -806
<< ndiffc >>
rect -275 430 -241 806
rect -17 430 17 806
rect 241 430 275 806
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect -275 -806 -241 -430
rect -17 -806 17 -430
rect 241 -806 275 -430
<< psubdiff >>
rect -389 958 -293 992
rect 293 958 389 992
rect -389 896 -355 958
rect 355 896 389 958
rect -389 -958 -355 -896
rect 355 -958 389 -896
rect -389 -992 -293 -958
rect 293 -992 389 -958
<< psubdiffcont >>
rect -293 958 293 992
rect -389 -896 -355 896
rect 355 -896 389 896
rect -293 -992 293 -958
<< poly >>
rect -229 890 -29 906
rect -229 856 -213 890
rect -45 856 -29 890
rect -229 818 -29 856
rect 29 890 229 906
rect 29 856 45 890
rect 213 856 229 890
rect 29 818 229 856
rect -229 380 -29 418
rect -229 346 -213 380
rect -45 346 -29 380
rect -229 330 -29 346
rect 29 380 229 418
rect 29 346 45 380
rect 213 346 229 380
rect 29 330 229 346
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect -229 -346 -29 -330
rect -229 -380 -213 -346
rect -45 -380 -29 -346
rect -229 -418 -29 -380
rect 29 -346 229 -330
rect 29 -380 45 -346
rect 213 -380 229 -346
rect 29 -418 229 -380
rect -229 -856 -29 -818
rect -229 -890 -213 -856
rect -45 -890 -29 -856
rect -229 -906 -29 -890
rect 29 -856 229 -818
rect 29 -890 45 -856
rect 213 -890 229 -856
rect 29 -906 229 -890
<< polycont >>
rect -213 856 -45 890
rect 45 856 213 890
rect -213 346 -45 380
rect 45 346 213 380
rect -213 238 -45 272
rect 45 238 213 272
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect -213 -380 -45 -346
rect 45 -380 213 -346
rect -213 -890 -45 -856
rect 45 -890 213 -856
<< locali >>
rect -389 958 -293 992
rect 293 958 389 992
rect -389 896 -355 958
rect 355 896 389 958
rect -229 856 -213 890
rect -45 856 -29 890
rect 29 856 45 890
rect 213 856 229 890
rect -275 806 -241 822
rect -275 414 -241 430
rect -17 806 17 822
rect -17 414 17 430
rect 241 806 275 822
rect 241 414 275 430
rect -229 346 -213 380
rect -45 346 -29 380
rect 29 346 45 380
rect 213 346 229 380
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect -229 -380 -213 -346
rect -45 -380 -29 -346
rect 29 -380 45 -346
rect 213 -380 229 -346
rect -275 -430 -241 -414
rect -275 -822 -241 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 241 -430 275 -414
rect 241 -822 275 -806
rect -229 -890 -213 -856
rect -45 -890 -29 -856
rect 29 -890 45 -856
rect 213 -890 229 -856
rect -389 -958 -355 -896
rect 355 -958 389 -896
rect -389 -992 -293 -958
rect 293 -992 389 -958
<< viali >>
rect -213 856 -45 890
rect 45 856 213 890
rect -275 430 -241 806
rect -17 430 17 806
rect 241 430 275 806
rect -213 346 -45 380
rect 45 346 213 380
rect -213 238 -45 272
rect 45 238 213 272
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect -213 -380 -45 -346
rect 45 -380 213 -346
rect -275 -806 -241 -430
rect -17 -806 17 -430
rect 241 -806 275 -430
rect -213 -890 -45 -856
rect 45 -890 213 -856
<< metal1 >>
rect -225 890 -33 896
rect -225 856 -213 890
rect -45 856 -33 890
rect -225 850 -33 856
rect 33 890 225 896
rect 33 856 45 890
rect 213 856 225 890
rect 33 850 225 856
rect -281 806 -235 818
rect -281 430 -275 806
rect -241 430 -235 806
rect -281 418 -235 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 235 806 281 818
rect 235 430 241 806
rect 275 430 281 806
rect 235 418 281 430
rect -225 380 -33 386
rect -225 346 -213 380
rect -45 346 -33 380
rect -225 340 -33 346
rect 33 380 225 386
rect 33 346 45 380
rect 213 346 225 380
rect 33 340 225 346
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
rect -225 -346 -33 -340
rect -225 -380 -213 -346
rect -45 -380 -33 -346
rect -225 -386 -33 -380
rect 33 -346 225 -340
rect 33 -380 45 -346
rect 213 -380 225 -346
rect 33 -386 225 -380
rect -281 -430 -235 -418
rect -281 -806 -275 -430
rect -241 -806 -235 -430
rect -281 -818 -235 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 235 -430 281 -418
rect 235 -806 241 -430
rect 275 -806 281 -430
rect 235 -818 281 -806
rect -225 -856 -33 -850
rect -225 -890 -213 -856
rect -45 -890 -33 -856
rect -225 -896 -33 -890
rect 33 -856 225 -850
rect 33 -890 45 -856
rect 213 -890 225 -856
rect 33 -896 225 -890
<< properties >>
string FIXED_BBOX -372 -975 372 975
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 1 m 3 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
