magic
tech sky130A
magscale 1 2
timestamp 1684930430
<< dnwell >>
rect 2776 3372 5220 5860
<< nwell >>
rect 2696 5654 5300 5940
rect 2696 3578 2982 5654
rect 5014 3578 5300 5654
rect 2696 3292 5300 3578
<< nsubdiff >>
rect 2733 5883 5263 5903
rect 2733 5849 2813 5883
rect 5183 5849 5263 5883
rect 2733 5829 5263 5849
rect 2733 5823 2807 5829
rect 2733 3409 2753 5823
rect 2787 3409 2807 5823
rect 2733 3403 2807 3409
rect 5189 5823 5263 5829
rect 5189 3409 5209 5823
rect 5243 3409 5263 5823
rect 5189 3403 5263 3409
rect 2733 3383 5263 3403
rect 2733 3349 2813 3383
rect 5183 3349 5263 3383
rect 2733 3329 5263 3349
<< nsubdiffcont >>
rect 2813 5849 5183 5883
rect 2753 3409 2787 5823
rect 5209 3409 5243 5823
rect 2813 3349 5183 3383
<< locali >>
rect 2753 5849 2813 5883
rect 5183 5849 5243 5883
rect 2753 5823 2787 5849
rect 5209 5823 5243 5849
rect 4100 4780 4160 4980
rect 3060 4460 3160 4560
rect 3060 3820 3160 3920
rect 4248 3636 4400 4984
rect 4240 3616 4416 3636
rect 2753 3383 2787 3409
rect 5209 3383 5243 3409
rect 2753 3349 2813 3383
rect 5183 3349 5243 3383
rect 3036 3340 3864 3349
<< viali >>
rect 3320 880 3600 1000
<< metal1 >>
rect 3180 4840 4264 4948
rect 3240 4808 3288 4840
rect 3432 4808 3480 4840
rect 3624 4808 3672 4840
rect 3816 4808 3856 4840
rect 4008 4808 4048 4840
rect 3226 4628 3236 4808
rect 3288 4628 3298 4808
rect 3418 4628 3428 4808
rect 3480 4628 3490 4808
rect 3610 4628 3620 4808
rect 3672 4628 3682 4808
rect 3802 4628 3812 4808
rect 3864 4628 3874 4808
rect 3994 4628 4004 4808
rect 4056 4628 4066 4808
rect 3816 4612 3856 4628
rect 4008 4600 4048 4628
rect 3130 4408 3140 4588
rect 3192 4408 3202 4588
rect 3322 4408 3332 4588
rect 3384 4408 3394 4588
rect 3514 4408 3524 4588
rect 3576 4408 3586 4588
rect 3706 4408 3716 4588
rect 3768 4408 3778 4588
rect 3898 4408 3908 4588
rect 3960 4408 3970 4588
rect 4090 4408 4100 4588
rect 4152 4408 4162 4588
rect 4192 4376 4264 4840
rect 3276 4220 4824 4376
rect 3226 4012 3236 4192
rect 3288 4012 3298 4192
rect 3418 4012 3428 4192
rect 3480 4012 3490 4192
rect 3610 4012 3620 4192
rect 3672 4012 3682 4192
rect 3802 4012 3812 4192
rect 3864 4012 3874 4192
rect 3994 4012 4004 4192
rect 4056 4012 4066 4192
rect 3130 3788 3140 3968
rect 3192 3788 3202 3968
rect 3322 3788 3332 3968
rect 3384 3788 3394 3968
rect 3514 3788 3524 3968
rect 3576 3788 3586 3968
rect 3706 3788 3716 3968
rect 3768 3788 3778 3968
rect 3898 3788 3908 3968
rect 3960 3788 3970 3968
rect 4090 3788 4100 3968
rect 4152 3788 4162 3968
rect 4196 3760 4264 4220
rect 3176 3652 4264 3760
rect 4564 3088 4700 3768
rect 3144 3004 3192 3088
rect 3336 3004 3384 3028
rect 3528 3004 3576 3024
rect 3720 3004 3768 3028
rect 3868 3004 4700 3088
rect 3144 2872 3192 2972
rect 3336 2884 3384 2972
rect 3528 2880 3576 2972
rect 3720 2884 3768 2972
rect 3224 2532 3300 2596
rect 3416 2528 3492 2592
rect 3608 2524 3684 2588
rect 3308 1000 3612 1006
rect 3308 880 3320 1000
rect 3600 880 3612 1000
rect 3308 874 3612 880
<< via1 >>
rect 3236 4628 3288 4808
rect 3428 4628 3480 4808
rect 3620 4628 3672 4808
rect 3812 4628 3864 4808
rect 4004 4628 4056 4808
rect 3140 4408 3192 4588
rect 3332 4408 3384 4588
rect 3524 4408 3576 4588
rect 3716 4408 3768 4588
rect 3908 4408 3960 4588
rect 4100 4408 4152 4588
rect 3236 4012 3288 4192
rect 3428 4012 3480 4192
rect 3620 4012 3672 4192
rect 3812 4012 3864 4192
rect 4004 4012 4056 4192
rect 3140 3788 3192 3968
rect 3332 3788 3384 3968
rect 3524 3788 3576 3968
rect 3716 3788 3768 3968
rect 3908 3788 3960 3968
rect 4100 3788 4152 3968
rect 3320 880 3600 1000
<< metal2 >>
rect 3236 4884 4060 4900
rect 3236 4808 3520 4884
rect 3852 4808 4060 4884
rect 3288 4640 3428 4808
rect 3236 4618 3288 4628
rect 3480 4652 3520 4808
rect 3480 4640 3620 4652
rect 3428 4618 3480 4628
rect 3672 4640 3812 4652
rect 3620 4618 3672 4628
rect 3864 4640 4004 4808
rect 3812 4618 3864 4628
rect 4056 4640 4060 4808
rect 4004 4618 4056 4628
rect 3140 4588 3192 4598
rect 3072 4568 3140 4578
rect 3332 4588 3384 4598
rect 3192 4568 3332 4580
rect 3524 4588 3576 4598
rect 3384 4568 3524 4580
rect 3404 4408 3524 4568
rect 3716 4588 3768 4598
rect 3576 4408 3716 4580
rect 3908 4588 3960 4598
rect 3768 4408 3908 4580
rect 4100 4588 4152 4598
rect 3960 4408 4100 4580
rect 3404 4336 4152 4408
rect 3072 4326 4152 4336
rect 3140 4320 4152 4326
rect 3236 4264 4056 4280
rect 3236 4192 3520 4264
rect 3852 4192 4056 4264
rect 3288 4020 3428 4192
rect 3236 4002 3288 4012
rect 3480 4032 3520 4192
rect 3480 4020 3620 4032
rect 3428 4002 3480 4012
rect 3672 4020 3812 4032
rect 3620 4002 3672 4012
rect 3864 4020 4004 4192
rect 3812 4002 3864 4012
rect 4004 4002 4056 4012
rect 3140 3968 3192 3978
rect 3072 3944 3140 3954
rect 3332 3968 3384 3978
rect 3192 3944 3332 3960
rect 3524 3968 3576 3978
rect 3384 3944 3524 3960
rect 3404 3788 3524 3944
rect 3716 3968 3768 3978
rect 3576 3788 3716 3960
rect 3908 3968 3960 3978
rect 3768 3788 3908 3960
rect 4100 3968 4152 3978
rect 3960 3788 4100 3960
rect 3404 3712 4152 3788
rect 3072 3702 4152 3712
rect 3140 3700 4152 3702
rect 3252 2708 3640 2718
rect 3252 2206 3640 2216
rect 3140 1000 3900 1260
rect 3140 920 3320 1000
rect 3600 920 3900 1000
rect 3320 870 3600 880
<< via2 >>
rect 3520 4808 3852 4884
rect 3520 4652 3620 4808
rect 3620 4652 3672 4808
rect 3672 4652 3812 4808
rect 3812 4652 3852 4808
rect 3072 4408 3140 4568
rect 3140 4408 3192 4568
rect 3192 4408 3332 4568
rect 3332 4408 3384 4568
rect 3384 4408 3404 4568
rect 3072 4336 3404 4408
rect 3520 4192 3852 4264
rect 3520 4032 3620 4192
rect 3620 4032 3672 4192
rect 3672 4032 3812 4192
rect 3812 4032 3852 4192
rect 3072 3788 3140 3944
rect 3140 3788 3192 3944
rect 3192 3788 3332 3944
rect 3332 3788 3384 3944
rect 3384 3788 3404 3944
rect 3072 3712 3404 3788
rect 3252 2216 3640 2708
<< metal3 >>
rect 3508 4884 3876 5064
rect 3508 4652 3520 4884
rect 3852 4652 3876 4884
rect 3056 4568 3420 4580
rect 3056 4336 3072 4568
rect 3404 4336 3420 4568
rect 3056 3944 3420 4336
rect 3508 4264 3876 4652
rect 3508 4032 3520 4264
rect 3852 4032 3876 4264
rect 3508 4016 3876 4032
rect 3056 3712 3072 3944
rect 3404 3712 3420 3944
rect 3056 2713 3420 3712
rect 3056 2708 3650 2713
rect 3056 2216 3252 2708
rect 3640 2216 3650 2708
rect 3056 2212 3650 2216
rect 3242 2211 3650 2212
use outd_curm  outd_curm_0
timestamp 1683888831
transform 1 0 3040 0 1 24
box -40 916 1002 3158
use sky130_fd_pr__nfet_01v8_lvt_CP5GGS  sky130_fd_pr__nfet_01v8_lvt_CP5GGS_0
timestamp 1683810998
transform 1 0 3647 0 1 4299
box -647 -719 647 719
use sky130_fd_pr__nfet_01v8_lvt_L8NDKD#0  sky130_fd_pr__nfet_01v8_lvt_L8NDKD_0
timestamp 1683810998
transform 0 -1 4650 1 0 4576
box -996 -310 996 310
<< end >>
