magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< psubdiff >>
rect 1800 -9000 2200 -8976
rect 1800 -9424 2200 -9400
rect 3000 -9000 3400 -8976
rect 3000 -9424 3400 -9400
rect 4200 -9000 4600 -8976
rect 4200 -9424 4600 -9400
rect 5400 -9000 5800 -8976
rect 5400 -9424 5800 -9400
rect 6600 -9000 7000 -8976
rect 6600 -9424 7000 -9400
rect 7800 -9000 8200 -8976
rect 7800 -9424 8200 -9400
<< psubdiffcont >>
rect 1800 -9400 2200 -9000
rect 3000 -9400 3400 -9000
rect 4200 -9400 4600 -9000
rect 5400 -9400 5800 -9000
rect 6600 -9400 7000 -9000
rect 7800 -9400 8200 -9000
<< locali >>
rect 4554 2042 4556 2140
rect 4770 2042 4772 2140
rect 1736 1288 1872 1292
rect 1868 1204 1872 1288
rect 1736 1100 1872 1204
rect 4554 474 4772 2042
rect 1800 -9000 2200 -8984
rect 1800 -9416 2200 -9400
rect 3000 -9000 3400 -8984
rect 3000 -9416 3400 -9400
rect 4200 -9000 4600 -8984
rect 4200 -9416 4600 -9400
rect 5400 -9000 5800 -8984
rect 5400 -9416 5800 -9400
rect 6600 -9000 7000 -8984
rect 6600 -9416 7000 -9400
rect 7800 -9000 8200 -8984
rect 7800 -9416 8200 -9400
<< viali >>
rect 4556 2042 4770 2156
rect 1736 1204 1868 1288
rect 1800 -9400 2200 -9000
rect 3000 -9400 3400 -9000
rect 4200 -9400 4600 -9000
rect 5400 -9400 5800 -9000
rect 6600 -9400 7000 -9000
rect 7800 -9400 8200 -9000
<< metal1 >>
rect 5030 2260 5040 2700
rect 7220 2260 7230 2700
rect 4544 2156 4782 2162
rect 4544 2042 4556 2156
rect 4770 2042 4782 2156
rect 4544 2036 4782 2042
rect 916 1784 1152 1880
rect 1080 1324 1152 1784
rect 808 1168 1152 1324
rect 1080 704 1152 1168
rect 876 552 1152 704
rect 1080 84 1152 552
rect 812 -68 1152 84
rect 1080 -532 1152 -68
rect 864 -688 1152 -532
rect 1080 -1148 1152 -688
rect 816 -1304 1152 -1148
rect 1080 -1768 1152 -1304
rect 900 -1920 1152 -1768
rect 1080 -2384 1152 -1920
rect 852 -2540 1152 -2384
rect 1080 -3004 1152 -2540
rect 860 -3160 1152 -3004
rect 1080 -3620 1152 -3160
rect 844 -3716 1152 -3620
rect 1220 1080 1230 1880
rect 1724 1288 1880 1294
rect 1724 1204 1736 1288
rect 1868 1204 1880 1288
rect 1724 1198 1880 1204
rect 1220 976 1620 1080
rect 1220 496 1230 976
rect 3664 852 3768 1088
rect 4048 852 4058 1088
rect 5034 1024 5044 1460
rect 7216 1024 7226 1460
rect 1220 340 1736 496
rect 1220 -140 1230 340
rect 3648 308 3768 544
rect 4048 308 4058 544
rect 4628 56 4736 208
rect 1220 -244 1664 -140
rect 3648 -244 3768 -8
rect 4048 -244 4058 -8
rect 4490 -116 4500 56
rect 4724 -116 4736 56
rect 1220 -3716 1230 -244
rect 4628 -468 4736 -116
rect 4790 -304 4800 44
rect 4856 -304 4866 44
rect 1284 -620 1632 -532
rect 3188 -620 3232 -532
rect 1284 -1084 1432 -620
rect 4628 -672 4736 -616
rect 4486 -844 4496 -672
rect 4720 -844 4736 -672
rect 1284 -1240 1756 -1084
rect 1284 -1700 1432 -1240
rect 4628 -1288 4736 -844
rect 4790 -1072 4800 -816
rect 4860 -1072 4870 -816
rect 4628 -1496 4736 -1432
rect 4490 -1668 4500 -1496
rect 4724 -1668 4736 -1496
rect 1284 -1796 1796 -1700
rect 1284 -1916 1484 -1796
rect 1284 -2068 1440 -1916
rect 1704 -2068 1714 -1916
rect 1284 -2088 1712 -2068
rect 4628 -2108 4736 -1668
rect 4786 -1912 4796 -1656
rect 4856 -1912 4866 -1656
rect -2996 -3840 -2424 -3812
rect -2996 -4008 -2960 -3840
rect -2448 -4008 -2424 -3840
rect -2996 -4444 -2424 -4008
rect -432 -3992 1420 -3980
rect -432 -4444 1456 -3992
rect -3240 -4976 1456 -4444
rect -3240 -4980 1420 -4976
rect 1788 -9000 2212 -8994
rect 1788 -9400 1800 -9000
rect 2200 -9400 2212 -9000
rect 1788 -9406 2212 -9400
rect 2988 -9000 3412 -8994
rect 2988 -9400 3000 -9000
rect 3400 -9400 3412 -9000
rect 2988 -9406 3412 -9400
rect 4188 -9000 4612 -8994
rect 4188 -9400 4200 -9000
rect 4600 -9400 4612 -9000
rect 4188 -9406 4612 -9400
rect 5388 -9000 5812 -8994
rect 5388 -9400 5400 -9000
rect 5800 -9400 5812 -9000
rect 5388 -9406 5812 -9400
rect 6588 -9000 7012 -8994
rect 6588 -9400 6600 -9000
rect 7000 -9400 7012 -9000
rect 6588 -9406 7012 -9400
rect 7788 -9000 8212 -8994
rect 7788 -9400 7800 -9000
rect 8200 -9400 8212 -9000
rect 7788 -9406 8212 -9400
<< via1 >>
rect 5040 2260 7220 2700
rect 4556 2042 4770 2156
rect 1152 -3716 1220 1880
rect 1736 1204 1868 1288
rect 3768 852 4048 1088
rect 5044 1024 7216 1460
rect 3768 308 4048 544
rect 3768 -244 4048 -8
rect 4500 -116 4724 56
rect 4800 -304 4856 44
rect 4496 -844 4720 -672
rect 4800 -1072 4860 -816
rect 4500 -1668 4724 -1496
rect 1440 -2068 1704 -1916
rect 4796 -1912 4856 -1656
rect -2960 -4008 -2448 -3840
rect 1800 -9400 2200 -9000
rect 3000 -9400 3400 -9000
rect 4200 -9400 4600 -9000
rect 5400 -9400 5800 -9000
rect 6600 -9400 7000 -9000
rect 7800 -9400 8200 -9000
<< metal2 >>
rect 5040 2700 7220 2710
rect 5040 2250 7220 2260
rect 4556 2156 4770 2166
rect 4556 2032 4770 2042
rect 1152 1880 1220 1890
rect 1112 -3716 1152 1880
rect 1220 -2108 1396 1880
rect 5044 1460 7216 1470
rect 1736 1288 1868 1298
rect 1736 1194 1868 1204
rect 3768 1088 4048 1098
rect 1484 1016 2456 1026
rect 1484 762 2456 772
rect 4048 852 4272 1088
rect 5044 1014 7216 1024
rect 2576 692 3668 702
rect 2576 438 3668 448
rect 3768 544 4272 852
rect 1484 384 2456 394
rect 1484 130 2456 140
rect 4048 340 4272 544
rect 4048 308 7076 340
rect 3768 232 7076 308
rect 2576 64 3668 74
rect 2576 -190 3668 -180
rect 3768 -8 4272 232
rect 4924 230 5216 232
rect 6008 172 6932 182
rect 4048 -172 4272 -8
rect 4500 56 4724 66
rect 4500 -126 4724 -116
rect 4800 44 4856 54
rect 4048 -244 4800 -172
rect 3768 -304 4800 -244
rect 5036 -68 6008 160
rect 5036 -78 6932 -68
rect 5036 -88 6816 -78
rect 6984 -168 7076 232
rect 6984 -172 7364 -168
rect 4856 -304 7364 -172
rect 3768 -420 7364 -304
rect 2580 -568 3664 -558
rect 2580 -814 3664 -804
rect 1476 -888 2460 -878
rect 1476 -1138 2460 -1128
rect 3768 -992 4376 -420
rect 4932 -582 5224 -420
rect 5800 -582 6092 -420
rect 6736 -578 7364 -420
rect 6008 -648 6932 -638
rect 4496 -672 4720 -662
rect 4496 -854 4720 -844
rect 4800 -816 4860 -806
rect 3768 -1072 4800 -992
rect 5036 -888 6008 -660
rect 5036 -898 6932 -888
rect 5036 -908 6816 -898
rect 7000 -992 7364 -578
rect 4860 -1072 7364 -992
rect 2580 -1188 3664 -1178
rect 2580 -1434 3664 -1424
rect 3768 -1240 7364 -1072
rect 1476 -1508 2460 -1498
rect 1476 -1758 2460 -1748
rect 3768 -1812 4376 -1240
rect 4932 -1402 5224 -1240
rect 5800 -1402 6092 -1240
rect 6736 -1402 7364 -1240
rect 6008 -1476 6932 -1466
rect 4500 -1496 4724 -1486
rect 4500 -1678 4724 -1668
rect 4796 -1656 4856 -1646
rect 1440 -1916 1704 -1906
rect 3768 -1912 4796 -1812
rect 5036 -1716 6008 -1480
rect 5036 -1726 6932 -1716
rect 5036 -1728 6816 -1726
rect 7000 -1812 7364 -1402
rect 4856 -1912 7364 -1812
rect 3768 -2000 7364 -1912
rect 1440 -2078 1704 -2068
rect 1740 -2060 7364 -2000
rect 1740 -2108 4376 -2060
rect 1220 -2544 4376 -2108
rect 4932 -2214 5224 -2060
rect 5800 -2214 6092 -2060
rect 6736 -2218 7364 -2060
rect 1220 -3716 1396 -2544
rect 1652 -2792 1764 -2544
rect 1944 -2772 2056 -2544
rect 2296 -2772 2408 -2544
rect 2660 -2772 2772 -2544
rect 2952 -2768 3064 -2544
rect 2952 -2772 3020 -2768
rect 3216 -2772 3328 -2544
rect 3464 -2772 3580 -2544
rect 3824 -2748 3932 -2544
rect 4024 -2748 4116 -2544
rect 4216 -2744 4376 -2544
rect 3468 -2776 3580 -2772
rect 7000 -2780 7364 -2218
rect 1152 -3726 1220 -3716
rect -2960 -3840 -2448 -3830
rect -2960 -4018 -2448 -4008
rect 1800 -9000 2200 -8990
rect 1800 -9410 2200 -9400
rect 3000 -9000 3400 -8990
rect 3000 -9410 3400 -9400
rect 4200 -9000 4600 -8990
rect 4200 -9410 4600 -9400
rect 5400 -9000 5800 -8990
rect 5400 -9410 5800 -9400
rect 6600 -9000 7000 -8990
rect 6600 -9410 7000 -9400
rect 7800 -9000 8200 -8990
rect 7800 -9410 8200 -9400
<< via2 >>
rect 5040 2260 7220 2700
rect 4556 2042 4770 2156
rect 1736 1204 1868 1288
rect 1484 772 2456 1016
rect 5044 1024 7216 1460
rect 2576 448 3668 692
rect 1484 140 2456 384
rect 2576 -180 3668 64
rect 4500 -116 4724 56
rect 6008 -68 6932 172
rect 2580 -804 3664 -568
rect 1476 -1128 2460 -888
rect 4496 -844 4720 -672
rect 6008 -888 6932 -648
rect 2580 -1424 3664 -1188
rect 1476 -1748 2460 -1508
rect 4500 -1668 4724 -1496
rect 1440 -2068 1704 -1916
rect 6008 -1716 6932 -1476
rect -2960 -4008 -2448 -3840
rect 1800 -9400 2200 -9000
rect 3000 -9400 3400 -9000
rect 4200 -9400 4600 -9000
rect 5400 -9400 5800 -9000
rect 6600 -9400 7000 -9000
rect 7800 -9400 8200 -9000
<< metal3 >>
rect -4448 3240 -1560 3244
rect -4448 2700 7420 3240
rect -4448 2320 5040 2700
rect -4448 2280 -1780 2320
rect -4448 1932 -3320 2280
rect -1720 2260 5040 2320
rect 7220 2260 7420 2700
rect -1720 2156 7420 2260
rect -1720 2042 4556 2156
rect 4770 2042 7420 2156
rect -1720 2040 7420 2042
rect 1460 1300 2480 2040
rect 4546 2037 4780 2040
rect 5034 1460 7226 1465
rect 1472 1288 2472 1300
rect 1472 1204 1736 1288
rect 1868 1204 2472 1288
rect -910 280 -900 1160
rect -60 280 -50 1160
rect 1472 1016 2472 1204
rect 5034 1024 5044 1460
rect 7216 1024 7296 1460
rect 5034 1019 7296 1024
rect 1472 772 1484 1016
rect 2456 772 2472 1016
rect 1472 384 2472 772
rect 5996 736 7296 1019
rect 1472 140 1484 384
rect 2456 140 2472 384
rect 1472 128 2472 140
rect 2564 692 3684 708
rect 2564 448 2576 692
rect 3668 448 3684 692
rect 2564 64 3684 448
rect 2564 -180 2576 64
rect 3668 32 3684 64
rect 5992 172 7296 736
rect 4490 56 4734 61
rect 4490 32 4500 56
rect 3668 -116 4500 32
rect 4724 28 4734 56
rect 4724 -116 4860 28
rect 3668 -180 4860 -116
rect 2564 -468 4860 -180
rect 2564 -568 3684 -468
rect 2564 -804 2580 -568
rect 3664 -804 3684 -568
rect 1016 -888 2476 -872
rect 1016 -1128 1476 -888
rect 2460 -1128 2476 -888
rect 1016 -1508 2476 -1128
rect 2564 -1188 3684 -804
rect 2564 -1424 2580 -1188
rect 3664 -1424 3684 -1188
rect 2564 -1444 3684 -1424
rect 4432 -672 4860 -468
rect 4432 -844 4496 -672
rect 4720 -844 4860 -672
rect -922 -1960 10 -1580
rect 1016 -1748 1476 -1508
rect 2460 -1748 2476 -1508
rect 4432 -1496 4860 -844
rect 4432 -1668 4500 -1496
rect 4724 -1668 4860 -1496
rect 5992 -68 6008 172
rect 6932 -68 7296 172
rect 5992 -648 7296 -68
rect 5992 -888 6008 -648
rect 6932 -888 7296 -648
rect 5992 -1476 7296 -888
rect 4490 -1673 4734 -1668
rect 5992 -1716 6008 -1476
rect 6932 -1716 7296 -1476
rect 5992 -1732 7296 -1716
rect 1016 -1764 2476 -1748
rect 1430 -1916 1714 -1911
rect -922 -2312 -900 -1960
rect -910 -2840 -900 -2312
rect -60 -2312 10 -1960
rect 1188 -2068 1440 -1916
rect 1704 -2068 1714 -1916
rect 1188 -2073 1714 -2068
rect 1188 -2108 1704 -2073
rect -60 -2840 -50 -2312
rect -2996 -3840 -2424 -3812
rect -2996 -4008 -2960 -3840
rect -2448 -4008 -2424 -3840
rect -1760 -3920 -560 -3800
rect -2996 -4460 -2424 -4008
rect -900 -4120 -560 -3920
rect 1188 -3988 1472 -2108
rect 1016 -4256 1472 -3988
rect 1790 -9000 2210 -8995
rect 1790 -9400 1800 -9000
rect 2200 -9400 2210 -9000
rect 1790 -9405 2210 -9400
rect 2990 -9000 3410 -8995
rect 2990 -9400 3000 -9000
rect 3400 -9400 3410 -9000
rect 2990 -9405 3410 -9400
rect 4190 -9000 4610 -8995
rect 4190 -9400 4200 -9000
rect 4600 -9400 4610 -9000
rect 4190 -9405 4610 -9400
rect 5390 -9000 5810 -8995
rect 5390 -9400 5400 -9000
rect 5800 -9400 5810 -9000
rect 5390 -9405 5810 -9400
rect 6590 -9000 7010 -8995
rect 6590 -9400 6600 -9000
rect 7000 -9400 7010 -9000
rect 6590 -9405 7010 -9400
rect 7790 -9000 8210 -8995
rect 7790 -9400 7800 -9000
rect 8200 -9400 8210 -9000
rect 7790 -9405 8210 -9400
<< via3 >>
rect -900 280 -60 1160
rect -900 -2840 -60 -1960
rect 1800 -9400 2200 -9000
rect 3000 -9400 3400 -9000
rect 4200 -9400 4600 -9000
rect 5400 -9400 5800 -9000
rect 6600 -9400 7000 -9000
rect 7800 -9400 8200 -9000
<< metal4 >>
rect -1860 1160 20 1200
rect -1860 280 -900 1160
rect -60 280 20 1160
rect -1860 220 20 280
rect -1880 -1960 0 -1900
rect -1880 -2840 -900 -1960
rect -60 -2840 0 -1960
rect -1880 -2880 0 -2840
rect -3440 -4720 -2020 -2980
rect -3440 -4800 -240 -4720
rect -3460 -5800 -240 -4800
rect -3460 -7940 -3340 -5800
rect -3460 -8300 -300 -7940
rect -3460 -9000 8480 -8300
rect -3460 -9400 1800 -9000
rect 2200 -9400 3000 -9000
rect 3400 -9400 4200 -9000
rect 4600 -9400 5400 -9000
rect 5800 -9400 6600 -9000
rect 7000 -9400 7800 -9000
rect 8200 -9400 8480 -9000
rect -3460 -9640 8480 -9400
use sky130_fd_pr__cap_mim_m3_1_2YC3NK#0  sky130_fd_pr__cap_mim_m3_1_2YC3NK_0
timestamp 1686659968
transform -1 0 -2878 0 -1 -508
box -1686 -3040 1686 3040
use sky130_fd_pr__cap_mim_m3_1_6FAAF3  sky130_fd_pr__cap_mim_m3_1_6FAAF3_1
timestamp 1686659968
transform 0 -1 360 1 0 -6574
box -2686 -1040 2686 1040
use sky130_fd_pr__cap_mim_m3_1_N3CXMH  sky130_fd_pr__cap_mim_m3_1_N3CXMH_0
timestamp 1686659968
transform -1 0 -2854 0 -1 -6240
box -1686 -2040 1686 2040
use sky130_fd_pr__res_xhigh_po_1p41_HK6UT6  sky130_fd_pr__res_xhigh_po_1p41_HK6UT6_0
timestamp 1686659968
transform 1 0 6132 0 1 1858
box -1252 -998 1252 998
use tia_casc  tia_casc_0
timestamp 1686659968
transform 1 0 -5880 0 1 -280
box 4800 -3520 7054 2244
use tia_currm  tia_currm_0
timestamp 1686659968
transform 1 0 4026 0 1 -540
box -2646 -8320 4424 -2144
use tia_inv  tia_inv_0
timestamp 1686659968
transform 1 0 -940 0 1 -1120
box 2300 -760 4622 2274
use tia_m1  tia_m1_0
timestamp 1686659968
transform 1 0 3100 0 1 -160
box 1400 -2320 4260 740
<< labels >>
rlabel metal3 -4130 2670 -3760 3010 1 VP
port 1 n
<< end >>
