magic
tech sky130A
magscale 1 2
timestamp 1687207894
<< metal1 >>
rect 41190 39800 41200 42800
rect 44800 42400 110200 42800
rect 44800 39800 107600 42400
rect 110000 39800 110200 42400
rect 34800 33200 35000 37800
rect 36200 33200 41200 37800
rect 44800 33200 44810 37800
rect 107800 32600 110200 39800
rect 37590 29800 37600 32600
rect 40000 30000 46000 32600
rect 47600 30000 47610 32600
rect 40000 29800 40010 30000
rect 107800 28200 108000 32600
rect 110000 28200 110200 32600
rect 86800 19200 90600 19600
rect 86590 17800 86600 19000
rect 87000 17800 88200 19000
rect 102390 18200 102400 19200
rect 103000 18200 104600 19200
rect 36590 10200 36600 13400
rect 40200 10200 46000 13400
rect 49600 10200 49610 13400
rect 87200 12600 88200 17800
rect 62000 11400 88200 12600
rect 62000 -1000 63000 11400
rect 49600 -1600 63000 -1000
rect 77700 9300 87400 10700
rect 88800 9300 88810 10700
rect 103200 9800 104600 18200
rect 45590 -2200 45600 -2000
rect 36590 -5000 36600 -2200
rect 40200 -5000 45600 -2200
rect 48200 -5000 48210 -2000
rect 49600 -6600 50200 -1600
rect 77700 -2300 78900 9300
rect 103200 8200 108000 9800
rect 49590 -6800 49600 -6600
rect 50200 -6800 50210 -6600
rect 78400 -8200 78900 -2300
rect 78990 -6400 79000 -6000
rect 79200 -6400 79210 -6000
rect 78400 -8600 78700 -8200
rect 79000 -8600 79010 -8200
rect 106600 -18400 108000 8200
rect 105800 -19700 108000 -18400
rect 36590 -24400 36600 -21200
rect 40200 -24400 45600 -21200
rect 48400 -24400 48410 -21200
rect 105800 -26600 107200 -19700
rect 62100 -27600 107200 -26600
rect 62100 -37100 62900 -27600
rect 50200 -37800 62900 -37100
rect 78000 -35300 107000 -35200
rect 78000 -36900 105900 -35300
rect 107100 -36900 107110 -35300
rect 78000 -37000 107000 -36900
rect 78000 -37800 78800 -37000
rect 36590 -40600 36600 -38000
rect 40200 -40600 45400 -38000
rect 49500 -40600 49510 -38000
rect 50200 -42200 50900 -37800
rect 49500 -42500 50900 -42200
rect 49490 -42800 49500 -42500
rect 49900 -42700 50900 -42500
rect 49900 -42800 49910 -42700
rect 78400 -43200 78800 -37800
rect 79390 -38800 79400 -37400
rect 82600 -38800 82610 -37400
rect 78990 -42500 79000 -42100
rect 79200 -42500 79210 -42100
rect 78400 -43600 79000 -43200
rect 78600 -43800 79000 -43600
rect 78590 -44400 78600 -43800
rect 79000 -44400 79010 -43800
<< via1 >>
rect 41200 39800 44800 42800
rect 107600 39800 110000 42400
rect 35000 33200 36200 37800
rect 41200 33200 44800 37800
rect 37600 29800 40000 32600
rect 46000 30000 47600 32600
rect 108000 28200 110000 32600
rect 86600 17800 87000 19000
rect 102400 18200 103000 19200
rect 36600 10200 40200 13400
rect 46000 10200 49600 13400
rect 87400 9300 88800 10700
rect 36600 -5000 40200 -2200
rect 45600 -5000 48200 -2000
rect 49600 -6800 50200 -6600
rect 79000 -6400 79200 -6000
rect 78700 -8600 79000 -8200
rect 36600 -24400 40200 -21200
rect 45600 -24400 48400 -21200
rect 105900 -36900 107100 -35300
rect 36600 -40600 40200 -38000
rect 45400 -40600 49500 -38000
rect 49500 -42800 49900 -42500
rect 79400 -38800 82600 -37400
rect 79000 -42500 79200 -42100
rect 78600 -44400 79000 -43800
<< metal2 >>
rect 41200 42800 44800 42810
rect 44800 42400 110200 42800
rect 44800 39800 107600 42400
rect 110000 39800 110200 42400
rect 41200 39790 44800 39800
rect 107600 39790 110200 39800
rect 35000 37800 36200 37810
rect 41200 37800 44800 37810
rect 34800 33200 35000 37800
rect 36200 33200 41200 37800
rect 35000 33190 36200 33200
rect 41200 33190 44800 33200
rect 37600 32600 40000 32610
rect 46000 32600 47600 32610
rect 40000 30000 46000 32600
rect 46000 29990 47600 30000
rect 107800 32600 110200 39790
rect 37600 29790 40000 29800
rect 107800 28200 108000 32600
rect 110000 28200 110200 32600
rect 108000 28190 110000 28200
rect 87400 23800 88800 23810
rect 86600 19000 87000 19010
rect 86600 17790 87000 17800
rect 36600 13400 40200 13410
rect 46000 13400 49600 13410
rect 40200 10200 46000 13400
rect 36600 10190 40200 10200
rect 46000 10190 49600 10200
rect 87400 10700 88800 22400
rect 102600 23400 103200 23410
rect 103200 22400 104600 23400
rect 102600 22390 104600 22400
rect 102400 19200 103000 19210
rect 102400 18190 103000 18200
rect 87400 9290 88800 9300
rect 103200 9800 104600 22390
rect 34200 9000 35800 9010
rect 50600 8800 52000 8810
rect 35800 7400 50600 8800
rect 103200 8200 108000 9800
rect 34200 7390 35800 7400
rect 50600 7390 52000 7400
rect 34200 6200 35800 6210
rect 35800 4600 47000 6000
rect 34200 4590 35800 4600
rect 45600 2800 47000 4600
rect 51000 2800 52400 2810
rect 45600 1400 51000 2800
rect 51000 1390 52400 1400
rect 43000 600 44600 610
rect 54600 600 56200 610
rect 44600 -600 54600 600
rect 43000 -610 44600 -600
rect 54600 -610 56200 -600
rect 45600 -2000 48200 -1990
rect 36600 -2200 40200 -2190
rect 40200 -5000 45600 -2200
rect 48200 -4600 53200 -2000
rect 36600 -5010 40200 -5000
rect 45600 -5010 48200 -5000
rect 59800 -5600 60600 -5590
rect 59800 -6410 60600 -6400
rect 73200 -5600 74000 -5590
rect 73200 -6410 74000 -6400
rect 79000 -6000 79200 -5990
rect 79000 -6410 79200 -6400
rect 49600 -6600 50200 -6590
rect 49600 -6810 50200 -6800
rect 78700 -8200 79000 -8190
rect 78700 -8610 79000 -8600
rect 106600 -18400 108000 8200
rect 105800 -19700 108000 -18400
rect 36600 -21200 40200 -21190
rect 45600 -21200 48400 -21190
rect 40200 -24400 45600 -21200
rect 36600 -24410 40200 -24400
rect 45600 -24410 48400 -24400
rect 34700 -26800 35900 -26790
rect 45800 -26800 47000 -26790
rect 35900 -28200 45800 -26800
rect 47000 -28200 47200 -26800
rect 34700 -28210 35900 -28200
rect 45800 -28210 47000 -28200
rect 34200 -31800 35800 -31790
rect 45400 -31800 47200 -31790
rect 35800 -34000 45400 -31800
rect 34200 -34010 35800 -34000
rect 45400 -34010 47200 -34000
rect 42400 -34500 44800 -34490
rect 54800 -34500 56600 -34490
rect 44800 -36300 54800 -34500
rect 42400 -36310 44800 -36300
rect 54800 -36310 56600 -36300
rect 105800 -35300 107200 -19700
rect 105800 -36900 105900 -35300
rect 107100 -36900 107200 -35300
rect 105800 -37000 107200 -36900
rect 79400 -37400 82600 -37390
rect 36600 -38000 40200 -37990
rect 45400 -38000 49500 -37990
rect 40200 -40600 45400 -38000
rect 49500 -40600 53100 -38000
rect 79400 -38810 82600 -38800
rect 36600 -40610 40200 -40600
rect 45400 -40610 49500 -40600
rect 59800 -41600 60200 -41590
rect 59800 -42410 60200 -42400
rect 73300 -41600 73700 -41590
rect 73300 -42410 73700 -42400
rect 79000 -42100 79200 -42090
rect 49500 -42500 49900 -42490
rect 79000 -42510 79200 -42500
rect 49500 -42810 49900 -42800
rect 78600 -43800 79000 -43790
rect 78600 -44410 79000 -44400
<< via2 >>
rect 41200 39800 44800 42800
rect 107600 39800 110000 42400
rect 35000 33200 36200 37800
rect 41200 33200 44800 37800
rect 37600 29800 40000 32600
rect 46000 30000 47600 32600
rect 108000 28200 110000 32600
rect 87400 22400 88800 23800
rect 86600 17800 87000 19000
rect 36600 10200 40200 13400
rect 46000 10200 49600 13400
rect 102600 22400 103200 23400
rect 102400 18200 103000 19200
rect 34200 7400 35800 9000
rect 50600 7400 52000 8800
rect 34200 4600 35800 6200
rect 51000 1400 52400 2800
rect 43000 -600 44600 600
rect 54600 -600 56200 600
rect 36600 -5000 40200 -2200
rect 45600 -5000 48200 -2000
rect 59800 -6400 60600 -5600
rect 73200 -6400 74000 -5600
rect 79000 -6400 79200 -6000
rect 78700 -8600 79000 -8200
rect 36600 -24400 40200 -21200
rect 45600 -24400 48400 -21200
rect 34700 -28200 35900 -26800
rect 45800 -28200 47000 -26800
rect 34200 -34000 35800 -31800
rect 45400 -34000 47200 -31800
rect 42400 -36300 44800 -34500
rect 54800 -36300 56600 -34500
rect 36600 -40600 40200 -38000
rect 45400 -40600 49500 -38000
rect 79400 -38800 82600 -37400
rect 59800 -42400 60200 -41600
rect 73300 -42400 73700 -41600
rect 79000 -42500 79200 -42100
rect 78600 -44400 79000 -43800
<< metal3 >>
rect 33780 42800 35140 42940
rect 41190 42800 44810 42805
rect 33780 38400 36600 42800
rect 40200 38400 40210 42800
rect 41190 39800 41200 42800
rect 44800 42400 112200 42800
rect 44800 39800 107600 42400
rect 110000 39800 112200 42400
rect 41190 39795 44810 39800
rect 107590 39795 112200 39800
rect 33780 38140 35140 38400
rect 34080 37805 35100 37840
rect 34080 37800 36210 37805
rect 34080 33200 35000 37800
rect 36200 33200 36210 37800
rect 34990 33195 36210 33200
rect 33800 32800 35160 32900
rect 36600 32800 40200 38400
rect 41200 37805 44800 39795
rect 108800 38200 112200 39795
rect 41190 37800 44810 37805
rect 41190 33200 41200 37800
rect 44800 33200 44810 37800
rect 104590 33200 104600 37800
rect 107400 33200 111800 37800
rect 41190 33195 44810 33200
rect 33800 32600 40200 32800
rect 33800 28200 36600 32600
rect 40200 28200 40210 32600
rect 33800 28100 35160 28200
rect 33800 16960 35800 17000
rect 33600 11940 35800 16960
rect 36600 13405 40200 28200
rect 41200 17000 44800 33195
rect 45990 32600 47610 32605
rect 45990 30000 46000 32600
rect 47600 30000 47610 32600
rect 45990 29995 47610 30000
rect 87390 23800 88810 23805
rect 87390 22400 87400 23800
rect 88800 22400 88810 23800
rect 87390 22395 88810 22400
rect 102590 23400 103210 23405
rect 102590 22400 102600 23400
rect 103200 22400 103210 23400
rect 102590 22395 103210 22400
rect 102390 19200 103010 19205
rect 86590 19000 87010 19005
rect 73000 18200 74200 18600
rect 73000 17400 73400 18200
rect 86590 17800 86600 19000
rect 87000 17800 87010 19000
rect 102390 18200 102400 19200
rect 103000 18200 103010 19200
rect 102390 18195 103010 18200
rect 64200 17000 73400 17400
rect 74190 17000 74200 17800
rect 75400 17000 75410 17800
rect 86590 17795 87010 17800
rect 89990 17000 90000 17800
rect 91200 17000 91210 17800
rect 41200 14000 49400 17000
rect 50400 14000 50410 17000
rect 34200 9005 35800 11940
rect 36590 13400 40210 13405
rect 36590 10200 36600 13400
rect 40200 10200 40210 13400
rect 36590 10195 40210 10200
rect 34190 9000 35810 9005
rect 34190 7400 34200 9000
rect 35800 7400 35810 9000
rect 34190 7395 35810 7400
rect 34190 6200 35810 6205
rect 34190 4600 34200 6200
rect 35800 4600 35810 6200
rect 34190 4595 35810 4600
rect 34200 -4000 35800 4595
rect 36600 -2195 40200 10195
rect 41200 600 44800 14000
rect 45990 13400 49610 13405
rect 74200 13400 75400 17000
rect 90000 13400 91200 17000
rect 104600 13400 107400 33200
rect 110520 32800 112240 32820
rect 107800 32600 112240 32800
rect 107800 28200 108000 32600
rect 110000 28200 112240 32600
rect 107990 28195 110010 28200
rect 110520 28100 112240 28200
rect 111720 15800 112380 17100
rect 109990 13800 110000 15800
rect 111400 13800 112380 15800
rect 45990 10200 46000 13400
rect 49600 11200 107400 13400
rect 111720 12100 112380 13800
rect 49600 10200 59400 11200
rect 79000 11000 107400 11200
rect 45990 10195 49610 10200
rect 50590 8800 52010 8805
rect 50590 7400 50600 8800
rect 52000 7400 52010 8800
rect 50590 7395 52010 7400
rect 50990 2800 52410 2805
rect 50990 1400 51000 2800
rect 52400 1400 52410 2800
rect 50990 1395 52410 1400
rect 79000 800 82200 11000
rect 41200 -600 43000 600
rect 44600 -600 44800 600
rect 34000 -4020 35800 -4000
rect 33580 -9000 35800 -4020
rect 36590 -2200 40210 -2195
rect 36590 -5000 36600 -2200
rect 40200 -5000 40210 -2200
rect 36590 -5005 40210 -5000
rect 33580 -9040 34260 -9000
rect 36600 -21195 40200 -5005
rect 41200 -15200 44800 -600
rect 54590 600 56210 605
rect 54590 -600 54600 600
rect 56200 -600 56210 600
rect 79000 -600 106200 800
rect 54590 -605 56210 -600
rect 45590 -2000 48210 -1995
rect 78990 -2000 79000 -600
rect 106200 -2000 106210 -600
rect 45590 -5000 45600 -2000
rect 48200 -4600 53200 -2000
rect 58190 -3800 58200 -2000
rect 59200 -3800 59210 -2000
rect 79000 -2200 106200 -2000
rect 48200 -5000 48210 -4600
rect 45590 -5005 48210 -5000
rect 59790 -5600 60610 -5595
rect 59790 -6400 59800 -5600
rect 60600 -6400 60610 -5600
rect 59790 -6405 60610 -6400
rect 73190 -5600 74010 -5595
rect 73190 -6400 73200 -5600
rect 74000 -6400 74010 -5600
rect 77000 -5995 79000 -5800
rect 77000 -6000 79210 -5995
rect 77000 -6200 79000 -6000
rect 78800 -6400 79000 -6200
rect 79200 -6400 79210 -6000
rect 73190 -6405 74010 -6400
rect 78990 -6405 79210 -6400
rect 111640 -7100 112300 -3860
rect 78690 -8200 79010 -8195
rect 77990 -8400 78000 -8200
rect 78200 -8400 78210 -8200
rect 78690 -8600 78700 -8200
rect 79000 -8600 79010 -8200
rect 109990 -8600 110000 -7100
rect 111100 -8600 112300 -7100
rect 78690 -8605 79010 -8600
rect 111640 -8860 112300 -8600
rect 80790 -10000 80800 -9700
rect 81400 -10000 81410 -9700
rect 41200 -19000 50400 -15200
rect 76800 -19000 83200 -15600
rect 36590 -21200 40210 -21195
rect 36590 -24400 36600 -21200
rect 40200 -24400 40210 -21200
rect 36590 -24405 40210 -24400
rect 33620 -25700 34300 -25020
rect 33620 -26795 35900 -25700
rect 33620 -26800 35910 -26795
rect 33620 -28200 34700 -26800
rect 35900 -28200 35910 -26800
rect 33620 -28205 35910 -28200
rect 33620 -29200 35900 -28205
rect 33620 -30040 34300 -29200
rect 34190 -31800 35810 -31795
rect 34190 -34000 34200 -31800
rect 35800 -34000 35810 -31800
rect 34190 -34005 35810 -34000
rect 34200 -46000 35800 -34005
rect 36600 -37995 40200 -24405
rect 41200 -34495 44800 -19000
rect 45590 -21200 48410 -21195
rect 45590 -24400 45600 -21200
rect 48400 -23200 82600 -21200
rect 48400 -24300 54700 -23200
rect 56600 -24300 82600 -23200
rect 48400 -24400 82600 -24300
rect 45590 -24405 48410 -24400
rect 50590 -26500 50600 -26400
rect 45800 -26795 50600 -26500
rect 45790 -26800 50600 -26795
rect 45790 -28200 45800 -26800
rect 47000 -28200 50600 -26800
rect 45790 -28205 47010 -28200
rect 50590 -28400 50600 -28200
rect 52600 -28400 52610 -26400
rect 54700 -27900 56600 -24400
rect 79200 -27500 105000 -24400
rect 45390 -31800 47210 -31795
rect 45390 -34000 45400 -31800
rect 47200 -34000 47400 -31800
rect 45390 -34005 47400 -34000
rect 41200 -34500 44810 -34495
rect 41200 -36300 42400 -34500
rect 44800 -36300 44810 -34500
rect 45400 -34700 47400 -34005
rect 50590 -34700 50600 -34400
rect 45400 -36200 50600 -34700
rect 50590 -36300 50600 -36200
rect 52600 -36300 52610 -34400
rect 54790 -34500 56610 -34495
rect 54790 -36300 54800 -34500
rect 56600 -36300 56610 -34500
rect 41200 -36305 44810 -36300
rect 54790 -36305 56610 -36300
rect 36590 -38000 40210 -37995
rect 36590 -40600 36600 -38000
rect 40200 -40600 40210 -38000
rect 36590 -40605 40210 -40600
rect 33900 -46040 34200 -46000
rect 33600 -47800 34200 -46040
rect 35800 -47800 35810 -46000
rect 33600 -51060 35500 -47800
rect 33900 -51100 35500 -51060
rect 36600 -62200 40200 -40605
rect 41200 -51200 44800 -36305
rect 79300 -37395 82600 -27500
rect 79300 -37400 82610 -37395
rect 45390 -38000 49510 -37995
rect 45390 -40600 45400 -38000
rect 49500 -38100 58310 -38000
rect 49500 -39000 57600 -38100
rect 58600 -39000 58610 -38100
rect 79300 -38300 79400 -37400
rect 79390 -38800 79400 -38300
rect 82600 -38800 82610 -37400
rect 101800 -38000 105000 -27500
rect 111700 -27800 112360 -24940
rect 107990 -29800 108000 -27800
rect 110200 -29800 112360 -27800
rect 111700 -29940 112360 -29800
rect 79390 -38805 82610 -38800
rect 49500 -39600 58310 -39000
rect 101790 -39400 101800 -38000
rect 105000 -38400 105010 -38000
rect 105000 -38800 105100 -38400
rect 105000 -39400 105010 -38800
rect 49500 -40600 58300 -39600
rect 45390 -40605 49510 -40600
rect 59790 -41600 60210 -41595
rect 59790 -42400 59800 -41600
rect 60200 -42400 60210 -41600
rect 59790 -42405 60210 -42400
rect 73290 -41600 73710 -41595
rect 73290 -42400 73300 -41600
rect 73700 -42400 73710 -41600
rect 76900 -42095 79100 -41900
rect 76900 -42100 79210 -42095
rect 76900 -42300 79000 -42100
rect 73290 -42405 73710 -42400
rect 78900 -42500 79000 -42300
rect 79200 -42500 79210 -42100
rect 78990 -42505 79210 -42500
rect 78590 -43000 78600 -42800
rect 78800 -43000 78810 -42800
rect 78600 -43400 78800 -43000
rect 78200 -43600 78800 -43400
rect 78200 -44000 78400 -43600
rect 78000 -44600 78400 -44000
rect 78590 -43800 79010 -43795
rect 78590 -44400 78600 -43800
rect 79000 -44400 79010 -43800
rect 78590 -44405 79010 -44400
rect 80790 -46000 80800 -45800
rect 81400 -46000 81410 -45800
rect 111720 -46200 112380 -45940
rect 107990 -49000 108000 -46200
rect 110200 -49000 112380 -46200
rect 111720 -50940 112380 -49000
rect 50100 -51200 50300 -51100
rect 41200 -51400 50300 -51200
rect 41200 -55000 50200 -51400
rect 76000 -54900 83300 -51700
rect 41200 -62200 44800 -55000
<< via3 >>
rect 36600 38400 40200 42800
rect 41200 39800 44800 42800
rect 107600 39800 110000 42400
rect 41200 33200 44800 37800
rect 104600 33200 107400 37800
rect 36600 29800 37600 32600
rect 37600 29800 40000 32600
rect 40000 29800 40200 32600
rect 36600 28200 40200 29800
rect 46000 30000 47600 32600
rect 87400 22400 88800 23800
rect 102600 22400 103200 23400
rect 86600 17800 87000 19000
rect 102400 18200 103000 19200
rect 74200 17000 75400 17800
rect 90000 17000 91200 17800
rect 49400 14000 50400 17000
rect 36600 10200 40200 13400
rect 108000 28400 110000 32600
rect 110000 13800 111400 15800
rect 46000 10200 49600 13400
rect 50600 7400 52000 8800
rect 51000 1400 52400 2800
rect 43000 -600 44600 600
rect 36600 -5000 40200 -2200
rect 54600 -600 56200 600
rect 79000 -2000 106200 -600
rect 45600 -3800 48200 -2000
rect 58200 -3800 59200 -2000
rect 59800 -6400 60600 -5600
rect 73200 -6400 74000 -5600
rect 78000 -8400 78200 -8200
rect 78700 -8600 79000 -8200
rect 110000 -8600 111100 -7100
rect 80800 -10000 81400 -9700
rect 36600 -24400 40200 -21200
rect 34200 -34000 35800 -31800
rect 45600 -24400 48400 -21200
rect 54700 -24300 56600 -23200
rect 50600 -28400 52600 -26400
rect 42400 -36300 44800 -34500
rect 50600 -36300 52600 -34400
rect 54800 -36300 56600 -34500
rect 36600 -40600 40200 -38000
rect 34200 -47800 35800 -46000
rect 45400 -40600 49500 -38000
rect 57600 -39000 58600 -38100
rect 79400 -38800 82600 -37400
rect 108000 -29800 110200 -27800
rect 101800 -39400 105000 -38000
rect 59800 -42400 60200 -41600
rect 73300 -42400 73700 -41600
rect 78600 -43000 78800 -42800
rect 78600 -44400 79000 -43800
rect 80800 -46000 81400 -45800
rect 108000 -49000 110200 -46200
<< metal4 >>
rect 36599 42800 40201 42801
rect 36599 38400 36600 42800
rect 40200 38400 40201 42800
rect 41199 42800 44801 42801
rect 41199 39800 41200 42800
rect 44800 42400 110200 42800
rect 44800 39800 107600 42400
rect 110000 39800 110200 42400
rect 41199 39799 44801 39800
rect 107599 39799 110200 39800
rect 36599 38399 40201 38400
rect 36600 32601 40200 38399
rect 41200 37801 44800 39799
rect 41199 37800 44801 37801
rect 41199 33200 41200 37800
rect 44800 33200 44801 37800
rect 104599 37800 107401 37801
rect 41199 33199 44801 33200
rect 45800 35400 55400 37400
rect 36599 32600 40201 32601
rect 36599 28200 36600 32600
rect 40200 28200 40201 32600
rect 36599 28199 40201 28200
rect 36600 13401 40200 28199
rect 41200 17000 44800 33199
rect 45800 32600 48000 35400
rect 104599 33200 104600 37800
rect 107400 33200 107401 37800
rect 104599 33199 107401 33200
rect 45800 30000 46000 32600
rect 47600 30000 48000 32600
rect 45999 29999 47601 30000
rect 87399 23800 88801 23801
rect 86800 22400 87400 23800
rect 88800 22400 88801 23800
rect 87399 22399 88801 22400
rect 102599 23400 103201 23401
rect 102599 22400 102600 23400
rect 103200 22400 103201 23400
rect 102599 22399 103201 22400
rect 102399 19200 103001 19201
rect 86599 19000 87001 19001
rect 74199 17800 75401 17801
rect 49399 17000 50401 17001
rect 41200 14000 49400 17000
rect 50400 14000 50401 17000
rect 74199 17000 74200 17800
rect 75400 17000 75401 17800
rect 86599 17800 86600 19000
rect 87000 17800 87001 19000
rect 102399 18200 102400 19200
rect 103000 18200 103001 19200
rect 102399 18199 103001 18200
rect 86599 17799 87001 17800
rect 89999 17800 91201 17801
rect 74199 16999 75401 17000
rect 89999 17000 90000 17800
rect 91200 17000 91201 17800
rect 89999 16999 91201 17000
rect 36599 13400 40201 13401
rect 36599 10200 36600 13400
rect 40200 10200 40201 13400
rect 36599 10199 40201 10200
rect 36600 -2199 40200 10199
rect 41200 600 44800 14000
rect 49399 13999 50401 14000
rect 45999 13400 49601 13401
rect 74200 13400 75400 16999
rect 90000 13400 91200 16999
rect 104600 13400 107400 33199
rect 107800 32600 110200 39799
rect 107800 28400 108000 32600
rect 110000 28400 110200 32600
rect 107999 28399 110001 28400
rect 109999 15800 111401 15801
rect 45999 10200 46000 13400
rect 49600 11200 107400 13400
rect 49600 10200 59400 11200
rect 79000 11000 107400 11200
rect 108200 13800 110000 15800
rect 111400 13800 111401 15800
rect 108200 13799 111401 13800
rect 45999 10199 49601 10200
rect 50599 8800 52001 8801
rect 50599 7400 50600 8800
rect 52000 7400 52001 8800
rect 54600 8400 56600 10200
rect 59800 9800 74200 10800
rect 50599 7399 52001 7400
rect 59800 5200 61200 9800
rect 49200 3600 54400 4600
rect 50999 2800 52401 2801
rect 50999 1400 51000 2800
rect 52400 1400 52401 2800
rect 53400 2800 54400 3600
rect 59200 3200 61200 5200
rect 53400 1800 60800 2800
rect 50999 1399 52401 1400
rect 51000 800 52400 1399
rect 41200 -600 43000 600
rect 44600 -600 44800 600
rect 36599 -2200 40201 -2199
rect 36599 -5000 36600 -2200
rect 40200 -5000 40201 -2200
rect 36599 -5001 40201 -5000
rect 36600 -21199 40200 -5001
rect 41200 -15200 44800 -600
rect 54599 600 56201 601
rect 54599 -600 54600 600
rect 56200 -600 56201 600
rect 54599 -601 56201 -600
rect 45599 -2000 48201 -1999
rect 58199 -2000 59201 -1999
rect 45599 -3800 45600 -2000
rect 48200 -3800 58200 -2000
rect 59200 -3800 59201 -2000
rect 45599 -3801 48201 -3800
rect 58199 -3801 59201 -3800
rect 59800 -5599 60800 1800
rect 73200 -5599 74200 9800
rect 79000 800 82200 11000
rect 79000 -599 106200 800
rect 78999 -600 106201 -599
rect 78999 -2000 79000 -600
rect 106200 -2000 106201 -600
rect 78999 -2001 106201 -2000
rect 79000 -2200 106200 -2001
rect 59799 -5600 60800 -5599
rect 59799 -6400 59800 -5600
rect 60600 -6400 60800 -5600
rect 59799 -6401 60800 -6400
rect 73199 -5600 74200 -5599
rect 108200 -5600 110000 13799
rect 73199 -6400 73200 -5600
rect 74000 -6400 74200 -5600
rect 73199 -6401 74001 -6400
rect 59800 -6600 60800 -6401
rect 106400 -6600 110000 -5600
rect 77200 -7100 77900 -6800
rect 78400 -7000 82600 -6800
rect 77999 -8200 78201 -8199
rect 78400 -8200 78600 -7000
rect 109999 -7100 111101 -7099
rect 77999 -8400 78000 -8200
rect 78200 -8400 78600 -8200
rect 78699 -8200 79001 -8199
rect 77999 -8401 78201 -8400
rect 78699 -8600 78700 -8200
rect 79000 -8600 81200 -8200
rect 106400 -8600 110000 -7100
rect 111100 -8600 111101 -7100
rect 78699 -8601 79001 -8600
rect 80800 -9699 81200 -8600
rect 109999 -8601 111101 -8600
rect 80799 -9700 81401 -9699
rect 80799 -10000 80800 -9700
rect 81400 -10000 81401 -9700
rect 80799 -10001 81401 -10000
rect 41200 -19000 50400 -15200
rect 76800 -19000 83200 -15600
rect 36599 -21200 40201 -21199
rect 36599 -24400 36600 -21200
rect 40200 -24400 40201 -21200
rect 36599 -24401 40201 -24400
rect 34199 -31800 35801 -31799
rect 34199 -34000 34200 -31800
rect 35800 -34000 35801 -31800
rect 34199 -34001 35801 -34000
rect 34200 -45999 35800 -34001
rect 36600 -37999 40200 -24401
rect 41200 -34499 44800 -19000
rect 45599 -21200 48401 -21199
rect 45599 -24400 45600 -21200
rect 48400 -23200 82600 -21200
rect 48400 -24300 54700 -23200
rect 56600 -24300 82600 -23200
rect 48400 -24400 82600 -24300
rect 45599 -24401 48401 -24400
rect 50599 -26400 52601 -26399
rect 50599 -28400 50600 -26400
rect 52600 -28400 52601 -26400
rect 54700 -27900 56600 -24400
rect 59800 -26400 74200 -25200
rect 50599 -28401 52601 -28400
rect 59800 -30400 61000 -26400
rect 49700 -32300 51700 -31400
rect 50700 -33000 51700 -32300
rect 58400 -32400 61000 -30400
rect 50700 -33900 60800 -33000
rect 50599 -34400 52601 -34399
rect 41200 -34500 44801 -34499
rect 41200 -36300 42400 -34500
rect 44800 -36300 44801 -34500
rect 41200 -36301 44801 -36300
rect 50599 -36300 50600 -34400
rect 52600 -36300 52601 -34400
rect 50599 -36301 52601 -36300
rect 54799 -34500 56601 -34499
rect 54799 -36300 54800 -34500
rect 56600 -36300 56601 -34500
rect 54799 -36301 56601 -36300
rect 36599 -38000 40201 -37999
rect 36599 -40600 36600 -38000
rect 40200 -40600 40201 -38000
rect 36599 -40601 40201 -40600
rect 34199 -46000 35801 -45999
rect 34199 -47800 34200 -46000
rect 35800 -47800 35801 -46000
rect 34199 -47801 35801 -47800
rect 36600 -62200 40200 -40601
rect 41200 -51200 44800 -36301
rect 45399 -38000 49501 -37999
rect 45399 -40600 45400 -38000
rect 49500 -38099 58600 -38000
rect 49500 -38100 58601 -38099
rect 49500 -39000 57600 -38100
rect 58600 -39000 58601 -38100
rect 49500 -39001 58601 -39000
rect 49500 -39600 58600 -39001
rect 49500 -40600 49501 -39600
rect 45399 -40601 49501 -40600
rect 59700 -41600 60800 -33900
rect 59700 -42300 59800 -41600
rect 59799 -42400 59800 -42300
rect 60200 -42300 60800 -41600
rect 73200 -41600 74200 -26400
rect 79200 -27500 105000 -24400
rect 79300 -37399 82600 -27500
rect 79300 -37400 82601 -37399
rect 79300 -38300 79400 -37400
rect 79399 -38800 79400 -38300
rect 82600 -38800 82601 -37400
rect 101800 -37999 105000 -27500
rect 107999 -27800 110201 -27799
rect 107999 -29800 108000 -27800
rect 110200 -29800 110201 -27800
rect 107999 -29801 110201 -29800
rect 79399 -38801 82601 -38800
rect 101799 -38000 105001 -37999
rect 101799 -39400 101800 -38000
rect 105000 -38400 105001 -38000
rect 105000 -38800 105100 -38400
rect 105000 -39400 105001 -38800
rect 101799 -39401 105001 -39400
rect 108000 -41600 110200 -29801
rect 60200 -42400 60201 -42300
rect 73200 -42400 73300 -41600
rect 73700 -42400 74200 -41600
rect 59799 -42401 60201 -42400
rect 73299 -42401 73701 -42400
rect 106400 -42600 110200 -41600
rect 78599 -42800 78801 -42799
rect 77300 -43100 77900 -42800
rect 78599 -43000 78600 -42800
rect 78800 -43000 82600 -42800
rect 78599 -43001 78801 -43000
rect 78599 -43800 79001 -43799
rect 78599 -44400 78600 -43800
rect 79000 -44400 81400 -43800
rect 106400 -44200 110200 -43000
rect 78599 -44401 79001 -44400
rect 80800 -45799 81400 -44400
rect 80799 -45800 81401 -45799
rect 80799 -46000 80800 -45800
rect 81400 -46000 81401 -45800
rect 80799 -46001 81401 -46000
rect 108000 -46199 110200 -44200
rect 107999 -46200 110201 -46199
rect 107999 -49000 108000 -46200
rect 110200 -49000 110201 -46200
rect 107999 -49001 110201 -49000
rect 41200 -55000 50200 -51200
rect 76000 -54900 83300 -51700
rect 41200 -62200 44800 -55000
<< metal5 >>
rect 50600 6800 52600 7200
rect 50600 5600 56200 6800
rect 49800 3200 50400 5200
rect 51000 1200 52600 5200
rect 55200 3200 56200 5600
rect 56800 3200 57400 5200
rect 50900 -28900 52600 -28100
rect 50900 -29900 56600 -28900
rect 49800 -32400 50000 -30400
rect 50600 -32400 52600 -30400
rect 55700 -32400 56600 -29900
rect 57200 -32400 57400 -30400
rect 50800 -34700 52600 -32400
rect 50400 3200 51000 5200
rect 56200 3200 56800 5200
rect 50000 -32400 50600 -30400
rect 56600 -32400 57200 -30400
use bias2_top  bias2_top_0 ~/code/hibpm-sky130a-tapeout/mag/bias
timestamp 1686510802
transform 1 0 74160 0 1 18200
box -160 -4200 12860 21010
use bias2_top_s  bias2_top_s_0 ~/code/hibpm-sky130a-tapeout/mag/bias
timestamp 1686327621
transform 1 0 89960 0 1 18200
box 40 -4200 12860 21010
use exp  exp_0 ~/code/hibpm-sky130a-tapeout/mag/experiment
timestamp 1686846378
transform 1 0 49024 0 1 -32176
box -1624 -4624 10424 5824
use exp  exp_1
timestamp 1686846378
transform 1 0 49024 0 1 3424
box -1624 -4624 10424 5824
use isource  isource_0 ~/code/hibpm-sky130a-tapeout/mag/isource
timestamp 1684166381
transform 1 0 49308 0 1 19900
box -308 -5900 23140 17576
use outd_50ohm_hg  outd_50ohm_hg_0 ~/code/hibpm-sky130a-tapeout/mag/outd_50Ohm
timestamp 1687207134
transform 1 0 89522 0 1 -46420
box -10522 -8580 17040 8520
use outd_50ohm_hg  outd_50ohm_hg_1
timestamp 1687207134
transform 1 0 89522 0 1 -10420
box -10522 -8580 17040 8520
use tia_top  tia_top_0 ~/code/hibpm-sky130a-tapeout/mag/tiaA
timestamp 1686667164
transform 1 0 52628 0 1 -50920
box -3628 -4080 25704 24280
use tia_top  tia_top_1
timestamp 1686667164
transform 1 0 52628 0 1 -14920
box -3628 -4080 25704 24280
<< labels >>
rlabel metal3 34000 28320 35060 32600 1 VDD
port 2 n
rlabel metal3 34220 33440 34880 37380 1 VSS
rlabel metal3 110520 28100 112240 32820 1 VSS
rlabel space 110540 33240 111840 37760 1 VDD
rlabel metal3 33800 -8200 35100 -4900 1 In_ref1
port 3 n
rlabel metal3 34000 12800 35300 16100 1 In1
port 4 n
rlabel metal3 34000 -50500 35000 -48200 1 In_ref2
port 5 n
rlabel metal3 33900 -28300 34500 -26300 1 In2
port 6 n
rlabel metal3 111400 -48600 112200 -46800 1 Out_P2
port 11 n
rlabel metal3 111200 -29600 112000 -28000 1 Out_N2
port 12 n
rlabel metal3 111600 -8400 112000 -7400 1 Out_P1
port 13 n
rlabel metal3 111600 14000 112200 15600 1 Out_N1
port 14 n
rlabel metal3 110600 38600 112000 42600 1 VSS
port 15 n
rlabel metal4 59700 -32000 60600 -30700 1 In2_e
rlabel metal4 53200 -33800 54100 -33300 1 In2_ref_r
rlabel metal4 53000 3900 53900 4400 1 In1_ref_r
rlabel metal4 59700 3700 60600 4200 1 In1_r
<< end >>
