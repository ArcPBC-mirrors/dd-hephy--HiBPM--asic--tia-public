magic
tech sky130A
magscale 1 2
timestamp 1684929745
<< metal3 >>
rect -1186 1612 1186 1640
rect -1186 -1612 1102 1612
rect 1166 -1612 1186 1612
rect -1186 -1640 1186 -1612
<< via3 >>
rect 1102 -1612 1166 1612
<< mimcap >>
rect -1146 1560 854 1600
rect -1146 -1560 -1106 1560
rect 814 -1560 854 1560
rect -1146 -1600 854 -1560
<< mimcapcontact >>
rect -1106 -1560 814 1560
<< metal4 >>
rect 1086 1612 1182 1628
rect -1107 1560 815 1561
rect -1107 -1560 -1106 1560
rect 814 -1560 815 1560
rect -1107 -1561 815 -1560
rect 1086 -1612 1102 1612
rect 1166 -1612 1182 1612
rect 1086 -1628 1182 -1612
<< properties >>
string FIXED_BBOX -1186 -1640 894 1640
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 16 val 329.88 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
