magic
tech sky130A
magscale 1 2
timestamp 1689781139
<< error_p >>
rect 36380 1091213 36382 1091297
rect 36464 1091172 36466 1091213
rect 122022 1091172 122024 1091297
rect 136822 1075313 136837 1075328
rect 136742 1075233 136757 1075248
rect 21647 1073352 21662 1073367
rect 21567 1073272 21582 1073287
rect 133389 1068693 133394 1068699
rect 136822 975313 136837 975328
rect 136742 975233 136757 975248
rect 21647 973352 21662 973367
rect 21567 973272 21582 973287
rect 133389 968693 133394 968699
rect 136822 875313 136837 875328
rect 136742 875233 136757 875248
rect 21647 873352 21662 873367
rect 21567 873272 21582 873287
rect 133389 868693 133394 868699
rect 136822 775313 136837 775328
rect 136742 775233 136757 775248
rect 21647 773352 21662 773367
rect 21567 773272 21582 773287
rect 133389 768693 133394 768699
rect 136822 675313 136837 675328
rect 136742 675233 136757 675248
rect 21647 673352 21662 673367
rect 21567 673272 21582 673287
rect 133389 668693 133394 668699
rect 136822 575313 136837 575328
rect 136742 575233 136757 575248
rect 21647 573352 21662 573367
rect 21567 573272 21582 573287
rect 133389 568693 133394 568699
rect 136822 475313 136837 475328
rect 136742 475233 136757 475248
rect 21647 473352 21662 473367
rect 21567 473272 21582 473287
rect 133389 468693 133394 468699
rect 136822 375313 136837 375328
rect 136742 375233 136757 375248
rect 21647 373352 21662 373367
rect 21567 373272 21582 373287
rect 133389 368693 133394 368699
rect 136822 275313 136837 275328
rect 136742 275233 136757 275248
rect 21647 273352 21662 273367
rect 21567 273272 21582 273287
rect 133389 268693 133394 268699
rect 36464 172387 36466 172512
rect 121938 172428 121940 172512
rect 122022 172387 122024 172428
rect 62058 171038 62114 171094
rect 63231 149964 63287 149988
use core4  core4_0
timestamp 1689778598
transform 1 0 6220 0 1 1038762
box 33200 -62200 112700 42900
use core4  core4_1
timestamp 1689778598
transform 1 0 6220 0 1 838800
box 33200 -62200 112700 42900
use core4  core4_2
timestamp 1689778598
transform 1 0 6220 0 1 938800
box 33200 -62200 112700 42900
use core4  core4_3
timestamp 1689778598
transform 1 0 6220 0 1 438800
box 33200 -62200 112700 42900
use core4  core4_4
timestamp 1689778598
transform 1 0 6220 0 1 338800
box 33200 -62200 112700 42900
use core4  core4_5
timestamp 1689778598
transform 1 0 6220 0 1 238800
box 33200 -62200 112700 42900
use core4  core4_6
timestamp 1689778598
transform 1 0 6220 0 1 538800
box 33200 -62200 112700 42900
use core4  core4_7
timestamp 1689778598
transform 1 0 6220 0 1 638600
box 33200 -62200 112700 42900
use core4  core4_8
timestamp 1689778598
transform 1 0 6220 0 1 738600
box 33200 -62200 112700 42900
use frame_modBC  frame_modBC_0 ~/code/hibpm-sky130a-tapeout/mag/frame
timestamp 1689779212
transform 1 0 6202 0 1 1038800
box -6000 -897800 152000 83800
<< end >>
