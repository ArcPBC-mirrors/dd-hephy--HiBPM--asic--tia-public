magic
tech sky130A
magscale 1 2
timestamp 1689861403
<< error_p >>
rect 53942 1116178 53946 1116194
rect 74942 1116178 74946 1116194
rect 95942 1116180 95944 1116194
rect 95944 1116178 95946 1116180
rect 116942 1116178 116946 1116194
rect 53946 1115958 53949 1116178
rect 74946 1115958 74949 1116178
rect 95946 1116137 95949 1116178
rect 116946 1115958 116949 1116178
rect 41189 1115909 41417 1115925
rect 62189 1115909 62417 1115925
rect 83189 1115909 83417 1115925
rect 104189 1115909 104417 1115925
rect 41186 1115898 41189 1115909
rect 62186 1115898 62189 1115909
rect 83186 1115898 83189 1115909
rect 104186 1115898 104189 1115909
rect 54206 1103442 54218 1103462
rect 75206 1103442 75218 1103462
rect 96206 1103442 96218 1103462
rect 117206 1103442 117218 1103462
rect 53982 1103435 54206 1103442
rect 74982 1103435 75206 1103442
rect 95982 1103435 96206 1103442
rect 116982 1103435 117206 1103442
rect 41455 1103182 41458 1103190
rect 62455 1103182 62458 1103190
rect 83455 1103182 83458 1103190
rect 104455 1103182 104458 1103190
rect 41458 1103166 41462 1103182
rect 62458 1103166 62462 1103182
rect 83458 1103166 83462 1103182
rect 104458 1103166 104462 1103182
rect 36380 1091213 36382 1091297
rect 36464 1091172 36466 1091213
rect 122022 1091172 122024 1091297
rect 19340 1080804 19360 1080816
rect 151500 1080813 151511 1080816
rect 19360 1080580 19367 1080804
rect 151511 1080585 151527 1080813
rect 6624 1080544 6844 1080547
rect 138784 1080544 139004 1080547
rect 6608 1080540 6624 1080544
rect 138768 1080540 138784 1080544
rect 19620 1068056 19636 1068060
rect 151780 1068056 151796 1068060
rect 19400 1068053 19620 1068056
rect 151560 1068053 151780 1068056
rect 6877 1067787 6893 1068015
rect 139037 1067796 139044 1068020
rect 6893 1067784 6904 1067787
rect 139044 1067784 139064 1067796
rect 19340 1060804 19360 1060816
rect 151500 1060813 151511 1060816
rect 19360 1060580 19367 1060804
rect 151511 1060585 151527 1060813
rect 6624 1060544 6844 1060547
rect 138784 1060544 139004 1060547
rect 6608 1060540 6624 1060544
rect 138768 1060540 138784 1060544
rect 19620 1048056 19636 1048060
rect 151780 1048056 151796 1048060
rect 19400 1048053 19620 1048056
rect 151560 1048053 151780 1048056
rect 6877 1047787 6893 1048015
rect 139037 1047796 139044 1048020
rect 6893 1047784 6904 1047787
rect 139044 1047784 139064 1047796
rect 19340 1040804 19360 1040816
rect 151500 1040813 151511 1040816
rect 19360 1040580 19367 1040804
rect 151511 1040585 151527 1040813
rect 6624 1040544 6844 1040547
rect 138784 1040544 139004 1040547
rect 6608 1040540 6624 1040544
rect 138768 1040540 138784 1040544
rect 19620 1028056 19636 1028060
rect 151780 1028056 151796 1028060
rect 19400 1028053 19620 1028056
rect 151560 1028053 151780 1028056
rect 6877 1027787 6893 1028015
rect 139037 1027796 139044 1028020
rect 6893 1027784 6904 1027787
rect 139044 1027784 139064 1027796
rect 19340 1020804 19360 1020816
rect 151500 1020813 151511 1020816
rect 19360 1020580 19367 1020804
rect 151511 1020585 151527 1020813
rect 6624 1020544 6844 1020547
rect 138784 1020544 139004 1020547
rect 6608 1020540 6624 1020544
rect 138768 1020540 138784 1020544
rect 19620 1008056 19636 1008060
rect 151780 1008056 151796 1008060
rect 19400 1008053 19620 1008056
rect 151560 1008053 151780 1008056
rect 6877 1007787 6893 1008015
rect 139037 1007796 139044 1008020
rect 6893 1007784 6904 1007787
rect 139044 1007784 139064 1007796
rect 19340 1000804 19360 1000816
rect 151500 1000813 151511 1000816
rect 19360 1000580 19367 1000804
rect 151511 1000585 151527 1000813
rect 6624 1000544 6844 1000547
rect 138784 1000544 139004 1000547
rect 6608 1000540 6624 1000544
rect 138768 1000540 138784 1000544
rect 19620 988056 19636 988060
rect 151780 988056 151796 988060
rect 19400 988053 19620 988056
rect 151560 988053 151780 988056
rect 6877 987787 6893 988015
rect 139037 987796 139044 988020
rect 6893 987784 6904 987787
rect 139044 987784 139064 987796
rect 19340 980804 19360 980816
rect 151500 980813 151511 980816
rect 19360 980580 19367 980804
rect 151511 980585 151527 980813
rect 6624 980544 6844 980547
rect 138784 980544 139004 980547
rect 6608 980540 6624 980544
rect 138768 980540 138784 980544
rect 19620 968056 19636 968060
rect 151780 968056 151796 968060
rect 19400 968053 19620 968056
rect 151560 968053 151780 968056
rect 6877 967787 6893 968015
rect 139037 967796 139044 968020
rect 6893 967784 6904 967787
rect 139044 967784 139064 967796
rect 19340 960804 19360 960816
rect 151500 960813 151511 960816
rect 19360 960580 19367 960804
rect 151511 960585 151527 960813
rect 6624 960544 6844 960547
rect 138784 960544 139004 960547
rect 6608 960540 6624 960544
rect 138768 960540 138784 960544
rect 19620 948056 19636 948060
rect 151780 948056 151796 948060
rect 19400 948053 19620 948056
rect 151560 948053 151780 948056
rect 6877 947787 6893 948015
rect 139037 947796 139044 948020
rect 6893 947784 6904 947787
rect 139044 947784 139064 947796
rect 19340 940804 19360 940816
rect 151500 940813 151511 940816
rect 19360 940580 19367 940804
rect 151511 940585 151527 940813
rect 6624 940544 6844 940547
rect 138784 940544 139004 940547
rect 6608 940540 6624 940544
rect 138768 940540 138784 940544
rect 19620 928056 19636 928060
rect 151780 928056 151796 928060
rect 19400 928053 19620 928056
rect 151560 928053 151780 928056
rect 6877 927787 6893 928015
rect 139037 927796 139044 928020
rect 6893 927784 6904 927787
rect 139044 927784 139064 927796
rect 19340 920804 19360 920816
rect 151500 920813 151511 920816
rect 19360 920580 19367 920804
rect 151511 920585 151527 920813
rect 6624 920544 6844 920547
rect 138784 920544 139004 920547
rect 6608 920540 6624 920544
rect 138768 920540 138784 920544
rect 19620 908056 19636 908060
rect 151780 908056 151796 908060
rect 19400 908053 19620 908056
rect 151560 908053 151780 908056
rect 6877 907787 6893 908015
rect 139037 907796 139044 908020
rect 6893 907784 6904 907787
rect 139044 907784 139064 907796
rect 19340 900804 19360 900816
rect 151500 900813 151511 900816
rect 19360 900580 19367 900804
rect 151511 900585 151527 900813
rect 6624 900544 6844 900547
rect 138784 900544 139004 900547
rect 6608 900540 6624 900544
rect 138768 900540 138784 900544
rect 19620 888056 19636 888060
rect 151780 888056 151796 888060
rect 19400 888053 19620 888056
rect 151560 888053 151780 888056
rect 6877 887787 6893 888015
rect 139037 887796 139044 888020
rect 6893 887784 6904 887787
rect 139044 887784 139064 887796
rect 19340 880804 19360 880816
rect 151500 880813 151511 880816
rect 19360 880580 19367 880804
rect 151511 880585 151527 880813
rect 6624 880544 6844 880547
rect 138784 880544 139004 880547
rect 6608 880540 6624 880544
rect 138768 880540 138784 880544
rect 19620 868056 19636 868060
rect 151780 868056 151796 868060
rect 19400 868053 19620 868056
rect 151560 868053 151780 868056
rect 6877 867787 6893 868015
rect 139037 867796 139044 868020
rect 6893 867784 6904 867787
rect 139044 867784 139064 867796
rect 19340 860804 19360 860816
rect 151500 860813 151511 860816
rect 19360 860580 19367 860804
rect 151511 860585 151527 860813
rect 6624 860544 6844 860547
rect 138784 860544 139004 860547
rect 6608 860540 6624 860544
rect 138768 860540 138784 860544
rect 19620 848056 19636 848060
rect 151780 848056 151796 848060
rect 19400 848053 19620 848056
rect 151560 848053 151780 848056
rect 6877 847787 6893 848015
rect 139037 847796 139044 848020
rect 6893 847784 6904 847787
rect 139044 847784 139064 847796
rect 19340 840804 19360 840816
rect 151500 840813 151511 840816
rect 19360 840580 19367 840804
rect 151511 840585 151527 840813
rect 6624 840544 6844 840547
rect 138784 840544 139004 840547
rect 6608 840540 6624 840544
rect 138768 840540 138784 840544
rect 19620 828056 19636 828060
rect 151780 828056 151796 828060
rect 19400 828053 19620 828056
rect 151560 828053 151780 828056
rect 6877 827787 6893 828015
rect 139037 827796 139044 828020
rect 6893 827784 6904 827787
rect 139044 827784 139064 827796
rect 19340 820804 19360 820816
rect 151500 820813 151511 820816
rect 19360 820580 19367 820804
rect 151511 820585 151527 820813
rect 6624 820544 6844 820547
rect 138784 820544 139004 820547
rect 6608 820540 6624 820544
rect 138768 820540 138784 820544
rect 19620 808056 19636 808060
rect 151780 808056 151796 808060
rect 19400 808053 19620 808056
rect 151560 808053 151780 808056
rect 6877 807787 6893 808015
rect 139037 807796 139044 808020
rect 6893 807784 6904 807787
rect 139044 807784 139064 807796
rect 19340 800804 19360 800816
rect 151500 800813 151511 800816
rect 19360 800580 19367 800804
rect 151511 800585 151527 800813
rect 6624 800544 6844 800547
rect 138784 800544 139004 800547
rect 6608 800540 6624 800544
rect 138768 800540 138784 800544
rect 19620 788056 19636 788060
rect 151780 788056 151796 788060
rect 19400 788053 19620 788056
rect 151560 788053 151780 788056
rect 6877 787787 6893 788015
rect 139037 787796 139044 788020
rect 6893 787784 6904 787787
rect 139044 787784 139064 787796
rect 19340 780804 19360 780816
rect 151500 780813 151511 780816
rect 19360 780580 19367 780804
rect 151511 780585 151527 780813
rect 6624 780544 6844 780547
rect 138784 780544 139004 780547
rect 6608 780540 6624 780544
rect 138768 780540 138784 780544
rect 19620 768056 19636 768060
rect 151780 768056 151796 768060
rect 19400 768053 19620 768056
rect 151560 768053 151780 768056
rect 6877 767787 6893 768015
rect 139037 767796 139044 768020
rect 6893 767784 6904 767787
rect 139044 767784 139064 767796
rect 19340 760804 19360 760816
rect 151500 760813 151511 760816
rect 19360 760580 19367 760804
rect 151511 760585 151527 760813
rect 6624 760544 6844 760547
rect 138784 760544 139004 760547
rect 6608 760540 6624 760544
rect 138768 760540 138784 760544
rect 19620 748056 19636 748060
rect 151780 748056 151796 748060
rect 19400 748053 19620 748056
rect 151560 748053 151780 748056
rect 6877 747787 6893 748015
rect 139037 747796 139044 748020
rect 6893 747784 6904 747787
rect 139044 747784 139064 747796
rect 19340 740804 19360 740816
rect 151500 740813 151511 740816
rect 19360 740580 19367 740804
rect 151511 740585 151527 740813
rect 6624 740544 6844 740547
rect 138784 740544 139004 740547
rect 6608 740540 6624 740544
rect 138768 740540 138784 740544
rect 19620 728056 19636 728060
rect 151780 728056 151796 728060
rect 19400 728053 19620 728056
rect 151560 728053 151780 728056
rect 6877 727787 6893 728015
rect 139037 727796 139044 728020
rect 6893 727784 6904 727787
rect 139044 727784 139064 727796
rect 19340 720804 19360 720816
rect 151500 720813 151511 720816
rect 19360 720580 19367 720804
rect 151511 720585 151527 720813
rect 6624 720544 6844 720547
rect 138784 720544 139004 720547
rect 6608 720540 6624 720544
rect 138768 720540 138784 720544
rect 19620 708056 19636 708060
rect 151780 708056 151796 708060
rect 19400 708053 19620 708056
rect 151560 708053 151780 708056
rect 6877 707787 6893 708015
rect 139037 707796 139044 708020
rect 6893 707784 6904 707787
rect 139044 707784 139064 707796
rect 19340 700804 19360 700816
rect 151500 700813 151511 700816
rect 19360 700580 19367 700804
rect 151511 700585 151527 700813
rect 6624 700544 6844 700547
rect 138784 700544 139004 700547
rect 6608 700540 6624 700544
rect 138768 700540 138784 700544
rect 19620 688056 19636 688060
rect 151780 688056 151796 688060
rect 19400 688053 19620 688056
rect 151560 688053 151780 688056
rect 6877 687787 6893 688015
rect 139037 687796 139044 688020
rect 6893 687784 6904 687787
rect 139044 687784 139064 687796
rect 19340 680804 19360 680816
rect 151500 680813 151511 680816
rect 19360 680580 19367 680804
rect 151511 680585 151527 680813
rect 6624 680544 6844 680547
rect 138784 680544 139004 680547
rect 6608 680540 6624 680544
rect 138768 680540 138784 680544
rect 19620 668056 19636 668060
rect 151780 668056 151796 668060
rect 19400 668053 19620 668056
rect 151560 668053 151780 668056
rect 6877 667787 6893 668015
rect 139037 667796 139044 668020
rect 6893 667784 6904 667787
rect 139044 667784 139064 667796
rect 19340 660804 19360 660816
rect 151500 660813 151511 660816
rect 19360 660580 19367 660804
rect 151511 660585 151527 660813
rect 6624 660544 6844 660547
rect 138784 660544 139004 660547
rect 6608 660540 6624 660544
rect 138768 660540 138784 660544
rect 19620 648056 19636 648060
rect 151780 648056 151796 648060
rect 19400 648053 19620 648056
rect 151560 648053 151780 648056
rect 6877 647787 6893 648015
rect 139037 647796 139044 648020
rect 6893 647784 6904 647787
rect 139044 647784 139064 647796
rect 19340 640804 19360 640816
rect 151500 640813 151511 640816
rect 19360 640580 19367 640804
rect 151511 640585 151527 640813
rect 6624 640544 6844 640547
rect 138784 640544 139004 640547
rect 6608 640540 6624 640544
rect 138768 640540 138784 640544
rect 19620 628056 19636 628060
rect 151780 628056 151796 628060
rect 19400 628053 19620 628056
rect 151560 628053 151780 628056
rect 6877 627787 6893 628015
rect 139037 627796 139044 628020
rect 6893 627784 6904 627787
rect 139044 627784 139064 627796
rect 19340 620804 19360 620816
rect 151500 620813 151511 620816
rect 19360 620580 19367 620804
rect 151511 620585 151527 620813
rect 6624 620544 6844 620547
rect 138784 620544 139004 620547
rect 6608 620540 6624 620544
rect 138768 620540 138784 620544
rect 19620 608056 19636 608060
rect 151780 608056 151796 608060
rect 19400 608053 19620 608056
rect 151560 608053 151780 608056
rect 6877 607787 6893 608015
rect 139037 607796 139044 608020
rect 6893 607784 6904 607787
rect 139044 607784 139064 607796
rect 19340 600804 19360 600816
rect 151500 600813 151511 600816
rect 19360 600580 19367 600804
rect 151511 600585 151527 600813
rect 6624 600544 6844 600547
rect 138784 600544 139004 600547
rect 6608 600540 6624 600544
rect 138768 600540 138784 600544
rect 19620 588056 19636 588060
rect 151780 588056 151796 588060
rect 19400 588053 19620 588056
rect 151560 588053 151780 588056
rect 6877 587787 6893 588015
rect 139037 587796 139044 588020
rect 6893 587784 6904 587787
rect 139044 587784 139064 587796
rect 19340 580804 19360 580816
rect 151500 580813 151511 580816
rect 19360 580580 19367 580804
rect 151511 580585 151527 580813
rect 6624 580544 6844 580547
rect 138784 580544 139004 580547
rect 6608 580540 6624 580544
rect 138768 580540 138784 580544
rect 19620 568056 19636 568060
rect 151780 568056 151796 568060
rect 19400 568053 19620 568056
rect 151560 568053 151780 568056
rect 6877 567787 6893 568015
rect 139037 567796 139044 568020
rect 6893 567784 6904 567787
rect 139044 567784 139064 567796
rect 19340 560804 19360 560816
rect 151500 560813 151511 560816
rect 19360 560580 19367 560804
rect 151511 560585 151527 560813
rect 6624 560544 6844 560547
rect 138784 560544 139004 560547
rect 6608 560540 6624 560544
rect 138768 560540 138784 560544
rect 19620 548056 19636 548060
rect 151780 548056 151796 548060
rect 19400 548053 19620 548056
rect 151560 548053 151780 548056
rect 6877 547787 6893 548015
rect 139037 547796 139044 548020
rect 6893 547784 6904 547787
rect 139044 547784 139064 547796
rect 19340 540804 19360 540816
rect 151500 540813 151511 540816
rect 19360 540580 19367 540804
rect 151511 540585 151527 540813
rect 6624 540544 6844 540547
rect 138784 540544 139004 540547
rect 6608 540540 6624 540544
rect 138768 540540 138784 540544
rect 19620 528056 19636 528060
rect 151780 528056 151796 528060
rect 19400 528053 19620 528056
rect 151560 528053 151780 528056
rect 6877 527787 6893 528015
rect 139037 527796 139044 528020
rect 6893 527784 6904 527787
rect 139044 527784 139064 527796
rect 19340 520804 19360 520816
rect 151500 520813 151511 520816
rect 19360 520580 19367 520804
rect 151511 520585 151527 520813
rect 6624 520544 6844 520547
rect 138784 520544 139004 520547
rect 6608 520540 6624 520544
rect 138768 520540 138784 520544
rect 19620 508056 19636 508060
rect 151780 508056 151796 508060
rect 19400 508053 19620 508056
rect 151560 508053 151780 508056
rect 6877 507787 6893 508015
rect 139037 507796 139044 508020
rect 6893 507784 6904 507787
rect 139044 507784 139064 507796
rect 19340 500804 19360 500816
rect 151500 500813 151511 500816
rect 19360 500580 19367 500804
rect 151511 500585 151527 500813
rect 6624 500544 6844 500547
rect 138784 500544 139004 500547
rect 6608 500540 6624 500544
rect 138768 500540 138784 500544
rect 19620 488056 19636 488060
rect 151780 488056 151796 488060
rect 19400 488053 19620 488056
rect 151560 488053 151780 488056
rect 6877 487787 6893 488015
rect 139037 487796 139044 488020
rect 6893 487784 6904 487787
rect 139044 487784 139064 487796
rect 19340 480804 19360 480816
rect 151500 480813 151511 480816
rect 19360 480580 19367 480804
rect 151511 480585 151527 480813
rect 6624 480544 6844 480547
rect 138784 480544 139004 480547
rect 6608 480540 6624 480544
rect 138768 480540 138784 480544
rect 19620 468056 19636 468060
rect 151780 468056 151796 468060
rect 19400 468053 19620 468056
rect 151560 468053 151780 468056
rect 6877 467787 6893 468015
rect 139037 467796 139044 468020
rect 6893 467784 6904 467787
rect 139044 467784 139064 467796
rect 19340 460804 19360 460816
rect 151500 460813 151511 460816
rect 19360 460580 19367 460804
rect 151511 460585 151527 460813
rect 6624 460544 6844 460547
rect 138784 460544 139004 460547
rect 6608 460540 6624 460544
rect 138768 460540 138784 460544
rect 19620 448056 19636 448060
rect 151780 448056 151796 448060
rect 19400 448053 19620 448056
rect 151560 448053 151780 448056
rect 6877 447787 6893 448015
rect 139037 447796 139044 448020
rect 6893 447784 6904 447787
rect 139044 447784 139064 447796
rect 19340 440804 19360 440816
rect 151500 440813 151511 440816
rect 19360 440580 19367 440804
rect 151511 440585 151527 440813
rect 6624 440544 6844 440547
rect 138784 440544 139004 440547
rect 6608 440540 6624 440544
rect 138768 440540 138784 440544
rect 19620 428056 19636 428060
rect 151780 428056 151796 428060
rect 19400 428053 19620 428056
rect 151560 428053 151780 428056
rect 6877 427787 6893 428015
rect 139037 427796 139044 428020
rect 6893 427784 6904 427787
rect 139044 427784 139064 427796
rect 19340 420804 19360 420816
rect 151500 420813 151511 420816
rect 19360 420580 19367 420804
rect 151511 420585 151527 420813
rect 6624 420544 6844 420547
rect 138784 420544 139004 420547
rect 6608 420540 6624 420544
rect 138768 420540 138784 420544
rect 19620 408056 19636 408060
rect 151780 408056 151796 408060
rect 19400 408053 19620 408056
rect 151560 408053 151780 408056
rect 6877 407787 6893 408015
rect 139037 407796 139044 408020
rect 6893 407784 6904 407787
rect 139044 407784 139064 407796
rect 19340 400804 19360 400816
rect 151500 400813 151511 400816
rect 19360 400580 19367 400804
rect 151511 400585 151527 400813
rect 6624 400544 6844 400547
rect 138784 400544 139004 400547
rect 6608 400540 6624 400544
rect 138768 400540 138784 400544
rect 19620 388056 19636 388060
rect 151780 388056 151796 388060
rect 19400 388053 19620 388056
rect 151560 388053 151780 388056
rect 6877 387787 6893 388015
rect 139037 387796 139044 388020
rect 6893 387784 6904 387787
rect 139044 387784 139064 387796
rect 19340 380804 19360 380816
rect 151500 380813 151511 380816
rect 19360 380580 19367 380804
rect 151511 380585 151527 380813
rect 6624 380544 6844 380547
rect 138784 380544 139004 380547
rect 6608 380540 6624 380544
rect 138768 380540 138784 380544
rect 19620 368056 19636 368060
rect 151780 368056 151796 368060
rect 19400 368053 19620 368056
rect 151560 368053 151780 368056
rect 6877 367787 6893 368015
rect 139037 367796 139044 368020
rect 6893 367784 6904 367787
rect 139044 367784 139064 367796
rect 19340 360804 19360 360816
rect 151500 360813 151511 360816
rect 19360 360580 19367 360804
rect 151511 360585 151527 360813
rect 6624 360544 6844 360547
rect 138784 360544 139004 360547
rect 6608 360540 6624 360544
rect 138768 360540 138784 360544
rect 19620 348056 19636 348060
rect 151780 348056 151796 348060
rect 19400 348053 19620 348056
rect 151560 348053 151780 348056
rect 6877 347787 6893 348015
rect 139037 347796 139044 348020
rect 6893 347784 6904 347787
rect 139044 347784 139064 347796
rect 19340 340804 19360 340816
rect 151500 340813 151511 340816
rect 19360 340580 19367 340804
rect 151511 340585 151527 340813
rect 6624 340544 6844 340547
rect 138784 340544 139004 340547
rect 6608 340540 6624 340544
rect 138768 340540 138784 340544
rect 19620 328056 19636 328060
rect 151780 328056 151796 328060
rect 19400 328053 19620 328056
rect 151560 328053 151780 328056
rect 6877 327787 6893 328015
rect 139037 327796 139044 328020
rect 6893 327784 6904 327787
rect 139044 327784 139064 327796
rect 19340 320804 19360 320816
rect 151500 320813 151511 320816
rect 19360 320580 19367 320804
rect 151511 320585 151527 320813
rect 6624 320544 6844 320547
rect 138784 320544 139004 320547
rect 6608 320540 6624 320544
rect 138768 320540 138784 320544
rect 19620 308056 19636 308060
rect 151780 308056 151796 308060
rect 19400 308053 19620 308056
rect 151560 308053 151780 308056
rect 6877 307787 6893 308015
rect 139037 307796 139044 308020
rect 6893 307784 6904 307787
rect 139044 307784 139064 307796
rect 19340 300804 19360 300816
rect 151500 300813 151511 300816
rect 19360 300580 19367 300804
rect 151511 300585 151527 300813
rect 6624 300544 6844 300547
rect 138784 300544 139004 300547
rect 6608 300540 6624 300544
rect 138768 300540 138784 300544
rect 19620 288056 19636 288060
rect 151780 288056 151796 288060
rect 19400 288053 19620 288056
rect 151560 288053 151780 288056
rect 6877 287787 6893 288015
rect 139037 287796 139044 288020
rect 6893 287784 6904 287787
rect 139044 287784 139064 287796
rect 19340 280804 19360 280816
rect 151500 280813 151511 280816
rect 19360 280580 19367 280804
rect 151511 280585 151527 280813
rect 6624 280544 6844 280547
rect 138784 280544 139004 280547
rect 6608 280540 6624 280544
rect 138768 280540 138784 280544
rect 19620 268056 19636 268060
rect 151780 268056 151796 268060
rect 19400 268053 19620 268056
rect 151560 268053 151780 268056
rect 6877 267787 6893 268015
rect 139037 267796 139044 268020
rect 6893 267784 6904 267787
rect 139044 267784 139064 267796
rect 19340 260804 19360 260816
rect 151500 260813 151511 260816
rect 19360 260580 19367 260804
rect 151511 260585 151527 260813
rect 6624 260544 6844 260547
rect 138784 260544 139004 260547
rect 6608 260540 6624 260544
rect 138768 260540 138784 260544
rect 19620 248056 19636 248060
rect 151780 248056 151796 248060
rect 19400 248053 19620 248056
rect 151560 248053 151780 248056
rect 6877 247787 6893 248015
rect 139037 247796 139044 248020
rect 6893 247784 6904 247787
rect 139044 247784 139064 247796
rect 19340 240804 19360 240816
rect 151500 240813 151511 240816
rect 19360 240580 19367 240804
rect 151511 240585 151527 240813
rect 6624 240544 6844 240547
rect 138784 240544 139004 240547
rect 6608 240540 6624 240544
rect 138768 240540 138784 240544
rect 19620 228056 19636 228060
rect 151780 228056 151796 228060
rect 19400 228053 19620 228056
rect 151560 228053 151780 228056
rect 6877 227787 6893 228015
rect 139037 227796 139044 228020
rect 6893 227784 6904 227787
rect 139044 227784 139064 227796
rect 19340 220804 19360 220816
rect 151500 220813 151511 220816
rect 19360 220580 19367 220804
rect 151511 220585 151527 220813
rect 6624 220544 6844 220547
rect 138784 220544 139004 220547
rect 6608 220540 6624 220544
rect 138768 220540 138784 220544
rect 19620 208056 19636 208060
rect 151780 208056 151796 208060
rect 19400 208053 19620 208056
rect 151560 208053 151780 208056
rect 6877 207787 6893 208015
rect 139037 207796 139044 208020
rect 6893 207784 6904 207787
rect 139044 207784 139064 207796
rect 19340 200804 19360 200816
rect 151500 200813 151511 200816
rect 19360 200580 19367 200804
rect 151511 200585 151527 200813
rect 6624 200544 6844 200547
rect 138784 200544 139004 200547
rect 6608 200540 6624 200544
rect 138768 200540 138784 200544
rect 19620 188056 19636 188060
rect 151780 188056 151796 188060
rect 19400 188053 19620 188056
rect 151560 188053 151780 188056
rect 6877 187787 6893 188015
rect 139037 187796 139044 188020
rect 6893 187784 6904 187787
rect 139044 187784 139064 187796
rect 36464 172387 36466 172512
rect 121938 172428 121940 172512
rect 122022 172387 122024 172428
rect 53942 160418 53946 160434
rect 74942 160418 74946 160434
rect 95942 160418 95946 160434
rect 116942 160418 116946 160434
rect 53946 160410 53949 160418
rect 74946 160410 74949 160418
rect 95946 160410 95949 160418
rect 116946 160410 116949 160418
rect 41198 160158 41422 160165
rect 62198 160158 62422 160165
rect 83198 160158 83422 160165
rect 104198 160158 104422 160165
rect 41186 160138 41198 160158
rect 62186 160138 62198 160158
rect 83186 160138 83198 160158
rect 104186 160138 104198 160158
rect 54215 147691 54218 147702
rect 75215 147691 75218 147702
rect 96215 147691 96218 147702
rect 117215 147691 117218 147702
rect 53987 147675 54215 147691
rect 74987 147675 75215 147691
rect 95987 147675 96215 147691
rect 116987 147675 117215 147691
rect 41455 147422 41458 147642
rect 62455 147422 62458 147463
rect 83455 147422 83458 147463
rect 104455 147422 104458 147642
rect 41458 147406 41462 147422
rect 62458 147420 62460 147422
rect 83458 147420 83460 147422
rect 62460 147406 62462 147420
rect 83460 147406 83462 147420
rect 104458 147406 104462 147422
use core4  core4_0
timestamp 1689861321
transform 1 0 6220 0 1 1038762
box 33200 -57200 112700 42900
use core4  core4_1
timestamp 1689861321
transform 1 0 6220 0 1 838800
box 33200 -57200 112700 42900
use core4  core4_2
timestamp 1689861321
transform 1 0 6220 0 1 938800
box 33200 -57200 112700 42900
use core4  core4_3
timestamp 1689861321
transform 1 0 6220 0 1 438800
box 33200 -57200 112700 42900
use core4  core4_4
timestamp 1689861321
transform 1 0 6220 0 1 338800
box 33200 -57200 112700 42900
use core4  core4_5
timestamp 1689861321
transform 1 0 6220 0 1 238800
box 33200 -57200 112700 42900
use core4  core4_6
timestamp 1689861321
transform 1 0 6220 0 1 538800
box 33200 -57200 112700 42900
use core4  core4_7
timestamp 1689861321
transform 1 0 6220 0 1 638600
box 33200 -57200 112700 42900
use core4  core4_8
timestamp 1689861321
transform 1 0 6220 0 1 738600
box 33200 -57200 112700 42900
use frame_modBC  frame_modBC_0 ~/code/hibpm-sky130a-tapeout/mag/frame
timestamp 1689775068
transform 1 0 6202 0 1 1038800
box -6000 -897800 152000 83800
<< end >>
