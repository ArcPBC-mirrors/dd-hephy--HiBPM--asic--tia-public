magic
tech sky130A
magscale 1 2
timestamp 1686667164
<< viali >>
rect 24360 5700 24580 5800
<< metal1 >>
rect 19540 19252 22096 19292
rect 19540 18996 21848 19252
rect 22068 18996 22096 19252
rect 19540 18960 22096 18996
rect 17222 18656 17232 18924
rect 17480 18656 17490 18924
rect 18182 18660 18192 18928
rect 18440 18660 18450 18928
rect 20234 18732 20244 18820
rect 20424 18732 20434 18820
rect 15156 15824 15968 15844
rect 15156 15716 15176 15824
rect 15348 15716 15968 15824
rect 15156 15696 15968 15716
rect 14276 13948 14532 13952
rect 14274 13844 14284 13948
rect 14416 13844 14532 13948
rect 14276 13840 14532 13844
rect 13872 13024 14068 13348
rect 15836 13228 15968 15696
rect 15836 13136 15848 13228
rect 15952 13136 15968 13228
rect 17240 13316 17404 18656
rect 21100 18100 21340 18120
rect 20770 17740 20780 18100
rect 21160 17740 21340 18100
rect 17240 13200 17260 13316
rect 17404 13200 17414 13316
rect 17240 13164 17404 13200
rect 15836 13124 15968 13136
rect 13872 12872 19380 13024
rect 11148 12796 11292 12800
rect 11148 12776 14500 12796
rect 11148 12676 14408 12776
rect 14484 12676 14500 12776
rect 11148 12664 14500 12676
rect 11148 11824 11292 12664
rect 1668 11652 11292 11824
rect 11404 12564 14168 12572
rect 11404 12412 14044 12564
rect 14192 12412 14202 12564
rect 11404 12404 14168 12412
rect -1380 4260 -1260 6000
rect 1668 4440 1800 11652
rect 11404 11564 11532 12404
rect 7124 11384 11532 11564
rect 7128 9092 7296 11384
rect 11404 11380 11532 11384
rect 11656 12196 14452 12212
rect 11656 12088 14340 12196
rect 14436 12088 14452 12196
rect 11656 12076 14452 12088
rect 10288 9700 11308 9712
rect 11656 9700 11804 12076
rect 10288 9500 11804 9700
rect 11656 9496 11804 9500
rect 1650 4320 1660 4440
rect 1820 4320 1830 4440
rect 1668 4284 1800 4320
rect -1380 4100 500 4260
rect 11540 4148 13600 4260
rect 11540 3672 11616 4148
rect 11784 3672 13600 4148
rect 14556 3748 14720 12872
rect 14804 12788 15192 12800
rect 14804 12780 15968 12788
rect 14804 12680 14824 12780
rect 14900 12772 15968 12780
rect 14900 12680 15848 12772
rect 15952 12680 15968 12772
rect 14804 12668 15968 12680
rect 14804 12664 15192 12668
rect 15004 11824 15124 12664
rect 15180 12476 17448 12512
rect 15180 12472 17256 12476
rect 15180 12364 15204 12472
rect 15300 12364 17256 12472
rect 15180 12360 17256 12364
rect 17400 12360 17448 12476
rect 15180 12344 17448 12360
rect 21100 12120 21340 17740
rect 21100 11880 25440 12120
rect 15000 11652 15124 11824
rect 15004 4440 15124 11652
rect 24330 8620 24340 9040
rect 24760 8620 24770 9040
rect 25220 8160 25440 11880
rect 24330 7740 24340 8160
rect 24760 7740 24770 8160
rect 25210 7740 25220 8160
rect 25640 7740 25650 8160
rect 24290 5920 24300 6480
rect 24600 5920 24610 6480
rect 24348 5800 24592 5806
rect 24348 5700 24360 5800
rect 24580 5700 24592 5800
rect 24348 5694 24592 5700
rect 14990 4320 15000 4440
rect 15130 4320 15140 4440
rect 15004 4264 15124 4320
rect 11540 3260 13600 3672
<< via1 >>
rect 21848 18996 22068 19252
rect 17232 18656 17480 18924
rect 18192 18660 18440 18928
rect 20244 18732 20424 18820
rect 15176 15716 15348 15824
rect 14284 13844 14416 13948
rect 15848 13136 15952 13228
rect 20780 17740 21160 18100
rect 17260 13200 17404 13316
rect 14408 12676 14484 12776
rect 14044 12412 14192 12564
rect 14340 12088 14436 12196
rect 1660 4320 1820 4440
rect 14824 12680 14900 12780
rect 15848 12680 15952 12772
rect 15204 12364 15300 12472
rect 17256 12360 17400 12476
rect 24340 8620 24760 9040
rect 24340 7740 24760 8160
rect 25220 7740 25640 8160
rect 24300 5920 24600 6480
rect 24360 5700 24580 5800
rect 15000 4320 15130 4440
<< metal2 >>
rect 21848 19252 22068 19262
rect 21848 18986 22068 18996
rect 17232 18924 17480 18934
rect 17232 18646 17480 18656
rect 18192 18928 18440 18938
rect 18440 18820 20436 18868
rect 18440 18732 20244 18820
rect 20424 18732 20436 18820
rect 18440 18708 20436 18732
rect 18192 18650 18440 18660
rect 20780 18100 21160 18110
rect 20780 17730 21160 17740
rect 15176 15824 15348 15834
rect 15176 15706 15348 15716
rect 14284 13948 14416 13958
rect 14276 13844 14284 13940
rect 14416 13844 14424 13940
rect 14036 13100 14204 13108
rect 14276 13100 14424 13844
rect 17260 13316 17408 13328
rect 14036 12996 14424 13100
rect -1200 12080 13840 12920
rect 14036 12564 14204 12996
rect 14276 12988 14424 12996
rect 15848 13228 15952 13240
rect 14400 12780 14920 12800
rect 14400 12776 14824 12780
rect 14400 12676 14408 12776
rect 14484 12680 14824 12776
rect 14900 12680 14920 12780
rect 14484 12676 14920 12680
rect 14400 12660 14920 12676
rect 15848 12772 15952 13136
rect 15848 12668 15952 12680
rect 17404 13200 17408 13316
rect 14036 12412 14044 12564
rect 14192 12412 14204 12564
rect 14036 12408 14204 12412
rect 15184 12472 15316 12496
rect 17260 12486 17408 13200
rect 14044 12402 14192 12408
rect 15184 12364 15204 12472
rect 15300 12364 15316 12472
rect 15184 12208 15316 12364
rect 17256 12476 17408 12486
rect 17400 12360 17408 12476
rect 17256 12350 17408 12360
rect 17260 12348 17408 12350
rect 14344 12206 15316 12208
rect -1200 11080 -260 12080
rect 3640 11600 13840 12080
rect 14340 12196 15316 12206
rect 14436 12108 15316 12196
rect 14436 12088 15292 12108
rect 14340 12084 15292 12088
rect 14340 12078 14436 12084
rect 3640 11480 24200 11600
rect -1200 10440 2400 11080
rect 11900 10440 15700 11120
rect 24020 10440 24200 11480
rect -1200 10300 24200 10440
rect 7200 8820 7560 9080
rect 20600 8840 20960 9100
rect 24340 9040 24760 9050
rect 24340 8610 24760 8620
rect -3060 8060 -2792 8252
rect 24340 8160 24760 8170
rect 24340 7730 24760 7740
rect 25220 8160 25640 8170
rect 25220 7730 25640 7740
rect 24300 6480 24600 6490
rect 24300 5910 24600 5920
rect 24360 5800 24580 5810
rect 5020 5460 5120 5780
rect 24360 5690 24580 5700
rect 1660 4440 1820 4450
rect 15000 4440 15130 4450
rect 1820 4420 1840 4430
rect 1820 4330 1840 4340
rect 1660 4310 1820 4320
rect 15000 4310 15130 4320
<< via2 >>
rect 21848 18996 22068 19252
rect 17232 18656 17480 18924
rect 18192 18660 18440 18928
rect 20780 17740 21160 18100
rect 15176 15716 15348 15824
rect -260 11480 3640 12080
rect -260 11120 24020 11480
rect -260 11080 11900 11120
rect 2400 10440 11900 11080
rect 15700 10440 24020 11120
rect 24340 8620 24760 9040
rect 24340 7740 24760 8160
rect 25220 7740 25640 8160
rect 24320 6120 24500 6360
rect 24360 5700 24580 5800
rect 1660 4340 1820 4420
rect 1820 4340 1840 4420
rect 15000 4320 15130 4440
<< metal3 >>
rect 9100 22920 23020 24280
rect 9120 12920 10600 22920
rect 21812 19252 23020 22920
rect 21812 18996 21848 19252
rect 22068 18996 23020 19252
rect 17222 18924 17490 18929
rect 17222 18656 17232 18924
rect 17480 18656 17490 18924
rect 17222 18651 17490 18656
rect 18182 18928 18450 18933
rect 18182 18660 18192 18928
rect 18440 18660 18450 18928
rect 18182 18655 18450 18660
rect 20770 18100 21170 18105
rect 20770 17740 20780 18100
rect 21160 17740 21170 18100
rect 20770 17735 21170 17740
rect 15166 15824 15358 15829
rect 15166 15716 15176 15824
rect 15348 15716 15358 15824
rect 15166 15711 15358 15716
rect -1200 12300 13840 12920
rect 19530 12740 19540 13120
rect 20000 12740 20010 13120
rect -1220 12080 16700 12300
rect -1220 11080 -260 12080
rect 3640 11620 16700 12080
rect 21812 11620 23020 18996
rect 3640 11480 24180 11620
rect -1220 10440 2400 11080
rect 11900 10440 15700 11120
rect 24020 10440 24180 11480
rect -1220 10280 24180 10440
rect 23800 9040 24800 9100
rect 23800 8660 24340 9040
rect 24330 8620 24340 8660
rect 24760 8660 24800 9040
rect 24760 8620 24770 8660
rect 24330 8615 24770 8620
rect 24330 8160 24770 8165
rect 24330 7740 24340 8160
rect 24760 7740 24770 8160
rect 24330 7735 24770 7740
rect 25210 8160 25650 8165
rect 25210 7740 25220 8160
rect 25640 7740 25650 8160
rect 25210 7735 25650 7740
rect 24980 6380 25560 6860
rect 24300 6360 25560 6380
rect 24300 6120 24320 6360
rect 24500 6340 25560 6360
rect 24500 6120 24980 6340
rect 24300 6100 24980 6120
rect 24350 5800 24590 5805
rect 24350 5700 24360 5800
rect 24580 5700 24590 5800
rect 24350 5695 24590 5700
rect 14990 4440 15140 4445
rect 1650 4420 1850 4425
rect 1650 4340 1660 4420
rect 1840 4340 1850 4420
rect 1650 4335 1850 4340
rect 14990 4320 15000 4440
rect 15130 4320 15140 4440
rect 14990 4315 15140 4320
rect -3250 -3680 -3240 -1280
rect 25320 -3680 25330 -1280
<< via3 >>
rect 17232 18656 17480 18924
rect 18192 18660 18440 18928
rect 19540 12740 20000 13120
rect 24340 8620 24760 9040
rect 24340 7740 24760 8160
rect 25220 7740 25640 8160
rect 24360 5700 24580 5800
rect -3240 -3680 25320 -1280
<< metal4 >>
rect 17480 18860 17520 18940
rect 18160 18928 18200 18940
rect 18160 18860 18192 18928
rect 17480 18680 18192 18860
rect 17480 18620 17520 18680
rect 18160 18660 18192 18680
rect 18160 18620 18200 18660
rect 11100 13140 18756 13760
rect 11100 13120 20040 13140
rect 11100 13012 19540 13120
rect 11096 12800 19540 13012
rect 11096 12664 14804 12800
rect 15192 12740 19540 12800
rect 20000 12740 20040 13120
rect 15192 12720 20040 12740
rect 15192 12664 18756 12720
rect 11096 12504 18756 12664
rect 11096 12500 16052 12504
rect 11096 12496 12280 12500
rect 12600 12496 13692 12500
rect 12600 10420 13560 12496
rect 24340 8500 24760 8580
rect 24340 8200 24760 8280
rect 24800 7740 24880 8160
rect 25100 7740 25180 8160
rect 24480 5801 25400 6040
rect 24359 5800 25400 5801
rect 24359 5700 24360 5800
rect 24580 5700 25400 5800
rect 24359 5699 25400 5700
rect -1700 -200 -1300 200
rect 24480 -200 25400 5699
rect -3628 -1280 25400 -200
rect -3628 -3680 -3240 -1280
rect 25320 -3680 25400 -1280
rect -3628 -4080 25400 -3680
<< via4 >>
rect 16980 18924 17480 19040
rect 16980 18656 17232 18924
rect 17232 18656 17480 18924
rect 18200 18928 18700 19040
rect 16980 18540 17480 18656
rect 18200 18660 18440 18928
rect 18440 18660 18700 18928
rect 18200 18540 18700 18660
rect 24300 9040 24800 9080
rect 24300 8620 24340 9040
rect 24340 8620 24760 9040
rect 24760 8620 24800 9040
rect 24300 8580 24800 8620
rect 24300 8160 24800 8200
rect 25180 8160 25680 8200
rect 24300 7740 24340 8160
rect 24340 7740 24760 8160
rect 24760 7740 24800 8160
rect 25180 7740 25220 8160
rect 25220 7740 25640 8160
rect 25640 7740 25680 8160
rect 24300 7700 24800 7740
rect 25180 7700 25680 7740
<< metal5 >>
rect 16956 19040 17504 19064
rect 16956 18540 16980 19040
rect 17480 18540 17504 19040
rect 16956 18516 17504 18540
rect 18176 19040 18724 19064
rect 18176 18540 18200 19040
rect 18700 18540 18724 19040
rect 18176 18516 18724 18540
rect 24276 9080 24824 9104
rect 24276 8580 24300 9080
rect 24800 8580 24824 9080
rect 24276 8556 24824 8580
rect 24276 8200 24824 8224
rect 24276 7700 24300 8200
rect 24800 7700 24824 8200
rect 24276 7676 24824 7700
rect 25156 8200 25704 8224
rect 25156 7700 25180 8200
rect 25680 7700 25704 8200
rect 25156 7676 25704 7700
use curr_filter  curr_filter_0
timestamp 1686659968
transform 1 0 -4440 0 1 -255
box 1140 -145 3180 8460
use sky130_fd_pr__cap_mim_m3_1_65KGHP  sky130_fd_pr__cap_mim_m3_1_65KGHP_0
timestamp 1685031707
transform 0 -1 24920 1 0 6466
box -686 -240 686 240
use sky130_fd_pr__res_xhigh_po_0p69_L5PD5X  sky130_fd_pr__res_xhigh_po_0p69_L5PD5X_0
timestamp 1685031707
transform 1 0 24535 0 1 6958
box -235 -1198 235 1198
use tia_bias  tia_bias_1
timestamp 1686659968
transform 1 0 10920 0 1 19376
box -120 -6836 10684 4104
use tia_core  tia_core_0
timestamp 1686659968
transform 1 0 16764 0 1 8240
box -4564 -9640 8480 3244
use tia_core  tia_core_1
timestamp 1686659968
transform 1 0 3364 0 1 8240
box -4564 -9640 8480 3244
use tia_outfilter  tia_outfilter_0
timestamp 1686659968
transform 1 0 19416 0 1 14810
box -2364 -3030 1784 4366
<< labels >>
rlabel metal1 25260 8460 25420 8660 1 Filter_out_1
port 1 n
rlabel metal4 24380 8240 24700 8260 1 Filter_in_2
port 3 n
rlabel metal3 24140 8780 24200 9040 1 Out_2
port 2 n
rlabel metal4 -2980 -2820 -2320 -2080 1 VN
port 4 n
rlabel metal2 7220 8840 7540 9060 1 Input_ref
port 5 n
rlabel metal2 20620 8860 20940 9080 1 Input
port 6 n
rlabel metal2 -1060 10880 -860 11260 1 VP
port 7 n
rlabel metal2 -3028 8212 -2816 8244 1 I_Bias1
port 8 n
rlabel metal3 25280 6380 25520 6800 1 Ref_out
port 9 n
<< end >>
