magic
tech sky130A
magscale 1 2
timestamp 1683557511
<< nwell >>
rect -11173 2281 -6907 3463
rect -6653 2281 -2387 3463
rect -2133 2281 2133 3463
rect 2387 2281 6653 3463
rect 6907 2281 11173 3463
rect -11173 845 -6907 2027
rect -6653 845 -2387 2027
rect -2133 845 2133 2027
rect 2387 845 6653 2027
rect 6907 845 11173 2027
rect -11173 -591 -6907 591
rect -6653 -591 -2387 591
rect -2133 -591 2133 591
rect 2387 -591 6653 591
rect 6907 -591 11173 591
rect -11173 -2027 -6907 -845
rect -6653 -2027 -2387 -845
rect -2133 -2027 2133 -845
rect 2387 -2027 6653 -845
rect 6907 -2027 11173 -845
rect -11173 -3463 -6907 -2281
rect -6653 -3463 -2387 -2281
rect -2133 -3463 2133 -2281
rect 2387 -3463 6653 -2281
rect 6907 -3463 11173 -2281
<< pwell >>
rect -11283 3463 11283 3573
rect -11283 2281 -11173 3463
rect -6907 2281 -6653 3463
rect -2387 2281 -2133 3463
rect 2133 2281 2387 3463
rect 6653 2281 6907 3463
rect 11173 2281 11283 3463
rect -11283 2027 11283 2281
rect -11283 845 -11173 2027
rect -6907 845 -6653 2027
rect -2387 845 -2133 2027
rect 2133 845 2387 2027
rect 6653 845 6907 2027
rect 11173 845 11283 2027
rect -11283 591 11283 845
rect -11283 -591 -11173 591
rect -6907 -591 -6653 591
rect -2387 -591 -2133 591
rect 2133 -591 2387 591
rect 6653 -591 6907 591
rect 11173 -591 11283 591
rect -11283 -845 11283 -591
rect -11283 -2027 -11173 -845
rect -6907 -2027 -6653 -845
rect -2387 -2027 -2133 -845
rect 2133 -2027 2387 -845
rect 6653 -2027 6907 -845
rect 11173 -2027 11283 -845
rect -11283 -2281 11283 -2027
rect -11283 -3463 -11173 -2281
rect -6907 -3463 -6653 -2281
rect -2387 -3463 -2133 -2281
rect 2133 -3463 2387 -2281
rect 6653 -3463 6907 -2281
rect 11173 -3463 11283 -2281
rect -11283 -3573 11283 -3463
<< varactor >>
rect -11040 2372 -7040 3372
rect -6520 2372 -2520 3372
rect -2000 2372 2000 3372
rect 2520 2372 6520 3372
rect 7040 2372 11040 3372
rect -11040 936 -7040 1936
rect -6520 936 -2520 1936
rect -2000 936 2000 1936
rect 2520 936 6520 1936
rect 7040 936 11040 1936
rect -11040 -500 -7040 500
rect -6520 -500 -2520 500
rect -2000 -500 2000 500
rect 2520 -500 6520 500
rect 7040 -500 11040 500
rect -11040 -1936 -7040 -936
rect -6520 -1936 -2520 -936
rect -2000 -1936 2000 -936
rect 2520 -1936 6520 -936
rect 7040 -1936 11040 -936
rect -11040 -3372 -7040 -2372
rect -6520 -3372 -2520 -2372
rect -2000 -3372 2000 -2372
rect 2520 -3372 6520 -2372
rect 7040 -3372 11040 -2372
<< psubdiff >>
rect -11247 3503 -11151 3537
rect 11151 3503 11247 3537
rect -11247 3441 -11213 3503
rect 11213 3441 11247 3503
rect -11247 -3503 -11213 -3441
rect 11213 -3503 11247 -3441
rect -11247 -3537 -11151 -3503
rect 11151 -3537 11247 -3503
<< nsubdiff >>
rect -11137 3348 -11040 3372
rect -11137 2396 -11125 3348
rect -11091 2396 -11040 3348
rect -11137 2372 -11040 2396
rect -7040 3348 -6943 3372
rect -7040 2396 -6989 3348
rect -6955 2396 -6943 3348
rect -7040 2372 -6943 2396
rect -6617 3348 -6520 3372
rect -6617 2396 -6605 3348
rect -6571 2396 -6520 3348
rect -6617 2372 -6520 2396
rect -2520 3348 -2423 3372
rect -2520 2396 -2469 3348
rect -2435 2396 -2423 3348
rect -2520 2372 -2423 2396
rect -2097 3348 -2000 3372
rect -2097 2396 -2085 3348
rect -2051 2396 -2000 3348
rect -2097 2372 -2000 2396
rect 2000 3348 2097 3372
rect 2000 2396 2051 3348
rect 2085 2396 2097 3348
rect 2000 2372 2097 2396
rect 2423 3348 2520 3372
rect 2423 2396 2435 3348
rect 2469 2396 2520 3348
rect 2423 2372 2520 2396
rect 6520 3348 6617 3372
rect 6520 2396 6571 3348
rect 6605 2396 6617 3348
rect 6520 2372 6617 2396
rect 6943 3348 7040 3372
rect 6943 2396 6955 3348
rect 6989 2396 7040 3348
rect 6943 2372 7040 2396
rect 11040 3348 11137 3372
rect 11040 2396 11091 3348
rect 11125 2396 11137 3348
rect 11040 2372 11137 2396
rect -11137 1912 -11040 1936
rect -11137 960 -11125 1912
rect -11091 960 -11040 1912
rect -11137 936 -11040 960
rect -7040 1912 -6943 1936
rect -7040 960 -6989 1912
rect -6955 960 -6943 1912
rect -7040 936 -6943 960
rect -6617 1912 -6520 1936
rect -6617 960 -6605 1912
rect -6571 960 -6520 1912
rect -6617 936 -6520 960
rect -2520 1912 -2423 1936
rect -2520 960 -2469 1912
rect -2435 960 -2423 1912
rect -2520 936 -2423 960
rect -2097 1912 -2000 1936
rect -2097 960 -2085 1912
rect -2051 960 -2000 1912
rect -2097 936 -2000 960
rect 2000 1912 2097 1936
rect 2000 960 2051 1912
rect 2085 960 2097 1912
rect 2000 936 2097 960
rect 2423 1912 2520 1936
rect 2423 960 2435 1912
rect 2469 960 2520 1912
rect 2423 936 2520 960
rect 6520 1912 6617 1936
rect 6520 960 6571 1912
rect 6605 960 6617 1912
rect 6520 936 6617 960
rect 6943 1912 7040 1936
rect 6943 960 6955 1912
rect 6989 960 7040 1912
rect 6943 936 7040 960
rect 11040 1912 11137 1936
rect 11040 960 11091 1912
rect 11125 960 11137 1912
rect 11040 936 11137 960
rect -11137 476 -11040 500
rect -11137 -476 -11125 476
rect -11091 -476 -11040 476
rect -11137 -500 -11040 -476
rect -7040 476 -6943 500
rect -7040 -476 -6989 476
rect -6955 -476 -6943 476
rect -7040 -500 -6943 -476
rect -6617 476 -6520 500
rect -6617 -476 -6605 476
rect -6571 -476 -6520 476
rect -6617 -500 -6520 -476
rect -2520 476 -2423 500
rect -2520 -476 -2469 476
rect -2435 -476 -2423 476
rect -2520 -500 -2423 -476
rect -2097 476 -2000 500
rect -2097 -476 -2085 476
rect -2051 -476 -2000 476
rect -2097 -500 -2000 -476
rect 2000 476 2097 500
rect 2000 -476 2051 476
rect 2085 -476 2097 476
rect 2000 -500 2097 -476
rect 2423 476 2520 500
rect 2423 -476 2435 476
rect 2469 -476 2520 476
rect 2423 -500 2520 -476
rect 6520 476 6617 500
rect 6520 -476 6571 476
rect 6605 -476 6617 476
rect 6520 -500 6617 -476
rect 6943 476 7040 500
rect 6943 -476 6955 476
rect 6989 -476 7040 476
rect 6943 -500 7040 -476
rect 11040 476 11137 500
rect 11040 -476 11091 476
rect 11125 -476 11137 476
rect 11040 -500 11137 -476
rect -11137 -960 -11040 -936
rect -11137 -1912 -11125 -960
rect -11091 -1912 -11040 -960
rect -11137 -1936 -11040 -1912
rect -7040 -960 -6943 -936
rect -7040 -1912 -6989 -960
rect -6955 -1912 -6943 -960
rect -7040 -1936 -6943 -1912
rect -6617 -960 -6520 -936
rect -6617 -1912 -6605 -960
rect -6571 -1912 -6520 -960
rect -6617 -1936 -6520 -1912
rect -2520 -960 -2423 -936
rect -2520 -1912 -2469 -960
rect -2435 -1912 -2423 -960
rect -2520 -1936 -2423 -1912
rect -2097 -960 -2000 -936
rect -2097 -1912 -2085 -960
rect -2051 -1912 -2000 -960
rect -2097 -1936 -2000 -1912
rect 2000 -960 2097 -936
rect 2000 -1912 2051 -960
rect 2085 -1912 2097 -960
rect 2000 -1936 2097 -1912
rect 2423 -960 2520 -936
rect 2423 -1912 2435 -960
rect 2469 -1912 2520 -960
rect 2423 -1936 2520 -1912
rect 6520 -960 6617 -936
rect 6520 -1912 6571 -960
rect 6605 -1912 6617 -960
rect 6520 -1936 6617 -1912
rect 6943 -960 7040 -936
rect 6943 -1912 6955 -960
rect 6989 -1912 7040 -960
rect 6943 -1936 7040 -1912
rect 11040 -960 11137 -936
rect 11040 -1912 11091 -960
rect 11125 -1912 11137 -960
rect 11040 -1936 11137 -1912
rect -11137 -2396 -11040 -2372
rect -11137 -3348 -11125 -2396
rect -11091 -3348 -11040 -2396
rect -11137 -3372 -11040 -3348
rect -7040 -2396 -6943 -2372
rect -7040 -3348 -6989 -2396
rect -6955 -3348 -6943 -2396
rect -7040 -3372 -6943 -3348
rect -6617 -2396 -6520 -2372
rect -6617 -3348 -6605 -2396
rect -6571 -3348 -6520 -2396
rect -6617 -3372 -6520 -3348
rect -2520 -2396 -2423 -2372
rect -2520 -3348 -2469 -2396
rect -2435 -3348 -2423 -2396
rect -2520 -3372 -2423 -3348
rect -2097 -2396 -2000 -2372
rect -2097 -3348 -2085 -2396
rect -2051 -3348 -2000 -2396
rect -2097 -3372 -2000 -3348
rect 2000 -2396 2097 -2372
rect 2000 -3348 2051 -2396
rect 2085 -3348 2097 -2396
rect 2000 -3372 2097 -3348
rect 2423 -2396 2520 -2372
rect 2423 -3348 2435 -2396
rect 2469 -3348 2520 -2396
rect 2423 -3372 2520 -3348
rect 6520 -2396 6617 -2372
rect 6520 -3348 6571 -2396
rect 6605 -3348 6617 -2396
rect 6520 -3372 6617 -3348
rect 6943 -2396 7040 -2372
rect 6943 -3348 6955 -2396
rect 6989 -3348 7040 -2396
rect 6943 -3372 7040 -3348
rect 11040 -2396 11137 -2372
rect 11040 -3348 11091 -2396
rect 11125 -3348 11137 -2396
rect 11040 -3372 11137 -3348
<< psubdiffcont >>
rect -11151 3503 11151 3537
rect -11247 -3441 -11213 3441
rect 11213 -3441 11247 3441
rect -11151 -3537 11151 -3503
<< nsubdiffcont >>
rect -11125 2396 -11091 3348
rect -6989 2396 -6955 3348
rect -6605 2396 -6571 3348
rect -2469 2396 -2435 3348
rect -2085 2396 -2051 3348
rect 2051 2396 2085 3348
rect 2435 2396 2469 3348
rect 6571 2396 6605 3348
rect 6955 2396 6989 3348
rect 11091 2396 11125 3348
rect -11125 960 -11091 1912
rect -6989 960 -6955 1912
rect -6605 960 -6571 1912
rect -2469 960 -2435 1912
rect -2085 960 -2051 1912
rect 2051 960 2085 1912
rect 2435 960 2469 1912
rect 6571 960 6605 1912
rect 6955 960 6989 1912
rect 11091 960 11125 1912
rect -11125 -476 -11091 476
rect -6989 -476 -6955 476
rect -6605 -476 -6571 476
rect -2469 -476 -2435 476
rect -2085 -476 -2051 476
rect 2051 -476 2085 476
rect 2435 -476 2469 476
rect 6571 -476 6605 476
rect 6955 -476 6989 476
rect 11091 -476 11125 476
rect -11125 -1912 -11091 -960
rect -6989 -1912 -6955 -960
rect -6605 -1912 -6571 -960
rect -2469 -1912 -2435 -960
rect -2085 -1912 -2051 -960
rect 2051 -1912 2085 -960
rect 2435 -1912 2469 -960
rect 6571 -1912 6605 -960
rect 6955 -1912 6989 -960
rect 11091 -1912 11125 -960
rect -11125 -3348 -11091 -2396
rect -6989 -3348 -6955 -2396
rect -6605 -3348 -6571 -2396
rect -2469 -3348 -2435 -2396
rect -2085 -3348 -2051 -2396
rect 2051 -3348 2085 -2396
rect 2435 -3348 2469 -2396
rect 6571 -3348 6605 -2396
rect 6955 -3348 6989 -2396
rect 11091 -3348 11125 -2396
<< poly >>
rect -11040 3444 -7040 3460
rect -11040 3410 -11024 3444
rect -7056 3410 -7040 3444
rect -11040 3372 -7040 3410
rect -6520 3444 -2520 3460
rect -6520 3410 -6504 3444
rect -2536 3410 -2520 3444
rect -6520 3372 -2520 3410
rect -2000 3444 2000 3460
rect -2000 3410 -1984 3444
rect 1984 3410 2000 3444
rect -2000 3372 2000 3410
rect 2520 3444 6520 3460
rect 2520 3410 2536 3444
rect 6504 3410 6520 3444
rect 2520 3372 6520 3410
rect 7040 3444 11040 3460
rect 7040 3410 7056 3444
rect 11024 3410 11040 3444
rect 7040 3372 11040 3410
rect -11040 2334 -7040 2372
rect -11040 2300 -11024 2334
rect -7056 2300 -7040 2334
rect -11040 2284 -7040 2300
rect -6520 2334 -2520 2372
rect -6520 2300 -6504 2334
rect -2536 2300 -2520 2334
rect -6520 2284 -2520 2300
rect -2000 2334 2000 2372
rect -2000 2300 -1984 2334
rect 1984 2300 2000 2334
rect -2000 2284 2000 2300
rect 2520 2334 6520 2372
rect 2520 2300 2536 2334
rect 6504 2300 6520 2334
rect 2520 2284 6520 2300
rect 7040 2334 11040 2372
rect 7040 2300 7056 2334
rect 11024 2300 11040 2334
rect 7040 2284 11040 2300
rect -11040 2008 -7040 2024
rect -11040 1974 -11024 2008
rect -7056 1974 -7040 2008
rect -11040 1936 -7040 1974
rect -6520 2008 -2520 2024
rect -6520 1974 -6504 2008
rect -2536 1974 -2520 2008
rect -6520 1936 -2520 1974
rect -2000 2008 2000 2024
rect -2000 1974 -1984 2008
rect 1984 1974 2000 2008
rect -2000 1936 2000 1974
rect 2520 2008 6520 2024
rect 2520 1974 2536 2008
rect 6504 1974 6520 2008
rect 2520 1936 6520 1974
rect 7040 2008 11040 2024
rect 7040 1974 7056 2008
rect 11024 1974 11040 2008
rect 7040 1936 11040 1974
rect -11040 898 -7040 936
rect -11040 864 -11024 898
rect -7056 864 -7040 898
rect -11040 848 -7040 864
rect -6520 898 -2520 936
rect -6520 864 -6504 898
rect -2536 864 -2520 898
rect -6520 848 -2520 864
rect -2000 898 2000 936
rect -2000 864 -1984 898
rect 1984 864 2000 898
rect -2000 848 2000 864
rect 2520 898 6520 936
rect 2520 864 2536 898
rect 6504 864 6520 898
rect 2520 848 6520 864
rect 7040 898 11040 936
rect 7040 864 7056 898
rect 11024 864 11040 898
rect 7040 848 11040 864
rect -11040 572 -7040 588
rect -11040 538 -11024 572
rect -7056 538 -7040 572
rect -11040 500 -7040 538
rect -6520 572 -2520 588
rect -6520 538 -6504 572
rect -2536 538 -2520 572
rect -6520 500 -2520 538
rect -2000 572 2000 588
rect -2000 538 -1984 572
rect 1984 538 2000 572
rect -2000 500 2000 538
rect 2520 572 6520 588
rect 2520 538 2536 572
rect 6504 538 6520 572
rect 2520 500 6520 538
rect 7040 572 11040 588
rect 7040 538 7056 572
rect 11024 538 11040 572
rect 7040 500 11040 538
rect -11040 -538 -7040 -500
rect -11040 -572 -11024 -538
rect -7056 -572 -7040 -538
rect -11040 -588 -7040 -572
rect -6520 -538 -2520 -500
rect -6520 -572 -6504 -538
rect -2536 -572 -2520 -538
rect -6520 -588 -2520 -572
rect -2000 -538 2000 -500
rect -2000 -572 -1984 -538
rect 1984 -572 2000 -538
rect -2000 -588 2000 -572
rect 2520 -538 6520 -500
rect 2520 -572 2536 -538
rect 6504 -572 6520 -538
rect 2520 -588 6520 -572
rect 7040 -538 11040 -500
rect 7040 -572 7056 -538
rect 11024 -572 11040 -538
rect 7040 -588 11040 -572
rect -11040 -864 -7040 -848
rect -11040 -898 -11024 -864
rect -7056 -898 -7040 -864
rect -11040 -936 -7040 -898
rect -6520 -864 -2520 -848
rect -6520 -898 -6504 -864
rect -2536 -898 -2520 -864
rect -6520 -936 -2520 -898
rect -2000 -864 2000 -848
rect -2000 -898 -1984 -864
rect 1984 -898 2000 -864
rect -2000 -936 2000 -898
rect 2520 -864 6520 -848
rect 2520 -898 2536 -864
rect 6504 -898 6520 -864
rect 2520 -936 6520 -898
rect 7040 -864 11040 -848
rect 7040 -898 7056 -864
rect 11024 -898 11040 -864
rect 7040 -936 11040 -898
rect -11040 -1974 -7040 -1936
rect -11040 -2008 -11024 -1974
rect -7056 -2008 -7040 -1974
rect -11040 -2024 -7040 -2008
rect -6520 -1974 -2520 -1936
rect -6520 -2008 -6504 -1974
rect -2536 -2008 -2520 -1974
rect -6520 -2024 -2520 -2008
rect -2000 -1974 2000 -1936
rect -2000 -2008 -1984 -1974
rect 1984 -2008 2000 -1974
rect -2000 -2024 2000 -2008
rect 2520 -1974 6520 -1936
rect 2520 -2008 2536 -1974
rect 6504 -2008 6520 -1974
rect 2520 -2024 6520 -2008
rect 7040 -1974 11040 -1936
rect 7040 -2008 7056 -1974
rect 11024 -2008 11040 -1974
rect 7040 -2024 11040 -2008
rect -11040 -2300 -7040 -2284
rect -11040 -2334 -11024 -2300
rect -7056 -2334 -7040 -2300
rect -11040 -2372 -7040 -2334
rect -6520 -2300 -2520 -2284
rect -6520 -2334 -6504 -2300
rect -2536 -2334 -2520 -2300
rect -6520 -2372 -2520 -2334
rect -2000 -2300 2000 -2284
rect -2000 -2334 -1984 -2300
rect 1984 -2334 2000 -2300
rect -2000 -2372 2000 -2334
rect 2520 -2300 6520 -2284
rect 2520 -2334 2536 -2300
rect 6504 -2334 6520 -2300
rect 2520 -2372 6520 -2334
rect 7040 -2300 11040 -2284
rect 7040 -2334 7056 -2300
rect 11024 -2334 11040 -2300
rect 7040 -2372 11040 -2334
rect -11040 -3410 -7040 -3372
rect -11040 -3444 -11024 -3410
rect -7056 -3444 -7040 -3410
rect -11040 -3460 -7040 -3444
rect -6520 -3410 -2520 -3372
rect -6520 -3444 -6504 -3410
rect -2536 -3444 -2520 -3410
rect -6520 -3460 -2520 -3444
rect -2000 -3410 2000 -3372
rect -2000 -3444 -1984 -3410
rect 1984 -3444 2000 -3410
rect -2000 -3460 2000 -3444
rect 2520 -3410 6520 -3372
rect 2520 -3444 2536 -3410
rect 6504 -3444 6520 -3410
rect 2520 -3460 6520 -3444
rect 7040 -3410 11040 -3372
rect 7040 -3444 7056 -3410
rect 11024 -3444 11040 -3410
rect 7040 -3460 11040 -3444
<< polycont >>
rect -11024 3410 -7056 3444
rect -6504 3410 -2536 3444
rect -1984 3410 1984 3444
rect 2536 3410 6504 3444
rect 7056 3410 11024 3444
rect -11024 2300 -7056 2334
rect -6504 2300 -2536 2334
rect -1984 2300 1984 2334
rect 2536 2300 6504 2334
rect 7056 2300 11024 2334
rect -11024 1974 -7056 2008
rect -6504 1974 -2536 2008
rect -1984 1974 1984 2008
rect 2536 1974 6504 2008
rect 7056 1974 11024 2008
rect -11024 864 -7056 898
rect -6504 864 -2536 898
rect -1984 864 1984 898
rect 2536 864 6504 898
rect 7056 864 11024 898
rect -11024 538 -7056 572
rect -6504 538 -2536 572
rect -1984 538 1984 572
rect 2536 538 6504 572
rect 7056 538 11024 572
rect -11024 -572 -7056 -538
rect -6504 -572 -2536 -538
rect -1984 -572 1984 -538
rect 2536 -572 6504 -538
rect 7056 -572 11024 -538
rect -11024 -898 -7056 -864
rect -6504 -898 -2536 -864
rect -1984 -898 1984 -864
rect 2536 -898 6504 -864
rect 7056 -898 11024 -864
rect -11024 -2008 -7056 -1974
rect -6504 -2008 -2536 -1974
rect -1984 -2008 1984 -1974
rect 2536 -2008 6504 -1974
rect 7056 -2008 11024 -1974
rect -11024 -2334 -7056 -2300
rect -6504 -2334 -2536 -2300
rect -1984 -2334 1984 -2300
rect 2536 -2334 6504 -2300
rect 7056 -2334 11024 -2300
rect -11024 -3444 -7056 -3410
rect -6504 -3444 -2536 -3410
rect -1984 -3444 1984 -3410
rect 2536 -3444 6504 -3410
rect 7056 -3444 11024 -3410
<< locali >>
rect -11247 3503 -11151 3537
rect 11151 3503 11247 3537
rect -11247 3441 -11213 3503
rect -11040 3410 -11024 3444
rect -7056 3410 -7040 3444
rect -6520 3410 -6504 3444
rect -2536 3410 -2520 3444
rect -2000 3410 -1984 3444
rect 1984 3410 2000 3444
rect 2520 3410 2536 3444
rect 6504 3410 6520 3444
rect 7040 3410 7056 3444
rect 11024 3410 11040 3444
rect 11213 3441 11247 3503
rect -11125 3348 -11091 3364
rect -11125 2380 -11091 2396
rect -6989 3348 -6955 3364
rect -6989 2380 -6955 2396
rect -6605 3348 -6571 3364
rect -6605 2380 -6571 2396
rect -2469 3348 -2435 3364
rect -2469 2380 -2435 2396
rect -2085 3348 -2051 3364
rect -2085 2380 -2051 2396
rect 2051 3348 2085 3364
rect 2051 2380 2085 2396
rect 2435 3348 2469 3364
rect 2435 2380 2469 2396
rect 6571 3348 6605 3364
rect 6571 2380 6605 2396
rect 6955 3348 6989 3364
rect 6955 2380 6989 2396
rect 11091 3348 11125 3364
rect 11091 2380 11125 2396
rect -11040 2300 -11024 2334
rect -7056 2300 -7040 2334
rect -6520 2300 -6504 2334
rect -2536 2300 -2520 2334
rect -2000 2300 -1984 2334
rect 1984 2300 2000 2334
rect 2520 2300 2536 2334
rect 6504 2300 6520 2334
rect 7040 2300 7056 2334
rect 11024 2300 11040 2334
rect -11040 1974 -11024 2008
rect -7056 1974 -7040 2008
rect -6520 1974 -6504 2008
rect -2536 1974 -2520 2008
rect -2000 1974 -1984 2008
rect 1984 1974 2000 2008
rect 2520 1974 2536 2008
rect 6504 1974 6520 2008
rect 7040 1974 7056 2008
rect 11024 1974 11040 2008
rect -11125 1912 -11091 1928
rect -11125 944 -11091 960
rect -6989 1912 -6955 1928
rect -6989 944 -6955 960
rect -6605 1912 -6571 1928
rect -6605 944 -6571 960
rect -2469 1912 -2435 1928
rect -2469 944 -2435 960
rect -2085 1912 -2051 1928
rect -2085 944 -2051 960
rect 2051 1912 2085 1928
rect 2051 944 2085 960
rect 2435 1912 2469 1928
rect 2435 944 2469 960
rect 6571 1912 6605 1928
rect 6571 944 6605 960
rect 6955 1912 6989 1928
rect 6955 944 6989 960
rect 11091 1912 11125 1928
rect 11091 944 11125 960
rect -11040 864 -11024 898
rect -7056 864 -7040 898
rect -6520 864 -6504 898
rect -2536 864 -2520 898
rect -2000 864 -1984 898
rect 1984 864 2000 898
rect 2520 864 2536 898
rect 6504 864 6520 898
rect 7040 864 7056 898
rect 11024 864 11040 898
rect -11040 538 -11024 572
rect -7056 538 -7040 572
rect -6520 538 -6504 572
rect -2536 538 -2520 572
rect -2000 538 -1984 572
rect 1984 538 2000 572
rect 2520 538 2536 572
rect 6504 538 6520 572
rect 7040 538 7056 572
rect 11024 538 11040 572
rect -11125 476 -11091 492
rect -11125 -492 -11091 -476
rect -6989 476 -6955 492
rect -6989 -492 -6955 -476
rect -6605 476 -6571 492
rect -6605 -492 -6571 -476
rect -2469 476 -2435 492
rect -2469 -492 -2435 -476
rect -2085 476 -2051 492
rect -2085 -492 -2051 -476
rect 2051 476 2085 492
rect 2051 -492 2085 -476
rect 2435 476 2469 492
rect 2435 -492 2469 -476
rect 6571 476 6605 492
rect 6571 -492 6605 -476
rect 6955 476 6989 492
rect 6955 -492 6989 -476
rect 11091 476 11125 492
rect 11091 -492 11125 -476
rect -11040 -572 -11024 -538
rect -7056 -572 -7040 -538
rect -6520 -572 -6504 -538
rect -2536 -572 -2520 -538
rect -2000 -572 -1984 -538
rect 1984 -572 2000 -538
rect 2520 -572 2536 -538
rect 6504 -572 6520 -538
rect 7040 -572 7056 -538
rect 11024 -572 11040 -538
rect -11040 -898 -11024 -864
rect -7056 -898 -7040 -864
rect -6520 -898 -6504 -864
rect -2536 -898 -2520 -864
rect -2000 -898 -1984 -864
rect 1984 -898 2000 -864
rect 2520 -898 2536 -864
rect 6504 -898 6520 -864
rect 7040 -898 7056 -864
rect 11024 -898 11040 -864
rect -11125 -960 -11091 -944
rect -11125 -1928 -11091 -1912
rect -6989 -960 -6955 -944
rect -6989 -1928 -6955 -1912
rect -6605 -960 -6571 -944
rect -6605 -1928 -6571 -1912
rect -2469 -960 -2435 -944
rect -2469 -1928 -2435 -1912
rect -2085 -960 -2051 -944
rect -2085 -1928 -2051 -1912
rect 2051 -960 2085 -944
rect 2051 -1928 2085 -1912
rect 2435 -960 2469 -944
rect 2435 -1928 2469 -1912
rect 6571 -960 6605 -944
rect 6571 -1928 6605 -1912
rect 6955 -960 6989 -944
rect 6955 -1928 6989 -1912
rect 11091 -960 11125 -944
rect 11091 -1928 11125 -1912
rect -11040 -2008 -11024 -1974
rect -7056 -2008 -7040 -1974
rect -6520 -2008 -6504 -1974
rect -2536 -2008 -2520 -1974
rect -2000 -2008 -1984 -1974
rect 1984 -2008 2000 -1974
rect 2520 -2008 2536 -1974
rect 6504 -2008 6520 -1974
rect 7040 -2008 7056 -1974
rect 11024 -2008 11040 -1974
rect -11040 -2334 -11024 -2300
rect -7056 -2334 -7040 -2300
rect -6520 -2334 -6504 -2300
rect -2536 -2334 -2520 -2300
rect -2000 -2334 -1984 -2300
rect 1984 -2334 2000 -2300
rect 2520 -2334 2536 -2300
rect 6504 -2334 6520 -2300
rect 7040 -2334 7056 -2300
rect 11024 -2334 11040 -2300
rect -11125 -2396 -11091 -2380
rect -11125 -3364 -11091 -3348
rect -6989 -2396 -6955 -2380
rect -6989 -3364 -6955 -3348
rect -6605 -2396 -6571 -2380
rect -6605 -3364 -6571 -3348
rect -2469 -2396 -2435 -2380
rect -2469 -3364 -2435 -3348
rect -2085 -2396 -2051 -2380
rect -2085 -3364 -2051 -3348
rect 2051 -2396 2085 -2380
rect 2051 -3364 2085 -3348
rect 2435 -2396 2469 -2380
rect 2435 -3364 2469 -3348
rect 6571 -2396 6605 -2380
rect 6571 -3364 6605 -3348
rect 6955 -2396 6989 -2380
rect 6955 -3364 6989 -3348
rect 11091 -2396 11125 -2380
rect 11091 -3364 11125 -3348
rect -11247 -3503 -11213 -3441
rect -11040 -3444 -11024 -3410
rect -7056 -3444 -7040 -3410
rect -6520 -3444 -6504 -3410
rect -2536 -3444 -2520 -3410
rect -2000 -3444 -1984 -3410
rect 1984 -3444 2000 -3410
rect 2520 -3444 2536 -3410
rect 6504 -3444 6520 -3410
rect 7040 -3444 7056 -3410
rect 11024 -3444 11040 -3410
rect 11213 -3503 11247 -3441
rect -11247 -3537 -11151 -3503
rect 11151 -3537 11247 -3503
<< viali >>
rect -11024 3410 -7056 3444
rect -6504 3410 -2536 3444
rect -1984 3410 1984 3444
rect 2536 3410 6504 3444
rect 7056 3410 11024 3444
rect -11125 2396 -11091 3348
rect -6989 2396 -6955 3348
rect -6605 2396 -6571 3348
rect -2469 2396 -2435 3348
rect -2085 2396 -2051 3348
rect 2051 2396 2085 3348
rect 2435 2396 2469 3348
rect 6571 2396 6605 3348
rect 6955 2396 6989 3348
rect 11091 2396 11125 3348
rect -11024 2300 -7056 2334
rect -6504 2300 -2536 2334
rect -1984 2300 1984 2334
rect 2536 2300 6504 2334
rect 7056 2300 11024 2334
rect -11024 1974 -7056 2008
rect -6504 1974 -2536 2008
rect -1984 1974 1984 2008
rect 2536 1974 6504 2008
rect 7056 1974 11024 2008
rect -11125 960 -11091 1912
rect -6989 960 -6955 1912
rect -6605 960 -6571 1912
rect -2469 960 -2435 1912
rect -2085 960 -2051 1912
rect 2051 960 2085 1912
rect 2435 960 2469 1912
rect 6571 960 6605 1912
rect 6955 960 6989 1912
rect 11091 960 11125 1912
rect -11024 864 -7056 898
rect -6504 864 -2536 898
rect -1984 864 1984 898
rect 2536 864 6504 898
rect 7056 864 11024 898
rect -11024 538 -7056 572
rect -6504 538 -2536 572
rect -1984 538 1984 572
rect 2536 538 6504 572
rect 7056 538 11024 572
rect -11125 -476 -11091 476
rect -6989 -476 -6955 476
rect -6605 -476 -6571 476
rect -2469 -476 -2435 476
rect -2085 -476 -2051 476
rect 2051 -476 2085 476
rect 2435 -476 2469 476
rect 6571 -476 6605 476
rect 6955 -476 6989 476
rect 11091 -476 11125 476
rect -11024 -572 -7056 -538
rect -6504 -572 -2536 -538
rect -1984 -572 1984 -538
rect 2536 -572 6504 -538
rect 7056 -572 11024 -538
rect -11024 -898 -7056 -864
rect -6504 -898 -2536 -864
rect -1984 -898 1984 -864
rect 2536 -898 6504 -864
rect 7056 -898 11024 -864
rect -11125 -1912 -11091 -960
rect -6989 -1912 -6955 -960
rect -6605 -1912 -6571 -960
rect -2469 -1912 -2435 -960
rect -2085 -1912 -2051 -960
rect 2051 -1912 2085 -960
rect 2435 -1912 2469 -960
rect 6571 -1912 6605 -960
rect 6955 -1912 6989 -960
rect 11091 -1912 11125 -960
rect -11024 -2008 -7056 -1974
rect -6504 -2008 -2536 -1974
rect -1984 -2008 1984 -1974
rect 2536 -2008 6504 -1974
rect 7056 -2008 11024 -1974
rect -11024 -2334 -7056 -2300
rect -6504 -2334 -2536 -2300
rect -1984 -2334 1984 -2300
rect 2536 -2334 6504 -2300
rect 7056 -2334 11024 -2300
rect -11125 -3348 -11091 -2396
rect -6989 -3348 -6955 -2396
rect -6605 -3348 -6571 -2396
rect -2469 -3348 -2435 -2396
rect -2085 -3348 -2051 -2396
rect 2051 -3348 2085 -2396
rect 2435 -3348 2469 -2396
rect 6571 -3348 6605 -2396
rect 6955 -3348 6989 -2396
rect 11091 -3348 11125 -2396
rect -11024 -3444 -7056 -3410
rect -6504 -3444 -2536 -3410
rect -1984 -3444 1984 -3410
rect 2536 -3444 6504 -3410
rect 7056 -3444 11024 -3410
<< metal1 >>
rect -11036 3444 -7044 3450
rect -11036 3410 -11024 3444
rect -7056 3410 -7044 3444
rect -11036 3404 -7044 3410
rect -6516 3444 -2524 3450
rect -6516 3410 -6504 3444
rect -2536 3410 -2524 3444
rect -6516 3404 -2524 3410
rect -1996 3444 1996 3450
rect -1996 3410 -1984 3444
rect 1984 3410 1996 3444
rect -1996 3404 1996 3410
rect 2524 3444 6516 3450
rect 2524 3410 2536 3444
rect 6504 3410 6516 3444
rect 2524 3404 6516 3410
rect 7044 3444 11036 3450
rect 7044 3410 7056 3444
rect 11024 3410 11036 3444
rect 7044 3404 11036 3410
rect -11131 3348 -11085 3360
rect -6995 3348 -6949 3360
rect -11131 2396 -11125 3348
rect -11091 2396 -6989 3348
rect -6955 2396 -6949 3348
rect -11131 2384 -11085 2396
rect -6995 2384 -6949 2396
rect -6611 3348 -6565 3360
rect -2475 3348 -2429 3360
rect -6611 2396 -6605 3348
rect -6571 2396 -2469 3348
rect -2435 2396 -2429 3348
rect -6611 2384 -6565 2396
rect -2475 2384 -2429 2396
rect -2091 3348 -2045 3360
rect 2045 3348 2091 3360
rect -2091 2396 -2085 3348
rect -2051 2396 2051 3348
rect 2085 2396 2091 3348
rect -2091 2384 -2045 2396
rect 2045 2384 2091 2396
rect 2429 3348 2475 3360
rect 6565 3348 6611 3360
rect 2429 2396 2435 3348
rect 2469 2396 6571 3348
rect 6605 2396 6611 3348
rect 2429 2384 2475 2396
rect 6565 2384 6611 2396
rect 6949 3348 6995 3360
rect 11085 3348 11131 3360
rect 6949 2396 6955 3348
rect 6989 2396 11091 3348
rect 11125 2396 11131 3348
rect 6949 2384 6995 2396
rect 11085 2384 11131 2396
rect -11036 2334 -7044 2340
rect -11036 2300 -11024 2334
rect -7056 2300 -7044 2334
rect -11036 2294 -7044 2300
rect -6516 2334 -2524 2340
rect -6516 2300 -6504 2334
rect -2536 2300 -2524 2334
rect -6516 2294 -2524 2300
rect -1996 2334 1996 2340
rect -1996 2300 -1984 2334
rect 1984 2300 1996 2334
rect -1996 2294 1996 2300
rect 2524 2334 6516 2340
rect 2524 2300 2536 2334
rect 6504 2300 6516 2334
rect 2524 2294 6516 2300
rect 7044 2334 11036 2340
rect 7044 2300 7056 2334
rect 11024 2300 11036 2334
rect 7044 2294 11036 2300
rect -11036 2008 -7044 2014
rect -11036 1974 -11024 2008
rect -7056 1974 -7044 2008
rect -11036 1968 -7044 1974
rect -6516 2008 -2524 2014
rect -6516 1974 -6504 2008
rect -2536 1974 -2524 2008
rect -6516 1968 -2524 1974
rect -1996 2008 1996 2014
rect -1996 1974 -1984 2008
rect 1984 1974 1996 2008
rect -1996 1968 1996 1974
rect 2524 2008 6516 2014
rect 2524 1974 2536 2008
rect 6504 1974 6516 2008
rect 2524 1968 6516 1974
rect 7044 2008 11036 2014
rect 7044 1974 7056 2008
rect 11024 1974 11036 2008
rect 7044 1968 11036 1974
rect -11131 1912 -11085 1924
rect -6995 1912 -6949 1924
rect -11131 960 -11125 1912
rect -11091 960 -6989 1912
rect -6955 960 -6949 1912
rect -11131 948 -11085 960
rect -6995 948 -6949 960
rect -6611 1912 -6565 1924
rect -2475 1912 -2429 1924
rect -6611 960 -6605 1912
rect -6571 960 -2469 1912
rect -2435 960 -2429 1912
rect -6611 948 -6565 960
rect -2475 948 -2429 960
rect -2091 1912 -2045 1924
rect 2045 1912 2091 1924
rect -2091 960 -2085 1912
rect -2051 960 2051 1912
rect 2085 960 2091 1912
rect -2091 948 -2045 960
rect 2045 948 2091 960
rect 2429 1912 2475 1924
rect 6565 1912 6611 1924
rect 2429 960 2435 1912
rect 2469 960 6571 1912
rect 6605 960 6611 1912
rect 2429 948 2475 960
rect 6565 948 6611 960
rect 6949 1912 6995 1924
rect 11085 1912 11131 1924
rect 6949 960 6955 1912
rect 6989 960 11091 1912
rect 11125 960 11131 1912
rect 6949 948 6995 960
rect 11085 948 11131 960
rect -11036 898 -7044 904
rect -11036 864 -11024 898
rect -7056 864 -7044 898
rect -11036 858 -7044 864
rect -6516 898 -2524 904
rect -6516 864 -6504 898
rect -2536 864 -2524 898
rect -6516 858 -2524 864
rect -1996 898 1996 904
rect -1996 864 -1984 898
rect 1984 864 1996 898
rect -1996 858 1996 864
rect 2524 898 6516 904
rect 2524 864 2536 898
rect 6504 864 6516 898
rect 2524 858 6516 864
rect 7044 898 11036 904
rect 7044 864 7056 898
rect 11024 864 11036 898
rect 7044 858 11036 864
rect -11036 572 -7044 578
rect -11036 538 -11024 572
rect -7056 538 -7044 572
rect -11036 532 -7044 538
rect -6516 572 -2524 578
rect -6516 538 -6504 572
rect -2536 538 -2524 572
rect -6516 532 -2524 538
rect -1996 572 1996 578
rect -1996 538 -1984 572
rect 1984 538 1996 572
rect -1996 532 1996 538
rect 2524 572 6516 578
rect 2524 538 2536 572
rect 6504 538 6516 572
rect 2524 532 6516 538
rect 7044 572 11036 578
rect 7044 538 7056 572
rect 11024 538 11036 572
rect 7044 532 11036 538
rect -11131 476 -11085 488
rect -6995 476 -6949 488
rect -11131 -476 -11125 476
rect -11091 -476 -6989 476
rect -6955 -476 -6949 476
rect -11131 -488 -11085 -476
rect -6995 -488 -6949 -476
rect -6611 476 -6565 488
rect -2475 476 -2429 488
rect -6611 -476 -6605 476
rect -6571 -476 -2469 476
rect -2435 -476 -2429 476
rect -6611 -488 -6565 -476
rect -2475 -488 -2429 -476
rect -2091 476 -2045 488
rect 2045 476 2091 488
rect -2091 -476 -2085 476
rect -2051 -476 2051 476
rect 2085 -476 2091 476
rect -2091 -488 -2045 -476
rect 2045 -488 2091 -476
rect 2429 476 2475 488
rect 6565 476 6611 488
rect 2429 -476 2435 476
rect 2469 -476 6571 476
rect 6605 -476 6611 476
rect 2429 -488 2475 -476
rect 6565 -488 6611 -476
rect 6949 476 6995 488
rect 11085 476 11131 488
rect 6949 -476 6955 476
rect 6989 -476 11091 476
rect 11125 -476 11131 476
rect 6949 -488 6995 -476
rect 11085 -488 11131 -476
rect -11036 -538 -7044 -532
rect -11036 -572 -11024 -538
rect -7056 -572 -7044 -538
rect -11036 -578 -7044 -572
rect -6516 -538 -2524 -532
rect -6516 -572 -6504 -538
rect -2536 -572 -2524 -538
rect -6516 -578 -2524 -572
rect -1996 -538 1996 -532
rect -1996 -572 -1984 -538
rect 1984 -572 1996 -538
rect -1996 -578 1996 -572
rect 2524 -538 6516 -532
rect 2524 -572 2536 -538
rect 6504 -572 6516 -538
rect 2524 -578 6516 -572
rect 7044 -538 11036 -532
rect 7044 -572 7056 -538
rect 11024 -572 11036 -538
rect 7044 -578 11036 -572
rect -11036 -864 -7044 -858
rect -11036 -898 -11024 -864
rect -7056 -898 -7044 -864
rect -11036 -904 -7044 -898
rect -6516 -864 -2524 -858
rect -6516 -898 -6504 -864
rect -2536 -898 -2524 -864
rect -6516 -904 -2524 -898
rect -1996 -864 1996 -858
rect -1996 -898 -1984 -864
rect 1984 -898 1996 -864
rect -1996 -904 1996 -898
rect 2524 -864 6516 -858
rect 2524 -898 2536 -864
rect 6504 -898 6516 -864
rect 2524 -904 6516 -898
rect 7044 -864 11036 -858
rect 7044 -898 7056 -864
rect 11024 -898 11036 -864
rect 7044 -904 11036 -898
rect -11131 -960 -11085 -948
rect -6995 -960 -6949 -948
rect -11131 -1912 -11125 -960
rect -11091 -1912 -6989 -960
rect -6955 -1912 -6949 -960
rect -11131 -1924 -11085 -1912
rect -6995 -1924 -6949 -1912
rect -6611 -960 -6565 -948
rect -2475 -960 -2429 -948
rect -6611 -1912 -6605 -960
rect -6571 -1912 -2469 -960
rect -2435 -1912 -2429 -960
rect -6611 -1924 -6565 -1912
rect -2475 -1924 -2429 -1912
rect -2091 -960 -2045 -948
rect 2045 -960 2091 -948
rect -2091 -1912 -2085 -960
rect -2051 -1912 2051 -960
rect 2085 -1912 2091 -960
rect -2091 -1924 -2045 -1912
rect 2045 -1924 2091 -1912
rect 2429 -960 2475 -948
rect 6565 -960 6611 -948
rect 2429 -1912 2435 -960
rect 2469 -1912 6571 -960
rect 6605 -1912 6611 -960
rect 2429 -1924 2475 -1912
rect 6565 -1924 6611 -1912
rect 6949 -960 6995 -948
rect 11085 -960 11131 -948
rect 6949 -1912 6955 -960
rect 6989 -1912 11091 -960
rect 11125 -1912 11131 -960
rect 6949 -1924 6995 -1912
rect 11085 -1924 11131 -1912
rect -11036 -1974 -7044 -1968
rect -11036 -2008 -11024 -1974
rect -7056 -2008 -7044 -1974
rect -11036 -2014 -7044 -2008
rect -6516 -1974 -2524 -1968
rect -6516 -2008 -6504 -1974
rect -2536 -2008 -2524 -1974
rect -6516 -2014 -2524 -2008
rect -1996 -1974 1996 -1968
rect -1996 -2008 -1984 -1974
rect 1984 -2008 1996 -1974
rect -1996 -2014 1996 -2008
rect 2524 -1974 6516 -1968
rect 2524 -2008 2536 -1974
rect 6504 -2008 6516 -1974
rect 2524 -2014 6516 -2008
rect 7044 -1974 11036 -1968
rect 7044 -2008 7056 -1974
rect 11024 -2008 11036 -1974
rect 7044 -2014 11036 -2008
rect -11036 -2300 -7044 -2294
rect -11036 -2334 -11024 -2300
rect -7056 -2334 -7044 -2300
rect -11036 -2340 -7044 -2334
rect -6516 -2300 -2524 -2294
rect -6516 -2334 -6504 -2300
rect -2536 -2334 -2524 -2300
rect -6516 -2340 -2524 -2334
rect -1996 -2300 1996 -2294
rect -1996 -2334 -1984 -2300
rect 1984 -2334 1996 -2300
rect -1996 -2340 1996 -2334
rect 2524 -2300 6516 -2294
rect 2524 -2334 2536 -2300
rect 6504 -2334 6516 -2300
rect 2524 -2340 6516 -2334
rect 7044 -2300 11036 -2294
rect 7044 -2334 7056 -2300
rect 11024 -2334 11036 -2300
rect 7044 -2340 11036 -2334
rect -11131 -2396 -11085 -2384
rect -6995 -2396 -6949 -2384
rect -11131 -3348 -11125 -2396
rect -11091 -3348 -6989 -2396
rect -6955 -3348 -6949 -2396
rect -11131 -3360 -11085 -3348
rect -6995 -3360 -6949 -3348
rect -6611 -2396 -6565 -2384
rect -2475 -2396 -2429 -2384
rect -6611 -3348 -6605 -2396
rect -6571 -3348 -2469 -2396
rect -2435 -3348 -2429 -2396
rect -6611 -3360 -6565 -3348
rect -2475 -3360 -2429 -3348
rect -2091 -2396 -2045 -2384
rect 2045 -2396 2091 -2384
rect -2091 -3348 -2085 -2396
rect -2051 -3348 2051 -2396
rect 2085 -3348 2091 -2396
rect -2091 -3360 -2045 -3348
rect 2045 -3360 2091 -3348
rect 2429 -2396 2475 -2384
rect 6565 -2396 6611 -2384
rect 2429 -3348 2435 -2396
rect 2469 -3348 6571 -2396
rect 6605 -3348 6611 -2396
rect 2429 -3360 2475 -3348
rect 6565 -3360 6611 -3348
rect 6949 -2396 6995 -2384
rect 11085 -2396 11131 -2384
rect 6949 -3348 6955 -2396
rect 6989 -3348 11091 -2396
rect 11125 -3348 11131 -2396
rect 6949 -3360 6995 -3348
rect 11085 -3360 11131 -3348
rect -11036 -3410 -7044 -3404
rect -11036 -3444 -11024 -3410
rect -7056 -3444 -7044 -3410
rect -11036 -3450 -7044 -3444
rect -6516 -3410 -2524 -3404
rect -6516 -3444 -6504 -3410
rect -2536 -3444 -2524 -3410
rect -6516 -3450 -2524 -3444
rect -1996 -3410 1996 -3404
rect -1996 -3444 -1984 -3410
rect 1984 -3444 1996 -3410
rect -1996 -3450 1996 -3444
rect 2524 -3410 6516 -3404
rect 2524 -3444 2536 -3410
rect 6504 -3444 6516 -3410
rect 2524 -3450 6516 -3444
rect 7044 -3410 11036 -3404
rect 7044 -3444 7056 -3410
rect 11024 -3444 11036 -3410
rect 7044 -3450 11036 -3444
<< properties >>
string FIXED_BBOX -11230 -3520 11230 3520
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5 l 20 m 5 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
