magic
tech sky130A
magscale 1 2
timestamp 1684929745
<< pwell >>
rect -874 -1482 874 1482
<< psubdiff >>
rect -838 1412 -742 1446
rect 742 1412 838 1446
rect -838 1350 -804 1412
rect 804 1350 838 1412
rect -838 -1412 -804 -1350
rect 804 -1412 838 -1350
rect -838 -1446 -742 -1412
rect 742 -1446 838 -1412
<< psubdiffcont >>
rect -742 1412 742 1446
rect -838 -1350 -804 1350
rect 804 -1350 838 1350
rect -742 -1446 742 -1412
<< xpolycontact >>
rect -708 884 -426 1316
rect -708 52 -426 484
rect -330 884 -48 1316
rect -330 52 -48 484
rect 48 884 330 1316
rect 48 52 330 484
rect 426 884 708 1316
rect 426 52 708 484
rect -708 -484 -426 -52
rect -708 -1316 -426 -884
rect -330 -484 -48 -52
rect -330 -1316 -48 -884
rect 48 -484 330 -52
rect 48 -1316 330 -884
rect 426 -484 708 -52
rect 426 -1316 708 -884
<< xpolyres >>
rect -708 484 -426 884
rect -330 484 -48 884
rect 48 484 330 884
rect 426 484 708 884
rect -708 -884 -426 -484
rect -330 -884 -48 -484
rect 48 -884 330 -484
rect 426 -884 708 -484
<< locali >>
rect -838 1412 -742 1446
rect 742 1412 838 1446
rect -838 1350 -804 1412
rect 804 1350 838 1412
rect -838 -1412 -804 -1350
rect 804 -1412 838 -1350
rect -838 -1446 -742 -1412
rect 742 -1446 838 -1412
<< viali >>
rect -692 901 -442 1298
rect -314 901 -64 1298
rect 64 901 314 1298
rect 442 901 692 1298
rect -692 70 -442 467
rect -314 70 -64 467
rect 64 70 314 467
rect 442 70 692 467
rect -692 -467 -442 -70
rect -314 -467 -64 -70
rect 64 -467 314 -70
rect 442 -467 692 -70
rect -692 -1298 -442 -901
rect -314 -1298 -64 -901
rect 64 -1298 314 -901
rect 442 -1298 692 -901
<< metal1 >>
rect -698 1298 -436 1310
rect -698 901 -692 1298
rect -442 901 -436 1298
rect -698 889 -436 901
rect -320 1298 -58 1310
rect -320 901 -314 1298
rect -64 901 -58 1298
rect -320 889 -58 901
rect 58 1298 320 1310
rect 58 901 64 1298
rect 314 901 320 1298
rect 58 889 320 901
rect 436 1298 698 1310
rect 436 901 442 1298
rect 692 901 698 1298
rect 436 889 698 901
rect -698 467 -436 479
rect -698 70 -692 467
rect -442 70 -436 467
rect -698 58 -436 70
rect -320 467 -58 479
rect -320 70 -314 467
rect -64 70 -58 467
rect -320 58 -58 70
rect 58 467 320 479
rect 58 70 64 467
rect 314 70 320 467
rect 58 58 320 70
rect 436 467 698 479
rect 436 70 442 467
rect 692 70 698 467
rect 436 58 698 70
rect -698 -70 -436 -58
rect -698 -467 -692 -70
rect -442 -467 -436 -70
rect -698 -479 -436 -467
rect -320 -70 -58 -58
rect -320 -467 -314 -70
rect -64 -467 -58 -70
rect -320 -479 -58 -467
rect 58 -70 320 -58
rect 58 -467 64 -70
rect 314 -467 320 -70
rect 58 -479 320 -467
rect 436 -70 698 -58
rect 436 -467 442 -70
rect 692 -467 698 -70
rect 436 -479 698 -467
rect -698 -901 -436 -889
rect -698 -1298 -692 -901
rect -442 -1298 -436 -901
rect -698 -1310 -436 -1298
rect -320 -901 -58 -889
rect -320 -1298 -314 -901
rect -64 -1298 -58 -901
rect -320 -1310 -58 -1298
rect 58 -901 320 -889
rect 58 -1298 64 -901
rect 314 -1298 320 -901
rect 58 -1310 320 -1298
rect 436 -901 698 -889
rect 436 -1298 442 -901
rect 692 -1298 698 -901
rect 436 -1310 698 -1298
<< res1p41 >>
rect -710 482 -424 886
rect -332 482 -46 886
rect 46 482 332 886
rect 424 482 710 886
rect -710 -886 -424 -482
rect -332 -886 -46 -482
rect 46 -886 332 -482
rect 424 -886 710 -482
<< properties >>
string FIXED_BBOX -821 -1429 821 1429
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 2 m 2 nx 4 wmin 1.410 lmin 0.50 rho 2000 val 3.103k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
