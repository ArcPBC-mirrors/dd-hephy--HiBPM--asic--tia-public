magic
tech sky130A
magscale 1 2
timestamp 1683889268
<< pwell >>
rect -1600 3804 526 6768
rect 1200 3804 3326 6768
rect -1180 3000 114 3804
rect 1620 3000 2914 3804
rect 4284 3002 7498 5674
rect 7924 3002 11138 5674
rect 11904 3002 15118 5674
rect 15544 3002 18758 5674
rect 4084 3000 11234 3002
rect -1720 1420 -810 2842
rect -680 1420 230 2842
rect 360 1420 1270 2842
rect 1400 1420 2310 2842
rect 2440 1420 3350 2842
rect 4084 1580 4994 3000
rect 5124 1580 6034 3000
rect 6164 1580 7074 3000
rect 7204 1580 8114 3000
rect 8244 1580 9154 3000
rect 9284 1580 10194 3000
rect 10324 1580 11234 3000
rect 11704 3000 18854 3002
rect 11704 1580 12614 3000
rect 12744 1580 13654 3000
rect 13784 1580 14694 3000
rect 14824 1580 15734 3000
rect 15864 1580 16774 3000
rect 16904 1580 17814 3000
rect 17944 1580 18854 3000
rect -1720 600 3482 1420
rect 4084 760 11366 1580
rect 11704 760 18986 1580
rect -7550 -1282 -6256 156
rect -7550 -3102 -6640 -1680
rect -6210 -1850 -5590 142
rect 4084 -660 4994 760
rect 5124 -660 6034 760
rect 6164 -660 7074 760
rect 7204 -660 8114 760
rect 8244 -660 9154 760
rect 9284 -660 10194 760
rect 10324 -660 11234 760
rect 11704 -660 12614 760
rect 12744 -660 13654 760
rect 13784 -660 14694 760
rect 14824 -660 15734 760
rect 15864 -660 16774 760
rect 16904 -660 17814 760
rect 17944 -660 18854 760
rect 4084 -1480 11366 -660
rect 11704 -1480 18986 -660
rect 4084 -2900 4994 -1480
rect 5124 -2900 6034 -1480
rect 6164 -2900 7074 -1480
rect 7204 -2900 8114 -1480
rect 8244 -2900 9154 -1480
rect 11704 -2900 12614 -1480
rect 12744 -2900 13654 -1480
rect 13784 -2900 14694 -1480
rect 14824 -2900 15734 -1480
rect 15864 -2900 16774 -1480
rect -7550 -3922 -6508 -3102
rect 4084 -3720 9286 -2900
rect 11704 -3720 16906 -2900
<< nmoslvt >>
rect -980 3210 -950 3610
rect -884 3210 -854 3610
rect -788 3210 -758 3610
rect -692 3210 -662 3610
rect -596 3210 -566 3610
rect -500 3210 -470 3610
rect -404 3210 -374 3610
rect -308 3210 -278 3610
rect -212 3210 -182 3610
rect -116 3210 -86 3610
rect 1820 3210 1850 3610
rect 1916 3210 1946 3610
rect 2012 3210 2042 3610
rect 2108 3210 2138 3610
rect 2204 3210 2234 3610
rect 2300 3210 2330 3610
rect 2396 3210 2426 3610
rect 2492 3210 2522 3610
rect 2588 3210 2618 3610
rect 2684 3210 2714 3610
rect 4484 5064 4514 5464
rect 4580 5064 4610 5464
rect 4676 5064 4706 5464
rect 4772 5064 4802 5464
rect 4868 5064 4898 5464
rect 4964 5064 4994 5464
rect 5060 5064 5090 5464
rect 5156 5064 5186 5464
rect 5252 5064 5282 5464
rect 5348 5064 5378 5464
rect 5444 5064 5474 5464
rect 5540 5064 5570 5464
rect 5636 5064 5666 5464
rect 5732 5064 5762 5464
rect 5828 5064 5858 5464
rect 5924 5064 5954 5464
rect 6020 5064 6050 5464
rect 6116 5064 6146 5464
rect 6212 5064 6242 5464
rect 6308 5064 6338 5464
rect 6404 5064 6434 5464
rect 6500 5064 6530 5464
rect 6596 5064 6626 5464
rect 6692 5064 6722 5464
rect 6788 5064 6818 5464
rect 6884 5064 6914 5464
rect 6980 5064 7010 5464
rect 7076 5064 7106 5464
rect 7172 5064 7202 5464
rect 7268 5064 7298 5464
rect 4484 4446 4514 4846
rect 4580 4446 4610 4846
rect 4676 4446 4706 4846
rect 4772 4446 4802 4846
rect 4868 4446 4898 4846
rect 4964 4446 4994 4846
rect 5060 4446 5090 4846
rect 5156 4446 5186 4846
rect 5252 4446 5282 4846
rect 5348 4446 5378 4846
rect 5444 4446 5474 4846
rect 5540 4446 5570 4846
rect 5636 4446 5666 4846
rect 5732 4446 5762 4846
rect 5828 4446 5858 4846
rect 5924 4446 5954 4846
rect 6020 4446 6050 4846
rect 6116 4446 6146 4846
rect 6212 4446 6242 4846
rect 6308 4446 6338 4846
rect 6404 4446 6434 4846
rect 6500 4446 6530 4846
rect 6596 4446 6626 4846
rect 6692 4446 6722 4846
rect 6788 4446 6818 4846
rect 6884 4446 6914 4846
rect 6980 4446 7010 4846
rect 7076 4446 7106 4846
rect 7172 4446 7202 4846
rect 7268 4446 7298 4846
rect 4484 3828 4514 4228
rect 4580 3828 4610 4228
rect 4676 3828 4706 4228
rect 4772 3828 4802 4228
rect 4868 3828 4898 4228
rect 4964 3828 4994 4228
rect 5060 3828 5090 4228
rect 5156 3828 5186 4228
rect 5252 3828 5282 4228
rect 5348 3828 5378 4228
rect 5444 3828 5474 4228
rect 5540 3828 5570 4228
rect 5636 3828 5666 4228
rect 5732 3828 5762 4228
rect 5828 3828 5858 4228
rect 5924 3828 5954 4228
rect 6020 3828 6050 4228
rect 6116 3828 6146 4228
rect 6212 3828 6242 4228
rect 6308 3828 6338 4228
rect 6404 3828 6434 4228
rect 6500 3828 6530 4228
rect 6596 3828 6626 4228
rect 6692 3828 6722 4228
rect 6788 3828 6818 4228
rect 6884 3828 6914 4228
rect 6980 3828 7010 4228
rect 7076 3828 7106 4228
rect 7172 3828 7202 4228
rect 7268 3828 7298 4228
rect 4484 3210 4514 3610
rect 4580 3210 4610 3610
rect 4676 3210 4706 3610
rect 4772 3210 4802 3610
rect 4868 3210 4898 3610
rect 4964 3210 4994 3610
rect 5060 3210 5090 3610
rect 5156 3210 5186 3610
rect 5252 3210 5282 3610
rect 5348 3210 5378 3610
rect 5444 3210 5474 3610
rect 5540 3210 5570 3610
rect 5636 3210 5666 3610
rect 5732 3210 5762 3610
rect 5828 3210 5858 3610
rect 5924 3210 5954 3610
rect 6020 3210 6050 3610
rect 6116 3210 6146 3610
rect 6212 3210 6242 3610
rect 6308 3210 6338 3610
rect 6404 3210 6434 3610
rect 6500 3210 6530 3610
rect 6596 3210 6626 3610
rect 6692 3210 6722 3610
rect 6788 3210 6818 3610
rect 6884 3210 6914 3610
rect 6980 3210 7010 3610
rect 7076 3210 7106 3610
rect 7172 3210 7202 3610
rect 7268 3210 7298 3610
rect 8124 5064 8154 5464
rect 8220 5064 8250 5464
rect 8316 5064 8346 5464
rect 8412 5064 8442 5464
rect 8508 5064 8538 5464
rect 8604 5064 8634 5464
rect 8700 5064 8730 5464
rect 8796 5064 8826 5464
rect 8892 5064 8922 5464
rect 8988 5064 9018 5464
rect 9084 5064 9114 5464
rect 9180 5064 9210 5464
rect 9276 5064 9306 5464
rect 9372 5064 9402 5464
rect 9468 5064 9498 5464
rect 9564 5064 9594 5464
rect 9660 5064 9690 5464
rect 9756 5064 9786 5464
rect 9852 5064 9882 5464
rect 9948 5064 9978 5464
rect 10044 5064 10074 5464
rect 10140 5064 10170 5464
rect 10236 5064 10266 5464
rect 10332 5064 10362 5464
rect 10428 5064 10458 5464
rect 10524 5064 10554 5464
rect 10620 5064 10650 5464
rect 10716 5064 10746 5464
rect 10812 5064 10842 5464
rect 10908 5064 10938 5464
rect 8124 4446 8154 4846
rect 8220 4446 8250 4846
rect 8316 4446 8346 4846
rect 8412 4446 8442 4846
rect 8508 4446 8538 4846
rect 8604 4446 8634 4846
rect 8700 4446 8730 4846
rect 8796 4446 8826 4846
rect 8892 4446 8922 4846
rect 8988 4446 9018 4846
rect 9084 4446 9114 4846
rect 9180 4446 9210 4846
rect 9276 4446 9306 4846
rect 9372 4446 9402 4846
rect 9468 4446 9498 4846
rect 9564 4446 9594 4846
rect 9660 4446 9690 4846
rect 9756 4446 9786 4846
rect 9852 4446 9882 4846
rect 9948 4446 9978 4846
rect 10044 4446 10074 4846
rect 10140 4446 10170 4846
rect 10236 4446 10266 4846
rect 10332 4446 10362 4846
rect 10428 4446 10458 4846
rect 10524 4446 10554 4846
rect 10620 4446 10650 4846
rect 10716 4446 10746 4846
rect 10812 4446 10842 4846
rect 10908 4446 10938 4846
rect 8124 3828 8154 4228
rect 8220 3828 8250 4228
rect 8316 3828 8346 4228
rect 8412 3828 8442 4228
rect 8508 3828 8538 4228
rect 8604 3828 8634 4228
rect 8700 3828 8730 4228
rect 8796 3828 8826 4228
rect 8892 3828 8922 4228
rect 8988 3828 9018 4228
rect 9084 3828 9114 4228
rect 9180 3828 9210 4228
rect 9276 3828 9306 4228
rect 9372 3828 9402 4228
rect 9468 3828 9498 4228
rect 9564 3828 9594 4228
rect 9660 3828 9690 4228
rect 9756 3828 9786 4228
rect 9852 3828 9882 4228
rect 9948 3828 9978 4228
rect 10044 3828 10074 4228
rect 10140 3828 10170 4228
rect 10236 3828 10266 4228
rect 10332 3828 10362 4228
rect 10428 3828 10458 4228
rect 10524 3828 10554 4228
rect 10620 3828 10650 4228
rect 10716 3828 10746 4228
rect 10812 3828 10842 4228
rect 10908 3828 10938 4228
rect 8124 3210 8154 3610
rect 8220 3210 8250 3610
rect 8316 3210 8346 3610
rect 8412 3210 8442 3610
rect 8508 3210 8538 3610
rect 8604 3210 8634 3610
rect 8700 3210 8730 3610
rect 8796 3210 8826 3610
rect 8892 3210 8922 3610
rect 8988 3210 9018 3610
rect 9084 3210 9114 3610
rect 9180 3210 9210 3610
rect 9276 3210 9306 3610
rect 9372 3210 9402 3610
rect 9468 3210 9498 3610
rect 9564 3210 9594 3610
rect 9660 3210 9690 3610
rect 9756 3210 9786 3610
rect 9852 3210 9882 3610
rect 9948 3210 9978 3610
rect 10044 3210 10074 3610
rect 10140 3210 10170 3610
rect 10236 3210 10266 3610
rect 10332 3210 10362 3610
rect 10428 3210 10458 3610
rect 10524 3210 10554 3610
rect 10620 3210 10650 3610
rect 10716 3210 10746 3610
rect 10812 3210 10842 3610
rect 10908 3210 10938 3610
rect 12104 5064 12134 5464
rect 12200 5064 12230 5464
rect 12296 5064 12326 5464
rect 12392 5064 12422 5464
rect 12488 5064 12518 5464
rect 12584 5064 12614 5464
rect 12680 5064 12710 5464
rect 12776 5064 12806 5464
rect 12872 5064 12902 5464
rect 12968 5064 12998 5464
rect 13064 5064 13094 5464
rect 13160 5064 13190 5464
rect 13256 5064 13286 5464
rect 13352 5064 13382 5464
rect 13448 5064 13478 5464
rect 13544 5064 13574 5464
rect 13640 5064 13670 5464
rect 13736 5064 13766 5464
rect 13832 5064 13862 5464
rect 13928 5064 13958 5464
rect 14024 5064 14054 5464
rect 14120 5064 14150 5464
rect 14216 5064 14246 5464
rect 14312 5064 14342 5464
rect 14408 5064 14438 5464
rect 14504 5064 14534 5464
rect 14600 5064 14630 5464
rect 14696 5064 14726 5464
rect 14792 5064 14822 5464
rect 14888 5064 14918 5464
rect 12104 4446 12134 4846
rect 12200 4446 12230 4846
rect 12296 4446 12326 4846
rect 12392 4446 12422 4846
rect 12488 4446 12518 4846
rect 12584 4446 12614 4846
rect 12680 4446 12710 4846
rect 12776 4446 12806 4846
rect 12872 4446 12902 4846
rect 12968 4446 12998 4846
rect 13064 4446 13094 4846
rect 13160 4446 13190 4846
rect 13256 4446 13286 4846
rect 13352 4446 13382 4846
rect 13448 4446 13478 4846
rect 13544 4446 13574 4846
rect 13640 4446 13670 4846
rect 13736 4446 13766 4846
rect 13832 4446 13862 4846
rect 13928 4446 13958 4846
rect 14024 4446 14054 4846
rect 14120 4446 14150 4846
rect 14216 4446 14246 4846
rect 14312 4446 14342 4846
rect 14408 4446 14438 4846
rect 14504 4446 14534 4846
rect 14600 4446 14630 4846
rect 14696 4446 14726 4846
rect 14792 4446 14822 4846
rect 14888 4446 14918 4846
rect 12104 3828 12134 4228
rect 12200 3828 12230 4228
rect 12296 3828 12326 4228
rect 12392 3828 12422 4228
rect 12488 3828 12518 4228
rect 12584 3828 12614 4228
rect 12680 3828 12710 4228
rect 12776 3828 12806 4228
rect 12872 3828 12902 4228
rect 12968 3828 12998 4228
rect 13064 3828 13094 4228
rect 13160 3828 13190 4228
rect 13256 3828 13286 4228
rect 13352 3828 13382 4228
rect 13448 3828 13478 4228
rect 13544 3828 13574 4228
rect 13640 3828 13670 4228
rect 13736 3828 13766 4228
rect 13832 3828 13862 4228
rect 13928 3828 13958 4228
rect 14024 3828 14054 4228
rect 14120 3828 14150 4228
rect 14216 3828 14246 4228
rect 14312 3828 14342 4228
rect 14408 3828 14438 4228
rect 14504 3828 14534 4228
rect 14600 3828 14630 4228
rect 14696 3828 14726 4228
rect 14792 3828 14822 4228
rect 14888 3828 14918 4228
rect 12104 3210 12134 3610
rect 12200 3210 12230 3610
rect 12296 3210 12326 3610
rect 12392 3210 12422 3610
rect 12488 3210 12518 3610
rect 12584 3210 12614 3610
rect 12680 3210 12710 3610
rect 12776 3210 12806 3610
rect 12872 3210 12902 3610
rect 12968 3210 12998 3610
rect 13064 3210 13094 3610
rect 13160 3210 13190 3610
rect 13256 3210 13286 3610
rect 13352 3210 13382 3610
rect 13448 3210 13478 3610
rect 13544 3210 13574 3610
rect 13640 3210 13670 3610
rect 13736 3210 13766 3610
rect 13832 3210 13862 3610
rect 13928 3210 13958 3610
rect 14024 3210 14054 3610
rect 14120 3210 14150 3610
rect 14216 3210 14246 3610
rect 14312 3210 14342 3610
rect 14408 3210 14438 3610
rect 14504 3210 14534 3610
rect 14600 3210 14630 3610
rect 14696 3210 14726 3610
rect 14792 3210 14822 3610
rect 14888 3210 14918 3610
rect 15744 5064 15774 5464
rect 15840 5064 15870 5464
rect 15936 5064 15966 5464
rect 16032 5064 16062 5464
rect 16128 5064 16158 5464
rect 16224 5064 16254 5464
rect 16320 5064 16350 5464
rect 16416 5064 16446 5464
rect 16512 5064 16542 5464
rect 16608 5064 16638 5464
rect 16704 5064 16734 5464
rect 16800 5064 16830 5464
rect 16896 5064 16926 5464
rect 16992 5064 17022 5464
rect 17088 5064 17118 5464
rect 17184 5064 17214 5464
rect 17280 5064 17310 5464
rect 17376 5064 17406 5464
rect 17472 5064 17502 5464
rect 17568 5064 17598 5464
rect 17664 5064 17694 5464
rect 17760 5064 17790 5464
rect 17856 5064 17886 5464
rect 17952 5064 17982 5464
rect 18048 5064 18078 5464
rect 18144 5064 18174 5464
rect 18240 5064 18270 5464
rect 18336 5064 18366 5464
rect 18432 5064 18462 5464
rect 18528 5064 18558 5464
rect 15744 4446 15774 4846
rect 15840 4446 15870 4846
rect 15936 4446 15966 4846
rect 16032 4446 16062 4846
rect 16128 4446 16158 4846
rect 16224 4446 16254 4846
rect 16320 4446 16350 4846
rect 16416 4446 16446 4846
rect 16512 4446 16542 4846
rect 16608 4446 16638 4846
rect 16704 4446 16734 4846
rect 16800 4446 16830 4846
rect 16896 4446 16926 4846
rect 16992 4446 17022 4846
rect 17088 4446 17118 4846
rect 17184 4446 17214 4846
rect 17280 4446 17310 4846
rect 17376 4446 17406 4846
rect 17472 4446 17502 4846
rect 17568 4446 17598 4846
rect 17664 4446 17694 4846
rect 17760 4446 17790 4846
rect 17856 4446 17886 4846
rect 17952 4446 17982 4846
rect 18048 4446 18078 4846
rect 18144 4446 18174 4846
rect 18240 4446 18270 4846
rect 18336 4446 18366 4846
rect 18432 4446 18462 4846
rect 18528 4446 18558 4846
rect 15744 3828 15774 4228
rect 15840 3828 15870 4228
rect 15936 3828 15966 4228
rect 16032 3828 16062 4228
rect 16128 3828 16158 4228
rect 16224 3828 16254 4228
rect 16320 3828 16350 4228
rect 16416 3828 16446 4228
rect 16512 3828 16542 4228
rect 16608 3828 16638 4228
rect 16704 3828 16734 4228
rect 16800 3828 16830 4228
rect 16896 3828 16926 4228
rect 16992 3828 17022 4228
rect 17088 3828 17118 4228
rect 17184 3828 17214 4228
rect 17280 3828 17310 4228
rect 17376 3828 17406 4228
rect 17472 3828 17502 4228
rect 17568 3828 17598 4228
rect 17664 3828 17694 4228
rect 17760 3828 17790 4228
rect 17856 3828 17886 4228
rect 17952 3828 17982 4228
rect 18048 3828 18078 4228
rect 18144 3828 18174 4228
rect 18240 3828 18270 4228
rect 18336 3828 18366 4228
rect 18432 3828 18462 4228
rect 18528 3828 18558 4228
rect 15744 3210 15774 3610
rect 15840 3210 15870 3610
rect 15936 3210 15966 3610
rect 16032 3210 16062 3610
rect 16128 3210 16158 3610
rect 16224 3210 16254 3610
rect 16320 3210 16350 3610
rect 16416 3210 16446 3610
rect 16512 3210 16542 3610
rect 16608 3210 16638 3610
rect 16704 3210 16734 3610
rect 16800 3210 16830 3610
rect 16896 3210 16926 3610
rect 16992 3210 17022 3610
rect 17088 3210 17118 3610
rect 17184 3210 17214 3610
rect 17280 3210 17310 3610
rect 17376 3210 17406 3610
rect 17472 3210 17502 3610
rect 17568 3210 17598 3610
rect 17664 3210 17694 3610
rect 17760 3210 17790 3610
rect 17856 3210 17886 3610
rect 17952 3210 17982 3610
rect 18048 3210 18078 3610
rect 18144 3210 18174 3610
rect 18240 3210 18270 3610
rect 18336 3210 18366 3610
rect 18432 3210 18462 3610
rect 18528 3210 18558 3610
rect -1520 2232 -1490 2632
rect -1424 2232 -1394 2632
rect -1328 2232 -1298 2632
rect -1232 2232 -1202 2632
rect -1136 2232 -1106 2632
rect -1040 2232 -1010 2632
rect -1520 1614 -1490 2014
rect -1424 1614 -1394 2014
rect -1328 1614 -1298 2014
rect -1232 1614 -1202 2014
rect -1136 1614 -1106 2014
rect -1040 1614 -1010 2014
rect -480 2232 -450 2632
rect -384 2232 -354 2632
rect -288 2232 -258 2632
rect -192 2232 -162 2632
rect -96 2232 -66 2632
rect 0 2232 30 2632
rect -480 1614 -450 2014
rect -384 1614 -354 2014
rect -288 1614 -258 2014
rect -192 1614 -162 2014
rect -96 1614 -66 2014
rect 0 1614 30 2014
rect 560 2232 590 2632
rect 656 2232 686 2632
rect 752 2232 782 2632
rect 848 2232 878 2632
rect 944 2232 974 2632
rect 1040 2232 1070 2632
rect 560 1614 590 2014
rect 656 1614 686 2014
rect 752 1614 782 2014
rect 848 1614 878 2014
rect 944 1614 974 2014
rect 1040 1614 1070 2014
rect 1600 2232 1630 2632
rect 1696 2232 1726 2632
rect 1792 2232 1822 2632
rect 1888 2232 1918 2632
rect 1984 2232 2014 2632
rect 2080 2232 2110 2632
rect 1600 1614 1630 2014
rect 1696 1614 1726 2014
rect 1792 1614 1822 2014
rect 1888 1614 1918 2014
rect 1984 1614 2014 2014
rect 2080 1614 2110 2014
rect 2640 2232 2670 2632
rect 2736 2232 2766 2632
rect 2832 2232 2862 2632
rect 2928 2232 2958 2632
rect 3024 2232 3054 2632
rect 3120 2232 3150 2632
rect 2640 1614 2670 2014
rect 2736 1614 2766 2014
rect 2832 1614 2862 2014
rect 2928 1614 2958 2014
rect 3024 1614 3054 2014
rect 3120 1614 3150 2014
rect 4284 2392 4314 2792
rect 4380 2392 4410 2792
rect 4476 2392 4506 2792
rect 4572 2392 4602 2792
rect 4668 2392 4698 2792
rect 4764 2392 4794 2792
rect 4284 1774 4314 2174
rect 4380 1774 4410 2174
rect 4476 1774 4506 2174
rect 4572 1774 4602 2174
rect 4668 1774 4698 2174
rect 4764 1774 4794 2174
rect 5324 2392 5354 2792
rect 5420 2392 5450 2792
rect 5516 2392 5546 2792
rect 5612 2392 5642 2792
rect 5708 2392 5738 2792
rect 5804 2392 5834 2792
rect 5324 1774 5354 2174
rect 5420 1774 5450 2174
rect 5516 1774 5546 2174
rect 5612 1774 5642 2174
rect 5708 1774 5738 2174
rect 5804 1774 5834 2174
rect 6364 2392 6394 2792
rect 6460 2392 6490 2792
rect 6556 2392 6586 2792
rect 6652 2392 6682 2792
rect 6748 2392 6778 2792
rect 6844 2392 6874 2792
rect 6364 1774 6394 2174
rect 6460 1774 6490 2174
rect 6556 1774 6586 2174
rect 6652 1774 6682 2174
rect 6748 1774 6778 2174
rect 6844 1774 6874 2174
rect 7404 2392 7434 2792
rect 7500 2392 7530 2792
rect 7596 2392 7626 2792
rect 7692 2392 7722 2792
rect 7788 2392 7818 2792
rect 7884 2392 7914 2792
rect 7404 1774 7434 2174
rect 7500 1774 7530 2174
rect 7596 1774 7626 2174
rect 7692 1774 7722 2174
rect 7788 1774 7818 2174
rect 7884 1774 7914 2174
rect 8444 2392 8474 2792
rect 8540 2392 8570 2792
rect 8636 2392 8666 2792
rect 8732 2392 8762 2792
rect 8828 2392 8858 2792
rect 8924 2392 8954 2792
rect 8444 1774 8474 2174
rect 8540 1774 8570 2174
rect 8636 1774 8666 2174
rect 8732 1774 8762 2174
rect 8828 1774 8858 2174
rect 8924 1774 8954 2174
rect 9484 2392 9514 2792
rect 9580 2392 9610 2792
rect 9676 2392 9706 2792
rect 9772 2392 9802 2792
rect 9868 2392 9898 2792
rect 9964 2392 9994 2792
rect 9484 1774 9514 2174
rect 9580 1774 9610 2174
rect 9676 1774 9706 2174
rect 9772 1774 9802 2174
rect 9868 1774 9898 2174
rect 9964 1774 9994 2174
rect 10524 2392 10554 2792
rect 10620 2392 10650 2792
rect 10716 2392 10746 2792
rect 10812 2392 10842 2792
rect 10908 2392 10938 2792
rect 11004 2392 11034 2792
rect 10524 1774 10554 2174
rect 10620 1774 10650 2174
rect 10716 1774 10746 2174
rect 10812 1774 10842 2174
rect 10908 1774 10938 2174
rect 11004 1774 11034 2174
rect 11904 2392 11934 2792
rect 12000 2392 12030 2792
rect 12096 2392 12126 2792
rect 12192 2392 12222 2792
rect 12288 2392 12318 2792
rect 12384 2392 12414 2792
rect 11904 1774 11934 2174
rect 12000 1774 12030 2174
rect 12096 1774 12126 2174
rect 12192 1774 12222 2174
rect 12288 1774 12318 2174
rect 12384 1774 12414 2174
rect 12944 2392 12974 2792
rect 13040 2392 13070 2792
rect 13136 2392 13166 2792
rect 13232 2392 13262 2792
rect 13328 2392 13358 2792
rect 13424 2392 13454 2792
rect 12944 1774 12974 2174
rect 13040 1774 13070 2174
rect 13136 1774 13166 2174
rect 13232 1774 13262 2174
rect 13328 1774 13358 2174
rect 13424 1774 13454 2174
rect 13984 2392 14014 2792
rect 14080 2392 14110 2792
rect 14176 2392 14206 2792
rect 14272 2392 14302 2792
rect 14368 2392 14398 2792
rect 14464 2392 14494 2792
rect 13984 1774 14014 2174
rect 14080 1774 14110 2174
rect 14176 1774 14206 2174
rect 14272 1774 14302 2174
rect 14368 1774 14398 2174
rect 14464 1774 14494 2174
rect 15024 2392 15054 2792
rect 15120 2392 15150 2792
rect 15216 2392 15246 2792
rect 15312 2392 15342 2792
rect 15408 2392 15438 2792
rect 15504 2392 15534 2792
rect 15024 1774 15054 2174
rect 15120 1774 15150 2174
rect 15216 1774 15246 2174
rect 15312 1774 15342 2174
rect 15408 1774 15438 2174
rect 15504 1774 15534 2174
rect 16064 2392 16094 2792
rect 16160 2392 16190 2792
rect 16256 2392 16286 2792
rect 16352 2392 16382 2792
rect 16448 2392 16478 2792
rect 16544 2392 16574 2792
rect 16064 1774 16094 2174
rect 16160 1774 16190 2174
rect 16256 1774 16286 2174
rect 16352 1774 16382 2174
rect 16448 1774 16478 2174
rect 16544 1774 16574 2174
rect 17104 2392 17134 2792
rect 17200 2392 17230 2792
rect 17296 2392 17326 2792
rect 17392 2392 17422 2792
rect 17488 2392 17518 2792
rect 17584 2392 17614 2792
rect 17104 1774 17134 2174
rect 17200 1774 17230 2174
rect 17296 1774 17326 2174
rect 17392 1774 17422 2174
rect 17488 1774 17518 2174
rect 17584 1774 17614 2174
rect 18144 2392 18174 2792
rect 18240 2392 18270 2792
rect 18336 2392 18366 2792
rect 18432 2392 18462 2792
rect 18528 2392 18558 2792
rect 18624 2392 18654 2792
rect 18144 1774 18174 2174
rect 18240 1774 18270 2174
rect 18336 1774 18366 2174
rect 18432 1774 18462 2174
rect 18528 1774 18558 2174
rect 18624 1774 18654 2174
rect -1524 810 -1464 1210
rect -1406 810 -1346 1210
rect -1288 810 -1228 1210
rect -1170 810 -1110 1210
rect -1052 810 -992 1210
rect -934 810 -874 1210
rect -484 810 -424 1210
rect -366 810 -306 1210
rect -248 810 -188 1210
rect -130 810 -70 1210
rect -12 810 48 1210
rect 106 810 166 1210
rect 556 810 616 1210
rect 674 810 734 1210
rect 792 810 852 1210
rect 910 810 970 1210
rect 1028 810 1088 1210
rect 1146 810 1206 1210
rect 1596 810 1656 1210
rect 1714 810 1774 1210
rect 1832 810 1892 1210
rect 1950 810 2010 1210
rect 2068 810 2128 1210
rect 2186 810 2246 1210
rect 2636 810 2696 1210
rect 2754 810 2814 1210
rect 2872 810 2932 1210
rect 2990 810 3050 1210
rect 3108 810 3168 1210
rect 3226 810 3286 1210
rect 4280 970 4340 1370
rect 4398 970 4458 1370
rect 4516 970 4576 1370
rect 4634 970 4694 1370
rect 4752 970 4812 1370
rect 4870 970 4930 1370
rect 5320 970 5380 1370
rect 5438 970 5498 1370
rect 5556 970 5616 1370
rect 5674 970 5734 1370
rect 5792 970 5852 1370
rect 5910 970 5970 1370
rect 6360 970 6420 1370
rect 6478 970 6538 1370
rect 6596 970 6656 1370
rect 6714 970 6774 1370
rect 6832 970 6892 1370
rect 6950 970 7010 1370
rect 7400 970 7460 1370
rect 7518 970 7578 1370
rect 7636 970 7696 1370
rect 7754 970 7814 1370
rect 7872 970 7932 1370
rect 7990 970 8050 1370
rect 8440 970 8500 1370
rect 8558 970 8618 1370
rect 8676 970 8736 1370
rect 8794 970 8854 1370
rect 8912 970 8972 1370
rect 9030 970 9090 1370
rect 9480 970 9540 1370
rect 9598 970 9658 1370
rect 9716 970 9776 1370
rect 9834 970 9894 1370
rect 9952 970 10012 1370
rect 10070 970 10130 1370
rect 10520 970 10580 1370
rect 10638 970 10698 1370
rect 10756 970 10816 1370
rect 10874 970 10934 1370
rect 10992 970 11052 1370
rect 11110 970 11170 1370
rect 11900 970 11960 1370
rect 12018 970 12078 1370
rect 12136 970 12196 1370
rect 12254 970 12314 1370
rect 12372 970 12432 1370
rect 12490 970 12550 1370
rect 12940 970 13000 1370
rect 13058 970 13118 1370
rect 13176 970 13236 1370
rect 13294 970 13354 1370
rect 13412 970 13472 1370
rect 13530 970 13590 1370
rect 13980 970 14040 1370
rect 14098 970 14158 1370
rect 14216 970 14276 1370
rect 14334 970 14394 1370
rect 14452 970 14512 1370
rect 14570 970 14630 1370
rect 15020 970 15080 1370
rect 15138 970 15198 1370
rect 15256 970 15316 1370
rect 15374 970 15434 1370
rect 15492 970 15552 1370
rect 15610 970 15670 1370
rect 16060 970 16120 1370
rect 16178 970 16238 1370
rect 16296 970 16356 1370
rect 16414 970 16474 1370
rect 16532 970 16592 1370
rect 16650 970 16710 1370
rect 17100 970 17160 1370
rect 17218 970 17278 1370
rect 17336 970 17396 1370
rect 17454 970 17514 1370
rect 17572 970 17632 1370
rect 17690 970 17750 1370
rect 18140 970 18200 1370
rect 18258 970 18318 1370
rect 18376 970 18436 1370
rect 18494 970 18554 1370
rect 18612 970 18672 1370
rect 18730 970 18790 1370
rect -7350 -454 -7320 -54
rect -7254 -454 -7224 -54
rect -7158 -454 -7128 -54
rect -7062 -454 -7032 -54
rect -6966 -454 -6936 -54
rect -6870 -454 -6840 -54
rect -6774 -454 -6744 -54
rect -6678 -454 -6648 -54
rect -6582 -454 -6552 -54
rect -6486 -454 -6456 -54
rect -7350 -1072 -7320 -672
rect -7254 -1072 -7224 -672
rect -7158 -1072 -7128 -672
rect -7062 -1072 -7032 -672
rect -6966 -1072 -6936 -672
rect -6870 -1072 -6840 -672
rect -6774 -1072 -6744 -672
rect -6678 -1072 -6648 -672
rect -6582 -1072 -6552 -672
rect -6486 -1072 -6456 -672
rect -7350 -2290 -7320 -1890
rect -7254 -2290 -7224 -1890
rect -7158 -2290 -7128 -1890
rect -7062 -2290 -7032 -1890
rect -6966 -2290 -6936 -1890
rect -6870 -2290 -6840 -1890
rect -7350 -2908 -7320 -2508
rect -7254 -2908 -7224 -2508
rect -7158 -2908 -7128 -2508
rect -7062 -2908 -7032 -2508
rect -6966 -2908 -6936 -2508
rect -6870 -2908 -6840 -2508
rect -6000 -1654 -5800 -54
rect 4284 152 4314 552
rect 4380 152 4410 552
rect 4476 152 4506 552
rect 4572 152 4602 552
rect 4668 152 4698 552
rect 4764 152 4794 552
rect 4284 -466 4314 -66
rect 4380 -466 4410 -66
rect 4476 -466 4506 -66
rect 4572 -466 4602 -66
rect 4668 -466 4698 -66
rect 4764 -466 4794 -66
rect 5324 152 5354 552
rect 5420 152 5450 552
rect 5516 152 5546 552
rect 5612 152 5642 552
rect 5708 152 5738 552
rect 5804 152 5834 552
rect 5324 -466 5354 -66
rect 5420 -466 5450 -66
rect 5516 -466 5546 -66
rect 5612 -466 5642 -66
rect 5708 -466 5738 -66
rect 5804 -466 5834 -66
rect 6364 152 6394 552
rect 6460 152 6490 552
rect 6556 152 6586 552
rect 6652 152 6682 552
rect 6748 152 6778 552
rect 6844 152 6874 552
rect 6364 -466 6394 -66
rect 6460 -466 6490 -66
rect 6556 -466 6586 -66
rect 6652 -466 6682 -66
rect 6748 -466 6778 -66
rect 6844 -466 6874 -66
rect 7404 152 7434 552
rect 7500 152 7530 552
rect 7596 152 7626 552
rect 7692 152 7722 552
rect 7788 152 7818 552
rect 7884 152 7914 552
rect 7404 -466 7434 -66
rect 7500 -466 7530 -66
rect 7596 -466 7626 -66
rect 7692 -466 7722 -66
rect 7788 -466 7818 -66
rect 7884 -466 7914 -66
rect 8444 152 8474 552
rect 8540 152 8570 552
rect 8636 152 8666 552
rect 8732 152 8762 552
rect 8828 152 8858 552
rect 8924 152 8954 552
rect 8444 -466 8474 -66
rect 8540 -466 8570 -66
rect 8636 -466 8666 -66
rect 8732 -466 8762 -66
rect 8828 -466 8858 -66
rect 8924 -466 8954 -66
rect 9484 152 9514 552
rect 9580 152 9610 552
rect 9676 152 9706 552
rect 9772 152 9802 552
rect 9868 152 9898 552
rect 9964 152 9994 552
rect 9484 -466 9514 -66
rect 9580 -466 9610 -66
rect 9676 -466 9706 -66
rect 9772 -466 9802 -66
rect 9868 -466 9898 -66
rect 9964 -466 9994 -66
rect 10524 152 10554 552
rect 10620 152 10650 552
rect 10716 152 10746 552
rect 10812 152 10842 552
rect 10908 152 10938 552
rect 11004 152 11034 552
rect 10524 -466 10554 -66
rect 10620 -466 10650 -66
rect 10716 -466 10746 -66
rect 10812 -466 10842 -66
rect 10908 -466 10938 -66
rect 11004 -466 11034 -66
rect 11904 152 11934 552
rect 12000 152 12030 552
rect 12096 152 12126 552
rect 12192 152 12222 552
rect 12288 152 12318 552
rect 12384 152 12414 552
rect 11904 -466 11934 -66
rect 12000 -466 12030 -66
rect 12096 -466 12126 -66
rect 12192 -466 12222 -66
rect 12288 -466 12318 -66
rect 12384 -466 12414 -66
rect 12944 152 12974 552
rect 13040 152 13070 552
rect 13136 152 13166 552
rect 13232 152 13262 552
rect 13328 152 13358 552
rect 13424 152 13454 552
rect 12944 -466 12974 -66
rect 13040 -466 13070 -66
rect 13136 -466 13166 -66
rect 13232 -466 13262 -66
rect 13328 -466 13358 -66
rect 13424 -466 13454 -66
rect 13984 152 14014 552
rect 14080 152 14110 552
rect 14176 152 14206 552
rect 14272 152 14302 552
rect 14368 152 14398 552
rect 14464 152 14494 552
rect 13984 -466 14014 -66
rect 14080 -466 14110 -66
rect 14176 -466 14206 -66
rect 14272 -466 14302 -66
rect 14368 -466 14398 -66
rect 14464 -466 14494 -66
rect 15024 152 15054 552
rect 15120 152 15150 552
rect 15216 152 15246 552
rect 15312 152 15342 552
rect 15408 152 15438 552
rect 15504 152 15534 552
rect 15024 -466 15054 -66
rect 15120 -466 15150 -66
rect 15216 -466 15246 -66
rect 15312 -466 15342 -66
rect 15408 -466 15438 -66
rect 15504 -466 15534 -66
rect 16064 152 16094 552
rect 16160 152 16190 552
rect 16256 152 16286 552
rect 16352 152 16382 552
rect 16448 152 16478 552
rect 16544 152 16574 552
rect 16064 -466 16094 -66
rect 16160 -466 16190 -66
rect 16256 -466 16286 -66
rect 16352 -466 16382 -66
rect 16448 -466 16478 -66
rect 16544 -466 16574 -66
rect 17104 152 17134 552
rect 17200 152 17230 552
rect 17296 152 17326 552
rect 17392 152 17422 552
rect 17488 152 17518 552
rect 17584 152 17614 552
rect 17104 -466 17134 -66
rect 17200 -466 17230 -66
rect 17296 -466 17326 -66
rect 17392 -466 17422 -66
rect 17488 -466 17518 -66
rect 17584 -466 17614 -66
rect 18144 152 18174 552
rect 18240 152 18270 552
rect 18336 152 18366 552
rect 18432 152 18462 552
rect 18528 152 18558 552
rect 18624 152 18654 552
rect 18144 -466 18174 -66
rect 18240 -466 18270 -66
rect 18336 -466 18366 -66
rect 18432 -466 18462 -66
rect 18528 -466 18558 -66
rect 18624 -466 18654 -66
rect 4280 -1270 4340 -870
rect 4398 -1270 4458 -870
rect 4516 -1270 4576 -870
rect 4634 -1270 4694 -870
rect 4752 -1270 4812 -870
rect 4870 -1270 4930 -870
rect 5320 -1270 5380 -870
rect 5438 -1270 5498 -870
rect 5556 -1270 5616 -870
rect 5674 -1270 5734 -870
rect 5792 -1270 5852 -870
rect 5910 -1270 5970 -870
rect 6360 -1270 6420 -870
rect 6478 -1270 6538 -870
rect 6596 -1270 6656 -870
rect 6714 -1270 6774 -870
rect 6832 -1270 6892 -870
rect 6950 -1270 7010 -870
rect 7400 -1270 7460 -870
rect 7518 -1270 7578 -870
rect 7636 -1270 7696 -870
rect 7754 -1270 7814 -870
rect 7872 -1270 7932 -870
rect 7990 -1270 8050 -870
rect 8440 -1270 8500 -870
rect 8558 -1270 8618 -870
rect 8676 -1270 8736 -870
rect 8794 -1270 8854 -870
rect 8912 -1270 8972 -870
rect 9030 -1270 9090 -870
rect 9480 -1270 9540 -870
rect 9598 -1270 9658 -870
rect 9716 -1270 9776 -870
rect 9834 -1270 9894 -870
rect 9952 -1270 10012 -870
rect 10070 -1270 10130 -870
rect 10520 -1270 10580 -870
rect 10638 -1270 10698 -870
rect 10756 -1270 10816 -870
rect 10874 -1270 10934 -870
rect 10992 -1270 11052 -870
rect 11110 -1270 11170 -870
rect 11900 -1270 11960 -870
rect 12018 -1270 12078 -870
rect 12136 -1270 12196 -870
rect 12254 -1270 12314 -870
rect 12372 -1270 12432 -870
rect 12490 -1270 12550 -870
rect 12940 -1270 13000 -870
rect 13058 -1270 13118 -870
rect 13176 -1270 13236 -870
rect 13294 -1270 13354 -870
rect 13412 -1270 13472 -870
rect 13530 -1270 13590 -870
rect 13980 -1270 14040 -870
rect 14098 -1270 14158 -870
rect 14216 -1270 14276 -870
rect 14334 -1270 14394 -870
rect 14452 -1270 14512 -870
rect 14570 -1270 14630 -870
rect 15020 -1270 15080 -870
rect 15138 -1270 15198 -870
rect 15256 -1270 15316 -870
rect 15374 -1270 15434 -870
rect 15492 -1270 15552 -870
rect 15610 -1270 15670 -870
rect 16060 -1270 16120 -870
rect 16178 -1270 16238 -870
rect 16296 -1270 16356 -870
rect 16414 -1270 16474 -870
rect 16532 -1270 16592 -870
rect 16650 -1270 16710 -870
rect 17100 -1270 17160 -870
rect 17218 -1270 17278 -870
rect 17336 -1270 17396 -870
rect 17454 -1270 17514 -870
rect 17572 -1270 17632 -870
rect 17690 -1270 17750 -870
rect 18140 -1270 18200 -870
rect 18258 -1270 18318 -870
rect 18376 -1270 18436 -870
rect 18494 -1270 18554 -870
rect 18612 -1270 18672 -870
rect 18730 -1270 18790 -870
rect 4284 -2088 4314 -1688
rect 4380 -2088 4410 -1688
rect 4476 -2088 4506 -1688
rect 4572 -2088 4602 -1688
rect 4668 -2088 4698 -1688
rect 4764 -2088 4794 -1688
rect 4284 -2706 4314 -2306
rect 4380 -2706 4410 -2306
rect 4476 -2706 4506 -2306
rect 4572 -2706 4602 -2306
rect 4668 -2706 4698 -2306
rect 4764 -2706 4794 -2306
rect 5324 -2088 5354 -1688
rect 5420 -2088 5450 -1688
rect 5516 -2088 5546 -1688
rect 5612 -2088 5642 -1688
rect 5708 -2088 5738 -1688
rect 5804 -2088 5834 -1688
rect 5324 -2706 5354 -2306
rect 5420 -2706 5450 -2306
rect 5516 -2706 5546 -2306
rect 5612 -2706 5642 -2306
rect 5708 -2706 5738 -2306
rect 5804 -2706 5834 -2306
rect 6364 -2088 6394 -1688
rect 6460 -2088 6490 -1688
rect 6556 -2088 6586 -1688
rect 6652 -2088 6682 -1688
rect 6748 -2088 6778 -1688
rect 6844 -2088 6874 -1688
rect 6364 -2706 6394 -2306
rect 6460 -2706 6490 -2306
rect 6556 -2706 6586 -2306
rect 6652 -2706 6682 -2306
rect 6748 -2706 6778 -2306
rect 6844 -2706 6874 -2306
rect 7404 -2088 7434 -1688
rect 7500 -2088 7530 -1688
rect 7596 -2088 7626 -1688
rect 7692 -2088 7722 -1688
rect 7788 -2088 7818 -1688
rect 7884 -2088 7914 -1688
rect 7404 -2706 7434 -2306
rect 7500 -2706 7530 -2306
rect 7596 -2706 7626 -2306
rect 7692 -2706 7722 -2306
rect 7788 -2706 7818 -2306
rect 7884 -2706 7914 -2306
rect 8444 -2088 8474 -1688
rect 8540 -2088 8570 -1688
rect 8636 -2088 8666 -1688
rect 8732 -2088 8762 -1688
rect 8828 -2088 8858 -1688
rect 8924 -2088 8954 -1688
rect 8444 -2706 8474 -2306
rect 8540 -2706 8570 -2306
rect 8636 -2706 8666 -2306
rect 8732 -2706 8762 -2306
rect 8828 -2706 8858 -2306
rect 8924 -2706 8954 -2306
rect 11904 -2088 11934 -1688
rect 12000 -2088 12030 -1688
rect 12096 -2088 12126 -1688
rect 12192 -2088 12222 -1688
rect 12288 -2088 12318 -1688
rect 12384 -2088 12414 -1688
rect 11904 -2706 11934 -2306
rect 12000 -2706 12030 -2306
rect 12096 -2706 12126 -2306
rect 12192 -2706 12222 -2306
rect 12288 -2706 12318 -2306
rect 12384 -2706 12414 -2306
rect 12944 -2088 12974 -1688
rect 13040 -2088 13070 -1688
rect 13136 -2088 13166 -1688
rect 13232 -2088 13262 -1688
rect 13328 -2088 13358 -1688
rect 13424 -2088 13454 -1688
rect 12944 -2706 12974 -2306
rect 13040 -2706 13070 -2306
rect 13136 -2706 13166 -2306
rect 13232 -2706 13262 -2306
rect 13328 -2706 13358 -2306
rect 13424 -2706 13454 -2306
rect 13984 -2088 14014 -1688
rect 14080 -2088 14110 -1688
rect 14176 -2088 14206 -1688
rect 14272 -2088 14302 -1688
rect 14368 -2088 14398 -1688
rect 14464 -2088 14494 -1688
rect 13984 -2706 14014 -2306
rect 14080 -2706 14110 -2306
rect 14176 -2706 14206 -2306
rect 14272 -2706 14302 -2306
rect 14368 -2706 14398 -2306
rect 14464 -2706 14494 -2306
rect 15024 -2088 15054 -1688
rect 15120 -2088 15150 -1688
rect 15216 -2088 15246 -1688
rect 15312 -2088 15342 -1688
rect 15408 -2088 15438 -1688
rect 15504 -2088 15534 -1688
rect 15024 -2706 15054 -2306
rect 15120 -2706 15150 -2306
rect 15216 -2706 15246 -2306
rect 15312 -2706 15342 -2306
rect 15408 -2706 15438 -2306
rect 15504 -2706 15534 -2306
rect 16064 -2088 16094 -1688
rect 16160 -2088 16190 -1688
rect 16256 -2088 16286 -1688
rect 16352 -2088 16382 -1688
rect 16448 -2088 16478 -1688
rect 16544 -2088 16574 -1688
rect 16064 -2706 16094 -2306
rect 16160 -2706 16190 -2306
rect 16256 -2706 16286 -2306
rect 16352 -2706 16382 -2306
rect 16448 -2706 16478 -2306
rect 16544 -2706 16574 -2306
rect -7354 -3712 -7294 -3312
rect -7236 -3712 -7176 -3312
rect -7118 -3712 -7058 -3312
rect -7000 -3712 -6940 -3312
rect -6882 -3712 -6822 -3312
rect -6764 -3712 -6704 -3312
rect 4280 -3510 4340 -3110
rect 4398 -3510 4458 -3110
rect 4516 -3510 4576 -3110
rect 4634 -3510 4694 -3110
rect 4752 -3510 4812 -3110
rect 4870 -3510 4930 -3110
rect 5320 -3510 5380 -3110
rect 5438 -3510 5498 -3110
rect 5556 -3510 5616 -3110
rect 5674 -3510 5734 -3110
rect 5792 -3510 5852 -3110
rect 5910 -3510 5970 -3110
rect 6360 -3510 6420 -3110
rect 6478 -3510 6538 -3110
rect 6596 -3510 6656 -3110
rect 6714 -3510 6774 -3110
rect 6832 -3510 6892 -3110
rect 6950 -3510 7010 -3110
rect 7400 -3510 7460 -3110
rect 7518 -3510 7578 -3110
rect 7636 -3510 7696 -3110
rect 7754 -3510 7814 -3110
rect 7872 -3510 7932 -3110
rect 7990 -3510 8050 -3110
rect 8440 -3510 8500 -3110
rect 8558 -3510 8618 -3110
rect 8676 -3510 8736 -3110
rect 8794 -3510 8854 -3110
rect 8912 -3510 8972 -3110
rect 9030 -3510 9090 -3110
rect 11900 -3510 11960 -3110
rect 12018 -3510 12078 -3110
rect 12136 -3510 12196 -3110
rect 12254 -3510 12314 -3110
rect 12372 -3510 12432 -3110
rect 12490 -3510 12550 -3110
rect 12940 -3510 13000 -3110
rect 13058 -3510 13118 -3110
rect 13176 -3510 13236 -3110
rect 13294 -3510 13354 -3110
rect 13412 -3510 13472 -3110
rect 13530 -3510 13590 -3110
rect 13980 -3510 14040 -3110
rect 14098 -3510 14158 -3110
rect 14216 -3510 14276 -3110
rect 14334 -3510 14394 -3110
rect 14452 -3510 14512 -3110
rect 14570 -3510 14630 -3110
rect 15020 -3510 15080 -3110
rect 15138 -3510 15198 -3110
rect 15256 -3510 15316 -3110
rect 15374 -3510 15434 -3110
rect 15492 -3510 15552 -3110
rect 15610 -3510 15670 -3110
rect 16060 -3510 16120 -3110
rect 16178 -3510 16238 -3110
rect 16296 -3510 16356 -3110
rect 16414 -3510 16474 -3110
rect 16532 -3510 16592 -3110
rect 16650 -3510 16710 -3110
<< ndiff >>
rect -1042 3598 -980 3610
rect -1042 3222 -1030 3598
rect -996 3222 -980 3598
rect -1042 3210 -980 3222
rect -950 3598 -884 3610
rect -950 3222 -934 3598
rect -900 3222 -884 3598
rect -950 3210 -884 3222
rect -854 3598 -788 3610
rect -854 3222 -838 3598
rect -804 3222 -788 3598
rect -854 3210 -788 3222
rect -758 3598 -692 3610
rect -758 3222 -742 3598
rect -708 3222 -692 3598
rect -758 3210 -692 3222
rect -662 3598 -596 3610
rect -662 3222 -646 3598
rect -612 3222 -596 3598
rect -662 3210 -596 3222
rect -566 3598 -500 3610
rect -566 3222 -550 3598
rect -516 3222 -500 3598
rect -566 3210 -500 3222
rect -470 3598 -404 3610
rect -470 3222 -454 3598
rect -420 3222 -404 3598
rect -470 3210 -404 3222
rect -374 3598 -308 3610
rect -374 3222 -358 3598
rect -324 3222 -308 3598
rect -374 3210 -308 3222
rect -278 3598 -212 3610
rect -278 3222 -262 3598
rect -228 3222 -212 3598
rect -278 3210 -212 3222
rect -182 3598 -116 3610
rect -182 3222 -166 3598
rect -132 3222 -116 3598
rect -182 3210 -116 3222
rect -86 3598 -24 3610
rect -86 3222 -70 3598
rect -36 3222 -24 3598
rect -86 3210 -24 3222
rect 1758 3598 1820 3610
rect 1758 3222 1770 3598
rect 1804 3222 1820 3598
rect 1758 3210 1820 3222
rect 1850 3598 1916 3610
rect 1850 3222 1866 3598
rect 1900 3222 1916 3598
rect 1850 3210 1916 3222
rect 1946 3598 2012 3610
rect 1946 3222 1962 3598
rect 1996 3222 2012 3598
rect 1946 3210 2012 3222
rect 2042 3598 2108 3610
rect 2042 3222 2058 3598
rect 2092 3222 2108 3598
rect 2042 3210 2108 3222
rect 2138 3598 2204 3610
rect 2138 3222 2154 3598
rect 2188 3222 2204 3598
rect 2138 3210 2204 3222
rect 2234 3598 2300 3610
rect 2234 3222 2250 3598
rect 2284 3222 2300 3598
rect 2234 3210 2300 3222
rect 2330 3598 2396 3610
rect 2330 3222 2346 3598
rect 2380 3222 2396 3598
rect 2330 3210 2396 3222
rect 2426 3598 2492 3610
rect 2426 3222 2442 3598
rect 2476 3222 2492 3598
rect 2426 3210 2492 3222
rect 2522 3598 2588 3610
rect 2522 3222 2538 3598
rect 2572 3222 2588 3598
rect 2522 3210 2588 3222
rect 2618 3598 2684 3610
rect 2618 3222 2634 3598
rect 2668 3222 2684 3598
rect 2618 3210 2684 3222
rect 2714 3598 2776 3610
rect 2714 3222 2730 3598
rect 2764 3222 2776 3598
rect 2714 3210 2776 3222
rect 4422 5452 4484 5464
rect 4422 5076 4434 5452
rect 4468 5076 4484 5452
rect 4422 5064 4484 5076
rect 4514 5452 4580 5464
rect 4514 5076 4530 5452
rect 4564 5076 4580 5452
rect 4514 5064 4580 5076
rect 4610 5452 4676 5464
rect 4610 5076 4626 5452
rect 4660 5076 4676 5452
rect 4610 5064 4676 5076
rect 4706 5452 4772 5464
rect 4706 5076 4722 5452
rect 4756 5076 4772 5452
rect 4706 5064 4772 5076
rect 4802 5452 4868 5464
rect 4802 5076 4818 5452
rect 4852 5076 4868 5452
rect 4802 5064 4868 5076
rect 4898 5452 4964 5464
rect 4898 5076 4914 5452
rect 4948 5076 4964 5452
rect 4898 5064 4964 5076
rect 4994 5452 5060 5464
rect 4994 5076 5010 5452
rect 5044 5076 5060 5452
rect 4994 5064 5060 5076
rect 5090 5452 5156 5464
rect 5090 5076 5106 5452
rect 5140 5076 5156 5452
rect 5090 5064 5156 5076
rect 5186 5452 5252 5464
rect 5186 5076 5202 5452
rect 5236 5076 5252 5452
rect 5186 5064 5252 5076
rect 5282 5452 5348 5464
rect 5282 5076 5298 5452
rect 5332 5076 5348 5452
rect 5282 5064 5348 5076
rect 5378 5452 5444 5464
rect 5378 5076 5394 5452
rect 5428 5076 5444 5452
rect 5378 5064 5444 5076
rect 5474 5452 5540 5464
rect 5474 5076 5490 5452
rect 5524 5076 5540 5452
rect 5474 5064 5540 5076
rect 5570 5452 5636 5464
rect 5570 5076 5586 5452
rect 5620 5076 5636 5452
rect 5570 5064 5636 5076
rect 5666 5452 5732 5464
rect 5666 5076 5682 5452
rect 5716 5076 5732 5452
rect 5666 5064 5732 5076
rect 5762 5452 5828 5464
rect 5762 5076 5778 5452
rect 5812 5076 5828 5452
rect 5762 5064 5828 5076
rect 5858 5452 5924 5464
rect 5858 5076 5874 5452
rect 5908 5076 5924 5452
rect 5858 5064 5924 5076
rect 5954 5452 6020 5464
rect 5954 5076 5970 5452
rect 6004 5076 6020 5452
rect 5954 5064 6020 5076
rect 6050 5452 6116 5464
rect 6050 5076 6066 5452
rect 6100 5076 6116 5452
rect 6050 5064 6116 5076
rect 6146 5452 6212 5464
rect 6146 5076 6162 5452
rect 6196 5076 6212 5452
rect 6146 5064 6212 5076
rect 6242 5452 6308 5464
rect 6242 5076 6258 5452
rect 6292 5076 6308 5452
rect 6242 5064 6308 5076
rect 6338 5452 6404 5464
rect 6338 5076 6354 5452
rect 6388 5076 6404 5452
rect 6338 5064 6404 5076
rect 6434 5452 6500 5464
rect 6434 5076 6450 5452
rect 6484 5076 6500 5452
rect 6434 5064 6500 5076
rect 6530 5452 6596 5464
rect 6530 5076 6546 5452
rect 6580 5076 6596 5452
rect 6530 5064 6596 5076
rect 6626 5452 6692 5464
rect 6626 5076 6642 5452
rect 6676 5076 6692 5452
rect 6626 5064 6692 5076
rect 6722 5452 6788 5464
rect 6722 5076 6738 5452
rect 6772 5076 6788 5452
rect 6722 5064 6788 5076
rect 6818 5452 6884 5464
rect 6818 5076 6834 5452
rect 6868 5076 6884 5452
rect 6818 5064 6884 5076
rect 6914 5452 6980 5464
rect 6914 5076 6930 5452
rect 6964 5076 6980 5452
rect 6914 5064 6980 5076
rect 7010 5452 7076 5464
rect 7010 5076 7026 5452
rect 7060 5076 7076 5452
rect 7010 5064 7076 5076
rect 7106 5452 7172 5464
rect 7106 5076 7122 5452
rect 7156 5076 7172 5452
rect 7106 5064 7172 5076
rect 7202 5452 7268 5464
rect 7202 5076 7218 5452
rect 7252 5076 7268 5452
rect 7202 5064 7268 5076
rect 7298 5452 7360 5464
rect 7298 5076 7314 5452
rect 7348 5076 7360 5452
rect 7298 5064 7360 5076
rect 4422 4834 4484 4846
rect 4422 4458 4434 4834
rect 4468 4458 4484 4834
rect 4422 4446 4484 4458
rect 4514 4834 4580 4846
rect 4514 4458 4530 4834
rect 4564 4458 4580 4834
rect 4514 4446 4580 4458
rect 4610 4834 4676 4846
rect 4610 4458 4626 4834
rect 4660 4458 4676 4834
rect 4610 4446 4676 4458
rect 4706 4834 4772 4846
rect 4706 4458 4722 4834
rect 4756 4458 4772 4834
rect 4706 4446 4772 4458
rect 4802 4834 4868 4846
rect 4802 4458 4818 4834
rect 4852 4458 4868 4834
rect 4802 4446 4868 4458
rect 4898 4834 4964 4846
rect 4898 4458 4914 4834
rect 4948 4458 4964 4834
rect 4898 4446 4964 4458
rect 4994 4834 5060 4846
rect 4994 4458 5010 4834
rect 5044 4458 5060 4834
rect 4994 4446 5060 4458
rect 5090 4834 5156 4846
rect 5090 4458 5106 4834
rect 5140 4458 5156 4834
rect 5090 4446 5156 4458
rect 5186 4834 5252 4846
rect 5186 4458 5202 4834
rect 5236 4458 5252 4834
rect 5186 4446 5252 4458
rect 5282 4834 5348 4846
rect 5282 4458 5298 4834
rect 5332 4458 5348 4834
rect 5282 4446 5348 4458
rect 5378 4834 5444 4846
rect 5378 4458 5394 4834
rect 5428 4458 5444 4834
rect 5378 4446 5444 4458
rect 5474 4834 5540 4846
rect 5474 4458 5490 4834
rect 5524 4458 5540 4834
rect 5474 4446 5540 4458
rect 5570 4834 5636 4846
rect 5570 4458 5586 4834
rect 5620 4458 5636 4834
rect 5570 4446 5636 4458
rect 5666 4834 5732 4846
rect 5666 4458 5682 4834
rect 5716 4458 5732 4834
rect 5666 4446 5732 4458
rect 5762 4834 5828 4846
rect 5762 4458 5778 4834
rect 5812 4458 5828 4834
rect 5762 4446 5828 4458
rect 5858 4834 5924 4846
rect 5858 4458 5874 4834
rect 5908 4458 5924 4834
rect 5858 4446 5924 4458
rect 5954 4834 6020 4846
rect 5954 4458 5970 4834
rect 6004 4458 6020 4834
rect 5954 4446 6020 4458
rect 6050 4834 6116 4846
rect 6050 4458 6066 4834
rect 6100 4458 6116 4834
rect 6050 4446 6116 4458
rect 6146 4834 6212 4846
rect 6146 4458 6162 4834
rect 6196 4458 6212 4834
rect 6146 4446 6212 4458
rect 6242 4834 6308 4846
rect 6242 4458 6258 4834
rect 6292 4458 6308 4834
rect 6242 4446 6308 4458
rect 6338 4834 6404 4846
rect 6338 4458 6354 4834
rect 6388 4458 6404 4834
rect 6338 4446 6404 4458
rect 6434 4834 6500 4846
rect 6434 4458 6450 4834
rect 6484 4458 6500 4834
rect 6434 4446 6500 4458
rect 6530 4834 6596 4846
rect 6530 4458 6546 4834
rect 6580 4458 6596 4834
rect 6530 4446 6596 4458
rect 6626 4834 6692 4846
rect 6626 4458 6642 4834
rect 6676 4458 6692 4834
rect 6626 4446 6692 4458
rect 6722 4834 6788 4846
rect 6722 4458 6738 4834
rect 6772 4458 6788 4834
rect 6722 4446 6788 4458
rect 6818 4834 6884 4846
rect 6818 4458 6834 4834
rect 6868 4458 6884 4834
rect 6818 4446 6884 4458
rect 6914 4834 6980 4846
rect 6914 4458 6930 4834
rect 6964 4458 6980 4834
rect 6914 4446 6980 4458
rect 7010 4834 7076 4846
rect 7010 4458 7026 4834
rect 7060 4458 7076 4834
rect 7010 4446 7076 4458
rect 7106 4834 7172 4846
rect 7106 4458 7122 4834
rect 7156 4458 7172 4834
rect 7106 4446 7172 4458
rect 7202 4834 7268 4846
rect 7202 4458 7218 4834
rect 7252 4458 7268 4834
rect 7202 4446 7268 4458
rect 7298 4834 7360 4846
rect 7298 4458 7314 4834
rect 7348 4458 7360 4834
rect 7298 4446 7360 4458
rect 4422 4216 4484 4228
rect 4422 3840 4434 4216
rect 4468 3840 4484 4216
rect 4422 3828 4484 3840
rect 4514 4216 4580 4228
rect 4514 3840 4530 4216
rect 4564 3840 4580 4216
rect 4514 3828 4580 3840
rect 4610 4216 4676 4228
rect 4610 3840 4626 4216
rect 4660 3840 4676 4216
rect 4610 3828 4676 3840
rect 4706 4216 4772 4228
rect 4706 3840 4722 4216
rect 4756 3840 4772 4216
rect 4706 3828 4772 3840
rect 4802 4216 4868 4228
rect 4802 3840 4818 4216
rect 4852 3840 4868 4216
rect 4802 3828 4868 3840
rect 4898 4216 4964 4228
rect 4898 3840 4914 4216
rect 4948 3840 4964 4216
rect 4898 3828 4964 3840
rect 4994 4216 5060 4228
rect 4994 3840 5010 4216
rect 5044 3840 5060 4216
rect 4994 3828 5060 3840
rect 5090 4216 5156 4228
rect 5090 3840 5106 4216
rect 5140 3840 5156 4216
rect 5090 3828 5156 3840
rect 5186 4216 5252 4228
rect 5186 3840 5202 4216
rect 5236 3840 5252 4216
rect 5186 3828 5252 3840
rect 5282 4216 5348 4228
rect 5282 3840 5298 4216
rect 5332 3840 5348 4216
rect 5282 3828 5348 3840
rect 5378 4216 5444 4228
rect 5378 3840 5394 4216
rect 5428 3840 5444 4216
rect 5378 3828 5444 3840
rect 5474 4216 5540 4228
rect 5474 3840 5490 4216
rect 5524 3840 5540 4216
rect 5474 3828 5540 3840
rect 5570 4216 5636 4228
rect 5570 3840 5586 4216
rect 5620 3840 5636 4216
rect 5570 3828 5636 3840
rect 5666 4216 5732 4228
rect 5666 3840 5682 4216
rect 5716 3840 5732 4216
rect 5666 3828 5732 3840
rect 5762 4216 5828 4228
rect 5762 3840 5778 4216
rect 5812 3840 5828 4216
rect 5762 3828 5828 3840
rect 5858 4216 5924 4228
rect 5858 3840 5874 4216
rect 5908 3840 5924 4216
rect 5858 3828 5924 3840
rect 5954 4216 6020 4228
rect 5954 3840 5970 4216
rect 6004 3840 6020 4216
rect 5954 3828 6020 3840
rect 6050 4216 6116 4228
rect 6050 3840 6066 4216
rect 6100 3840 6116 4216
rect 6050 3828 6116 3840
rect 6146 4216 6212 4228
rect 6146 3840 6162 4216
rect 6196 3840 6212 4216
rect 6146 3828 6212 3840
rect 6242 4216 6308 4228
rect 6242 3840 6258 4216
rect 6292 3840 6308 4216
rect 6242 3828 6308 3840
rect 6338 4216 6404 4228
rect 6338 3840 6354 4216
rect 6388 3840 6404 4216
rect 6338 3828 6404 3840
rect 6434 4216 6500 4228
rect 6434 3840 6450 4216
rect 6484 3840 6500 4216
rect 6434 3828 6500 3840
rect 6530 4216 6596 4228
rect 6530 3840 6546 4216
rect 6580 3840 6596 4216
rect 6530 3828 6596 3840
rect 6626 4216 6692 4228
rect 6626 3840 6642 4216
rect 6676 3840 6692 4216
rect 6626 3828 6692 3840
rect 6722 4216 6788 4228
rect 6722 3840 6738 4216
rect 6772 3840 6788 4216
rect 6722 3828 6788 3840
rect 6818 4216 6884 4228
rect 6818 3840 6834 4216
rect 6868 3840 6884 4216
rect 6818 3828 6884 3840
rect 6914 4216 6980 4228
rect 6914 3840 6930 4216
rect 6964 3840 6980 4216
rect 6914 3828 6980 3840
rect 7010 4216 7076 4228
rect 7010 3840 7026 4216
rect 7060 3840 7076 4216
rect 7010 3828 7076 3840
rect 7106 4216 7172 4228
rect 7106 3840 7122 4216
rect 7156 3840 7172 4216
rect 7106 3828 7172 3840
rect 7202 4216 7268 4228
rect 7202 3840 7218 4216
rect 7252 3840 7268 4216
rect 7202 3828 7268 3840
rect 7298 4216 7360 4228
rect 7298 3840 7314 4216
rect 7348 3840 7360 4216
rect 7298 3828 7360 3840
rect 4422 3598 4484 3610
rect 4422 3222 4434 3598
rect 4468 3222 4484 3598
rect 4422 3210 4484 3222
rect 4514 3598 4580 3610
rect 4514 3222 4530 3598
rect 4564 3222 4580 3598
rect 4514 3210 4580 3222
rect 4610 3598 4676 3610
rect 4610 3222 4626 3598
rect 4660 3222 4676 3598
rect 4610 3210 4676 3222
rect 4706 3598 4772 3610
rect 4706 3222 4722 3598
rect 4756 3222 4772 3598
rect 4706 3210 4772 3222
rect 4802 3598 4868 3610
rect 4802 3222 4818 3598
rect 4852 3222 4868 3598
rect 4802 3210 4868 3222
rect 4898 3598 4964 3610
rect 4898 3222 4914 3598
rect 4948 3222 4964 3598
rect 4898 3210 4964 3222
rect 4994 3598 5060 3610
rect 4994 3222 5010 3598
rect 5044 3222 5060 3598
rect 4994 3210 5060 3222
rect 5090 3598 5156 3610
rect 5090 3222 5106 3598
rect 5140 3222 5156 3598
rect 5090 3210 5156 3222
rect 5186 3598 5252 3610
rect 5186 3222 5202 3598
rect 5236 3222 5252 3598
rect 5186 3210 5252 3222
rect 5282 3598 5348 3610
rect 5282 3222 5298 3598
rect 5332 3222 5348 3598
rect 5282 3210 5348 3222
rect 5378 3598 5444 3610
rect 5378 3222 5394 3598
rect 5428 3222 5444 3598
rect 5378 3210 5444 3222
rect 5474 3598 5540 3610
rect 5474 3222 5490 3598
rect 5524 3222 5540 3598
rect 5474 3210 5540 3222
rect 5570 3598 5636 3610
rect 5570 3222 5586 3598
rect 5620 3222 5636 3598
rect 5570 3210 5636 3222
rect 5666 3598 5732 3610
rect 5666 3222 5682 3598
rect 5716 3222 5732 3598
rect 5666 3210 5732 3222
rect 5762 3598 5828 3610
rect 5762 3222 5778 3598
rect 5812 3222 5828 3598
rect 5762 3210 5828 3222
rect 5858 3598 5924 3610
rect 5858 3222 5874 3598
rect 5908 3222 5924 3598
rect 5858 3210 5924 3222
rect 5954 3598 6020 3610
rect 5954 3222 5970 3598
rect 6004 3222 6020 3598
rect 5954 3210 6020 3222
rect 6050 3598 6116 3610
rect 6050 3222 6066 3598
rect 6100 3222 6116 3598
rect 6050 3210 6116 3222
rect 6146 3598 6212 3610
rect 6146 3222 6162 3598
rect 6196 3222 6212 3598
rect 6146 3210 6212 3222
rect 6242 3598 6308 3610
rect 6242 3222 6258 3598
rect 6292 3222 6308 3598
rect 6242 3210 6308 3222
rect 6338 3598 6404 3610
rect 6338 3222 6354 3598
rect 6388 3222 6404 3598
rect 6338 3210 6404 3222
rect 6434 3598 6500 3610
rect 6434 3222 6450 3598
rect 6484 3222 6500 3598
rect 6434 3210 6500 3222
rect 6530 3598 6596 3610
rect 6530 3222 6546 3598
rect 6580 3222 6596 3598
rect 6530 3210 6596 3222
rect 6626 3598 6692 3610
rect 6626 3222 6642 3598
rect 6676 3222 6692 3598
rect 6626 3210 6692 3222
rect 6722 3598 6788 3610
rect 6722 3222 6738 3598
rect 6772 3222 6788 3598
rect 6722 3210 6788 3222
rect 6818 3598 6884 3610
rect 6818 3222 6834 3598
rect 6868 3222 6884 3598
rect 6818 3210 6884 3222
rect 6914 3598 6980 3610
rect 6914 3222 6930 3598
rect 6964 3222 6980 3598
rect 6914 3210 6980 3222
rect 7010 3598 7076 3610
rect 7010 3222 7026 3598
rect 7060 3222 7076 3598
rect 7010 3210 7076 3222
rect 7106 3598 7172 3610
rect 7106 3222 7122 3598
rect 7156 3222 7172 3598
rect 7106 3210 7172 3222
rect 7202 3598 7268 3610
rect 7202 3222 7218 3598
rect 7252 3222 7268 3598
rect 7202 3210 7268 3222
rect 7298 3598 7360 3610
rect 7298 3222 7314 3598
rect 7348 3222 7360 3598
rect 7298 3210 7360 3222
rect 8062 5452 8124 5464
rect 8062 5076 8074 5452
rect 8108 5076 8124 5452
rect 8062 5064 8124 5076
rect 8154 5452 8220 5464
rect 8154 5076 8170 5452
rect 8204 5076 8220 5452
rect 8154 5064 8220 5076
rect 8250 5452 8316 5464
rect 8250 5076 8266 5452
rect 8300 5076 8316 5452
rect 8250 5064 8316 5076
rect 8346 5452 8412 5464
rect 8346 5076 8362 5452
rect 8396 5076 8412 5452
rect 8346 5064 8412 5076
rect 8442 5452 8508 5464
rect 8442 5076 8458 5452
rect 8492 5076 8508 5452
rect 8442 5064 8508 5076
rect 8538 5452 8604 5464
rect 8538 5076 8554 5452
rect 8588 5076 8604 5452
rect 8538 5064 8604 5076
rect 8634 5452 8700 5464
rect 8634 5076 8650 5452
rect 8684 5076 8700 5452
rect 8634 5064 8700 5076
rect 8730 5452 8796 5464
rect 8730 5076 8746 5452
rect 8780 5076 8796 5452
rect 8730 5064 8796 5076
rect 8826 5452 8892 5464
rect 8826 5076 8842 5452
rect 8876 5076 8892 5452
rect 8826 5064 8892 5076
rect 8922 5452 8988 5464
rect 8922 5076 8938 5452
rect 8972 5076 8988 5452
rect 8922 5064 8988 5076
rect 9018 5452 9084 5464
rect 9018 5076 9034 5452
rect 9068 5076 9084 5452
rect 9018 5064 9084 5076
rect 9114 5452 9180 5464
rect 9114 5076 9130 5452
rect 9164 5076 9180 5452
rect 9114 5064 9180 5076
rect 9210 5452 9276 5464
rect 9210 5076 9226 5452
rect 9260 5076 9276 5452
rect 9210 5064 9276 5076
rect 9306 5452 9372 5464
rect 9306 5076 9322 5452
rect 9356 5076 9372 5452
rect 9306 5064 9372 5076
rect 9402 5452 9468 5464
rect 9402 5076 9418 5452
rect 9452 5076 9468 5452
rect 9402 5064 9468 5076
rect 9498 5452 9564 5464
rect 9498 5076 9514 5452
rect 9548 5076 9564 5452
rect 9498 5064 9564 5076
rect 9594 5452 9660 5464
rect 9594 5076 9610 5452
rect 9644 5076 9660 5452
rect 9594 5064 9660 5076
rect 9690 5452 9756 5464
rect 9690 5076 9706 5452
rect 9740 5076 9756 5452
rect 9690 5064 9756 5076
rect 9786 5452 9852 5464
rect 9786 5076 9802 5452
rect 9836 5076 9852 5452
rect 9786 5064 9852 5076
rect 9882 5452 9948 5464
rect 9882 5076 9898 5452
rect 9932 5076 9948 5452
rect 9882 5064 9948 5076
rect 9978 5452 10044 5464
rect 9978 5076 9994 5452
rect 10028 5076 10044 5452
rect 9978 5064 10044 5076
rect 10074 5452 10140 5464
rect 10074 5076 10090 5452
rect 10124 5076 10140 5452
rect 10074 5064 10140 5076
rect 10170 5452 10236 5464
rect 10170 5076 10186 5452
rect 10220 5076 10236 5452
rect 10170 5064 10236 5076
rect 10266 5452 10332 5464
rect 10266 5076 10282 5452
rect 10316 5076 10332 5452
rect 10266 5064 10332 5076
rect 10362 5452 10428 5464
rect 10362 5076 10378 5452
rect 10412 5076 10428 5452
rect 10362 5064 10428 5076
rect 10458 5452 10524 5464
rect 10458 5076 10474 5452
rect 10508 5076 10524 5452
rect 10458 5064 10524 5076
rect 10554 5452 10620 5464
rect 10554 5076 10570 5452
rect 10604 5076 10620 5452
rect 10554 5064 10620 5076
rect 10650 5452 10716 5464
rect 10650 5076 10666 5452
rect 10700 5076 10716 5452
rect 10650 5064 10716 5076
rect 10746 5452 10812 5464
rect 10746 5076 10762 5452
rect 10796 5076 10812 5452
rect 10746 5064 10812 5076
rect 10842 5452 10908 5464
rect 10842 5076 10858 5452
rect 10892 5076 10908 5452
rect 10842 5064 10908 5076
rect 10938 5452 11000 5464
rect 10938 5076 10954 5452
rect 10988 5076 11000 5452
rect 10938 5064 11000 5076
rect 8062 4834 8124 4846
rect 8062 4458 8074 4834
rect 8108 4458 8124 4834
rect 8062 4446 8124 4458
rect 8154 4834 8220 4846
rect 8154 4458 8170 4834
rect 8204 4458 8220 4834
rect 8154 4446 8220 4458
rect 8250 4834 8316 4846
rect 8250 4458 8266 4834
rect 8300 4458 8316 4834
rect 8250 4446 8316 4458
rect 8346 4834 8412 4846
rect 8346 4458 8362 4834
rect 8396 4458 8412 4834
rect 8346 4446 8412 4458
rect 8442 4834 8508 4846
rect 8442 4458 8458 4834
rect 8492 4458 8508 4834
rect 8442 4446 8508 4458
rect 8538 4834 8604 4846
rect 8538 4458 8554 4834
rect 8588 4458 8604 4834
rect 8538 4446 8604 4458
rect 8634 4834 8700 4846
rect 8634 4458 8650 4834
rect 8684 4458 8700 4834
rect 8634 4446 8700 4458
rect 8730 4834 8796 4846
rect 8730 4458 8746 4834
rect 8780 4458 8796 4834
rect 8730 4446 8796 4458
rect 8826 4834 8892 4846
rect 8826 4458 8842 4834
rect 8876 4458 8892 4834
rect 8826 4446 8892 4458
rect 8922 4834 8988 4846
rect 8922 4458 8938 4834
rect 8972 4458 8988 4834
rect 8922 4446 8988 4458
rect 9018 4834 9084 4846
rect 9018 4458 9034 4834
rect 9068 4458 9084 4834
rect 9018 4446 9084 4458
rect 9114 4834 9180 4846
rect 9114 4458 9130 4834
rect 9164 4458 9180 4834
rect 9114 4446 9180 4458
rect 9210 4834 9276 4846
rect 9210 4458 9226 4834
rect 9260 4458 9276 4834
rect 9210 4446 9276 4458
rect 9306 4834 9372 4846
rect 9306 4458 9322 4834
rect 9356 4458 9372 4834
rect 9306 4446 9372 4458
rect 9402 4834 9468 4846
rect 9402 4458 9418 4834
rect 9452 4458 9468 4834
rect 9402 4446 9468 4458
rect 9498 4834 9564 4846
rect 9498 4458 9514 4834
rect 9548 4458 9564 4834
rect 9498 4446 9564 4458
rect 9594 4834 9660 4846
rect 9594 4458 9610 4834
rect 9644 4458 9660 4834
rect 9594 4446 9660 4458
rect 9690 4834 9756 4846
rect 9690 4458 9706 4834
rect 9740 4458 9756 4834
rect 9690 4446 9756 4458
rect 9786 4834 9852 4846
rect 9786 4458 9802 4834
rect 9836 4458 9852 4834
rect 9786 4446 9852 4458
rect 9882 4834 9948 4846
rect 9882 4458 9898 4834
rect 9932 4458 9948 4834
rect 9882 4446 9948 4458
rect 9978 4834 10044 4846
rect 9978 4458 9994 4834
rect 10028 4458 10044 4834
rect 9978 4446 10044 4458
rect 10074 4834 10140 4846
rect 10074 4458 10090 4834
rect 10124 4458 10140 4834
rect 10074 4446 10140 4458
rect 10170 4834 10236 4846
rect 10170 4458 10186 4834
rect 10220 4458 10236 4834
rect 10170 4446 10236 4458
rect 10266 4834 10332 4846
rect 10266 4458 10282 4834
rect 10316 4458 10332 4834
rect 10266 4446 10332 4458
rect 10362 4834 10428 4846
rect 10362 4458 10378 4834
rect 10412 4458 10428 4834
rect 10362 4446 10428 4458
rect 10458 4834 10524 4846
rect 10458 4458 10474 4834
rect 10508 4458 10524 4834
rect 10458 4446 10524 4458
rect 10554 4834 10620 4846
rect 10554 4458 10570 4834
rect 10604 4458 10620 4834
rect 10554 4446 10620 4458
rect 10650 4834 10716 4846
rect 10650 4458 10666 4834
rect 10700 4458 10716 4834
rect 10650 4446 10716 4458
rect 10746 4834 10812 4846
rect 10746 4458 10762 4834
rect 10796 4458 10812 4834
rect 10746 4446 10812 4458
rect 10842 4834 10908 4846
rect 10842 4458 10858 4834
rect 10892 4458 10908 4834
rect 10842 4446 10908 4458
rect 10938 4834 11000 4846
rect 10938 4458 10954 4834
rect 10988 4458 11000 4834
rect 10938 4446 11000 4458
rect 8062 4216 8124 4228
rect 8062 3840 8074 4216
rect 8108 3840 8124 4216
rect 8062 3828 8124 3840
rect 8154 4216 8220 4228
rect 8154 3840 8170 4216
rect 8204 3840 8220 4216
rect 8154 3828 8220 3840
rect 8250 4216 8316 4228
rect 8250 3840 8266 4216
rect 8300 3840 8316 4216
rect 8250 3828 8316 3840
rect 8346 4216 8412 4228
rect 8346 3840 8362 4216
rect 8396 3840 8412 4216
rect 8346 3828 8412 3840
rect 8442 4216 8508 4228
rect 8442 3840 8458 4216
rect 8492 3840 8508 4216
rect 8442 3828 8508 3840
rect 8538 4216 8604 4228
rect 8538 3840 8554 4216
rect 8588 3840 8604 4216
rect 8538 3828 8604 3840
rect 8634 4216 8700 4228
rect 8634 3840 8650 4216
rect 8684 3840 8700 4216
rect 8634 3828 8700 3840
rect 8730 4216 8796 4228
rect 8730 3840 8746 4216
rect 8780 3840 8796 4216
rect 8730 3828 8796 3840
rect 8826 4216 8892 4228
rect 8826 3840 8842 4216
rect 8876 3840 8892 4216
rect 8826 3828 8892 3840
rect 8922 4216 8988 4228
rect 8922 3840 8938 4216
rect 8972 3840 8988 4216
rect 8922 3828 8988 3840
rect 9018 4216 9084 4228
rect 9018 3840 9034 4216
rect 9068 3840 9084 4216
rect 9018 3828 9084 3840
rect 9114 4216 9180 4228
rect 9114 3840 9130 4216
rect 9164 3840 9180 4216
rect 9114 3828 9180 3840
rect 9210 4216 9276 4228
rect 9210 3840 9226 4216
rect 9260 3840 9276 4216
rect 9210 3828 9276 3840
rect 9306 4216 9372 4228
rect 9306 3840 9322 4216
rect 9356 3840 9372 4216
rect 9306 3828 9372 3840
rect 9402 4216 9468 4228
rect 9402 3840 9418 4216
rect 9452 3840 9468 4216
rect 9402 3828 9468 3840
rect 9498 4216 9564 4228
rect 9498 3840 9514 4216
rect 9548 3840 9564 4216
rect 9498 3828 9564 3840
rect 9594 4216 9660 4228
rect 9594 3840 9610 4216
rect 9644 3840 9660 4216
rect 9594 3828 9660 3840
rect 9690 4216 9756 4228
rect 9690 3840 9706 4216
rect 9740 3840 9756 4216
rect 9690 3828 9756 3840
rect 9786 4216 9852 4228
rect 9786 3840 9802 4216
rect 9836 3840 9852 4216
rect 9786 3828 9852 3840
rect 9882 4216 9948 4228
rect 9882 3840 9898 4216
rect 9932 3840 9948 4216
rect 9882 3828 9948 3840
rect 9978 4216 10044 4228
rect 9978 3840 9994 4216
rect 10028 3840 10044 4216
rect 9978 3828 10044 3840
rect 10074 4216 10140 4228
rect 10074 3840 10090 4216
rect 10124 3840 10140 4216
rect 10074 3828 10140 3840
rect 10170 4216 10236 4228
rect 10170 3840 10186 4216
rect 10220 3840 10236 4216
rect 10170 3828 10236 3840
rect 10266 4216 10332 4228
rect 10266 3840 10282 4216
rect 10316 3840 10332 4216
rect 10266 3828 10332 3840
rect 10362 4216 10428 4228
rect 10362 3840 10378 4216
rect 10412 3840 10428 4216
rect 10362 3828 10428 3840
rect 10458 4216 10524 4228
rect 10458 3840 10474 4216
rect 10508 3840 10524 4216
rect 10458 3828 10524 3840
rect 10554 4216 10620 4228
rect 10554 3840 10570 4216
rect 10604 3840 10620 4216
rect 10554 3828 10620 3840
rect 10650 4216 10716 4228
rect 10650 3840 10666 4216
rect 10700 3840 10716 4216
rect 10650 3828 10716 3840
rect 10746 4216 10812 4228
rect 10746 3840 10762 4216
rect 10796 3840 10812 4216
rect 10746 3828 10812 3840
rect 10842 4216 10908 4228
rect 10842 3840 10858 4216
rect 10892 3840 10908 4216
rect 10842 3828 10908 3840
rect 10938 4216 11000 4228
rect 10938 3840 10954 4216
rect 10988 3840 11000 4216
rect 10938 3828 11000 3840
rect 8062 3598 8124 3610
rect 8062 3222 8074 3598
rect 8108 3222 8124 3598
rect 8062 3210 8124 3222
rect 8154 3598 8220 3610
rect 8154 3222 8170 3598
rect 8204 3222 8220 3598
rect 8154 3210 8220 3222
rect 8250 3598 8316 3610
rect 8250 3222 8266 3598
rect 8300 3222 8316 3598
rect 8250 3210 8316 3222
rect 8346 3598 8412 3610
rect 8346 3222 8362 3598
rect 8396 3222 8412 3598
rect 8346 3210 8412 3222
rect 8442 3598 8508 3610
rect 8442 3222 8458 3598
rect 8492 3222 8508 3598
rect 8442 3210 8508 3222
rect 8538 3598 8604 3610
rect 8538 3222 8554 3598
rect 8588 3222 8604 3598
rect 8538 3210 8604 3222
rect 8634 3598 8700 3610
rect 8634 3222 8650 3598
rect 8684 3222 8700 3598
rect 8634 3210 8700 3222
rect 8730 3598 8796 3610
rect 8730 3222 8746 3598
rect 8780 3222 8796 3598
rect 8730 3210 8796 3222
rect 8826 3598 8892 3610
rect 8826 3222 8842 3598
rect 8876 3222 8892 3598
rect 8826 3210 8892 3222
rect 8922 3598 8988 3610
rect 8922 3222 8938 3598
rect 8972 3222 8988 3598
rect 8922 3210 8988 3222
rect 9018 3598 9084 3610
rect 9018 3222 9034 3598
rect 9068 3222 9084 3598
rect 9018 3210 9084 3222
rect 9114 3598 9180 3610
rect 9114 3222 9130 3598
rect 9164 3222 9180 3598
rect 9114 3210 9180 3222
rect 9210 3598 9276 3610
rect 9210 3222 9226 3598
rect 9260 3222 9276 3598
rect 9210 3210 9276 3222
rect 9306 3598 9372 3610
rect 9306 3222 9322 3598
rect 9356 3222 9372 3598
rect 9306 3210 9372 3222
rect 9402 3598 9468 3610
rect 9402 3222 9418 3598
rect 9452 3222 9468 3598
rect 9402 3210 9468 3222
rect 9498 3598 9564 3610
rect 9498 3222 9514 3598
rect 9548 3222 9564 3598
rect 9498 3210 9564 3222
rect 9594 3598 9660 3610
rect 9594 3222 9610 3598
rect 9644 3222 9660 3598
rect 9594 3210 9660 3222
rect 9690 3598 9756 3610
rect 9690 3222 9706 3598
rect 9740 3222 9756 3598
rect 9690 3210 9756 3222
rect 9786 3598 9852 3610
rect 9786 3222 9802 3598
rect 9836 3222 9852 3598
rect 9786 3210 9852 3222
rect 9882 3598 9948 3610
rect 9882 3222 9898 3598
rect 9932 3222 9948 3598
rect 9882 3210 9948 3222
rect 9978 3598 10044 3610
rect 9978 3222 9994 3598
rect 10028 3222 10044 3598
rect 9978 3210 10044 3222
rect 10074 3598 10140 3610
rect 10074 3222 10090 3598
rect 10124 3222 10140 3598
rect 10074 3210 10140 3222
rect 10170 3598 10236 3610
rect 10170 3222 10186 3598
rect 10220 3222 10236 3598
rect 10170 3210 10236 3222
rect 10266 3598 10332 3610
rect 10266 3222 10282 3598
rect 10316 3222 10332 3598
rect 10266 3210 10332 3222
rect 10362 3598 10428 3610
rect 10362 3222 10378 3598
rect 10412 3222 10428 3598
rect 10362 3210 10428 3222
rect 10458 3598 10524 3610
rect 10458 3222 10474 3598
rect 10508 3222 10524 3598
rect 10458 3210 10524 3222
rect 10554 3598 10620 3610
rect 10554 3222 10570 3598
rect 10604 3222 10620 3598
rect 10554 3210 10620 3222
rect 10650 3598 10716 3610
rect 10650 3222 10666 3598
rect 10700 3222 10716 3598
rect 10650 3210 10716 3222
rect 10746 3598 10812 3610
rect 10746 3222 10762 3598
rect 10796 3222 10812 3598
rect 10746 3210 10812 3222
rect 10842 3598 10908 3610
rect 10842 3222 10858 3598
rect 10892 3222 10908 3598
rect 10842 3210 10908 3222
rect 10938 3598 11000 3610
rect 10938 3222 10954 3598
rect 10988 3222 11000 3598
rect 10938 3210 11000 3222
rect 12042 5452 12104 5464
rect 12042 5076 12054 5452
rect 12088 5076 12104 5452
rect 12042 5064 12104 5076
rect 12134 5452 12200 5464
rect 12134 5076 12150 5452
rect 12184 5076 12200 5452
rect 12134 5064 12200 5076
rect 12230 5452 12296 5464
rect 12230 5076 12246 5452
rect 12280 5076 12296 5452
rect 12230 5064 12296 5076
rect 12326 5452 12392 5464
rect 12326 5076 12342 5452
rect 12376 5076 12392 5452
rect 12326 5064 12392 5076
rect 12422 5452 12488 5464
rect 12422 5076 12438 5452
rect 12472 5076 12488 5452
rect 12422 5064 12488 5076
rect 12518 5452 12584 5464
rect 12518 5076 12534 5452
rect 12568 5076 12584 5452
rect 12518 5064 12584 5076
rect 12614 5452 12680 5464
rect 12614 5076 12630 5452
rect 12664 5076 12680 5452
rect 12614 5064 12680 5076
rect 12710 5452 12776 5464
rect 12710 5076 12726 5452
rect 12760 5076 12776 5452
rect 12710 5064 12776 5076
rect 12806 5452 12872 5464
rect 12806 5076 12822 5452
rect 12856 5076 12872 5452
rect 12806 5064 12872 5076
rect 12902 5452 12968 5464
rect 12902 5076 12918 5452
rect 12952 5076 12968 5452
rect 12902 5064 12968 5076
rect 12998 5452 13064 5464
rect 12998 5076 13014 5452
rect 13048 5076 13064 5452
rect 12998 5064 13064 5076
rect 13094 5452 13160 5464
rect 13094 5076 13110 5452
rect 13144 5076 13160 5452
rect 13094 5064 13160 5076
rect 13190 5452 13256 5464
rect 13190 5076 13206 5452
rect 13240 5076 13256 5452
rect 13190 5064 13256 5076
rect 13286 5452 13352 5464
rect 13286 5076 13302 5452
rect 13336 5076 13352 5452
rect 13286 5064 13352 5076
rect 13382 5452 13448 5464
rect 13382 5076 13398 5452
rect 13432 5076 13448 5452
rect 13382 5064 13448 5076
rect 13478 5452 13544 5464
rect 13478 5076 13494 5452
rect 13528 5076 13544 5452
rect 13478 5064 13544 5076
rect 13574 5452 13640 5464
rect 13574 5076 13590 5452
rect 13624 5076 13640 5452
rect 13574 5064 13640 5076
rect 13670 5452 13736 5464
rect 13670 5076 13686 5452
rect 13720 5076 13736 5452
rect 13670 5064 13736 5076
rect 13766 5452 13832 5464
rect 13766 5076 13782 5452
rect 13816 5076 13832 5452
rect 13766 5064 13832 5076
rect 13862 5452 13928 5464
rect 13862 5076 13878 5452
rect 13912 5076 13928 5452
rect 13862 5064 13928 5076
rect 13958 5452 14024 5464
rect 13958 5076 13974 5452
rect 14008 5076 14024 5452
rect 13958 5064 14024 5076
rect 14054 5452 14120 5464
rect 14054 5076 14070 5452
rect 14104 5076 14120 5452
rect 14054 5064 14120 5076
rect 14150 5452 14216 5464
rect 14150 5076 14166 5452
rect 14200 5076 14216 5452
rect 14150 5064 14216 5076
rect 14246 5452 14312 5464
rect 14246 5076 14262 5452
rect 14296 5076 14312 5452
rect 14246 5064 14312 5076
rect 14342 5452 14408 5464
rect 14342 5076 14358 5452
rect 14392 5076 14408 5452
rect 14342 5064 14408 5076
rect 14438 5452 14504 5464
rect 14438 5076 14454 5452
rect 14488 5076 14504 5452
rect 14438 5064 14504 5076
rect 14534 5452 14600 5464
rect 14534 5076 14550 5452
rect 14584 5076 14600 5452
rect 14534 5064 14600 5076
rect 14630 5452 14696 5464
rect 14630 5076 14646 5452
rect 14680 5076 14696 5452
rect 14630 5064 14696 5076
rect 14726 5452 14792 5464
rect 14726 5076 14742 5452
rect 14776 5076 14792 5452
rect 14726 5064 14792 5076
rect 14822 5452 14888 5464
rect 14822 5076 14838 5452
rect 14872 5076 14888 5452
rect 14822 5064 14888 5076
rect 14918 5452 14980 5464
rect 14918 5076 14934 5452
rect 14968 5076 14980 5452
rect 14918 5064 14980 5076
rect 12042 4834 12104 4846
rect 12042 4458 12054 4834
rect 12088 4458 12104 4834
rect 12042 4446 12104 4458
rect 12134 4834 12200 4846
rect 12134 4458 12150 4834
rect 12184 4458 12200 4834
rect 12134 4446 12200 4458
rect 12230 4834 12296 4846
rect 12230 4458 12246 4834
rect 12280 4458 12296 4834
rect 12230 4446 12296 4458
rect 12326 4834 12392 4846
rect 12326 4458 12342 4834
rect 12376 4458 12392 4834
rect 12326 4446 12392 4458
rect 12422 4834 12488 4846
rect 12422 4458 12438 4834
rect 12472 4458 12488 4834
rect 12422 4446 12488 4458
rect 12518 4834 12584 4846
rect 12518 4458 12534 4834
rect 12568 4458 12584 4834
rect 12518 4446 12584 4458
rect 12614 4834 12680 4846
rect 12614 4458 12630 4834
rect 12664 4458 12680 4834
rect 12614 4446 12680 4458
rect 12710 4834 12776 4846
rect 12710 4458 12726 4834
rect 12760 4458 12776 4834
rect 12710 4446 12776 4458
rect 12806 4834 12872 4846
rect 12806 4458 12822 4834
rect 12856 4458 12872 4834
rect 12806 4446 12872 4458
rect 12902 4834 12968 4846
rect 12902 4458 12918 4834
rect 12952 4458 12968 4834
rect 12902 4446 12968 4458
rect 12998 4834 13064 4846
rect 12998 4458 13014 4834
rect 13048 4458 13064 4834
rect 12998 4446 13064 4458
rect 13094 4834 13160 4846
rect 13094 4458 13110 4834
rect 13144 4458 13160 4834
rect 13094 4446 13160 4458
rect 13190 4834 13256 4846
rect 13190 4458 13206 4834
rect 13240 4458 13256 4834
rect 13190 4446 13256 4458
rect 13286 4834 13352 4846
rect 13286 4458 13302 4834
rect 13336 4458 13352 4834
rect 13286 4446 13352 4458
rect 13382 4834 13448 4846
rect 13382 4458 13398 4834
rect 13432 4458 13448 4834
rect 13382 4446 13448 4458
rect 13478 4834 13544 4846
rect 13478 4458 13494 4834
rect 13528 4458 13544 4834
rect 13478 4446 13544 4458
rect 13574 4834 13640 4846
rect 13574 4458 13590 4834
rect 13624 4458 13640 4834
rect 13574 4446 13640 4458
rect 13670 4834 13736 4846
rect 13670 4458 13686 4834
rect 13720 4458 13736 4834
rect 13670 4446 13736 4458
rect 13766 4834 13832 4846
rect 13766 4458 13782 4834
rect 13816 4458 13832 4834
rect 13766 4446 13832 4458
rect 13862 4834 13928 4846
rect 13862 4458 13878 4834
rect 13912 4458 13928 4834
rect 13862 4446 13928 4458
rect 13958 4834 14024 4846
rect 13958 4458 13974 4834
rect 14008 4458 14024 4834
rect 13958 4446 14024 4458
rect 14054 4834 14120 4846
rect 14054 4458 14070 4834
rect 14104 4458 14120 4834
rect 14054 4446 14120 4458
rect 14150 4834 14216 4846
rect 14150 4458 14166 4834
rect 14200 4458 14216 4834
rect 14150 4446 14216 4458
rect 14246 4834 14312 4846
rect 14246 4458 14262 4834
rect 14296 4458 14312 4834
rect 14246 4446 14312 4458
rect 14342 4834 14408 4846
rect 14342 4458 14358 4834
rect 14392 4458 14408 4834
rect 14342 4446 14408 4458
rect 14438 4834 14504 4846
rect 14438 4458 14454 4834
rect 14488 4458 14504 4834
rect 14438 4446 14504 4458
rect 14534 4834 14600 4846
rect 14534 4458 14550 4834
rect 14584 4458 14600 4834
rect 14534 4446 14600 4458
rect 14630 4834 14696 4846
rect 14630 4458 14646 4834
rect 14680 4458 14696 4834
rect 14630 4446 14696 4458
rect 14726 4834 14792 4846
rect 14726 4458 14742 4834
rect 14776 4458 14792 4834
rect 14726 4446 14792 4458
rect 14822 4834 14888 4846
rect 14822 4458 14838 4834
rect 14872 4458 14888 4834
rect 14822 4446 14888 4458
rect 14918 4834 14980 4846
rect 14918 4458 14934 4834
rect 14968 4458 14980 4834
rect 14918 4446 14980 4458
rect 12042 4216 12104 4228
rect 12042 3840 12054 4216
rect 12088 3840 12104 4216
rect 12042 3828 12104 3840
rect 12134 4216 12200 4228
rect 12134 3840 12150 4216
rect 12184 3840 12200 4216
rect 12134 3828 12200 3840
rect 12230 4216 12296 4228
rect 12230 3840 12246 4216
rect 12280 3840 12296 4216
rect 12230 3828 12296 3840
rect 12326 4216 12392 4228
rect 12326 3840 12342 4216
rect 12376 3840 12392 4216
rect 12326 3828 12392 3840
rect 12422 4216 12488 4228
rect 12422 3840 12438 4216
rect 12472 3840 12488 4216
rect 12422 3828 12488 3840
rect 12518 4216 12584 4228
rect 12518 3840 12534 4216
rect 12568 3840 12584 4216
rect 12518 3828 12584 3840
rect 12614 4216 12680 4228
rect 12614 3840 12630 4216
rect 12664 3840 12680 4216
rect 12614 3828 12680 3840
rect 12710 4216 12776 4228
rect 12710 3840 12726 4216
rect 12760 3840 12776 4216
rect 12710 3828 12776 3840
rect 12806 4216 12872 4228
rect 12806 3840 12822 4216
rect 12856 3840 12872 4216
rect 12806 3828 12872 3840
rect 12902 4216 12968 4228
rect 12902 3840 12918 4216
rect 12952 3840 12968 4216
rect 12902 3828 12968 3840
rect 12998 4216 13064 4228
rect 12998 3840 13014 4216
rect 13048 3840 13064 4216
rect 12998 3828 13064 3840
rect 13094 4216 13160 4228
rect 13094 3840 13110 4216
rect 13144 3840 13160 4216
rect 13094 3828 13160 3840
rect 13190 4216 13256 4228
rect 13190 3840 13206 4216
rect 13240 3840 13256 4216
rect 13190 3828 13256 3840
rect 13286 4216 13352 4228
rect 13286 3840 13302 4216
rect 13336 3840 13352 4216
rect 13286 3828 13352 3840
rect 13382 4216 13448 4228
rect 13382 3840 13398 4216
rect 13432 3840 13448 4216
rect 13382 3828 13448 3840
rect 13478 4216 13544 4228
rect 13478 3840 13494 4216
rect 13528 3840 13544 4216
rect 13478 3828 13544 3840
rect 13574 4216 13640 4228
rect 13574 3840 13590 4216
rect 13624 3840 13640 4216
rect 13574 3828 13640 3840
rect 13670 4216 13736 4228
rect 13670 3840 13686 4216
rect 13720 3840 13736 4216
rect 13670 3828 13736 3840
rect 13766 4216 13832 4228
rect 13766 3840 13782 4216
rect 13816 3840 13832 4216
rect 13766 3828 13832 3840
rect 13862 4216 13928 4228
rect 13862 3840 13878 4216
rect 13912 3840 13928 4216
rect 13862 3828 13928 3840
rect 13958 4216 14024 4228
rect 13958 3840 13974 4216
rect 14008 3840 14024 4216
rect 13958 3828 14024 3840
rect 14054 4216 14120 4228
rect 14054 3840 14070 4216
rect 14104 3840 14120 4216
rect 14054 3828 14120 3840
rect 14150 4216 14216 4228
rect 14150 3840 14166 4216
rect 14200 3840 14216 4216
rect 14150 3828 14216 3840
rect 14246 4216 14312 4228
rect 14246 3840 14262 4216
rect 14296 3840 14312 4216
rect 14246 3828 14312 3840
rect 14342 4216 14408 4228
rect 14342 3840 14358 4216
rect 14392 3840 14408 4216
rect 14342 3828 14408 3840
rect 14438 4216 14504 4228
rect 14438 3840 14454 4216
rect 14488 3840 14504 4216
rect 14438 3828 14504 3840
rect 14534 4216 14600 4228
rect 14534 3840 14550 4216
rect 14584 3840 14600 4216
rect 14534 3828 14600 3840
rect 14630 4216 14696 4228
rect 14630 3840 14646 4216
rect 14680 3840 14696 4216
rect 14630 3828 14696 3840
rect 14726 4216 14792 4228
rect 14726 3840 14742 4216
rect 14776 3840 14792 4216
rect 14726 3828 14792 3840
rect 14822 4216 14888 4228
rect 14822 3840 14838 4216
rect 14872 3840 14888 4216
rect 14822 3828 14888 3840
rect 14918 4216 14980 4228
rect 14918 3840 14934 4216
rect 14968 3840 14980 4216
rect 14918 3828 14980 3840
rect 12042 3598 12104 3610
rect 12042 3222 12054 3598
rect 12088 3222 12104 3598
rect 12042 3210 12104 3222
rect 12134 3598 12200 3610
rect 12134 3222 12150 3598
rect 12184 3222 12200 3598
rect 12134 3210 12200 3222
rect 12230 3598 12296 3610
rect 12230 3222 12246 3598
rect 12280 3222 12296 3598
rect 12230 3210 12296 3222
rect 12326 3598 12392 3610
rect 12326 3222 12342 3598
rect 12376 3222 12392 3598
rect 12326 3210 12392 3222
rect 12422 3598 12488 3610
rect 12422 3222 12438 3598
rect 12472 3222 12488 3598
rect 12422 3210 12488 3222
rect 12518 3598 12584 3610
rect 12518 3222 12534 3598
rect 12568 3222 12584 3598
rect 12518 3210 12584 3222
rect 12614 3598 12680 3610
rect 12614 3222 12630 3598
rect 12664 3222 12680 3598
rect 12614 3210 12680 3222
rect 12710 3598 12776 3610
rect 12710 3222 12726 3598
rect 12760 3222 12776 3598
rect 12710 3210 12776 3222
rect 12806 3598 12872 3610
rect 12806 3222 12822 3598
rect 12856 3222 12872 3598
rect 12806 3210 12872 3222
rect 12902 3598 12968 3610
rect 12902 3222 12918 3598
rect 12952 3222 12968 3598
rect 12902 3210 12968 3222
rect 12998 3598 13064 3610
rect 12998 3222 13014 3598
rect 13048 3222 13064 3598
rect 12998 3210 13064 3222
rect 13094 3598 13160 3610
rect 13094 3222 13110 3598
rect 13144 3222 13160 3598
rect 13094 3210 13160 3222
rect 13190 3598 13256 3610
rect 13190 3222 13206 3598
rect 13240 3222 13256 3598
rect 13190 3210 13256 3222
rect 13286 3598 13352 3610
rect 13286 3222 13302 3598
rect 13336 3222 13352 3598
rect 13286 3210 13352 3222
rect 13382 3598 13448 3610
rect 13382 3222 13398 3598
rect 13432 3222 13448 3598
rect 13382 3210 13448 3222
rect 13478 3598 13544 3610
rect 13478 3222 13494 3598
rect 13528 3222 13544 3598
rect 13478 3210 13544 3222
rect 13574 3598 13640 3610
rect 13574 3222 13590 3598
rect 13624 3222 13640 3598
rect 13574 3210 13640 3222
rect 13670 3598 13736 3610
rect 13670 3222 13686 3598
rect 13720 3222 13736 3598
rect 13670 3210 13736 3222
rect 13766 3598 13832 3610
rect 13766 3222 13782 3598
rect 13816 3222 13832 3598
rect 13766 3210 13832 3222
rect 13862 3598 13928 3610
rect 13862 3222 13878 3598
rect 13912 3222 13928 3598
rect 13862 3210 13928 3222
rect 13958 3598 14024 3610
rect 13958 3222 13974 3598
rect 14008 3222 14024 3598
rect 13958 3210 14024 3222
rect 14054 3598 14120 3610
rect 14054 3222 14070 3598
rect 14104 3222 14120 3598
rect 14054 3210 14120 3222
rect 14150 3598 14216 3610
rect 14150 3222 14166 3598
rect 14200 3222 14216 3598
rect 14150 3210 14216 3222
rect 14246 3598 14312 3610
rect 14246 3222 14262 3598
rect 14296 3222 14312 3598
rect 14246 3210 14312 3222
rect 14342 3598 14408 3610
rect 14342 3222 14358 3598
rect 14392 3222 14408 3598
rect 14342 3210 14408 3222
rect 14438 3598 14504 3610
rect 14438 3222 14454 3598
rect 14488 3222 14504 3598
rect 14438 3210 14504 3222
rect 14534 3598 14600 3610
rect 14534 3222 14550 3598
rect 14584 3222 14600 3598
rect 14534 3210 14600 3222
rect 14630 3598 14696 3610
rect 14630 3222 14646 3598
rect 14680 3222 14696 3598
rect 14630 3210 14696 3222
rect 14726 3598 14792 3610
rect 14726 3222 14742 3598
rect 14776 3222 14792 3598
rect 14726 3210 14792 3222
rect 14822 3598 14888 3610
rect 14822 3222 14838 3598
rect 14872 3222 14888 3598
rect 14822 3210 14888 3222
rect 14918 3598 14980 3610
rect 14918 3222 14934 3598
rect 14968 3222 14980 3598
rect 14918 3210 14980 3222
rect 15682 5452 15744 5464
rect 15682 5076 15694 5452
rect 15728 5076 15744 5452
rect 15682 5064 15744 5076
rect 15774 5452 15840 5464
rect 15774 5076 15790 5452
rect 15824 5076 15840 5452
rect 15774 5064 15840 5076
rect 15870 5452 15936 5464
rect 15870 5076 15886 5452
rect 15920 5076 15936 5452
rect 15870 5064 15936 5076
rect 15966 5452 16032 5464
rect 15966 5076 15982 5452
rect 16016 5076 16032 5452
rect 15966 5064 16032 5076
rect 16062 5452 16128 5464
rect 16062 5076 16078 5452
rect 16112 5076 16128 5452
rect 16062 5064 16128 5076
rect 16158 5452 16224 5464
rect 16158 5076 16174 5452
rect 16208 5076 16224 5452
rect 16158 5064 16224 5076
rect 16254 5452 16320 5464
rect 16254 5076 16270 5452
rect 16304 5076 16320 5452
rect 16254 5064 16320 5076
rect 16350 5452 16416 5464
rect 16350 5076 16366 5452
rect 16400 5076 16416 5452
rect 16350 5064 16416 5076
rect 16446 5452 16512 5464
rect 16446 5076 16462 5452
rect 16496 5076 16512 5452
rect 16446 5064 16512 5076
rect 16542 5452 16608 5464
rect 16542 5076 16558 5452
rect 16592 5076 16608 5452
rect 16542 5064 16608 5076
rect 16638 5452 16704 5464
rect 16638 5076 16654 5452
rect 16688 5076 16704 5452
rect 16638 5064 16704 5076
rect 16734 5452 16800 5464
rect 16734 5076 16750 5452
rect 16784 5076 16800 5452
rect 16734 5064 16800 5076
rect 16830 5452 16896 5464
rect 16830 5076 16846 5452
rect 16880 5076 16896 5452
rect 16830 5064 16896 5076
rect 16926 5452 16992 5464
rect 16926 5076 16942 5452
rect 16976 5076 16992 5452
rect 16926 5064 16992 5076
rect 17022 5452 17088 5464
rect 17022 5076 17038 5452
rect 17072 5076 17088 5452
rect 17022 5064 17088 5076
rect 17118 5452 17184 5464
rect 17118 5076 17134 5452
rect 17168 5076 17184 5452
rect 17118 5064 17184 5076
rect 17214 5452 17280 5464
rect 17214 5076 17230 5452
rect 17264 5076 17280 5452
rect 17214 5064 17280 5076
rect 17310 5452 17376 5464
rect 17310 5076 17326 5452
rect 17360 5076 17376 5452
rect 17310 5064 17376 5076
rect 17406 5452 17472 5464
rect 17406 5076 17422 5452
rect 17456 5076 17472 5452
rect 17406 5064 17472 5076
rect 17502 5452 17568 5464
rect 17502 5076 17518 5452
rect 17552 5076 17568 5452
rect 17502 5064 17568 5076
rect 17598 5452 17664 5464
rect 17598 5076 17614 5452
rect 17648 5076 17664 5452
rect 17598 5064 17664 5076
rect 17694 5452 17760 5464
rect 17694 5076 17710 5452
rect 17744 5076 17760 5452
rect 17694 5064 17760 5076
rect 17790 5452 17856 5464
rect 17790 5076 17806 5452
rect 17840 5076 17856 5452
rect 17790 5064 17856 5076
rect 17886 5452 17952 5464
rect 17886 5076 17902 5452
rect 17936 5076 17952 5452
rect 17886 5064 17952 5076
rect 17982 5452 18048 5464
rect 17982 5076 17998 5452
rect 18032 5076 18048 5452
rect 17982 5064 18048 5076
rect 18078 5452 18144 5464
rect 18078 5076 18094 5452
rect 18128 5076 18144 5452
rect 18078 5064 18144 5076
rect 18174 5452 18240 5464
rect 18174 5076 18190 5452
rect 18224 5076 18240 5452
rect 18174 5064 18240 5076
rect 18270 5452 18336 5464
rect 18270 5076 18286 5452
rect 18320 5076 18336 5452
rect 18270 5064 18336 5076
rect 18366 5452 18432 5464
rect 18366 5076 18382 5452
rect 18416 5076 18432 5452
rect 18366 5064 18432 5076
rect 18462 5452 18528 5464
rect 18462 5076 18478 5452
rect 18512 5076 18528 5452
rect 18462 5064 18528 5076
rect 18558 5452 18620 5464
rect 18558 5076 18574 5452
rect 18608 5076 18620 5452
rect 18558 5064 18620 5076
rect 15682 4834 15744 4846
rect 15682 4458 15694 4834
rect 15728 4458 15744 4834
rect 15682 4446 15744 4458
rect 15774 4834 15840 4846
rect 15774 4458 15790 4834
rect 15824 4458 15840 4834
rect 15774 4446 15840 4458
rect 15870 4834 15936 4846
rect 15870 4458 15886 4834
rect 15920 4458 15936 4834
rect 15870 4446 15936 4458
rect 15966 4834 16032 4846
rect 15966 4458 15982 4834
rect 16016 4458 16032 4834
rect 15966 4446 16032 4458
rect 16062 4834 16128 4846
rect 16062 4458 16078 4834
rect 16112 4458 16128 4834
rect 16062 4446 16128 4458
rect 16158 4834 16224 4846
rect 16158 4458 16174 4834
rect 16208 4458 16224 4834
rect 16158 4446 16224 4458
rect 16254 4834 16320 4846
rect 16254 4458 16270 4834
rect 16304 4458 16320 4834
rect 16254 4446 16320 4458
rect 16350 4834 16416 4846
rect 16350 4458 16366 4834
rect 16400 4458 16416 4834
rect 16350 4446 16416 4458
rect 16446 4834 16512 4846
rect 16446 4458 16462 4834
rect 16496 4458 16512 4834
rect 16446 4446 16512 4458
rect 16542 4834 16608 4846
rect 16542 4458 16558 4834
rect 16592 4458 16608 4834
rect 16542 4446 16608 4458
rect 16638 4834 16704 4846
rect 16638 4458 16654 4834
rect 16688 4458 16704 4834
rect 16638 4446 16704 4458
rect 16734 4834 16800 4846
rect 16734 4458 16750 4834
rect 16784 4458 16800 4834
rect 16734 4446 16800 4458
rect 16830 4834 16896 4846
rect 16830 4458 16846 4834
rect 16880 4458 16896 4834
rect 16830 4446 16896 4458
rect 16926 4834 16992 4846
rect 16926 4458 16942 4834
rect 16976 4458 16992 4834
rect 16926 4446 16992 4458
rect 17022 4834 17088 4846
rect 17022 4458 17038 4834
rect 17072 4458 17088 4834
rect 17022 4446 17088 4458
rect 17118 4834 17184 4846
rect 17118 4458 17134 4834
rect 17168 4458 17184 4834
rect 17118 4446 17184 4458
rect 17214 4834 17280 4846
rect 17214 4458 17230 4834
rect 17264 4458 17280 4834
rect 17214 4446 17280 4458
rect 17310 4834 17376 4846
rect 17310 4458 17326 4834
rect 17360 4458 17376 4834
rect 17310 4446 17376 4458
rect 17406 4834 17472 4846
rect 17406 4458 17422 4834
rect 17456 4458 17472 4834
rect 17406 4446 17472 4458
rect 17502 4834 17568 4846
rect 17502 4458 17518 4834
rect 17552 4458 17568 4834
rect 17502 4446 17568 4458
rect 17598 4834 17664 4846
rect 17598 4458 17614 4834
rect 17648 4458 17664 4834
rect 17598 4446 17664 4458
rect 17694 4834 17760 4846
rect 17694 4458 17710 4834
rect 17744 4458 17760 4834
rect 17694 4446 17760 4458
rect 17790 4834 17856 4846
rect 17790 4458 17806 4834
rect 17840 4458 17856 4834
rect 17790 4446 17856 4458
rect 17886 4834 17952 4846
rect 17886 4458 17902 4834
rect 17936 4458 17952 4834
rect 17886 4446 17952 4458
rect 17982 4834 18048 4846
rect 17982 4458 17998 4834
rect 18032 4458 18048 4834
rect 17982 4446 18048 4458
rect 18078 4834 18144 4846
rect 18078 4458 18094 4834
rect 18128 4458 18144 4834
rect 18078 4446 18144 4458
rect 18174 4834 18240 4846
rect 18174 4458 18190 4834
rect 18224 4458 18240 4834
rect 18174 4446 18240 4458
rect 18270 4834 18336 4846
rect 18270 4458 18286 4834
rect 18320 4458 18336 4834
rect 18270 4446 18336 4458
rect 18366 4834 18432 4846
rect 18366 4458 18382 4834
rect 18416 4458 18432 4834
rect 18366 4446 18432 4458
rect 18462 4834 18528 4846
rect 18462 4458 18478 4834
rect 18512 4458 18528 4834
rect 18462 4446 18528 4458
rect 18558 4834 18620 4846
rect 18558 4458 18574 4834
rect 18608 4458 18620 4834
rect 18558 4446 18620 4458
rect 15682 4216 15744 4228
rect 15682 3840 15694 4216
rect 15728 3840 15744 4216
rect 15682 3828 15744 3840
rect 15774 4216 15840 4228
rect 15774 3840 15790 4216
rect 15824 3840 15840 4216
rect 15774 3828 15840 3840
rect 15870 4216 15936 4228
rect 15870 3840 15886 4216
rect 15920 3840 15936 4216
rect 15870 3828 15936 3840
rect 15966 4216 16032 4228
rect 15966 3840 15982 4216
rect 16016 3840 16032 4216
rect 15966 3828 16032 3840
rect 16062 4216 16128 4228
rect 16062 3840 16078 4216
rect 16112 3840 16128 4216
rect 16062 3828 16128 3840
rect 16158 4216 16224 4228
rect 16158 3840 16174 4216
rect 16208 3840 16224 4216
rect 16158 3828 16224 3840
rect 16254 4216 16320 4228
rect 16254 3840 16270 4216
rect 16304 3840 16320 4216
rect 16254 3828 16320 3840
rect 16350 4216 16416 4228
rect 16350 3840 16366 4216
rect 16400 3840 16416 4216
rect 16350 3828 16416 3840
rect 16446 4216 16512 4228
rect 16446 3840 16462 4216
rect 16496 3840 16512 4216
rect 16446 3828 16512 3840
rect 16542 4216 16608 4228
rect 16542 3840 16558 4216
rect 16592 3840 16608 4216
rect 16542 3828 16608 3840
rect 16638 4216 16704 4228
rect 16638 3840 16654 4216
rect 16688 3840 16704 4216
rect 16638 3828 16704 3840
rect 16734 4216 16800 4228
rect 16734 3840 16750 4216
rect 16784 3840 16800 4216
rect 16734 3828 16800 3840
rect 16830 4216 16896 4228
rect 16830 3840 16846 4216
rect 16880 3840 16896 4216
rect 16830 3828 16896 3840
rect 16926 4216 16992 4228
rect 16926 3840 16942 4216
rect 16976 3840 16992 4216
rect 16926 3828 16992 3840
rect 17022 4216 17088 4228
rect 17022 3840 17038 4216
rect 17072 3840 17088 4216
rect 17022 3828 17088 3840
rect 17118 4216 17184 4228
rect 17118 3840 17134 4216
rect 17168 3840 17184 4216
rect 17118 3828 17184 3840
rect 17214 4216 17280 4228
rect 17214 3840 17230 4216
rect 17264 3840 17280 4216
rect 17214 3828 17280 3840
rect 17310 4216 17376 4228
rect 17310 3840 17326 4216
rect 17360 3840 17376 4216
rect 17310 3828 17376 3840
rect 17406 4216 17472 4228
rect 17406 3840 17422 4216
rect 17456 3840 17472 4216
rect 17406 3828 17472 3840
rect 17502 4216 17568 4228
rect 17502 3840 17518 4216
rect 17552 3840 17568 4216
rect 17502 3828 17568 3840
rect 17598 4216 17664 4228
rect 17598 3840 17614 4216
rect 17648 3840 17664 4216
rect 17598 3828 17664 3840
rect 17694 4216 17760 4228
rect 17694 3840 17710 4216
rect 17744 3840 17760 4216
rect 17694 3828 17760 3840
rect 17790 4216 17856 4228
rect 17790 3840 17806 4216
rect 17840 3840 17856 4216
rect 17790 3828 17856 3840
rect 17886 4216 17952 4228
rect 17886 3840 17902 4216
rect 17936 3840 17952 4216
rect 17886 3828 17952 3840
rect 17982 4216 18048 4228
rect 17982 3840 17998 4216
rect 18032 3840 18048 4216
rect 17982 3828 18048 3840
rect 18078 4216 18144 4228
rect 18078 3840 18094 4216
rect 18128 3840 18144 4216
rect 18078 3828 18144 3840
rect 18174 4216 18240 4228
rect 18174 3840 18190 4216
rect 18224 3840 18240 4216
rect 18174 3828 18240 3840
rect 18270 4216 18336 4228
rect 18270 3840 18286 4216
rect 18320 3840 18336 4216
rect 18270 3828 18336 3840
rect 18366 4216 18432 4228
rect 18366 3840 18382 4216
rect 18416 3840 18432 4216
rect 18366 3828 18432 3840
rect 18462 4216 18528 4228
rect 18462 3840 18478 4216
rect 18512 3840 18528 4216
rect 18462 3828 18528 3840
rect 18558 4216 18620 4228
rect 18558 3840 18574 4216
rect 18608 3840 18620 4216
rect 18558 3828 18620 3840
rect 15682 3598 15744 3610
rect 15682 3222 15694 3598
rect 15728 3222 15744 3598
rect 15682 3210 15744 3222
rect 15774 3598 15840 3610
rect 15774 3222 15790 3598
rect 15824 3222 15840 3598
rect 15774 3210 15840 3222
rect 15870 3598 15936 3610
rect 15870 3222 15886 3598
rect 15920 3222 15936 3598
rect 15870 3210 15936 3222
rect 15966 3598 16032 3610
rect 15966 3222 15982 3598
rect 16016 3222 16032 3598
rect 15966 3210 16032 3222
rect 16062 3598 16128 3610
rect 16062 3222 16078 3598
rect 16112 3222 16128 3598
rect 16062 3210 16128 3222
rect 16158 3598 16224 3610
rect 16158 3222 16174 3598
rect 16208 3222 16224 3598
rect 16158 3210 16224 3222
rect 16254 3598 16320 3610
rect 16254 3222 16270 3598
rect 16304 3222 16320 3598
rect 16254 3210 16320 3222
rect 16350 3598 16416 3610
rect 16350 3222 16366 3598
rect 16400 3222 16416 3598
rect 16350 3210 16416 3222
rect 16446 3598 16512 3610
rect 16446 3222 16462 3598
rect 16496 3222 16512 3598
rect 16446 3210 16512 3222
rect 16542 3598 16608 3610
rect 16542 3222 16558 3598
rect 16592 3222 16608 3598
rect 16542 3210 16608 3222
rect 16638 3598 16704 3610
rect 16638 3222 16654 3598
rect 16688 3222 16704 3598
rect 16638 3210 16704 3222
rect 16734 3598 16800 3610
rect 16734 3222 16750 3598
rect 16784 3222 16800 3598
rect 16734 3210 16800 3222
rect 16830 3598 16896 3610
rect 16830 3222 16846 3598
rect 16880 3222 16896 3598
rect 16830 3210 16896 3222
rect 16926 3598 16992 3610
rect 16926 3222 16942 3598
rect 16976 3222 16992 3598
rect 16926 3210 16992 3222
rect 17022 3598 17088 3610
rect 17022 3222 17038 3598
rect 17072 3222 17088 3598
rect 17022 3210 17088 3222
rect 17118 3598 17184 3610
rect 17118 3222 17134 3598
rect 17168 3222 17184 3598
rect 17118 3210 17184 3222
rect 17214 3598 17280 3610
rect 17214 3222 17230 3598
rect 17264 3222 17280 3598
rect 17214 3210 17280 3222
rect 17310 3598 17376 3610
rect 17310 3222 17326 3598
rect 17360 3222 17376 3598
rect 17310 3210 17376 3222
rect 17406 3598 17472 3610
rect 17406 3222 17422 3598
rect 17456 3222 17472 3598
rect 17406 3210 17472 3222
rect 17502 3598 17568 3610
rect 17502 3222 17518 3598
rect 17552 3222 17568 3598
rect 17502 3210 17568 3222
rect 17598 3598 17664 3610
rect 17598 3222 17614 3598
rect 17648 3222 17664 3598
rect 17598 3210 17664 3222
rect 17694 3598 17760 3610
rect 17694 3222 17710 3598
rect 17744 3222 17760 3598
rect 17694 3210 17760 3222
rect 17790 3598 17856 3610
rect 17790 3222 17806 3598
rect 17840 3222 17856 3598
rect 17790 3210 17856 3222
rect 17886 3598 17952 3610
rect 17886 3222 17902 3598
rect 17936 3222 17952 3598
rect 17886 3210 17952 3222
rect 17982 3598 18048 3610
rect 17982 3222 17998 3598
rect 18032 3222 18048 3598
rect 17982 3210 18048 3222
rect 18078 3598 18144 3610
rect 18078 3222 18094 3598
rect 18128 3222 18144 3598
rect 18078 3210 18144 3222
rect 18174 3598 18240 3610
rect 18174 3222 18190 3598
rect 18224 3222 18240 3598
rect 18174 3210 18240 3222
rect 18270 3598 18336 3610
rect 18270 3222 18286 3598
rect 18320 3222 18336 3598
rect 18270 3210 18336 3222
rect 18366 3598 18432 3610
rect 18366 3222 18382 3598
rect 18416 3222 18432 3598
rect 18366 3210 18432 3222
rect 18462 3598 18528 3610
rect 18462 3222 18478 3598
rect 18512 3222 18528 3598
rect 18462 3210 18528 3222
rect 18558 3598 18620 3610
rect 18558 3222 18574 3598
rect 18608 3222 18620 3598
rect 18558 3210 18620 3222
rect -1582 2620 -1520 2632
rect -1582 2244 -1570 2620
rect -1536 2244 -1520 2620
rect -1582 2232 -1520 2244
rect -1490 2620 -1424 2632
rect -1490 2244 -1474 2620
rect -1440 2244 -1424 2620
rect -1490 2232 -1424 2244
rect -1394 2620 -1328 2632
rect -1394 2244 -1378 2620
rect -1344 2244 -1328 2620
rect -1394 2232 -1328 2244
rect -1298 2620 -1232 2632
rect -1298 2244 -1282 2620
rect -1248 2244 -1232 2620
rect -1298 2232 -1232 2244
rect -1202 2620 -1136 2632
rect -1202 2244 -1186 2620
rect -1152 2244 -1136 2620
rect -1202 2232 -1136 2244
rect -1106 2620 -1040 2632
rect -1106 2244 -1090 2620
rect -1056 2244 -1040 2620
rect -1106 2232 -1040 2244
rect -1010 2620 -948 2632
rect -1010 2244 -994 2620
rect -960 2244 -948 2620
rect -1010 2232 -948 2244
rect -1582 2002 -1520 2014
rect -1582 1626 -1570 2002
rect -1536 1626 -1520 2002
rect -1582 1614 -1520 1626
rect -1490 2002 -1424 2014
rect -1490 1626 -1474 2002
rect -1440 1626 -1424 2002
rect -1490 1614 -1424 1626
rect -1394 2002 -1328 2014
rect -1394 1626 -1378 2002
rect -1344 1626 -1328 2002
rect -1394 1614 -1328 1626
rect -1298 2002 -1232 2014
rect -1298 1626 -1282 2002
rect -1248 1626 -1232 2002
rect -1298 1614 -1232 1626
rect -1202 2002 -1136 2014
rect -1202 1626 -1186 2002
rect -1152 1626 -1136 2002
rect -1202 1614 -1136 1626
rect -1106 2002 -1040 2014
rect -1106 1626 -1090 2002
rect -1056 1626 -1040 2002
rect -1106 1614 -1040 1626
rect -1010 2002 -948 2014
rect -1010 1626 -994 2002
rect -960 1626 -948 2002
rect -1010 1614 -948 1626
rect -542 2620 -480 2632
rect -542 2244 -530 2620
rect -496 2244 -480 2620
rect -542 2232 -480 2244
rect -450 2620 -384 2632
rect -450 2244 -434 2620
rect -400 2244 -384 2620
rect -450 2232 -384 2244
rect -354 2620 -288 2632
rect -354 2244 -338 2620
rect -304 2244 -288 2620
rect -354 2232 -288 2244
rect -258 2620 -192 2632
rect -258 2244 -242 2620
rect -208 2244 -192 2620
rect -258 2232 -192 2244
rect -162 2620 -96 2632
rect -162 2244 -146 2620
rect -112 2244 -96 2620
rect -162 2232 -96 2244
rect -66 2620 0 2632
rect -66 2244 -50 2620
rect -16 2244 0 2620
rect -66 2232 0 2244
rect 30 2620 92 2632
rect 30 2244 46 2620
rect 80 2244 92 2620
rect 30 2232 92 2244
rect -542 2002 -480 2014
rect -542 1626 -530 2002
rect -496 1626 -480 2002
rect -542 1614 -480 1626
rect -450 2002 -384 2014
rect -450 1626 -434 2002
rect -400 1626 -384 2002
rect -450 1614 -384 1626
rect -354 2002 -288 2014
rect -354 1626 -338 2002
rect -304 1626 -288 2002
rect -354 1614 -288 1626
rect -258 2002 -192 2014
rect -258 1626 -242 2002
rect -208 1626 -192 2002
rect -258 1614 -192 1626
rect -162 2002 -96 2014
rect -162 1626 -146 2002
rect -112 1626 -96 2002
rect -162 1614 -96 1626
rect -66 2002 0 2014
rect -66 1626 -50 2002
rect -16 1626 0 2002
rect -66 1614 0 1626
rect 30 2002 92 2014
rect 30 1626 46 2002
rect 80 1626 92 2002
rect 30 1614 92 1626
rect 498 2620 560 2632
rect 498 2244 510 2620
rect 544 2244 560 2620
rect 498 2232 560 2244
rect 590 2620 656 2632
rect 590 2244 606 2620
rect 640 2244 656 2620
rect 590 2232 656 2244
rect 686 2620 752 2632
rect 686 2244 702 2620
rect 736 2244 752 2620
rect 686 2232 752 2244
rect 782 2620 848 2632
rect 782 2244 798 2620
rect 832 2244 848 2620
rect 782 2232 848 2244
rect 878 2620 944 2632
rect 878 2244 894 2620
rect 928 2244 944 2620
rect 878 2232 944 2244
rect 974 2620 1040 2632
rect 974 2244 990 2620
rect 1024 2244 1040 2620
rect 974 2232 1040 2244
rect 1070 2620 1132 2632
rect 1070 2244 1086 2620
rect 1120 2244 1132 2620
rect 1070 2232 1132 2244
rect 498 2002 560 2014
rect 498 1626 510 2002
rect 544 1626 560 2002
rect 498 1614 560 1626
rect 590 2002 656 2014
rect 590 1626 606 2002
rect 640 1626 656 2002
rect 590 1614 656 1626
rect 686 2002 752 2014
rect 686 1626 702 2002
rect 736 1626 752 2002
rect 686 1614 752 1626
rect 782 2002 848 2014
rect 782 1626 798 2002
rect 832 1626 848 2002
rect 782 1614 848 1626
rect 878 2002 944 2014
rect 878 1626 894 2002
rect 928 1626 944 2002
rect 878 1614 944 1626
rect 974 2002 1040 2014
rect 974 1626 990 2002
rect 1024 1626 1040 2002
rect 974 1614 1040 1626
rect 1070 2002 1132 2014
rect 1070 1626 1086 2002
rect 1120 1626 1132 2002
rect 1070 1614 1132 1626
rect 1538 2620 1600 2632
rect 1538 2244 1550 2620
rect 1584 2244 1600 2620
rect 1538 2232 1600 2244
rect 1630 2620 1696 2632
rect 1630 2244 1646 2620
rect 1680 2244 1696 2620
rect 1630 2232 1696 2244
rect 1726 2620 1792 2632
rect 1726 2244 1742 2620
rect 1776 2244 1792 2620
rect 1726 2232 1792 2244
rect 1822 2620 1888 2632
rect 1822 2244 1838 2620
rect 1872 2244 1888 2620
rect 1822 2232 1888 2244
rect 1918 2620 1984 2632
rect 1918 2244 1934 2620
rect 1968 2244 1984 2620
rect 1918 2232 1984 2244
rect 2014 2620 2080 2632
rect 2014 2244 2030 2620
rect 2064 2244 2080 2620
rect 2014 2232 2080 2244
rect 2110 2620 2172 2632
rect 2110 2244 2126 2620
rect 2160 2244 2172 2620
rect 2110 2232 2172 2244
rect 1538 2002 1600 2014
rect 1538 1626 1550 2002
rect 1584 1626 1600 2002
rect 1538 1614 1600 1626
rect 1630 2002 1696 2014
rect 1630 1626 1646 2002
rect 1680 1626 1696 2002
rect 1630 1614 1696 1626
rect 1726 2002 1792 2014
rect 1726 1626 1742 2002
rect 1776 1626 1792 2002
rect 1726 1614 1792 1626
rect 1822 2002 1888 2014
rect 1822 1626 1838 2002
rect 1872 1626 1888 2002
rect 1822 1614 1888 1626
rect 1918 2002 1984 2014
rect 1918 1626 1934 2002
rect 1968 1626 1984 2002
rect 1918 1614 1984 1626
rect 2014 2002 2080 2014
rect 2014 1626 2030 2002
rect 2064 1626 2080 2002
rect 2014 1614 2080 1626
rect 2110 2002 2172 2014
rect 2110 1626 2126 2002
rect 2160 1626 2172 2002
rect 2110 1614 2172 1626
rect 2578 2620 2640 2632
rect 2578 2244 2590 2620
rect 2624 2244 2640 2620
rect 2578 2232 2640 2244
rect 2670 2620 2736 2632
rect 2670 2244 2686 2620
rect 2720 2244 2736 2620
rect 2670 2232 2736 2244
rect 2766 2620 2832 2632
rect 2766 2244 2782 2620
rect 2816 2244 2832 2620
rect 2766 2232 2832 2244
rect 2862 2620 2928 2632
rect 2862 2244 2878 2620
rect 2912 2244 2928 2620
rect 2862 2232 2928 2244
rect 2958 2620 3024 2632
rect 2958 2244 2974 2620
rect 3008 2244 3024 2620
rect 2958 2232 3024 2244
rect 3054 2620 3120 2632
rect 3054 2244 3070 2620
rect 3104 2244 3120 2620
rect 3054 2232 3120 2244
rect 3150 2620 3212 2632
rect 3150 2244 3166 2620
rect 3200 2244 3212 2620
rect 3150 2232 3212 2244
rect 2578 2002 2640 2014
rect 2578 1626 2590 2002
rect 2624 1626 2640 2002
rect 2578 1614 2640 1626
rect 2670 2002 2736 2014
rect 2670 1626 2686 2002
rect 2720 1626 2736 2002
rect 2670 1614 2736 1626
rect 2766 2002 2832 2014
rect 2766 1626 2782 2002
rect 2816 1626 2832 2002
rect 2766 1614 2832 1626
rect 2862 2002 2928 2014
rect 2862 1626 2878 2002
rect 2912 1626 2928 2002
rect 2862 1614 2928 1626
rect 2958 2002 3024 2014
rect 2958 1626 2974 2002
rect 3008 1626 3024 2002
rect 2958 1614 3024 1626
rect 3054 2002 3120 2014
rect 3054 1626 3070 2002
rect 3104 1626 3120 2002
rect 3054 1614 3120 1626
rect 3150 2002 3212 2014
rect 3150 1626 3166 2002
rect 3200 1626 3212 2002
rect 3150 1614 3212 1626
rect 4222 2780 4284 2792
rect 4222 2404 4234 2780
rect 4268 2404 4284 2780
rect 4222 2392 4284 2404
rect 4314 2780 4380 2792
rect 4314 2404 4330 2780
rect 4364 2404 4380 2780
rect 4314 2392 4380 2404
rect 4410 2780 4476 2792
rect 4410 2404 4426 2780
rect 4460 2404 4476 2780
rect 4410 2392 4476 2404
rect 4506 2780 4572 2792
rect 4506 2404 4522 2780
rect 4556 2404 4572 2780
rect 4506 2392 4572 2404
rect 4602 2780 4668 2792
rect 4602 2404 4618 2780
rect 4652 2404 4668 2780
rect 4602 2392 4668 2404
rect 4698 2780 4764 2792
rect 4698 2404 4714 2780
rect 4748 2404 4764 2780
rect 4698 2392 4764 2404
rect 4794 2780 4856 2792
rect 4794 2404 4810 2780
rect 4844 2404 4856 2780
rect 4794 2392 4856 2404
rect 4222 2162 4284 2174
rect 4222 1786 4234 2162
rect 4268 1786 4284 2162
rect 4222 1774 4284 1786
rect 4314 2162 4380 2174
rect 4314 1786 4330 2162
rect 4364 1786 4380 2162
rect 4314 1774 4380 1786
rect 4410 2162 4476 2174
rect 4410 1786 4426 2162
rect 4460 1786 4476 2162
rect 4410 1774 4476 1786
rect 4506 2162 4572 2174
rect 4506 1786 4522 2162
rect 4556 1786 4572 2162
rect 4506 1774 4572 1786
rect 4602 2162 4668 2174
rect 4602 1786 4618 2162
rect 4652 1786 4668 2162
rect 4602 1774 4668 1786
rect 4698 2162 4764 2174
rect 4698 1786 4714 2162
rect 4748 1786 4764 2162
rect 4698 1774 4764 1786
rect 4794 2162 4856 2174
rect 4794 1786 4810 2162
rect 4844 1786 4856 2162
rect 4794 1774 4856 1786
rect 5262 2780 5324 2792
rect 5262 2404 5274 2780
rect 5308 2404 5324 2780
rect 5262 2392 5324 2404
rect 5354 2780 5420 2792
rect 5354 2404 5370 2780
rect 5404 2404 5420 2780
rect 5354 2392 5420 2404
rect 5450 2780 5516 2792
rect 5450 2404 5466 2780
rect 5500 2404 5516 2780
rect 5450 2392 5516 2404
rect 5546 2780 5612 2792
rect 5546 2404 5562 2780
rect 5596 2404 5612 2780
rect 5546 2392 5612 2404
rect 5642 2780 5708 2792
rect 5642 2404 5658 2780
rect 5692 2404 5708 2780
rect 5642 2392 5708 2404
rect 5738 2780 5804 2792
rect 5738 2404 5754 2780
rect 5788 2404 5804 2780
rect 5738 2392 5804 2404
rect 5834 2780 5896 2792
rect 5834 2404 5850 2780
rect 5884 2404 5896 2780
rect 5834 2392 5896 2404
rect 5262 2162 5324 2174
rect 5262 1786 5274 2162
rect 5308 1786 5324 2162
rect 5262 1774 5324 1786
rect 5354 2162 5420 2174
rect 5354 1786 5370 2162
rect 5404 1786 5420 2162
rect 5354 1774 5420 1786
rect 5450 2162 5516 2174
rect 5450 1786 5466 2162
rect 5500 1786 5516 2162
rect 5450 1774 5516 1786
rect 5546 2162 5612 2174
rect 5546 1786 5562 2162
rect 5596 1786 5612 2162
rect 5546 1774 5612 1786
rect 5642 2162 5708 2174
rect 5642 1786 5658 2162
rect 5692 1786 5708 2162
rect 5642 1774 5708 1786
rect 5738 2162 5804 2174
rect 5738 1786 5754 2162
rect 5788 1786 5804 2162
rect 5738 1774 5804 1786
rect 5834 2162 5896 2174
rect 5834 1786 5850 2162
rect 5884 1786 5896 2162
rect 5834 1774 5896 1786
rect 6302 2780 6364 2792
rect 6302 2404 6314 2780
rect 6348 2404 6364 2780
rect 6302 2392 6364 2404
rect 6394 2780 6460 2792
rect 6394 2404 6410 2780
rect 6444 2404 6460 2780
rect 6394 2392 6460 2404
rect 6490 2780 6556 2792
rect 6490 2404 6506 2780
rect 6540 2404 6556 2780
rect 6490 2392 6556 2404
rect 6586 2780 6652 2792
rect 6586 2404 6602 2780
rect 6636 2404 6652 2780
rect 6586 2392 6652 2404
rect 6682 2780 6748 2792
rect 6682 2404 6698 2780
rect 6732 2404 6748 2780
rect 6682 2392 6748 2404
rect 6778 2780 6844 2792
rect 6778 2404 6794 2780
rect 6828 2404 6844 2780
rect 6778 2392 6844 2404
rect 6874 2780 6936 2792
rect 6874 2404 6890 2780
rect 6924 2404 6936 2780
rect 6874 2392 6936 2404
rect 6302 2162 6364 2174
rect 6302 1786 6314 2162
rect 6348 1786 6364 2162
rect 6302 1774 6364 1786
rect 6394 2162 6460 2174
rect 6394 1786 6410 2162
rect 6444 1786 6460 2162
rect 6394 1774 6460 1786
rect 6490 2162 6556 2174
rect 6490 1786 6506 2162
rect 6540 1786 6556 2162
rect 6490 1774 6556 1786
rect 6586 2162 6652 2174
rect 6586 1786 6602 2162
rect 6636 1786 6652 2162
rect 6586 1774 6652 1786
rect 6682 2162 6748 2174
rect 6682 1786 6698 2162
rect 6732 1786 6748 2162
rect 6682 1774 6748 1786
rect 6778 2162 6844 2174
rect 6778 1786 6794 2162
rect 6828 1786 6844 2162
rect 6778 1774 6844 1786
rect 6874 2162 6936 2174
rect 6874 1786 6890 2162
rect 6924 1786 6936 2162
rect 6874 1774 6936 1786
rect 7342 2780 7404 2792
rect 7342 2404 7354 2780
rect 7388 2404 7404 2780
rect 7342 2392 7404 2404
rect 7434 2780 7500 2792
rect 7434 2404 7450 2780
rect 7484 2404 7500 2780
rect 7434 2392 7500 2404
rect 7530 2780 7596 2792
rect 7530 2404 7546 2780
rect 7580 2404 7596 2780
rect 7530 2392 7596 2404
rect 7626 2780 7692 2792
rect 7626 2404 7642 2780
rect 7676 2404 7692 2780
rect 7626 2392 7692 2404
rect 7722 2780 7788 2792
rect 7722 2404 7738 2780
rect 7772 2404 7788 2780
rect 7722 2392 7788 2404
rect 7818 2780 7884 2792
rect 7818 2404 7834 2780
rect 7868 2404 7884 2780
rect 7818 2392 7884 2404
rect 7914 2780 7976 2792
rect 7914 2404 7930 2780
rect 7964 2404 7976 2780
rect 7914 2392 7976 2404
rect 7342 2162 7404 2174
rect 7342 1786 7354 2162
rect 7388 1786 7404 2162
rect 7342 1774 7404 1786
rect 7434 2162 7500 2174
rect 7434 1786 7450 2162
rect 7484 1786 7500 2162
rect 7434 1774 7500 1786
rect 7530 2162 7596 2174
rect 7530 1786 7546 2162
rect 7580 1786 7596 2162
rect 7530 1774 7596 1786
rect 7626 2162 7692 2174
rect 7626 1786 7642 2162
rect 7676 1786 7692 2162
rect 7626 1774 7692 1786
rect 7722 2162 7788 2174
rect 7722 1786 7738 2162
rect 7772 1786 7788 2162
rect 7722 1774 7788 1786
rect 7818 2162 7884 2174
rect 7818 1786 7834 2162
rect 7868 1786 7884 2162
rect 7818 1774 7884 1786
rect 7914 2162 7976 2174
rect 7914 1786 7930 2162
rect 7964 1786 7976 2162
rect 7914 1774 7976 1786
rect 8382 2780 8444 2792
rect 8382 2404 8394 2780
rect 8428 2404 8444 2780
rect 8382 2392 8444 2404
rect 8474 2780 8540 2792
rect 8474 2404 8490 2780
rect 8524 2404 8540 2780
rect 8474 2392 8540 2404
rect 8570 2780 8636 2792
rect 8570 2404 8586 2780
rect 8620 2404 8636 2780
rect 8570 2392 8636 2404
rect 8666 2780 8732 2792
rect 8666 2404 8682 2780
rect 8716 2404 8732 2780
rect 8666 2392 8732 2404
rect 8762 2780 8828 2792
rect 8762 2404 8778 2780
rect 8812 2404 8828 2780
rect 8762 2392 8828 2404
rect 8858 2780 8924 2792
rect 8858 2404 8874 2780
rect 8908 2404 8924 2780
rect 8858 2392 8924 2404
rect 8954 2780 9016 2792
rect 8954 2404 8970 2780
rect 9004 2404 9016 2780
rect 8954 2392 9016 2404
rect 8382 2162 8444 2174
rect 8382 1786 8394 2162
rect 8428 1786 8444 2162
rect 8382 1774 8444 1786
rect 8474 2162 8540 2174
rect 8474 1786 8490 2162
rect 8524 1786 8540 2162
rect 8474 1774 8540 1786
rect 8570 2162 8636 2174
rect 8570 1786 8586 2162
rect 8620 1786 8636 2162
rect 8570 1774 8636 1786
rect 8666 2162 8732 2174
rect 8666 1786 8682 2162
rect 8716 1786 8732 2162
rect 8666 1774 8732 1786
rect 8762 2162 8828 2174
rect 8762 1786 8778 2162
rect 8812 1786 8828 2162
rect 8762 1774 8828 1786
rect 8858 2162 8924 2174
rect 8858 1786 8874 2162
rect 8908 1786 8924 2162
rect 8858 1774 8924 1786
rect 8954 2162 9016 2174
rect 8954 1786 8970 2162
rect 9004 1786 9016 2162
rect 8954 1774 9016 1786
rect 9422 2780 9484 2792
rect 9422 2404 9434 2780
rect 9468 2404 9484 2780
rect 9422 2392 9484 2404
rect 9514 2780 9580 2792
rect 9514 2404 9530 2780
rect 9564 2404 9580 2780
rect 9514 2392 9580 2404
rect 9610 2780 9676 2792
rect 9610 2404 9626 2780
rect 9660 2404 9676 2780
rect 9610 2392 9676 2404
rect 9706 2780 9772 2792
rect 9706 2404 9722 2780
rect 9756 2404 9772 2780
rect 9706 2392 9772 2404
rect 9802 2780 9868 2792
rect 9802 2404 9818 2780
rect 9852 2404 9868 2780
rect 9802 2392 9868 2404
rect 9898 2780 9964 2792
rect 9898 2404 9914 2780
rect 9948 2404 9964 2780
rect 9898 2392 9964 2404
rect 9994 2780 10056 2792
rect 9994 2404 10010 2780
rect 10044 2404 10056 2780
rect 9994 2392 10056 2404
rect 9422 2162 9484 2174
rect 9422 1786 9434 2162
rect 9468 1786 9484 2162
rect 9422 1774 9484 1786
rect 9514 2162 9580 2174
rect 9514 1786 9530 2162
rect 9564 1786 9580 2162
rect 9514 1774 9580 1786
rect 9610 2162 9676 2174
rect 9610 1786 9626 2162
rect 9660 1786 9676 2162
rect 9610 1774 9676 1786
rect 9706 2162 9772 2174
rect 9706 1786 9722 2162
rect 9756 1786 9772 2162
rect 9706 1774 9772 1786
rect 9802 2162 9868 2174
rect 9802 1786 9818 2162
rect 9852 1786 9868 2162
rect 9802 1774 9868 1786
rect 9898 2162 9964 2174
rect 9898 1786 9914 2162
rect 9948 1786 9964 2162
rect 9898 1774 9964 1786
rect 9994 2162 10056 2174
rect 9994 1786 10010 2162
rect 10044 1786 10056 2162
rect 9994 1774 10056 1786
rect 10462 2780 10524 2792
rect 10462 2404 10474 2780
rect 10508 2404 10524 2780
rect 10462 2392 10524 2404
rect 10554 2780 10620 2792
rect 10554 2404 10570 2780
rect 10604 2404 10620 2780
rect 10554 2392 10620 2404
rect 10650 2780 10716 2792
rect 10650 2404 10666 2780
rect 10700 2404 10716 2780
rect 10650 2392 10716 2404
rect 10746 2780 10812 2792
rect 10746 2404 10762 2780
rect 10796 2404 10812 2780
rect 10746 2392 10812 2404
rect 10842 2780 10908 2792
rect 10842 2404 10858 2780
rect 10892 2404 10908 2780
rect 10842 2392 10908 2404
rect 10938 2780 11004 2792
rect 10938 2404 10954 2780
rect 10988 2404 11004 2780
rect 10938 2392 11004 2404
rect 11034 2780 11096 2792
rect 11034 2404 11050 2780
rect 11084 2404 11096 2780
rect 11034 2392 11096 2404
rect 10462 2162 10524 2174
rect 10462 1786 10474 2162
rect 10508 1786 10524 2162
rect 10462 1774 10524 1786
rect 10554 2162 10620 2174
rect 10554 1786 10570 2162
rect 10604 1786 10620 2162
rect 10554 1774 10620 1786
rect 10650 2162 10716 2174
rect 10650 1786 10666 2162
rect 10700 1786 10716 2162
rect 10650 1774 10716 1786
rect 10746 2162 10812 2174
rect 10746 1786 10762 2162
rect 10796 1786 10812 2162
rect 10746 1774 10812 1786
rect 10842 2162 10908 2174
rect 10842 1786 10858 2162
rect 10892 1786 10908 2162
rect 10842 1774 10908 1786
rect 10938 2162 11004 2174
rect 10938 1786 10954 2162
rect 10988 1786 11004 2162
rect 10938 1774 11004 1786
rect 11034 2162 11096 2174
rect 11034 1786 11050 2162
rect 11084 1786 11096 2162
rect 11034 1774 11096 1786
rect 11842 2780 11904 2792
rect 11842 2404 11854 2780
rect 11888 2404 11904 2780
rect 11842 2392 11904 2404
rect 11934 2780 12000 2792
rect 11934 2404 11950 2780
rect 11984 2404 12000 2780
rect 11934 2392 12000 2404
rect 12030 2780 12096 2792
rect 12030 2404 12046 2780
rect 12080 2404 12096 2780
rect 12030 2392 12096 2404
rect 12126 2780 12192 2792
rect 12126 2404 12142 2780
rect 12176 2404 12192 2780
rect 12126 2392 12192 2404
rect 12222 2780 12288 2792
rect 12222 2404 12238 2780
rect 12272 2404 12288 2780
rect 12222 2392 12288 2404
rect 12318 2780 12384 2792
rect 12318 2404 12334 2780
rect 12368 2404 12384 2780
rect 12318 2392 12384 2404
rect 12414 2780 12476 2792
rect 12414 2404 12430 2780
rect 12464 2404 12476 2780
rect 12414 2392 12476 2404
rect 11842 2162 11904 2174
rect 11842 1786 11854 2162
rect 11888 1786 11904 2162
rect 11842 1774 11904 1786
rect 11934 2162 12000 2174
rect 11934 1786 11950 2162
rect 11984 1786 12000 2162
rect 11934 1774 12000 1786
rect 12030 2162 12096 2174
rect 12030 1786 12046 2162
rect 12080 1786 12096 2162
rect 12030 1774 12096 1786
rect 12126 2162 12192 2174
rect 12126 1786 12142 2162
rect 12176 1786 12192 2162
rect 12126 1774 12192 1786
rect 12222 2162 12288 2174
rect 12222 1786 12238 2162
rect 12272 1786 12288 2162
rect 12222 1774 12288 1786
rect 12318 2162 12384 2174
rect 12318 1786 12334 2162
rect 12368 1786 12384 2162
rect 12318 1774 12384 1786
rect 12414 2162 12476 2174
rect 12414 1786 12430 2162
rect 12464 1786 12476 2162
rect 12414 1774 12476 1786
rect 12882 2780 12944 2792
rect 12882 2404 12894 2780
rect 12928 2404 12944 2780
rect 12882 2392 12944 2404
rect 12974 2780 13040 2792
rect 12974 2404 12990 2780
rect 13024 2404 13040 2780
rect 12974 2392 13040 2404
rect 13070 2780 13136 2792
rect 13070 2404 13086 2780
rect 13120 2404 13136 2780
rect 13070 2392 13136 2404
rect 13166 2780 13232 2792
rect 13166 2404 13182 2780
rect 13216 2404 13232 2780
rect 13166 2392 13232 2404
rect 13262 2780 13328 2792
rect 13262 2404 13278 2780
rect 13312 2404 13328 2780
rect 13262 2392 13328 2404
rect 13358 2780 13424 2792
rect 13358 2404 13374 2780
rect 13408 2404 13424 2780
rect 13358 2392 13424 2404
rect 13454 2780 13516 2792
rect 13454 2404 13470 2780
rect 13504 2404 13516 2780
rect 13454 2392 13516 2404
rect 12882 2162 12944 2174
rect 12882 1786 12894 2162
rect 12928 1786 12944 2162
rect 12882 1774 12944 1786
rect 12974 2162 13040 2174
rect 12974 1786 12990 2162
rect 13024 1786 13040 2162
rect 12974 1774 13040 1786
rect 13070 2162 13136 2174
rect 13070 1786 13086 2162
rect 13120 1786 13136 2162
rect 13070 1774 13136 1786
rect 13166 2162 13232 2174
rect 13166 1786 13182 2162
rect 13216 1786 13232 2162
rect 13166 1774 13232 1786
rect 13262 2162 13328 2174
rect 13262 1786 13278 2162
rect 13312 1786 13328 2162
rect 13262 1774 13328 1786
rect 13358 2162 13424 2174
rect 13358 1786 13374 2162
rect 13408 1786 13424 2162
rect 13358 1774 13424 1786
rect 13454 2162 13516 2174
rect 13454 1786 13470 2162
rect 13504 1786 13516 2162
rect 13454 1774 13516 1786
rect 13922 2780 13984 2792
rect 13922 2404 13934 2780
rect 13968 2404 13984 2780
rect 13922 2392 13984 2404
rect 14014 2780 14080 2792
rect 14014 2404 14030 2780
rect 14064 2404 14080 2780
rect 14014 2392 14080 2404
rect 14110 2780 14176 2792
rect 14110 2404 14126 2780
rect 14160 2404 14176 2780
rect 14110 2392 14176 2404
rect 14206 2780 14272 2792
rect 14206 2404 14222 2780
rect 14256 2404 14272 2780
rect 14206 2392 14272 2404
rect 14302 2780 14368 2792
rect 14302 2404 14318 2780
rect 14352 2404 14368 2780
rect 14302 2392 14368 2404
rect 14398 2780 14464 2792
rect 14398 2404 14414 2780
rect 14448 2404 14464 2780
rect 14398 2392 14464 2404
rect 14494 2780 14556 2792
rect 14494 2404 14510 2780
rect 14544 2404 14556 2780
rect 14494 2392 14556 2404
rect 13922 2162 13984 2174
rect 13922 1786 13934 2162
rect 13968 1786 13984 2162
rect 13922 1774 13984 1786
rect 14014 2162 14080 2174
rect 14014 1786 14030 2162
rect 14064 1786 14080 2162
rect 14014 1774 14080 1786
rect 14110 2162 14176 2174
rect 14110 1786 14126 2162
rect 14160 1786 14176 2162
rect 14110 1774 14176 1786
rect 14206 2162 14272 2174
rect 14206 1786 14222 2162
rect 14256 1786 14272 2162
rect 14206 1774 14272 1786
rect 14302 2162 14368 2174
rect 14302 1786 14318 2162
rect 14352 1786 14368 2162
rect 14302 1774 14368 1786
rect 14398 2162 14464 2174
rect 14398 1786 14414 2162
rect 14448 1786 14464 2162
rect 14398 1774 14464 1786
rect 14494 2162 14556 2174
rect 14494 1786 14510 2162
rect 14544 1786 14556 2162
rect 14494 1774 14556 1786
rect 14962 2780 15024 2792
rect 14962 2404 14974 2780
rect 15008 2404 15024 2780
rect 14962 2392 15024 2404
rect 15054 2780 15120 2792
rect 15054 2404 15070 2780
rect 15104 2404 15120 2780
rect 15054 2392 15120 2404
rect 15150 2780 15216 2792
rect 15150 2404 15166 2780
rect 15200 2404 15216 2780
rect 15150 2392 15216 2404
rect 15246 2780 15312 2792
rect 15246 2404 15262 2780
rect 15296 2404 15312 2780
rect 15246 2392 15312 2404
rect 15342 2780 15408 2792
rect 15342 2404 15358 2780
rect 15392 2404 15408 2780
rect 15342 2392 15408 2404
rect 15438 2780 15504 2792
rect 15438 2404 15454 2780
rect 15488 2404 15504 2780
rect 15438 2392 15504 2404
rect 15534 2780 15596 2792
rect 15534 2404 15550 2780
rect 15584 2404 15596 2780
rect 15534 2392 15596 2404
rect 14962 2162 15024 2174
rect 14962 1786 14974 2162
rect 15008 1786 15024 2162
rect 14962 1774 15024 1786
rect 15054 2162 15120 2174
rect 15054 1786 15070 2162
rect 15104 1786 15120 2162
rect 15054 1774 15120 1786
rect 15150 2162 15216 2174
rect 15150 1786 15166 2162
rect 15200 1786 15216 2162
rect 15150 1774 15216 1786
rect 15246 2162 15312 2174
rect 15246 1786 15262 2162
rect 15296 1786 15312 2162
rect 15246 1774 15312 1786
rect 15342 2162 15408 2174
rect 15342 1786 15358 2162
rect 15392 1786 15408 2162
rect 15342 1774 15408 1786
rect 15438 2162 15504 2174
rect 15438 1786 15454 2162
rect 15488 1786 15504 2162
rect 15438 1774 15504 1786
rect 15534 2162 15596 2174
rect 15534 1786 15550 2162
rect 15584 1786 15596 2162
rect 15534 1774 15596 1786
rect 16002 2780 16064 2792
rect 16002 2404 16014 2780
rect 16048 2404 16064 2780
rect 16002 2392 16064 2404
rect 16094 2780 16160 2792
rect 16094 2404 16110 2780
rect 16144 2404 16160 2780
rect 16094 2392 16160 2404
rect 16190 2780 16256 2792
rect 16190 2404 16206 2780
rect 16240 2404 16256 2780
rect 16190 2392 16256 2404
rect 16286 2780 16352 2792
rect 16286 2404 16302 2780
rect 16336 2404 16352 2780
rect 16286 2392 16352 2404
rect 16382 2780 16448 2792
rect 16382 2404 16398 2780
rect 16432 2404 16448 2780
rect 16382 2392 16448 2404
rect 16478 2780 16544 2792
rect 16478 2404 16494 2780
rect 16528 2404 16544 2780
rect 16478 2392 16544 2404
rect 16574 2780 16636 2792
rect 16574 2404 16590 2780
rect 16624 2404 16636 2780
rect 16574 2392 16636 2404
rect 16002 2162 16064 2174
rect 16002 1786 16014 2162
rect 16048 1786 16064 2162
rect 16002 1774 16064 1786
rect 16094 2162 16160 2174
rect 16094 1786 16110 2162
rect 16144 1786 16160 2162
rect 16094 1774 16160 1786
rect 16190 2162 16256 2174
rect 16190 1786 16206 2162
rect 16240 1786 16256 2162
rect 16190 1774 16256 1786
rect 16286 2162 16352 2174
rect 16286 1786 16302 2162
rect 16336 1786 16352 2162
rect 16286 1774 16352 1786
rect 16382 2162 16448 2174
rect 16382 1786 16398 2162
rect 16432 1786 16448 2162
rect 16382 1774 16448 1786
rect 16478 2162 16544 2174
rect 16478 1786 16494 2162
rect 16528 1786 16544 2162
rect 16478 1774 16544 1786
rect 16574 2162 16636 2174
rect 16574 1786 16590 2162
rect 16624 1786 16636 2162
rect 16574 1774 16636 1786
rect 17042 2780 17104 2792
rect 17042 2404 17054 2780
rect 17088 2404 17104 2780
rect 17042 2392 17104 2404
rect 17134 2780 17200 2792
rect 17134 2404 17150 2780
rect 17184 2404 17200 2780
rect 17134 2392 17200 2404
rect 17230 2780 17296 2792
rect 17230 2404 17246 2780
rect 17280 2404 17296 2780
rect 17230 2392 17296 2404
rect 17326 2780 17392 2792
rect 17326 2404 17342 2780
rect 17376 2404 17392 2780
rect 17326 2392 17392 2404
rect 17422 2780 17488 2792
rect 17422 2404 17438 2780
rect 17472 2404 17488 2780
rect 17422 2392 17488 2404
rect 17518 2780 17584 2792
rect 17518 2404 17534 2780
rect 17568 2404 17584 2780
rect 17518 2392 17584 2404
rect 17614 2780 17676 2792
rect 17614 2404 17630 2780
rect 17664 2404 17676 2780
rect 17614 2392 17676 2404
rect 17042 2162 17104 2174
rect 17042 1786 17054 2162
rect 17088 1786 17104 2162
rect 17042 1774 17104 1786
rect 17134 2162 17200 2174
rect 17134 1786 17150 2162
rect 17184 1786 17200 2162
rect 17134 1774 17200 1786
rect 17230 2162 17296 2174
rect 17230 1786 17246 2162
rect 17280 1786 17296 2162
rect 17230 1774 17296 1786
rect 17326 2162 17392 2174
rect 17326 1786 17342 2162
rect 17376 1786 17392 2162
rect 17326 1774 17392 1786
rect 17422 2162 17488 2174
rect 17422 1786 17438 2162
rect 17472 1786 17488 2162
rect 17422 1774 17488 1786
rect 17518 2162 17584 2174
rect 17518 1786 17534 2162
rect 17568 1786 17584 2162
rect 17518 1774 17584 1786
rect 17614 2162 17676 2174
rect 17614 1786 17630 2162
rect 17664 1786 17676 2162
rect 17614 1774 17676 1786
rect 18082 2780 18144 2792
rect 18082 2404 18094 2780
rect 18128 2404 18144 2780
rect 18082 2392 18144 2404
rect 18174 2780 18240 2792
rect 18174 2404 18190 2780
rect 18224 2404 18240 2780
rect 18174 2392 18240 2404
rect 18270 2780 18336 2792
rect 18270 2404 18286 2780
rect 18320 2404 18336 2780
rect 18270 2392 18336 2404
rect 18366 2780 18432 2792
rect 18366 2404 18382 2780
rect 18416 2404 18432 2780
rect 18366 2392 18432 2404
rect 18462 2780 18528 2792
rect 18462 2404 18478 2780
rect 18512 2404 18528 2780
rect 18462 2392 18528 2404
rect 18558 2780 18624 2792
rect 18558 2404 18574 2780
rect 18608 2404 18624 2780
rect 18558 2392 18624 2404
rect 18654 2780 18716 2792
rect 18654 2404 18670 2780
rect 18704 2404 18716 2780
rect 18654 2392 18716 2404
rect 18082 2162 18144 2174
rect 18082 1786 18094 2162
rect 18128 1786 18144 2162
rect 18082 1774 18144 1786
rect 18174 2162 18240 2174
rect 18174 1786 18190 2162
rect 18224 1786 18240 2162
rect 18174 1774 18240 1786
rect 18270 2162 18336 2174
rect 18270 1786 18286 2162
rect 18320 1786 18336 2162
rect 18270 1774 18336 1786
rect 18366 2162 18432 2174
rect 18366 1786 18382 2162
rect 18416 1786 18432 2162
rect 18366 1774 18432 1786
rect 18462 2162 18528 2174
rect 18462 1786 18478 2162
rect 18512 1786 18528 2162
rect 18462 1774 18528 1786
rect 18558 2162 18624 2174
rect 18558 1786 18574 2162
rect 18608 1786 18624 2162
rect 18558 1774 18624 1786
rect 18654 2162 18716 2174
rect 18654 1786 18670 2162
rect 18704 1786 18716 2162
rect 18654 1774 18716 1786
rect -1582 1198 -1524 1210
rect -1582 822 -1570 1198
rect -1536 822 -1524 1198
rect -1582 810 -1524 822
rect -1464 1198 -1406 1210
rect -1464 822 -1452 1198
rect -1418 822 -1406 1198
rect -1464 810 -1406 822
rect -1346 1198 -1288 1210
rect -1346 822 -1334 1198
rect -1300 822 -1288 1198
rect -1346 810 -1288 822
rect -1228 1198 -1170 1210
rect -1228 822 -1216 1198
rect -1182 822 -1170 1198
rect -1228 810 -1170 822
rect -1110 1198 -1052 1210
rect -1110 822 -1098 1198
rect -1064 822 -1052 1198
rect -1110 810 -1052 822
rect -992 1198 -934 1210
rect -992 822 -980 1198
rect -946 822 -934 1198
rect -992 810 -934 822
rect -874 1198 -816 1210
rect -874 822 -862 1198
rect -828 822 -816 1198
rect -874 810 -816 822
rect -542 1198 -484 1210
rect -542 822 -530 1198
rect -496 822 -484 1198
rect -542 810 -484 822
rect -424 1198 -366 1210
rect -424 822 -412 1198
rect -378 822 -366 1198
rect -424 810 -366 822
rect -306 1198 -248 1210
rect -306 822 -294 1198
rect -260 822 -248 1198
rect -306 810 -248 822
rect -188 1198 -130 1210
rect -188 822 -176 1198
rect -142 822 -130 1198
rect -188 810 -130 822
rect -70 1198 -12 1210
rect -70 822 -58 1198
rect -24 822 -12 1198
rect -70 810 -12 822
rect 48 1198 106 1210
rect 48 822 60 1198
rect 94 822 106 1198
rect 48 810 106 822
rect 166 1198 224 1210
rect 166 822 178 1198
rect 212 822 224 1198
rect 166 810 224 822
rect 498 1198 556 1210
rect 498 822 510 1198
rect 544 822 556 1198
rect 498 810 556 822
rect 616 1198 674 1210
rect 616 822 628 1198
rect 662 822 674 1198
rect 616 810 674 822
rect 734 1198 792 1210
rect 734 822 746 1198
rect 780 822 792 1198
rect 734 810 792 822
rect 852 1198 910 1210
rect 852 822 864 1198
rect 898 822 910 1198
rect 852 810 910 822
rect 970 1198 1028 1210
rect 970 822 982 1198
rect 1016 822 1028 1198
rect 970 810 1028 822
rect 1088 1198 1146 1210
rect 1088 822 1100 1198
rect 1134 822 1146 1198
rect 1088 810 1146 822
rect 1206 1198 1264 1210
rect 1206 822 1218 1198
rect 1252 822 1264 1198
rect 1206 810 1264 822
rect 1538 1198 1596 1210
rect 1538 822 1550 1198
rect 1584 822 1596 1198
rect 1538 810 1596 822
rect 1656 1198 1714 1210
rect 1656 822 1668 1198
rect 1702 822 1714 1198
rect 1656 810 1714 822
rect 1774 1198 1832 1210
rect 1774 822 1786 1198
rect 1820 822 1832 1198
rect 1774 810 1832 822
rect 1892 1198 1950 1210
rect 1892 822 1904 1198
rect 1938 822 1950 1198
rect 1892 810 1950 822
rect 2010 1198 2068 1210
rect 2010 822 2022 1198
rect 2056 822 2068 1198
rect 2010 810 2068 822
rect 2128 1198 2186 1210
rect 2128 822 2140 1198
rect 2174 822 2186 1198
rect 2128 810 2186 822
rect 2246 1198 2304 1210
rect 2246 822 2258 1198
rect 2292 822 2304 1198
rect 2246 810 2304 822
rect 2578 1198 2636 1210
rect 2578 822 2590 1198
rect 2624 822 2636 1198
rect 2578 810 2636 822
rect 2696 1198 2754 1210
rect 2696 822 2708 1198
rect 2742 822 2754 1198
rect 2696 810 2754 822
rect 2814 1198 2872 1210
rect 2814 822 2826 1198
rect 2860 822 2872 1198
rect 2814 810 2872 822
rect 2932 1198 2990 1210
rect 2932 822 2944 1198
rect 2978 822 2990 1198
rect 2932 810 2990 822
rect 3050 1198 3108 1210
rect 3050 822 3062 1198
rect 3096 822 3108 1198
rect 3050 810 3108 822
rect 3168 1198 3226 1210
rect 3168 822 3180 1198
rect 3214 822 3226 1198
rect 3168 810 3226 822
rect 3286 1198 3344 1210
rect 3286 822 3298 1198
rect 3332 822 3344 1198
rect 3286 810 3344 822
rect 4222 1358 4280 1370
rect 4222 982 4234 1358
rect 4268 982 4280 1358
rect 4222 970 4280 982
rect 4340 1358 4398 1370
rect 4340 982 4352 1358
rect 4386 982 4398 1358
rect 4340 970 4398 982
rect 4458 1358 4516 1370
rect 4458 982 4470 1358
rect 4504 982 4516 1358
rect 4458 970 4516 982
rect 4576 1358 4634 1370
rect 4576 982 4588 1358
rect 4622 982 4634 1358
rect 4576 970 4634 982
rect 4694 1358 4752 1370
rect 4694 982 4706 1358
rect 4740 982 4752 1358
rect 4694 970 4752 982
rect 4812 1358 4870 1370
rect 4812 982 4824 1358
rect 4858 982 4870 1358
rect 4812 970 4870 982
rect 4930 1358 4988 1370
rect 4930 982 4942 1358
rect 4976 982 4988 1358
rect 4930 970 4988 982
rect 5262 1358 5320 1370
rect 5262 982 5274 1358
rect 5308 982 5320 1358
rect 5262 970 5320 982
rect 5380 1358 5438 1370
rect 5380 982 5392 1358
rect 5426 982 5438 1358
rect 5380 970 5438 982
rect 5498 1358 5556 1370
rect 5498 982 5510 1358
rect 5544 982 5556 1358
rect 5498 970 5556 982
rect 5616 1358 5674 1370
rect 5616 982 5628 1358
rect 5662 982 5674 1358
rect 5616 970 5674 982
rect 5734 1358 5792 1370
rect 5734 982 5746 1358
rect 5780 982 5792 1358
rect 5734 970 5792 982
rect 5852 1358 5910 1370
rect 5852 982 5864 1358
rect 5898 982 5910 1358
rect 5852 970 5910 982
rect 5970 1358 6028 1370
rect 5970 982 5982 1358
rect 6016 982 6028 1358
rect 5970 970 6028 982
rect 6302 1358 6360 1370
rect 6302 982 6314 1358
rect 6348 982 6360 1358
rect 6302 970 6360 982
rect 6420 1358 6478 1370
rect 6420 982 6432 1358
rect 6466 982 6478 1358
rect 6420 970 6478 982
rect 6538 1358 6596 1370
rect 6538 982 6550 1358
rect 6584 982 6596 1358
rect 6538 970 6596 982
rect 6656 1358 6714 1370
rect 6656 982 6668 1358
rect 6702 982 6714 1358
rect 6656 970 6714 982
rect 6774 1358 6832 1370
rect 6774 982 6786 1358
rect 6820 982 6832 1358
rect 6774 970 6832 982
rect 6892 1358 6950 1370
rect 6892 982 6904 1358
rect 6938 982 6950 1358
rect 6892 970 6950 982
rect 7010 1358 7068 1370
rect 7010 982 7022 1358
rect 7056 982 7068 1358
rect 7010 970 7068 982
rect 7342 1358 7400 1370
rect 7342 982 7354 1358
rect 7388 982 7400 1358
rect 7342 970 7400 982
rect 7460 1358 7518 1370
rect 7460 982 7472 1358
rect 7506 982 7518 1358
rect 7460 970 7518 982
rect 7578 1358 7636 1370
rect 7578 982 7590 1358
rect 7624 982 7636 1358
rect 7578 970 7636 982
rect 7696 1358 7754 1370
rect 7696 982 7708 1358
rect 7742 982 7754 1358
rect 7696 970 7754 982
rect 7814 1358 7872 1370
rect 7814 982 7826 1358
rect 7860 982 7872 1358
rect 7814 970 7872 982
rect 7932 1358 7990 1370
rect 7932 982 7944 1358
rect 7978 982 7990 1358
rect 7932 970 7990 982
rect 8050 1358 8108 1370
rect 8050 982 8062 1358
rect 8096 982 8108 1358
rect 8050 970 8108 982
rect 8382 1358 8440 1370
rect 8382 982 8394 1358
rect 8428 982 8440 1358
rect 8382 970 8440 982
rect 8500 1358 8558 1370
rect 8500 982 8512 1358
rect 8546 982 8558 1358
rect 8500 970 8558 982
rect 8618 1358 8676 1370
rect 8618 982 8630 1358
rect 8664 982 8676 1358
rect 8618 970 8676 982
rect 8736 1358 8794 1370
rect 8736 982 8748 1358
rect 8782 982 8794 1358
rect 8736 970 8794 982
rect 8854 1358 8912 1370
rect 8854 982 8866 1358
rect 8900 982 8912 1358
rect 8854 970 8912 982
rect 8972 1358 9030 1370
rect 8972 982 8984 1358
rect 9018 982 9030 1358
rect 8972 970 9030 982
rect 9090 1358 9148 1370
rect 9090 982 9102 1358
rect 9136 982 9148 1358
rect 9090 970 9148 982
rect 9422 1358 9480 1370
rect 9422 982 9434 1358
rect 9468 982 9480 1358
rect 9422 970 9480 982
rect 9540 1358 9598 1370
rect 9540 982 9552 1358
rect 9586 982 9598 1358
rect 9540 970 9598 982
rect 9658 1358 9716 1370
rect 9658 982 9670 1358
rect 9704 982 9716 1358
rect 9658 970 9716 982
rect 9776 1358 9834 1370
rect 9776 982 9788 1358
rect 9822 982 9834 1358
rect 9776 970 9834 982
rect 9894 1358 9952 1370
rect 9894 982 9906 1358
rect 9940 982 9952 1358
rect 9894 970 9952 982
rect 10012 1358 10070 1370
rect 10012 982 10024 1358
rect 10058 982 10070 1358
rect 10012 970 10070 982
rect 10130 1358 10188 1370
rect 10130 982 10142 1358
rect 10176 982 10188 1358
rect 10130 970 10188 982
rect 10462 1358 10520 1370
rect 10462 982 10474 1358
rect 10508 982 10520 1358
rect 10462 970 10520 982
rect 10580 1358 10638 1370
rect 10580 982 10592 1358
rect 10626 982 10638 1358
rect 10580 970 10638 982
rect 10698 1358 10756 1370
rect 10698 982 10710 1358
rect 10744 982 10756 1358
rect 10698 970 10756 982
rect 10816 1358 10874 1370
rect 10816 982 10828 1358
rect 10862 982 10874 1358
rect 10816 970 10874 982
rect 10934 1358 10992 1370
rect 10934 982 10946 1358
rect 10980 982 10992 1358
rect 10934 970 10992 982
rect 11052 1358 11110 1370
rect 11052 982 11064 1358
rect 11098 982 11110 1358
rect 11052 970 11110 982
rect 11170 1358 11228 1370
rect 11170 982 11182 1358
rect 11216 982 11228 1358
rect 11170 970 11228 982
rect 11842 1358 11900 1370
rect 11842 982 11854 1358
rect 11888 982 11900 1358
rect 11842 970 11900 982
rect 11960 1358 12018 1370
rect 11960 982 11972 1358
rect 12006 982 12018 1358
rect 11960 970 12018 982
rect 12078 1358 12136 1370
rect 12078 982 12090 1358
rect 12124 982 12136 1358
rect 12078 970 12136 982
rect 12196 1358 12254 1370
rect 12196 982 12208 1358
rect 12242 982 12254 1358
rect 12196 970 12254 982
rect 12314 1358 12372 1370
rect 12314 982 12326 1358
rect 12360 982 12372 1358
rect 12314 970 12372 982
rect 12432 1358 12490 1370
rect 12432 982 12444 1358
rect 12478 982 12490 1358
rect 12432 970 12490 982
rect 12550 1358 12608 1370
rect 12550 982 12562 1358
rect 12596 982 12608 1358
rect 12550 970 12608 982
rect 12882 1358 12940 1370
rect 12882 982 12894 1358
rect 12928 982 12940 1358
rect 12882 970 12940 982
rect 13000 1358 13058 1370
rect 13000 982 13012 1358
rect 13046 982 13058 1358
rect 13000 970 13058 982
rect 13118 1358 13176 1370
rect 13118 982 13130 1358
rect 13164 982 13176 1358
rect 13118 970 13176 982
rect 13236 1358 13294 1370
rect 13236 982 13248 1358
rect 13282 982 13294 1358
rect 13236 970 13294 982
rect 13354 1358 13412 1370
rect 13354 982 13366 1358
rect 13400 982 13412 1358
rect 13354 970 13412 982
rect 13472 1358 13530 1370
rect 13472 982 13484 1358
rect 13518 982 13530 1358
rect 13472 970 13530 982
rect 13590 1358 13648 1370
rect 13590 982 13602 1358
rect 13636 982 13648 1358
rect 13590 970 13648 982
rect 13922 1358 13980 1370
rect 13922 982 13934 1358
rect 13968 982 13980 1358
rect 13922 970 13980 982
rect 14040 1358 14098 1370
rect 14040 982 14052 1358
rect 14086 982 14098 1358
rect 14040 970 14098 982
rect 14158 1358 14216 1370
rect 14158 982 14170 1358
rect 14204 982 14216 1358
rect 14158 970 14216 982
rect 14276 1358 14334 1370
rect 14276 982 14288 1358
rect 14322 982 14334 1358
rect 14276 970 14334 982
rect 14394 1358 14452 1370
rect 14394 982 14406 1358
rect 14440 982 14452 1358
rect 14394 970 14452 982
rect 14512 1358 14570 1370
rect 14512 982 14524 1358
rect 14558 982 14570 1358
rect 14512 970 14570 982
rect 14630 1358 14688 1370
rect 14630 982 14642 1358
rect 14676 982 14688 1358
rect 14630 970 14688 982
rect 14962 1358 15020 1370
rect 14962 982 14974 1358
rect 15008 982 15020 1358
rect 14962 970 15020 982
rect 15080 1358 15138 1370
rect 15080 982 15092 1358
rect 15126 982 15138 1358
rect 15080 970 15138 982
rect 15198 1358 15256 1370
rect 15198 982 15210 1358
rect 15244 982 15256 1358
rect 15198 970 15256 982
rect 15316 1358 15374 1370
rect 15316 982 15328 1358
rect 15362 982 15374 1358
rect 15316 970 15374 982
rect 15434 1358 15492 1370
rect 15434 982 15446 1358
rect 15480 982 15492 1358
rect 15434 970 15492 982
rect 15552 1358 15610 1370
rect 15552 982 15564 1358
rect 15598 982 15610 1358
rect 15552 970 15610 982
rect 15670 1358 15728 1370
rect 15670 982 15682 1358
rect 15716 982 15728 1358
rect 15670 970 15728 982
rect 16002 1358 16060 1370
rect 16002 982 16014 1358
rect 16048 982 16060 1358
rect 16002 970 16060 982
rect 16120 1358 16178 1370
rect 16120 982 16132 1358
rect 16166 982 16178 1358
rect 16120 970 16178 982
rect 16238 1358 16296 1370
rect 16238 982 16250 1358
rect 16284 982 16296 1358
rect 16238 970 16296 982
rect 16356 1358 16414 1370
rect 16356 982 16368 1358
rect 16402 982 16414 1358
rect 16356 970 16414 982
rect 16474 1358 16532 1370
rect 16474 982 16486 1358
rect 16520 982 16532 1358
rect 16474 970 16532 982
rect 16592 1358 16650 1370
rect 16592 982 16604 1358
rect 16638 982 16650 1358
rect 16592 970 16650 982
rect 16710 1358 16768 1370
rect 16710 982 16722 1358
rect 16756 982 16768 1358
rect 16710 970 16768 982
rect 17042 1358 17100 1370
rect 17042 982 17054 1358
rect 17088 982 17100 1358
rect 17042 970 17100 982
rect 17160 1358 17218 1370
rect 17160 982 17172 1358
rect 17206 982 17218 1358
rect 17160 970 17218 982
rect 17278 1358 17336 1370
rect 17278 982 17290 1358
rect 17324 982 17336 1358
rect 17278 970 17336 982
rect 17396 1358 17454 1370
rect 17396 982 17408 1358
rect 17442 982 17454 1358
rect 17396 970 17454 982
rect 17514 1358 17572 1370
rect 17514 982 17526 1358
rect 17560 982 17572 1358
rect 17514 970 17572 982
rect 17632 1358 17690 1370
rect 17632 982 17644 1358
rect 17678 982 17690 1358
rect 17632 970 17690 982
rect 17750 1358 17808 1370
rect 17750 982 17762 1358
rect 17796 982 17808 1358
rect 17750 970 17808 982
rect 18082 1358 18140 1370
rect 18082 982 18094 1358
rect 18128 982 18140 1358
rect 18082 970 18140 982
rect 18200 1358 18258 1370
rect 18200 982 18212 1358
rect 18246 982 18258 1358
rect 18200 970 18258 982
rect 18318 1358 18376 1370
rect 18318 982 18330 1358
rect 18364 982 18376 1358
rect 18318 970 18376 982
rect 18436 1358 18494 1370
rect 18436 982 18448 1358
rect 18482 982 18494 1358
rect 18436 970 18494 982
rect 18554 1358 18612 1370
rect 18554 982 18566 1358
rect 18600 982 18612 1358
rect 18554 970 18612 982
rect 18672 1358 18730 1370
rect 18672 982 18684 1358
rect 18718 982 18730 1358
rect 18672 970 18730 982
rect 18790 1358 18848 1370
rect 18790 982 18802 1358
rect 18836 982 18848 1358
rect 18790 970 18848 982
rect -7412 -66 -7350 -54
rect -7412 -442 -7400 -66
rect -7366 -442 -7350 -66
rect -7412 -454 -7350 -442
rect -7320 -66 -7254 -54
rect -7320 -442 -7304 -66
rect -7270 -442 -7254 -66
rect -7320 -454 -7254 -442
rect -7224 -66 -7158 -54
rect -7224 -442 -7208 -66
rect -7174 -442 -7158 -66
rect -7224 -454 -7158 -442
rect -7128 -66 -7062 -54
rect -7128 -442 -7112 -66
rect -7078 -442 -7062 -66
rect -7128 -454 -7062 -442
rect -7032 -66 -6966 -54
rect -7032 -442 -7016 -66
rect -6982 -442 -6966 -66
rect -7032 -454 -6966 -442
rect -6936 -66 -6870 -54
rect -6936 -442 -6920 -66
rect -6886 -442 -6870 -66
rect -6936 -454 -6870 -442
rect -6840 -66 -6774 -54
rect -6840 -442 -6824 -66
rect -6790 -442 -6774 -66
rect -6840 -454 -6774 -442
rect -6744 -66 -6678 -54
rect -6744 -442 -6728 -66
rect -6694 -442 -6678 -66
rect -6744 -454 -6678 -442
rect -6648 -66 -6582 -54
rect -6648 -442 -6632 -66
rect -6598 -442 -6582 -66
rect -6648 -454 -6582 -442
rect -6552 -66 -6486 -54
rect -6552 -442 -6536 -66
rect -6502 -442 -6486 -66
rect -6552 -454 -6486 -442
rect -6456 -66 -6394 -54
rect -6456 -442 -6440 -66
rect -6406 -442 -6394 -66
rect -6456 -454 -6394 -442
rect -7412 -684 -7350 -672
rect -7412 -1060 -7400 -684
rect -7366 -1060 -7350 -684
rect -7412 -1072 -7350 -1060
rect -7320 -684 -7254 -672
rect -7320 -1060 -7304 -684
rect -7270 -1060 -7254 -684
rect -7320 -1072 -7254 -1060
rect -7224 -684 -7158 -672
rect -7224 -1060 -7208 -684
rect -7174 -1060 -7158 -684
rect -7224 -1072 -7158 -1060
rect -7128 -684 -7062 -672
rect -7128 -1060 -7112 -684
rect -7078 -1060 -7062 -684
rect -7128 -1072 -7062 -1060
rect -7032 -684 -6966 -672
rect -7032 -1060 -7016 -684
rect -6982 -1060 -6966 -684
rect -7032 -1072 -6966 -1060
rect -6936 -684 -6870 -672
rect -6936 -1060 -6920 -684
rect -6886 -1060 -6870 -684
rect -6936 -1072 -6870 -1060
rect -6840 -684 -6774 -672
rect -6840 -1060 -6824 -684
rect -6790 -1060 -6774 -684
rect -6840 -1072 -6774 -1060
rect -6744 -684 -6678 -672
rect -6744 -1060 -6728 -684
rect -6694 -1060 -6678 -684
rect -6744 -1072 -6678 -1060
rect -6648 -684 -6582 -672
rect -6648 -1060 -6632 -684
rect -6598 -1060 -6582 -684
rect -6648 -1072 -6582 -1060
rect -6552 -684 -6486 -672
rect -6552 -1060 -6536 -684
rect -6502 -1060 -6486 -684
rect -6552 -1072 -6486 -1060
rect -6456 -684 -6394 -672
rect -6456 -1060 -6440 -684
rect -6406 -1060 -6394 -684
rect -6456 -1072 -6394 -1060
rect -7412 -1902 -7350 -1890
rect -7412 -2278 -7400 -1902
rect -7366 -2278 -7350 -1902
rect -7412 -2290 -7350 -2278
rect -7320 -1902 -7254 -1890
rect -7320 -2278 -7304 -1902
rect -7270 -2278 -7254 -1902
rect -7320 -2290 -7254 -2278
rect -7224 -1902 -7158 -1890
rect -7224 -2278 -7208 -1902
rect -7174 -2278 -7158 -1902
rect -7224 -2290 -7158 -2278
rect -7128 -1902 -7062 -1890
rect -7128 -2278 -7112 -1902
rect -7078 -2278 -7062 -1902
rect -7128 -2290 -7062 -2278
rect -7032 -1902 -6966 -1890
rect -7032 -2278 -7016 -1902
rect -6982 -2278 -6966 -1902
rect -7032 -2290 -6966 -2278
rect -6936 -1902 -6870 -1890
rect -6936 -2278 -6920 -1902
rect -6886 -2278 -6870 -1902
rect -6936 -2290 -6870 -2278
rect -6840 -1902 -6778 -1890
rect -6840 -2278 -6824 -1902
rect -6790 -2278 -6778 -1902
rect -6840 -2290 -6778 -2278
rect -7412 -2520 -7350 -2508
rect -7412 -2896 -7400 -2520
rect -7366 -2896 -7350 -2520
rect -7412 -2908 -7350 -2896
rect -7320 -2520 -7254 -2508
rect -7320 -2896 -7304 -2520
rect -7270 -2896 -7254 -2520
rect -7320 -2908 -7254 -2896
rect -7224 -2520 -7158 -2508
rect -7224 -2896 -7208 -2520
rect -7174 -2896 -7158 -2520
rect -7224 -2908 -7158 -2896
rect -7128 -2520 -7062 -2508
rect -7128 -2896 -7112 -2520
rect -7078 -2896 -7062 -2520
rect -7128 -2908 -7062 -2896
rect -7032 -2520 -6966 -2508
rect -7032 -2896 -7016 -2520
rect -6982 -2896 -6966 -2520
rect -7032 -2908 -6966 -2896
rect -6936 -2520 -6870 -2508
rect -6936 -2896 -6920 -2520
rect -6886 -2896 -6870 -2520
rect -6936 -2908 -6870 -2896
rect -6840 -2520 -6778 -2508
rect -6840 -2896 -6824 -2520
rect -6790 -2896 -6778 -2520
rect -6840 -2908 -6778 -2896
rect -6000 -8 -5800 4
rect -6000 -42 -5988 -8
rect -5812 -42 -5800 -8
rect -6000 -54 -5800 -42
rect -6000 -1666 -5800 -1654
rect -6000 -1700 -5988 -1666
rect -5812 -1700 -5800 -1666
rect -6000 -1712 -5800 -1700
rect 4222 540 4284 552
rect 4222 164 4234 540
rect 4268 164 4284 540
rect 4222 152 4284 164
rect 4314 540 4380 552
rect 4314 164 4330 540
rect 4364 164 4380 540
rect 4314 152 4380 164
rect 4410 540 4476 552
rect 4410 164 4426 540
rect 4460 164 4476 540
rect 4410 152 4476 164
rect 4506 540 4572 552
rect 4506 164 4522 540
rect 4556 164 4572 540
rect 4506 152 4572 164
rect 4602 540 4668 552
rect 4602 164 4618 540
rect 4652 164 4668 540
rect 4602 152 4668 164
rect 4698 540 4764 552
rect 4698 164 4714 540
rect 4748 164 4764 540
rect 4698 152 4764 164
rect 4794 540 4856 552
rect 4794 164 4810 540
rect 4844 164 4856 540
rect 4794 152 4856 164
rect 4222 -78 4284 -66
rect 4222 -454 4234 -78
rect 4268 -454 4284 -78
rect 4222 -466 4284 -454
rect 4314 -78 4380 -66
rect 4314 -454 4330 -78
rect 4364 -454 4380 -78
rect 4314 -466 4380 -454
rect 4410 -78 4476 -66
rect 4410 -454 4426 -78
rect 4460 -454 4476 -78
rect 4410 -466 4476 -454
rect 4506 -78 4572 -66
rect 4506 -454 4522 -78
rect 4556 -454 4572 -78
rect 4506 -466 4572 -454
rect 4602 -78 4668 -66
rect 4602 -454 4618 -78
rect 4652 -454 4668 -78
rect 4602 -466 4668 -454
rect 4698 -78 4764 -66
rect 4698 -454 4714 -78
rect 4748 -454 4764 -78
rect 4698 -466 4764 -454
rect 4794 -78 4856 -66
rect 4794 -454 4810 -78
rect 4844 -454 4856 -78
rect 4794 -466 4856 -454
rect 5262 540 5324 552
rect 5262 164 5274 540
rect 5308 164 5324 540
rect 5262 152 5324 164
rect 5354 540 5420 552
rect 5354 164 5370 540
rect 5404 164 5420 540
rect 5354 152 5420 164
rect 5450 540 5516 552
rect 5450 164 5466 540
rect 5500 164 5516 540
rect 5450 152 5516 164
rect 5546 540 5612 552
rect 5546 164 5562 540
rect 5596 164 5612 540
rect 5546 152 5612 164
rect 5642 540 5708 552
rect 5642 164 5658 540
rect 5692 164 5708 540
rect 5642 152 5708 164
rect 5738 540 5804 552
rect 5738 164 5754 540
rect 5788 164 5804 540
rect 5738 152 5804 164
rect 5834 540 5896 552
rect 5834 164 5850 540
rect 5884 164 5896 540
rect 5834 152 5896 164
rect 5262 -78 5324 -66
rect 5262 -454 5274 -78
rect 5308 -454 5324 -78
rect 5262 -466 5324 -454
rect 5354 -78 5420 -66
rect 5354 -454 5370 -78
rect 5404 -454 5420 -78
rect 5354 -466 5420 -454
rect 5450 -78 5516 -66
rect 5450 -454 5466 -78
rect 5500 -454 5516 -78
rect 5450 -466 5516 -454
rect 5546 -78 5612 -66
rect 5546 -454 5562 -78
rect 5596 -454 5612 -78
rect 5546 -466 5612 -454
rect 5642 -78 5708 -66
rect 5642 -454 5658 -78
rect 5692 -454 5708 -78
rect 5642 -466 5708 -454
rect 5738 -78 5804 -66
rect 5738 -454 5754 -78
rect 5788 -454 5804 -78
rect 5738 -466 5804 -454
rect 5834 -78 5896 -66
rect 5834 -454 5850 -78
rect 5884 -454 5896 -78
rect 5834 -466 5896 -454
rect 6302 540 6364 552
rect 6302 164 6314 540
rect 6348 164 6364 540
rect 6302 152 6364 164
rect 6394 540 6460 552
rect 6394 164 6410 540
rect 6444 164 6460 540
rect 6394 152 6460 164
rect 6490 540 6556 552
rect 6490 164 6506 540
rect 6540 164 6556 540
rect 6490 152 6556 164
rect 6586 540 6652 552
rect 6586 164 6602 540
rect 6636 164 6652 540
rect 6586 152 6652 164
rect 6682 540 6748 552
rect 6682 164 6698 540
rect 6732 164 6748 540
rect 6682 152 6748 164
rect 6778 540 6844 552
rect 6778 164 6794 540
rect 6828 164 6844 540
rect 6778 152 6844 164
rect 6874 540 6936 552
rect 6874 164 6890 540
rect 6924 164 6936 540
rect 6874 152 6936 164
rect 6302 -78 6364 -66
rect 6302 -454 6314 -78
rect 6348 -454 6364 -78
rect 6302 -466 6364 -454
rect 6394 -78 6460 -66
rect 6394 -454 6410 -78
rect 6444 -454 6460 -78
rect 6394 -466 6460 -454
rect 6490 -78 6556 -66
rect 6490 -454 6506 -78
rect 6540 -454 6556 -78
rect 6490 -466 6556 -454
rect 6586 -78 6652 -66
rect 6586 -454 6602 -78
rect 6636 -454 6652 -78
rect 6586 -466 6652 -454
rect 6682 -78 6748 -66
rect 6682 -454 6698 -78
rect 6732 -454 6748 -78
rect 6682 -466 6748 -454
rect 6778 -78 6844 -66
rect 6778 -454 6794 -78
rect 6828 -454 6844 -78
rect 6778 -466 6844 -454
rect 6874 -78 6936 -66
rect 6874 -454 6890 -78
rect 6924 -454 6936 -78
rect 6874 -466 6936 -454
rect 7342 540 7404 552
rect 7342 164 7354 540
rect 7388 164 7404 540
rect 7342 152 7404 164
rect 7434 540 7500 552
rect 7434 164 7450 540
rect 7484 164 7500 540
rect 7434 152 7500 164
rect 7530 540 7596 552
rect 7530 164 7546 540
rect 7580 164 7596 540
rect 7530 152 7596 164
rect 7626 540 7692 552
rect 7626 164 7642 540
rect 7676 164 7692 540
rect 7626 152 7692 164
rect 7722 540 7788 552
rect 7722 164 7738 540
rect 7772 164 7788 540
rect 7722 152 7788 164
rect 7818 540 7884 552
rect 7818 164 7834 540
rect 7868 164 7884 540
rect 7818 152 7884 164
rect 7914 540 7976 552
rect 7914 164 7930 540
rect 7964 164 7976 540
rect 7914 152 7976 164
rect 7342 -78 7404 -66
rect 7342 -454 7354 -78
rect 7388 -454 7404 -78
rect 7342 -466 7404 -454
rect 7434 -78 7500 -66
rect 7434 -454 7450 -78
rect 7484 -454 7500 -78
rect 7434 -466 7500 -454
rect 7530 -78 7596 -66
rect 7530 -454 7546 -78
rect 7580 -454 7596 -78
rect 7530 -466 7596 -454
rect 7626 -78 7692 -66
rect 7626 -454 7642 -78
rect 7676 -454 7692 -78
rect 7626 -466 7692 -454
rect 7722 -78 7788 -66
rect 7722 -454 7738 -78
rect 7772 -454 7788 -78
rect 7722 -466 7788 -454
rect 7818 -78 7884 -66
rect 7818 -454 7834 -78
rect 7868 -454 7884 -78
rect 7818 -466 7884 -454
rect 7914 -78 7976 -66
rect 7914 -454 7930 -78
rect 7964 -454 7976 -78
rect 7914 -466 7976 -454
rect 8382 540 8444 552
rect 8382 164 8394 540
rect 8428 164 8444 540
rect 8382 152 8444 164
rect 8474 540 8540 552
rect 8474 164 8490 540
rect 8524 164 8540 540
rect 8474 152 8540 164
rect 8570 540 8636 552
rect 8570 164 8586 540
rect 8620 164 8636 540
rect 8570 152 8636 164
rect 8666 540 8732 552
rect 8666 164 8682 540
rect 8716 164 8732 540
rect 8666 152 8732 164
rect 8762 540 8828 552
rect 8762 164 8778 540
rect 8812 164 8828 540
rect 8762 152 8828 164
rect 8858 540 8924 552
rect 8858 164 8874 540
rect 8908 164 8924 540
rect 8858 152 8924 164
rect 8954 540 9016 552
rect 8954 164 8970 540
rect 9004 164 9016 540
rect 8954 152 9016 164
rect 8382 -78 8444 -66
rect 8382 -454 8394 -78
rect 8428 -454 8444 -78
rect 8382 -466 8444 -454
rect 8474 -78 8540 -66
rect 8474 -454 8490 -78
rect 8524 -454 8540 -78
rect 8474 -466 8540 -454
rect 8570 -78 8636 -66
rect 8570 -454 8586 -78
rect 8620 -454 8636 -78
rect 8570 -466 8636 -454
rect 8666 -78 8732 -66
rect 8666 -454 8682 -78
rect 8716 -454 8732 -78
rect 8666 -466 8732 -454
rect 8762 -78 8828 -66
rect 8762 -454 8778 -78
rect 8812 -454 8828 -78
rect 8762 -466 8828 -454
rect 8858 -78 8924 -66
rect 8858 -454 8874 -78
rect 8908 -454 8924 -78
rect 8858 -466 8924 -454
rect 8954 -78 9016 -66
rect 8954 -454 8970 -78
rect 9004 -454 9016 -78
rect 8954 -466 9016 -454
rect 9422 540 9484 552
rect 9422 164 9434 540
rect 9468 164 9484 540
rect 9422 152 9484 164
rect 9514 540 9580 552
rect 9514 164 9530 540
rect 9564 164 9580 540
rect 9514 152 9580 164
rect 9610 540 9676 552
rect 9610 164 9626 540
rect 9660 164 9676 540
rect 9610 152 9676 164
rect 9706 540 9772 552
rect 9706 164 9722 540
rect 9756 164 9772 540
rect 9706 152 9772 164
rect 9802 540 9868 552
rect 9802 164 9818 540
rect 9852 164 9868 540
rect 9802 152 9868 164
rect 9898 540 9964 552
rect 9898 164 9914 540
rect 9948 164 9964 540
rect 9898 152 9964 164
rect 9994 540 10056 552
rect 9994 164 10010 540
rect 10044 164 10056 540
rect 9994 152 10056 164
rect 9422 -78 9484 -66
rect 9422 -454 9434 -78
rect 9468 -454 9484 -78
rect 9422 -466 9484 -454
rect 9514 -78 9580 -66
rect 9514 -454 9530 -78
rect 9564 -454 9580 -78
rect 9514 -466 9580 -454
rect 9610 -78 9676 -66
rect 9610 -454 9626 -78
rect 9660 -454 9676 -78
rect 9610 -466 9676 -454
rect 9706 -78 9772 -66
rect 9706 -454 9722 -78
rect 9756 -454 9772 -78
rect 9706 -466 9772 -454
rect 9802 -78 9868 -66
rect 9802 -454 9818 -78
rect 9852 -454 9868 -78
rect 9802 -466 9868 -454
rect 9898 -78 9964 -66
rect 9898 -454 9914 -78
rect 9948 -454 9964 -78
rect 9898 -466 9964 -454
rect 9994 -78 10056 -66
rect 9994 -454 10010 -78
rect 10044 -454 10056 -78
rect 9994 -466 10056 -454
rect 10462 540 10524 552
rect 10462 164 10474 540
rect 10508 164 10524 540
rect 10462 152 10524 164
rect 10554 540 10620 552
rect 10554 164 10570 540
rect 10604 164 10620 540
rect 10554 152 10620 164
rect 10650 540 10716 552
rect 10650 164 10666 540
rect 10700 164 10716 540
rect 10650 152 10716 164
rect 10746 540 10812 552
rect 10746 164 10762 540
rect 10796 164 10812 540
rect 10746 152 10812 164
rect 10842 540 10908 552
rect 10842 164 10858 540
rect 10892 164 10908 540
rect 10842 152 10908 164
rect 10938 540 11004 552
rect 10938 164 10954 540
rect 10988 164 11004 540
rect 10938 152 11004 164
rect 11034 540 11096 552
rect 11034 164 11050 540
rect 11084 164 11096 540
rect 11034 152 11096 164
rect 10462 -78 10524 -66
rect 10462 -454 10474 -78
rect 10508 -454 10524 -78
rect 10462 -466 10524 -454
rect 10554 -78 10620 -66
rect 10554 -454 10570 -78
rect 10604 -454 10620 -78
rect 10554 -466 10620 -454
rect 10650 -78 10716 -66
rect 10650 -454 10666 -78
rect 10700 -454 10716 -78
rect 10650 -466 10716 -454
rect 10746 -78 10812 -66
rect 10746 -454 10762 -78
rect 10796 -454 10812 -78
rect 10746 -466 10812 -454
rect 10842 -78 10908 -66
rect 10842 -454 10858 -78
rect 10892 -454 10908 -78
rect 10842 -466 10908 -454
rect 10938 -78 11004 -66
rect 10938 -454 10954 -78
rect 10988 -454 11004 -78
rect 10938 -466 11004 -454
rect 11034 -78 11096 -66
rect 11034 -454 11050 -78
rect 11084 -454 11096 -78
rect 11034 -466 11096 -454
rect 11842 540 11904 552
rect 11842 164 11854 540
rect 11888 164 11904 540
rect 11842 152 11904 164
rect 11934 540 12000 552
rect 11934 164 11950 540
rect 11984 164 12000 540
rect 11934 152 12000 164
rect 12030 540 12096 552
rect 12030 164 12046 540
rect 12080 164 12096 540
rect 12030 152 12096 164
rect 12126 540 12192 552
rect 12126 164 12142 540
rect 12176 164 12192 540
rect 12126 152 12192 164
rect 12222 540 12288 552
rect 12222 164 12238 540
rect 12272 164 12288 540
rect 12222 152 12288 164
rect 12318 540 12384 552
rect 12318 164 12334 540
rect 12368 164 12384 540
rect 12318 152 12384 164
rect 12414 540 12476 552
rect 12414 164 12430 540
rect 12464 164 12476 540
rect 12414 152 12476 164
rect 11842 -78 11904 -66
rect 11842 -454 11854 -78
rect 11888 -454 11904 -78
rect 11842 -466 11904 -454
rect 11934 -78 12000 -66
rect 11934 -454 11950 -78
rect 11984 -454 12000 -78
rect 11934 -466 12000 -454
rect 12030 -78 12096 -66
rect 12030 -454 12046 -78
rect 12080 -454 12096 -78
rect 12030 -466 12096 -454
rect 12126 -78 12192 -66
rect 12126 -454 12142 -78
rect 12176 -454 12192 -78
rect 12126 -466 12192 -454
rect 12222 -78 12288 -66
rect 12222 -454 12238 -78
rect 12272 -454 12288 -78
rect 12222 -466 12288 -454
rect 12318 -78 12384 -66
rect 12318 -454 12334 -78
rect 12368 -454 12384 -78
rect 12318 -466 12384 -454
rect 12414 -78 12476 -66
rect 12414 -454 12430 -78
rect 12464 -454 12476 -78
rect 12414 -466 12476 -454
rect 12882 540 12944 552
rect 12882 164 12894 540
rect 12928 164 12944 540
rect 12882 152 12944 164
rect 12974 540 13040 552
rect 12974 164 12990 540
rect 13024 164 13040 540
rect 12974 152 13040 164
rect 13070 540 13136 552
rect 13070 164 13086 540
rect 13120 164 13136 540
rect 13070 152 13136 164
rect 13166 540 13232 552
rect 13166 164 13182 540
rect 13216 164 13232 540
rect 13166 152 13232 164
rect 13262 540 13328 552
rect 13262 164 13278 540
rect 13312 164 13328 540
rect 13262 152 13328 164
rect 13358 540 13424 552
rect 13358 164 13374 540
rect 13408 164 13424 540
rect 13358 152 13424 164
rect 13454 540 13516 552
rect 13454 164 13470 540
rect 13504 164 13516 540
rect 13454 152 13516 164
rect 12882 -78 12944 -66
rect 12882 -454 12894 -78
rect 12928 -454 12944 -78
rect 12882 -466 12944 -454
rect 12974 -78 13040 -66
rect 12974 -454 12990 -78
rect 13024 -454 13040 -78
rect 12974 -466 13040 -454
rect 13070 -78 13136 -66
rect 13070 -454 13086 -78
rect 13120 -454 13136 -78
rect 13070 -466 13136 -454
rect 13166 -78 13232 -66
rect 13166 -454 13182 -78
rect 13216 -454 13232 -78
rect 13166 -466 13232 -454
rect 13262 -78 13328 -66
rect 13262 -454 13278 -78
rect 13312 -454 13328 -78
rect 13262 -466 13328 -454
rect 13358 -78 13424 -66
rect 13358 -454 13374 -78
rect 13408 -454 13424 -78
rect 13358 -466 13424 -454
rect 13454 -78 13516 -66
rect 13454 -454 13470 -78
rect 13504 -454 13516 -78
rect 13454 -466 13516 -454
rect 13922 540 13984 552
rect 13922 164 13934 540
rect 13968 164 13984 540
rect 13922 152 13984 164
rect 14014 540 14080 552
rect 14014 164 14030 540
rect 14064 164 14080 540
rect 14014 152 14080 164
rect 14110 540 14176 552
rect 14110 164 14126 540
rect 14160 164 14176 540
rect 14110 152 14176 164
rect 14206 540 14272 552
rect 14206 164 14222 540
rect 14256 164 14272 540
rect 14206 152 14272 164
rect 14302 540 14368 552
rect 14302 164 14318 540
rect 14352 164 14368 540
rect 14302 152 14368 164
rect 14398 540 14464 552
rect 14398 164 14414 540
rect 14448 164 14464 540
rect 14398 152 14464 164
rect 14494 540 14556 552
rect 14494 164 14510 540
rect 14544 164 14556 540
rect 14494 152 14556 164
rect 13922 -78 13984 -66
rect 13922 -454 13934 -78
rect 13968 -454 13984 -78
rect 13922 -466 13984 -454
rect 14014 -78 14080 -66
rect 14014 -454 14030 -78
rect 14064 -454 14080 -78
rect 14014 -466 14080 -454
rect 14110 -78 14176 -66
rect 14110 -454 14126 -78
rect 14160 -454 14176 -78
rect 14110 -466 14176 -454
rect 14206 -78 14272 -66
rect 14206 -454 14222 -78
rect 14256 -454 14272 -78
rect 14206 -466 14272 -454
rect 14302 -78 14368 -66
rect 14302 -454 14318 -78
rect 14352 -454 14368 -78
rect 14302 -466 14368 -454
rect 14398 -78 14464 -66
rect 14398 -454 14414 -78
rect 14448 -454 14464 -78
rect 14398 -466 14464 -454
rect 14494 -78 14556 -66
rect 14494 -454 14510 -78
rect 14544 -454 14556 -78
rect 14494 -466 14556 -454
rect 14962 540 15024 552
rect 14962 164 14974 540
rect 15008 164 15024 540
rect 14962 152 15024 164
rect 15054 540 15120 552
rect 15054 164 15070 540
rect 15104 164 15120 540
rect 15054 152 15120 164
rect 15150 540 15216 552
rect 15150 164 15166 540
rect 15200 164 15216 540
rect 15150 152 15216 164
rect 15246 540 15312 552
rect 15246 164 15262 540
rect 15296 164 15312 540
rect 15246 152 15312 164
rect 15342 540 15408 552
rect 15342 164 15358 540
rect 15392 164 15408 540
rect 15342 152 15408 164
rect 15438 540 15504 552
rect 15438 164 15454 540
rect 15488 164 15504 540
rect 15438 152 15504 164
rect 15534 540 15596 552
rect 15534 164 15550 540
rect 15584 164 15596 540
rect 15534 152 15596 164
rect 14962 -78 15024 -66
rect 14962 -454 14974 -78
rect 15008 -454 15024 -78
rect 14962 -466 15024 -454
rect 15054 -78 15120 -66
rect 15054 -454 15070 -78
rect 15104 -454 15120 -78
rect 15054 -466 15120 -454
rect 15150 -78 15216 -66
rect 15150 -454 15166 -78
rect 15200 -454 15216 -78
rect 15150 -466 15216 -454
rect 15246 -78 15312 -66
rect 15246 -454 15262 -78
rect 15296 -454 15312 -78
rect 15246 -466 15312 -454
rect 15342 -78 15408 -66
rect 15342 -454 15358 -78
rect 15392 -454 15408 -78
rect 15342 -466 15408 -454
rect 15438 -78 15504 -66
rect 15438 -454 15454 -78
rect 15488 -454 15504 -78
rect 15438 -466 15504 -454
rect 15534 -78 15596 -66
rect 15534 -454 15550 -78
rect 15584 -454 15596 -78
rect 15534 -466 15596 -454
rect 16002 540 16064 552
rect 16002 164 16014 540
rect 16048 164 16064 540
rect 16002 152 16064 164
rect 16094 540 16160 552
rect 16094 164 16110 540
rect 16144 164 16160 540
rect 16094 152 16160 164
rect 16190 540 16256 552
rect 16190 164 16206 540
rect 16240 164 16256 540
rect 16190 152 16256 164
rect 16286 540 16352 552
rect 16286 164 16302 540
rect 16336 164 16352 540
rect 16286 152 16352 164
rect 16382 540 16448 552
rect 16382 164 16398 540
rect 16432 164 16448 540
rect 16382 152 16448 164
rect 16478 540 16544 552
rect 16478 164 16494 540
rect 16528 164 16544 540
rect 16478 152 16544 164
rect 16574 540 16636 552
rect 16574 164 16590 540
rect 16624 164 16636 540
rect 16574 152 16636 164
rect 16002 -78 16064 -66
rect 16002 -454 16014 -78
rect 16048 -454 16064 -78
rect 16002 -466 16064 -454
rect 16094 -78 16160 -66
rect 16094 -454 16110 -78
rect 16144 -454 16160 -78
rect 16094 -466 16160 -454
rect 16190 -78 16256 -66
rect 16190 -454 16206 -78
rect 16240 -454 16256 -78
rect 16190 -466 16256 -454
rect 16286 -78 16352 -66
rect 16286 -454 16302 -78
rect 16336 -454 16352 -78
rect 16286 -466 16352 -454
rect 16382 -78 16448 -66
rect 16382 -454 16398 -78
rect 16432 -454 16448 -78
rect 16382 -466 16448 -454
rect 16478 -78 16544 -66
rect 16478 -454 16494 -78
rect 16528 -454 16544 -78
rect 16478 -466 16544 -454
rect 16574 -78 16636 -66
rect 16574 -454 16590 -78
rect 16624 -454 16636 -78
rect 16574 -466 16636 -454
rect 17042 540 17104 552
rect 17042 164 17054 540
rect 17088 164 17104 540
rect 17042 152 17104 164
rect 17134 540 17200 552
rect 17134 164 17150 540
rect 17184 164 17200 540
rect 17134 152 17200 164
rect 17230 540 17296 552
rect 17230 164 17246 540
rect 17280 164 17296 540
rect 17230 152 17296 164
rect 17326 540 17392 552
rect 17326 164 17342 540
rect 17376 164 17392 540
rect 17326 152 17392 164
rect 17422 540 17488 552
rect 17422 164 17438 540
rect 17472 164 17488 540
rect 17422 152 17488 164
rect 17518 540 17584 552
rect 17518 164 17534 540
rect 17568 164 17584 540
rect 17518 152 17584 164
rect 17614 540 17676 552
rect 17614 164 17630 540
rect 17664 164 17676 540
rect 17614 152 17676 164
rect 17042 -78 17104 -66
rect 17042 -454 17054 -78
rect 17088 -454 17104 -78
rect 17042 -466 17104 -454
rect 17134 -78 17200 -66
rect 17134 -454 17150 -78
rect 17184 -454 17200 -78
rect 17134 -466 17200 -454
rect 17230 -78 17296 -66
rect 17230 -454 17246 -78
rect 17280 -454 17296 -78
rect 17230 -466 17296 -454
rect 17326 -78 17392 -66
rect 17326 -454 17342 -78
rect 17376 -454 17392 -78
rect 17326 -466 17392 -454
rect 17422 -78 17488 -66
rect 17422 -454 17438 -78
rect 17472 -454 17488 -78
rect 17422 -466 17488 -454
rect 17518 -78 17584 -66
rect 17518 -454 17534 -78
rect 17568 -454 17584 -78
rect 17518 -466 17584 -454
rect 17614 -78 17676 -66
rect 17614 -454 17630 -78
rect 17664 -454 17676 -78
rect 17614 -466 17676 -454
rect 18082 540 18144 552
rect 18082 164 18094 540
rect 18128 164 18144 540
rect 18082 152 18144 164
rect 18174 540 18240 552
rect 18174 164 18190 540
rect 18224 164 18240 540
rect 18174 152 18240 164
rect 18270 540 18336 552
rect 18270 164 18286 540
rect 18320 164 18336 540
rect 18270 152 18336 164
rect 18366 540 18432 552
rect 18366 164 18382 540
rect 18416 164 18432 540
rect 18366 152 18432 164
rect 18462 540 18528 552
rect 18462 164 18478 540
rect 18512 164 18528 540
rect 18462 152 18528 164
rect 18558 540 18624 552
rect 18558 164 18574 540
rect 18608 164 18624 540
rect 18558 152 18624 164
rect 18654 540 18716 552
rect 18654 164 18670 540
rect 18704 164 18716 540
rect 18654 152 18716 164
rect 18082 -78 18144 -66
rect 18082 -454 18094 -78
rect 18128 -454 18144 -78
rect 18082 -466 18144 -454
rect 18174 -78 18240 -66
rect 18174 -454 18190 -78
rect 18224 -454 18240 -78
rect 18174 -466 18240 -454
rect 18270 -78 18336 -66
rect 18270 -454 18286 -78
rect 18320 -454 18336 -78
rect 18270 -466 18336 -454
rect 18366 -78 18432 -66
rect 18366 -454 18382 -78
rect 18416 -454 18432 -78
rect 18366 -466 18432 -454
rect 18462 -78 18528 -66
rect 18462 -454 18478 -78
rect 18512 -454 18528 -78
rect 18462 -466 18528 -454
rect 18558 -78 18624 -66
rect 18558 -454 18574 -78
rect 18608 -454 18624 -78
rect 18558 -466 18624 -454
rect 18654 -78 18716 -66
rect 18654 -454 18670 -78
rect 18704 -454 18716 -78
rect 18654 -466 18716 -454
rect 4222 -882 4280 -870
rect 4222 -1258 4234 -882
rect 4268 -1258 4280 -882
rect 4222 -1270 4280 -1258
rect 4340 -882 4398 -870
rect 4340 -1258 4352 -882
rect 4386 -1258 4398 -882
rect 4340 -1270 4398 -1258
rect 4458 -882 4516 -870
rect 4458 -1258 4470 -882
rect 4504 -1258 4516 -882
rect 4458 -1270 4516 -1258
rect 4576 -882 4634 -870
rect 4576 -1258 4588 -882
rect 4622 -1258 4634 -882
rect 4576 -1270 4634 -1258
rect 4694 -882 4752 -870
rect 4694 -1258 4706 -882
rect 4740 -1258 4752 -882
rect 4694 -1270 4752 -1258
rect 4812 -882 4870 -870
rect 4812 -1258 4824 -882
rect 4858 -1258 4870 -882
rect 4812 -1270 4870 -1258
rect 4930 -882 4988 -870
rect 4930 -1258 4942 -882
rect 4976 -1258 4988 -882
rect 4930 -1270 4988 -1258
rect 5262 -882 5320 -870
rect 5262 -1258 5274 -882
rect 5308 -1258 5320 -882
rect 5262 -1270 5320 -1258
rect 5380 -882 5438 -870
rect 5380 -1258 5392 -882
rect 5426 -1258 5438 -882
rect 5380 -1270 5438 -1258
rect 5498 -882 5556 -870
rect 5498 -1258 5510 -882
rect 5544 -1258 5556 -882
rect 5498 -1270 5556 -1258
rect 5616 -882 5674 -870
rect 5616 -1258 5628 -882
rect 5662 -1258 5674 -882
rect 5616 -1270 5674 -1258
rect 5734 -882 5792 -870
rect 5734 -1258 5746 -882
rect 5780 -1258 5792 -882
rect 5734 -1270 5792 -1258
rect 5852 -882 5910 -870
rect 5852 -1258 5864 -882
rect 5898 -1258 5910 -882
rect 5852 -1270 5910 -1258
rect 5970 -882 6028 -870
rect 5970 -1258 5982 -882
rect 6016 -1258 6028 -882
rect 5970 -1270 6028 -1258
rect 6302 -882 6360 -870
rect 6302 -1258 6314 -882
rect 6348 -1258 6360 -882
rect 6302 -1270 6360 -1258
rect 6420 -882 6478 -870
rect 6420 -1258 6432 -882
rect 6466 -1258 6478 -882
rect 6420 -1270 6478 -1258
rect 6538 -882 6596 -870
rect 6538 -1258 6550 -882
rect 6584 -1258 6596 -882
rect 6538 -1270 6596 -1258
rect 6656 -882 6714 -870
rect 6656 -1258 6668 -882
rect 6702 -1258 6714 -882
rect 6656 -1270 6714 -1258
rect 6774 -882 6832 -870
rect 6774 -1258 6786 -882
rect 6820 -1258 6832 -882
rect 6774 -1270 6832 -1258
rect 6892 -882 6950 -870
rect 6892 -1258 6904 -882
rect 6938 -1258 6950 -882
rect 6892 -1270 6950 -1258
rect 7010 -882 7068 -870
rect 7010 -1258 7022 -882
rect 7056 -1258 7068 -882
rect 7010 -1270 7068 -1258
rect 7342 -882 7400 -870
rect 7342 -1258 7354 -882
rect 7388 -1258 7400 -882
rect 7342 -1270 7400 -1258
rect 7460 -882 7518 -870
rect 7460 -1258 7472 -882
rect 7506 -1258 7518 -882
rect 7460 -1270 7518 -1258
rect 7578 -882 7636 -870
rect 7578 -1258 7590 -882
rect 7624 -1258 7636 -882
rect 7578 -1270 7636 -1258
rect 7696 -882 7754 -870
rect 7696 -1258 7708 -882
rect 7742 -1258 7754 -882
rect 7696 -1270 7754 -1258
rect 7814 -882 7872 -870
rect 7814 -1258 7826 -882
rect 7860 -1258 7872 -882
rect 7814 -1270 7872 -1258
rect 7932 -882 7990 -870
rect 7932 -1258 7944 -882
rect 7978 -1258 7990 -882
rect 7932 -1270 7990 -1258
rect 8050 -882 8108 -870
rect 8050 -1258 8062 -882
rect 8096 -1258 8108 -882
rect 8050 -1270 8108 -1258
rect 8382 -882 8440 -870
rect 8382 -1258 8394 -882
rect 8428 -1258 8440 -882
rect 8382 -1270 8440 -1258
rect 8500 -882 8558 -870
rect 8500 -1258 8512 -882
rect 8546 -1258 8558 -882
rect 8500 -1270 8558 -1258
rect 8618 -882 8676 -870
rect 8618 -1258 8630 -882
rect 8664 -1258 8676 -882
rect 8618 -1270 8676 -1258
rect 8736 -882 8794 -870
rect 8736 -1258 8748 -882
rect 8782 -1258 8794 -882
rect 8736 -1270 8794 -1258
rect 8854 -882 8912 -870
rect 8854 -1258 8866 -882
rect 8900 -1258 8912 -882
rect 8854 -1270 8912 -1258
rect 8972 -882 9030 -870
rect 8972 -1258 8984 -882
rect 9018 -1258 9030 -882
rect 8972 -1270 9030 -1258
rect 9090 -882 9148 -870
rect 9090 -1258 9102 -882
rect 9136 -1258 9148 -882
rect 9090 -1270 9148 -1258
rect 9422 -882 9480 -870
rect 9422 -1258 9434 -882
rect 9468 -1258 9480 -882
rect 9422 -1270 9480 -1258
rect 9540 -882 9598 -870
rect 9540 -1258 9552 -882
rect 9586 -1258 9598 -882
rect 9540 -1270 9598 -1258
rect 9658 -882 9716 -870
rect 9658 -1258 9670 -882
rect 9704 -1258 9716 -882
rect 9658 -1270 9716 -1258
rect 9776 -882 9834 -870
rect 9776 -1258 9788 -882
rect 9822 -1258 9834 -882
rect 9776 -1270 9834 -1258
rect 9894 -882 9952 -870
rect 9894 -1258 9906 -882
rect 9940 -1258 9952 -882
rect 9894 -1270 9952 -1258
rect 10012 -882 10070 -870
rect 10012 -1258 10024 -882
rect 10058 -1258 10070 -882
rect 10012 -1270 10070 -1258
rect 10130 -882 10188 -870
rect 10130 -1258 10142 -882
rect 10176 -1258 10188 -882
rect 10130 -1270 10188 -1258
rect 10462 -882 10520 -870
rect 10462 -1258 10474 -882
rect 10508 -1258 10520 -882
rect 10462 -1270 10520 -1258
rect 10580 -882 10638 -870
rect 10580 -1258 10592 -882
rect 10626 -1258 10638 -882
rect 10580 -1270 10638 -1258
rect 10698 -882 10756 -870
rect 10698 -1258 10710 -882
rect 10744 -1258 10756 -882
rect 10698 -1270 10756 -1258
rect 10816 -882 10874 -870
rect 10816 -1258 10828 -882
rect 10862 -1258 10874 -882
rect 10816 -1270 10874 -1258
rect 10934 -882 10992 -870
rect 10934 -1258 10946 -882
rect 10980 -1258 10992 -882
rect 10934 -1270 10992 -1258
rect 11052 -882 11110 -870
rect 11052 -1258 11064 -882
rect 11098 -1258 11110 -882
rect 11052 -1270 11110 -1258
rect 11170 -882 11228 -870
rect 11170 -1258 11182 -882
rect 11216 -1258 11228 -882
rect 11170 -1270 11228 -1258
rect 11842 -882 11900 -870
rect 11842 -1258 11854 -882
rect 11888 -1258 11900 -882
rect 11842 -1270 11900 -1258
rect 11960 -882 12018 -870
rect 11960 -1258 11972 -882
rect 12006 -1258 12018 -882
rect 11960 -1270 12018 -1258
rect 12078 -882 12136 -870
rect 12078 -1258 12090 -882
rect 12124 -1258 12136 -882
rect 12078 -1270 12136 -1258
rect 12196 -882 12254 -870
rect 12196 -1258 12208 -882
rect 12242 -1258 12254 -882
rect 12196 -1270 12254 -1258
rect 12314 -882 12372 -870
rect 12314 -1258 12326 -882
rect 12360 -1258 12372 -882
rect 12314 -1270 12372 -1258
rect 12432 -882 12490 -870
rect 12432 -1258 12444 -882
rect 12478 -1258 12490 -882
rect 12432 -1270 12490 -1258
rect 12550 -882 12608 -870
rect 12550 -1258 12562 -882
rect 12596 -1258 12608 -882
rect 12550 -1270 12608 -1258
rect 12882 -882 12940 -870
rect 12882 -1258 12894 -882
rect 12928 -1258 12940 -882
rect 12882 -1270 12940 -1258
rect 13000 -882 13058 -870
rect 13000 -1258 13012 -882
rect 13046 -1258 13058 -882
rect 13000 -1270 13058 -1258
rect 13118 -882 13176 -870
rect 13118 -1258 13130 -882
rect 13164 -1258 13176 -882
rect 13118 -1270 13176 -1258
rect 13236 -882 13294 -870
rect 13236 -1258 13248 -882
rect 13282 -1258 13294 -882
rect 13236 -1270 13294 -1258
rect 13354 -882 13412 -870
rect 13354 -1258 13366 -882
rect 13400 -1258 13412 -882
rect 13354 -1270 13412 -1258
rect 13472 -882 13530 -870
rect 13472 -1258 13484 -882
rect 13518 -1258 13530 -882
rect 13472 -1270 13530 -1258
rect 13590 -882 13648 -870
rect 13590 -1258 13602 -882
rect 13636 -1258 13648 -882
rect 13590 -1270 13648 -1258
rect 13922 -882 13980 -870
rect 13922 -1258 13934 -882
rect 13968 -1258 13980 -882
rect 13922 -1270 13980 -1258
rect 14040 -882 14098 -870
rect 14040 -1258 14052 -882
rect 14086 -1258 14098 -882
rect 14040 -1270 14098 -1258
rect 14158 -882 14216 -870
rect 14158 -1258 14170 -882
rect 14204 -1258 14216 -882
rect 14158 -1270 14216 -1258
rect 14276 -882 14334 -870
rect 14276 -1258 14288 -882
rect 14322 -1258 14334 -882
rect 14276 -1270 14334 -1258
rect 14394 -882 14452 -870
rect 14394 -1258 14406 -882
rect 14440 -1258 14452 -882
rect 14394 -1270 14452 -1258
rect 14512 -882 14570 -870
rect 14512 -1258 14524 -882
rect 14558 -1258 14570 -882
rect 14512 -1270 14570 -1258
rect 14630 -882 14688 -870
rect 14630 -1258 14642 -882
rect 14676 -1258 14688 -882
rect 14630 -1270 14688 -1258
rect 14962 -882 15020 -870
rect 14962 -1258 14974 -882
rect 15008 -1258 15020 -882
rect 14962 -1270 15020 -1258
rect 15080 -882 15138 -870
rect 15080 -1258 15092 -882
rect 15126 -1258 15138 -882
rect 15080 -1270 15138 -1258
rect 15198 -882 15256 -870
rect 15198 -1258 15210 -882
rect 15244 -1258 15256 -882
rect 15198 -1270 15256 -1258
rect 15316 -882 15374 -870
rect 15316 -1258 15328 -882
rect 15362 -1258 15374 -882
rect 15316 -1270 15374 -1258
rect 15434 -882 15492 -870
rect 15434 -1258 15446 -882
rect 15480 -1258 15492 -882
rect 15434 -1270 15492 -1258
rect 15552 -882 15610 -870
rect 15552 -1258 15564 -882
rect 15598 -1258 15610 -882
rect 15552 -1270 15610 -1258
rect 15670 -882 15728 -870
rect 15670 -1258 15682 -882
rect 15716 -1258 15728 -882
rect 15670 -1270 15728 -1258
rect 16002 -882 16060 -870
rect 16002 -1258 16014 -882
rect 16048 -1258 16060 -882
rect 16002 -1270 16060 -1258
rect 16120 -882 16178 -870
rect 16120 -1258 16132 -882
rect 16166 -1258 16178 -882
rect 16120 -1270 16178 -1258
rect 16238 -882 16296 -870
rect 16238 -1258 16250 -882
rect 16284 -1258 16296 -882
rect 16238 -1270 16296 -1258
rect 16356 -882 16414 -870
rect 16356 -1258 16368 -882
rect 16402 -1258 16414 -882
rect 16356 -1270 16414 -1258
rect 16474 -882 16532 -870
rect 16474 -1258 16486 -882
rect 16520 -1258 16532 -882
rect 16474 -1270 16532 -1258
rect 16592 -882 16650 -870
rect 16592 -1258 16604 -882
rect 16638 -1258 16650 -882
rect 16592 -1270 16650 -1258
rect 16710 -882 16768 -870
rect 16710 -1258 16722 -882
rect 16756 -1258 16768 -882
rect 16710 -1270 16768 -1258
rect 17042 -882 17100 -870
rect 17042 -1258 17054 -882
rect 17088 -1258 17100 -882
rect 17042 -1270 17100 -1258
rect 17160 -882 17218 -870
rect 17160 -1258 17172 -882
rect 17206 -1258 17218 -882
rect 17160 -1270 17218 -1258
rect 17278 -882 17336 -870
rect 17278 -1258 17290 -882
rect 17324 -1258 17336 -882
rect 17278 -1270 17336 -1258
rect 17396 -882 17454 -870
rect 17396 -1258 17408 -882
rect 17442 -1258 17454 -882
rect 17396 -1270 17454 -1258
rect 17514 -882 17572 -870
rect 17514 -1258 17526 -882
rect 17560 -1258 17572 -882
rect 17514 -1270 17572 -1258
rect 17632 -882 17690 -870
rect 17632 -1258 17644 -882
rect 17678 -1258 17690 -882
rect 17632 -1270 17690 -1258
rect 17750 -882 17808 -870
rect 17750 -1258 17762 -882
rect 17796 -1258 17808 -882
rect 17750 -1270 17808 -1258
rect 18082 -882 18140 -870
rect 18082 -1258 18094 -882
rect 18128 -1258 18140 -882
rect 18082 -1270 18140 -1258
rect 18200 -882 18258 -870
rect 18200 -1258 18212 -882
rect 18246 -1258 18258 -882
rect 18200 -1270 18258 -1258
rect 18318 -882 18376 -870
rect 18318 -1258 18330 -882
rect 18364 -1258 18376 -882
rect 18318 -1270 18376 -1258
rect 18436 -882 18494 -870
rect 18436 -1258 18448 -882
rect 18482 -1258 18494 -882
rect 18436 -1270 18494 -1258
rect 18554 -882 18612 -870
rect 18554 -1258 18566 -882
rect 18600 -1258 18612 -882
rect 18554 -1270 18612 -1258
rect 18672 -882 18730 -870
rect 18672 -1258 18684 -882
rect 18718 -1258 18730 -882
rect 18672 -1270 18730 -1258
rect 18790 -882 18848 -870
rect 18790 -1258 18802 -882
rect 18836 -1258 18848 -882
rect 18790 -1270 18848 -1258
rect 4222 -1700 4284 -1688
rect 4222 -2076 4234 -1700
rect 4268 -2076 4284 -1700
rect 4222 -2088 4284 -2076
rect 4314 -1700 4380 -1688
rect 4314 -2076 4330 -1700
rect 4364 -2076 4380 -1700
rect 4314 -2088 4380 -2076
rect 4410 -1700 4476 -1688
rect 4410 -2076 4426 -1700
rect 4460 -2076 4476 -1700
rect 4410 -2088 4476 -2076
rect 4506 -1700 4572 -1688
rect 4506 -2076 4522 -1700
rect 4556 -2076 4572 -1700
rect 4506 -2088 4572 -2076
rect 4602 -1700 4668 -1688
rect 4602 -2076 4618 -1700
rect 4652 -2076 4668 -1700
rect 4602 -2088 4668 -2076
rect 4698 -1700 4764 -1688
rect 4698 -2076 4714 -1700
rect 4748 -2076 4764 -1700
rect 4698 -2088 4764 -2076
rect 4794 -1700 4856 -1688
rect 4794 -2076 4810 -1700
rect 4844 -2076 4856 -1700
rect 4794 -2088 4856 -2076
rect 4222 -2318 4284 -2306
rect 4222 -2694 4234 -2318
rect 4268 -2694 4284 -2318
rect 4222 -2706 4284 -2694
rect 4314 -2318 4380 -2306
rect 4314 -2694 4330 -2318
rect 4364 -2694 4380 -2318
rect 4314 -2706 4380 -2694
rect 4410 -2318 4476 -2306
rect 4410 -2694 4426 -2318
rect 4460 -2694 4476 -2318
rect 4410 -2706 4476 -2694
rect 4506 -2318 4572 -2306
rect 4506 -2694 4522 -2318
rect 4556 -2694 4572 -2318
rect 4506 -2706 4572 -2694
rect 4602 -2318 4668 -2306
rect 4602 -2694 4618 -2318
rect 4652 -2694 4668 -2318
rect 4602 -2706 4668 -2694
rect 4698 -2318 4764 -2306
rect 4698 -2694 4714 -2318
rect 4748 -2694 4764 -2318
rect 4698 -2706 4764 -2694
rect 4794 -2318 4856 -2306
rect 4794 -2694 4810 -2318
rect 4844 -2694 4856 -2318
rect 4794 -2706 4856 -2694
rect 5262 -1700 5324 -1688
rect 5262 -2076 5274 -1700
rect 5308 -2076 5324 -1700
rect 5262 -2088 5324 -2076
rect 5354 -1700 5420 -1688
rect 5354 -2076 5370 -1700
rect 5404 -2076 5420 -1700
rect 5354 -2088 5420 -2076
rect 5450 -1700 5516 -1688
rect 5450 -2076 5466 -1700
rect 5500 -2076 5516 -1700
rect 5450 -2088 5516 -2076
rect 5546 -1700 5612 -1688
rect 5546 -2076 5562 -1700
rect 5596 -2076 5612 -1700
rect 5546 -2088 5612 -2076
rect 5642 -1700 5708 -1688
rect 5642 -2076 5658 -1700
rect 5692 -2076 5708 -1700
rect 5642 -2088 5708 -2076
rect 5738 -1700 5804 -1688
rect 5738 -2076 5754 -1700
rect 5788 -2076 5804 -1700
rect 5738 -2088 5804 -2076
rect 5834 -1700 5896 -1688
rect 5834 -2076 5850 -1700
rect 5884 -2076 5896 -1700
rect 5834 -2088 5896 -2076
rect 5262 -2318 5324 -2306
rect 5262 -2694 5274 -2318
rect 5308 -2694 5324 -2318
rect 5262 -2706 5324 -2694
rect 5354 -2318 5420 -2306
rect 5354 -2694 5370 -2318
rect 5404 -2694 5420 -2318
rect 5354 -2706 5420 -2694
rect 5450 -2318 5516 -2306
rect 5450 -2694 5466 -2318
rect 5500 -2694 5516 -2318
rect 5450 -2706 5516 -2694
rect 5546 -2318 5612 -2306
rect 5546 -2694 5562 -2318
rect 5596 -2694 5612 -2318
rect 5546 -2706 5612 -2694
rect 5642 -2318 5708 -2306
rect 5642 -2694 5658 -2318
rect 5692 -2694 5708 -2318
rect 5642 -2706 5708 -2694
rect 5738 -2318 5804 -2306
rect 5738 -2694 5754 -2318
rect 5788 -2694 5804 -2318
rect 5738 -2706 5804 -2694
rect 5834 -2318 5896 -2306
rect 5834 -2694 5850 -2318
rect 5884 -2694 5896 -2318
rect 5834 -2706 5896 -2694
rect 6302 -1700 6364 -1688
rect 6302 -2076 6314 -1700
rect 6348 -2076 6364 -1700
rect 6302 -2088 6364 -2076
rect 6394 -1700 6460 -1688
rect 6394 -2076 6410 -1700
rect 6444 -2076 6460 -1700
rect 6394 -2088 6460 -2076
rect 6490 -1700 6556 -1688
rect 6490 -2076 6506 -1700
rect 6540 -2076 6556 -1700
rect 6490 -2088 6556 -2076
rect 6586 -1700 6652 -1688
rect 6586 -2076 6602 -1700
rect 6636 -2076 6652 -1700
rect 6586 -2088 6652 -2076
rect 6682 -1700 6748 -1688
rect 6682 -2076 6698 -1700
rect 6732 -2076 6748 -1700
rect 6682 -2088 6748 -2076
rect 6778 -1700 6844 -1688
rect 6778 -2076 6794 -1700
rect 6828 -2076 6844 -1700
rect 6778 -2088 6844 -2076
rect 6874 -1700 6936 -1688
rect 6874 -2076 6890 -1700
rect 6924 -2076 6936 -1700
rect 6874 -2088 6936 -2076
rect 6302 -2318 6364 -2306
rect 6302 -2694 6314 -2318
rect 6348 -2694 6364 -2318
rect 6302 -2706 6364 -2694
rect 6394 -2318 6460 -2306
rect 6394 -2694 6410 -2318
rect 6444 -2694 6460 -2318
rect 6394 -2706 6460 -2694
rect 6490 -2318 6556 -2306
rect 6490 -2694 6506 -2318
rect 6540 -2694 6556 -2318
rect 6490 -2706 6556 -2694
rect 6586 -2318 6652 -2306
rect 6586 -2694 6602 -2318
rect 6636 -2694 6652 -2318
rect 6586 -2706 6652 -2694
rect 6682 -2318 6748 -2306
rect 6682 -2694 6698 -2318
rect 6732 -2694 6748 -2318
rect 6682 -2706 6748 -2694
rect 6778 -2318 6844 -2306
rect 6778 -2694 6794 -2318
rect 6828 -2694 6844 -2318
rect 6778 -2706 6844 -2694
rect 6874 -2318 6936 -2306
rect 6874 -2694 6890 -2318
rect 6924 -2694 6936 -2318
rect 6874 -2706 6936 -2694
rect 7342 -1700 7404 -1688
rect 7342 -2076 7354 -1700
rect 7388 -2076 7404 -1700
rect 7342 -2088 7404 -2076
rect 7434 -1700 7500 -1688
rect 7434 -2076 7450 -1700
rect 7484 -2076 7500 -1700
rect 7434 -2088 7500 -2076
rect 7530 -1700 7596 -1688
rect 7530 -2076 7546 -1700
rect 7580 -2076 7596 -1700
rect 7530 -2088 7596 -2076
rect 7626 -1700 7692 -1688
rect 7626 -2076 7642 -1700
rect 7676 -2076 7692 -1700
rect 7626 -2088 7692 -2076
rect 7722 -1700 7788 -1688
rect 7722 -2076 7738 -1700
rect 7772 -2076 7788 -1700
rect 7722 -2088 7788 -2076
rect 7818 -1700 7884 -1688
rect 7818 -2076 7834 -1700
rect 7868 -2076 7884 -1700
rect 7818 -2088 7884 -2076
rect 7914 -1700 7976 -1688
rect 7914 -2076 7930 -1700
rect 7964 -2076 7976 -1700
rect 7914 -2088 7976 -2076
rect 7342 -2318 7404 -2306
rect 7342 -2694 7354 -2318
rect 7388 -2694 7404 -2318
rect 7342 -2706 7404 -2694
rect 7434 -2318 7500 -2306
rect 7434 -2694 7450 -2318
rect 7484 -2694 7500 -2318
rect 7434 -2706 7500 -2694
rect 7530 -2318 7596 -2306
rect 7530 -2694 7546 -2318
rect 7580 -2694 7596 -2318
rect 7530 -2706 7596 -2694
rect 7626 -2318 7692 -2306
rect 7626 -2694 7642 -2318
rect 7676 -2694 7692 -2318
rect 7626 -2706 7692 -2694
rect 7722 -2318 7788 -2306
rect 7722 -2694 7738 -2318
rect 7772 -2694 7788 -2318
rect 7722 -2706 7788 -2694
rect 7818 -2318 7884 -2306
rect 7818 -2694 7834 -2318
rect 7868 -2694 7884 -2318
rect 7818 -2706 7884 -2694
rect 7914 -2318 7976 -2306
rect 7914 -2694 7930 -2318
rect 7964 -2694 7976 -2318
rect 7914 -2706 7976 -2694
rect 8382 -1700 8444 -1688
rect 8382 -2076 8394 -1700
rect 8428 -2076 8444 -1700
rect 8382 -2088 8444 -2076
rect 8474 -1700 8540 -1688
rect 8474 -2076 8490 -1700
rect 8524 -2076 8540 -1700
rect 8474 -2088 8540 -2076
rect 8570 -1700 8636 -1688
rect 8570 -2076 8586 -1700
rect 8620 -2076 8636 -1700
rect 8570 -2088 8636 -2076
rect 8666 -1700 8732 -1688
rect 8666 -2076 8682 -1700
rect 8716 -2076 8732 -1700
rect 8666 -2088 8732 -2076
rect 8762 -1700 8828 -1688
rect 8762 -2076 8778 -1700
rect 8812 -2076 8828 -1700
rect 8762 -2088 8828 -2076
rect 8858 -1700 8924 -1688
rect 8858 -2076 8874 -1700
rect 8908 -2076 8924 -1700
rect 8858 -2088 8924 -2076
rect 8954 -1700 9016 -1688
rect 8954 -2076 8970 -1700
rect 9004 -2076 9016 -1700
rect 8954 -2088 9016 -2076
rect 8382 -2318 8444 -2306
rect 8382 -2694 8394 -2318
rect 8428 -2694 8444 -2318
rect 8382 -2706 8444 -2694
rect 8474 -2318 8540 -2306
rect 8474 -2694 8490 -2318
rect 8524 -2694 8540 -2318
rect 8474 -2706 8540 -2694
rect 8570 -2318 8636 -2306
rect 8570 -2694 8586 -2318
rect 8620 -2694 8636 -2318
rect 8570 -2706 8636 -2694
rect 8666 -2318 8732 -2306
rect 8666 -2694 8682 -2318
rect 8716 -2694 8732 -2318
rect 8666 -2706 8732 -2694
rect 8762 -2318 8828 -2306
rect 8762 -2694 8778 -2318
rect 8812 -2694 8828 -2318
rect 8762 -2706 8828 -2694
rect 8858 -2318 8924 -2306
rect 8858 -2694 8874 -2318
rect 8908 -2694 8924 -2318
rect 8858 -2706 8924 -2694
rect 8954 -2318 9016 -2306
rect 8954 -2694 8970 -2318
rect 9004 -2694 9016 -2318
rect 8954 -2706 9016 -2694
rect 11842 -1700 11904 -1688
rect 11842 -2076 11854 -1700
rect 11888 -2076 11904 -1700
rect 11842 -2088 11904 -2076
rect 11934 -1700 12000 -1688
rect 11934 -2076 11950 -1700
rect 11984 -2076 12000 -1700
rect 11934 -2088 12000 -2076
rect 12030 -1700 12096 -1688
rect 12030 -2076 12046 -1700
rect 12080 -2076 12096 -1700
rect 12030 -2088 12096 -2076
rect 12126 -1700 12192 -1688
rect 12126 -2076 12142 -1700
rect 12176 -2076 12192 -1700
rect 12126 -2088 12192 -2076
rect 12222 -1700 12288 -1688
rect 12222 -2076 12238 -1700
rect 12272 -2076 12288 -1700
rect 12222 -2088 12288 -2076
rect 12318 -1700 12384 -1688
rect 12318 -2076 12334 -1700
rect 12368 -2076 12384 -1700
rect 12318 -2088 12384 -2076
rect 12414 -1700 12476 -1688
rect 12414 -2076 12430 -1700
rect 12464 -2076 12476 -1700
rect 12414 -2088 12476 -2076
rect 11842 -2318 11904 -2306
rect 11842 -2694 11854 -2318
rect 11888 -2694 11904 -2318
rect 11842 -2706 11904 -2694
rect 11934 -2318 12000 -2306
rect 11934 -2694 11950 -2318
rect 11984 -2694 12000 -2318
rect 11934 -2706 12000 -2694
rect 12030 -2318 12096 -2306
rect 12030 -2694 12046 -2318
rect 12080 -2694 12096 -2318
rect 12030 -2706 12096 -2694
rect 12126 -2318 12192 -2306
rect 12126 -2694 12142 -2318
rect 12176 -2694 12192 -2318
rect 12126 -2706 12192 -2694
rect 12222 -2318 12288 -2306
rect 12222 -2694 12238 -2318
rect 12272 -2694 12288 -2318
rect 12222 -2706 12288 -2694
rect 12318 -2318 12384 -2306
rect 12318 -2694 12334 -2318
rect 12368 -2694 12384 -2318
rect 12318 -2706 12384 -2694
rect 12414 -2318 12476 -2306
rect 12414 -2694 12430 -2318
rect 12464 -2694 12476 -2318
rect 12414 -2706 12476 -2694
rect 12882 -1700 12944 -1688
rect 12882 -2076 12894 -1700
rect 12928 -2076 12944 -1700
rect 12882 -2088 12944 -2076
rect 12974 -1700 13040 -1688
rect 12974 -2076 12990 -1700
rect 13024 -2076 13040 -1700
rect 12974 -2088 13040 -2076
rect 13070 -1700 13136 -1688
rect 13070 -2076 13086 -1700
rect 13120 -2076 13136 -1700
rect 13070 -2088 13136 -2076
rect 13166 -1700 13232 -1688
rect 13166 -2076 13182 -1700
rect 13216 -2076 13232 -1700
rect 13166 -2088 13232 -2076
rect 13262 -1700 13328 -1688
rect 13262 -2076 13278 -1700
rect 13312 -2076 13328 -1700
rect 13262 -2088 13328 -2076
rect 13358 -1700 13424 -1688
rect 13358 -2076 13374 -1700
rect 13408 -2076 13424 -1700
rect 13358 -2088 13424 -2076
rect 13454 -1700 13516 -1688
rect 13454 -2076 13470 -1700
rect 13504 -2076 13516 -1700
rect 13454 -2088 13516 -2076
rect 12882 -2318 12944 -2306
rect 12882 -2694 12894 -2318
rect 12928 -2694 12944 -2318
rect 12882 -2706 12944 -2694
rect 12974 -2318 13040 -2306
rect 12974 -2694 12990 -2318
rect 13024 -2694 13040 -2318
rect 12974 -2706 13040 -2694
rect 13070 -2318 13136 -2306
rect 13070 -2694 13086 -2318
rect 13120 -2694 13136 -2318
rect 13070 -2706 13136 -2694
rect 13166 -2318 13232 -2306
rect 13166 -2694 13182 -2318
rect 13216 -2694 13232 -2318
rect 13166 -2706 13232 -2694
rect 13262 -2318 13328 -2306
rect 13262 -2694 13278 -2318
rect 13312 -2694 13328 -2318
rect 13262 -2706 13328 -2694
rect 13358 -2318 13424 -2306
rect 13358 -2694 13374 -2318
rect 13408 -2694 13424 -2318
rect 13358 -2706 13424 -2694
rect 13454 -2318 13516 -2306
rect 13454 -2694 13470 -2318
rect 13504 -2694 13516 -2318
rect 13454 -2706 13516 -2694
rect 13922 -1700 13984 -1688
rect 13922 -2076 13934 -1700
rect 13968 -2076 13984 -1700
rect 13922 -2088 13984 -2076
rect 14014 -1700 14080 -1688
rect 14014 -2076 14030 -1700
rect 14064 -2076 14080 -1700
rect 14014 -2088 14080 -2076
rect 14110 -1700 14176 -1688
rect 14110 -2076 14126 -1700
rect 14160 -2076 14176 -1700
rect 14110 -2088 14176 -2076
rect 14206 -1700 14272 -1688
rect 14206 -2076 14222 -1700
rect 14256 -2076 14272 -1700
rect 14206 -2088 14272 -2076
rect 14302 -1700 14368 -1688
rect 14302 -2076 14318 -1700
rect 14352 -2076 14368 -1700
rect 14302 -2088 14368 -2076
rect 14398 -1700 14464 -1688
rect 14398 -2076 14414 -1700
rect 14448 -2076 14464 -1700
rect 14398 -2088 14464 -2076
rect 14494 -1700 14556 -1688
rect 14494 -2076 14510 -1700
rect 14544 -2076 14556 -1700
rect 14494 -2088 14556 -2076
rect 13922 -2318 13984 -2306
rect 13922 -2694 13934 -2318
rect 13968 -2694 13984 -2318
rect 13922 -2706 13984 -2694
rect 14014 -2318 14080 -2306
rect 14014 -2694 14030 -2318
rect 14064 -2694 14080 -2318
rect 14014 -2706 14080 -2694
rect 14110 -2318 14176 -2306
rect 14110 -2694 14126 -2318
rect 14160 -2694 14176 -2318
rect 14110 -2706 14176 -2694
rect 14206 -2318 14272 -2306
rect 14206 -2694 14222 -2318
rect 14256 -2694 14272 -2318
rect 14206 -2706 14272 -2694
rect 14302 -2318 14368 -2306
rect 14302 -2694 14318 -2318
rect 14352 -2694 14368 -2318
rect 14302 -2706 14368 -2694
rect 14398 -2318 14464 -2306
rect 14398 -2694 14414 -2318
rect 14448 -2694 14464 -2318
rect 14398 -2706 14464 -2694
rect 14494 -2318 14556 -2306
rect 14494 -2694 14510 -2318
rect 14544 -2694 14556 -2318
rect 14494 -2706 14556 -2694
rect 14962 -1700 15024 -1688
rect 14962 -2076 14974 -1700
rect 15008 -2076 15024 -1700
rect 14962 -2088 15024 -2076
rect 15054 -1700 15120 -1688
rect 15054 -2076 15070 -1700
rect 15104 -2076 15120 -1700
rect 15054 -2088 15120 -2076
rect 15150 -1700 15216 -1688
rect 15150 -2076 15166 -1700
rect 15200 -2076 15216 -1700
rect 15150 -2088 15216 -2076
rect 15246 -1700 15312 -1688
rect 15246 -2076 15262 -1700
rect 15296 -2076 15312 -1700
rect 15246 -2088 15312 -2076
rect 15342 -1700 15408 -1688
rect 15342 -2076 15358 -1700
rect 15392 -2076 15408 -1700
rect 15342 -2088 15408 -2076
rect 15438 -1700 15504 -1688
rect 15438 -2076 15454 -1700
rect 15488 -2076 15504 -1700
rect 15438 -2088 15504 -2076
rect 15534 -1700 15596 -1688
rect 15534 -2076 15550 -1700
rect 15584 -2076 15596 -1700
rect 15534 -2088 15596 -2076
rect 14962 -2318 15024 -2306
rect 14962 -2694 14974 -2318
rect 15008 -2694 15024 -2318
rect 14962 -2706 15024 -2694
rect 15054 -2318 15120 -2306
rect 15054 -2694 15070 -2318
rect 15104 -2694 15120 -2318
rect 15054 -2706 15120 -2694
rect 15150 -2318 15216 -2306
rect 15150 -2694 15166 -2318
rect 15200 -2694 15216 -2318
rect 15150 -2706 15216 -2694
rect 15246 -2318 15312 -2306
rect 15246 -2694 15262 -2318
rect 15296 -2694 15312 -2318
rect 15246 -2706 15312 -2694
rect 15342 -2318 15408 -2306
rect 15342 -2694 15358 -2318
rect 15392 -2694 15408 -2318
rect 15342 -2706 15408 -2694
rect 15438 -2318 15504 -2306
rect 15438 -2694 15454 -2318
rect 15488 -2694 15504 -2318
rect 15438 -2706 15504 -2694
rect 15534 -2318 15596 -2306
rect 15534 -2694 15550 -2318
rect 15584 -2694 15596 -2318
rect 15534 -2706 15596 -2694
rect 16002 -1700 16064 -1688
rect 16002 -2076 16014 -1700
rect 16048 -2076 16064 -1700
rect 16002 -2088 16064 -2076
rect 16094 -1700 16160 -1688
rect 16094 -2076 16110 -1700
rect 16144 -2076 16160 -1700
rect 16094 -2088 16160 -2076
rect 16190 -1700 16256 -1688
rect 16190 -2076 16206 -1700
rect 16240 -2076 16256 -1700
rect 16190 -2088 16256 -2076
rect 16286 -1700 16352 -1688
rect 16286 -2076 16302 -1700
rect 16336 -2076 16352 -1700
rect 16286 -2088 16352 -2076
rect 16382 -1700 16448 -1688
rect 16382 -2076 16398 -1700
rect 16432 -2076 16448 -1700
rect 16382 -2088 16448 -2076
rect 16478 -1700 16544 -1688
rect 16478 -2076 16494 -1700
rect 16528 -2076 16544 -1700
rect 16478 -2088 16544 -2076
rect 16574 -1700 16636 -1688
rect 16574 -2076 16590 -1700
rect 16624 -2076 16636 -1700
rect 16574 -2088 16636 -2076
rect 16002 -2318 16064 -2306
rect 16002 -2694 16014 -2318
rect 16048 -2694 16064 -2318
rect 16002 -2706 16064 -2694
rect 16094 -2318 16160 -2306
rect 16094 -2694 16110 -2318
rect 16144 -2694 16160 -2318
rect 16094 -2706 16160 -2694
rect 16190 -2318 16256 -2306
rect 16190 -2694 16206 -2318
rect 16240 -2694 16256 -2318
rect 16190 -2706 16256 -2694
rect 16286 -2318 16352 -2306
rect 16286 -2694 16302 -2318
rect 16336 -2694 16352 -2318
rect 16286 -2706 16352 -2694
rect 16382 -2318 16448 -2306
rect 16382 -2694 16398 -2318
rect 16432 -2694 16448 -2318
rect 16382 -2706 16448 -2694
rect 16478 -2318 16544 -2306
rect 16478 -2694 16494 -2318
rect 16528 -2694 16544 -2318
rect 16478 -2706 16544 -2694
rect 16574 -2318 16636 -2306
rect 16574 -2694 16590 -2318
rect 16624 -2694 16636 -2318
rect 16574 -2706 16636 -2694
rect -7412 -3324 -7354 -3312
rect -7412 -3700 -7400 -3324
rect -7366 -3700 -7354 -3324
rect -7412 -3712 -7354 -3700
rect -7294 -3324 -7236 -3312
rect -7294 -3700 -7282 -3324
rect -7248 -3700 -7236 -3324
rect -7294 -3712 -7236 -3700
rect -7176 -3324 -7118 -3312
rect -7176 -3700 -7164 -3324
rect -7130 -3700 -7118 -3324
rect -7176 -3712 -7118 -3700
rect -7058 -3324 -7000 -3312
rect -7058 -3700 -7046 -3324
rect -7012 -3700 -7000 -3324
rect -7058 -3712 -7000 -3700
rect -6940 -3324 -6882 -3312
rect -6940 -3700 -6928 -3324
rect -6894 -3700 -6882 -3324
rect -6940 -3712 -6882 -3700
rect -6822 -3324 -6764 -3312
rect -6822 -3700 -6810 -3324
rect -6776 -3700 -6764 -3324
rect -6822 -3712 -6764 -3700
rect -6704 -3324 -6646 -3312
rect -6704 -3700 -6692 -3324
rect -6658 -3700 -6646 -3324
rect -6704 -3712 -6646 -3700
rect 4222 -3122 4280 -3110
rect 4222 -3498 4234 -3122
rect 4268 -3498 4280 -3122
rect 4222 -3510 4280 -3498
rect 4340 -3122 4398 -3110
rect 4340 -3498 4352 -3122
rect 4386 -3498 4398 -3122
rect 4340 -3510 4398 -3498
rect 4458 -3122 4516 -3110
rect 4458 -3498 4470 -3122
rect 4504 -3498 4516 -3122
rect 4458 -3510 4516 -3498
rect 4576 -3122 4634 -3110
rect 4576 -3498 4588 -3122
rect 4622 -3498 4634 -3122
rect 4576 -3510 4634 -3498
rect 4694 -3122 4752 -3110
rect 4694 -3498 4706 -3122
rect 4740 -3498 4752 -3122
rect 4694 -3510 4752 -3498
rect 4812 -3122 4870 -3110
rect 4812 -3498 4824 -3122
rect 4858 -3498 4870 -3122
rect 4812 -3510 4870 -3498
rect 4930 -3122 4988 -3110
rect 4930 -3498 4942 -3122
rect 4976 -3498 4988 -3122
rect 4930 -3510 4988 -3498
rect 5262 -3122 5320 -3110
rect 5262 -3498 5274 -3122
rect 5308 -3498 5320 -3122
rect 5262 -3510 5320 -3498
rect 5380 -3122 5438 -3110
rect 5380 -3498 5392 -3122
rect 5426 -3498 5438 -3122
rect 5380 -3510 5438 -3498
rect 5498 -3122 5556 -3110
rect 5498 -3498 5510 -3122
rect 5544 -3498 5556 -3122
rect 5498 -3510 5556 -3498
rect 5616 -3122 5674 -3110
rect 5616 -3498 5628 -3122
rect 5662 -3498 5674 -3122
rect 5616 -3510 5674 -3498
rect 5734 -3122 5792 -3110
rect 5734 -3498 5746 -3122
rect 5780 -3498 5792 -3122
rect 5734 -3510 5792 -3498
rect 5852 -3122 5910 -3110
rect 5852 -3498 5864 -3122
rect 5898 -3498 5910 -3122
rect 5852 -3510 5910 -3498
rect 5970 -3122 6028 -3110
rect 5970 -3498 5982 -3122
rect 6016 -3498 6028 -3122
rect 5970 -3510 6028 -3498
rect 6302 -3122 6360 -3110
rect 6302 -3498 6314 -3122
rect 6348 -3498 6360 -3122
rect 6302 -3510 6360 -3498
rect 6420 -3122 6478 -3110
rect 6420 -3498 6432 -3122
rect 6466 -3498 6478 -3122
rect 6420 -3510 6478 -3498
rect 6538 -3122 6596 -3110
rect 6538 -3498 6550 -3122
rect 6584 -3498 6596 -3122
rect 6538 -3510 6596 -3498
rect 6656 -3122 6714 -3110
rect 6656 -3498 6668 -3122
rect 6702 -3498 6714 -3122
rect 6656 -3510 6714 -3498
rect 6774 -3122 6832 -3110
rect 6774 -3498 6786 -3122
rect 6820 -3498 6832 -3122
rect 6774 -3510 6832 -3498
rect 6892 -3122 6950 -3110
rect 6892 -3498 6904 -3122
rect 6938 -3498 6950 -3122
rect 6892 -3510 6950 -3498
rect 7010 -3122 7068 -3110
rect 7010 -3498 7022 -3122
rect 7056 -3498 7068 -3122
rect 7010 -3510 7068 -3498
rect 7342 -3122 7400 -3110
rect 7342 -3498 7354 -3122
rect 7388 -3498 7400 -3122
rect 7342 -3510 7400 -3498
rect 7460 -3122 7518 -3110
rect 7460 -3498 7472 -3122
rect 7506 -3498 7518 -3122
rect 7460 -3510 7518 -3498
rect 7578 -3122 7636 -3110
rect 7578 -3498 7590 -3122
rect 7624 -3498 7636 -3122
rect 7578 -3510 7636 -3498
rect 7696 -3122 7754 -3110
rect 7696 -3498 7708 -3122
rect 7742 -3498 7754 -3122
rect 7696 -3510 7754 -3498
rect 7814 -3122 7872 -3110
rect 7814 -3498 7826 -3122
rect 7860 -3498 7872 -3122
rect 7814 -3510 7872 -3498
rect 7932 -3122 7990 -3110
rect 7932 -3498 7944 -3122
rect 7978 -3498 7990 -3122
rect 7932 -3510 7990 -3498
rect 8050 -3122 8108 -3110
rect 8050 -3498 8062 -3122
rect 8096 -3498 8108 -3122
rect 8050 -3510 8108 -3498
rect 8382 -3122 8440 -3110
rect 8382 -3498 8394 -3122
rect 8428 -3498 8440 -3122
rect 8382 -3510 8440 -3498
rect 8500 -3122 8558 -3110
rect 8500 -3498 8512 -3122
rect 8546 -3498 8558 -3122
rect 8500 -3510 8558 -3498
rect 8618 -3122 8676 -3110
rect 8618 -3498 8630 -3122
rect 8664 -3498 8676 -3122
rect 8618 -3510 8676 -3498
rect 8736 -3122 8794 -3110
rect 8736 -3498 8748 -3122
rect 8782 -3498 8794 -3122
rect 8736 -3510 8794 -3498
rect 8854 -3122 8912 -3110
rect 8854 -3498 8866 -3122
rect 8900 -3498 8912 -3122
rect 8854 -3510 8912 -3498
rect 8972 -3122 9030 -3110
rect 8972 -3498 8984 -3122
rect 9018 -3498 9030 -3122
rect 8972 -3510 9030 -3498
rect 9090 -3122 9148 -3110
rect 9090 -3498 9102 -3122
rect 9136 -3498 9148 -3122
rect 9090 -3510 9148 -3498
rect 11842 -3122 11900 -3110
rect 11842 -3498 11854 -3122
rect 11888 -3498 11900 -3122
rect 11842 -3510 11900 -3498
rect 11960 -3122 12018 -3110
rect 11960 -3498 11972 -3122
rect 12006 -3498 12018 -3122
rect 11960 -3510 12018 -3498
rect 12078 -3122 12136 -3110
rect 12078 -3498 12090 -3122
rect 12124 -3498 12136 -3122
rect 12078 -3510 12136 -3498
rect 12196 -3122 12254 -3110
rect 12196 -3498 12208 -3122
rect 12242 -3498 12254 -3122
rect 12196 -3510 12254 -3498
rect 12314 -3122 12372 -3110
rect 12314 -3498 12326 -3122
rect 12360 -3498 12372 -3122
rect 12314 -3510 12372 -3498
rect 12432 -3122 12490 -3110
rect 12432 -3498 12444 -3122
rect 12478 -3498 12490 -3122
rect 12432 -3510 12490 -3498
rect 12550 -3122 12608 -3110
rect 12550 -3498 12562 -3122
rect 12596 -3498 12608 -3122
rect 12550 -3510 12608 -3498
rect 12882 -3122 12940 -3110
rect 12882 -3498 12894 -3122
rect 12928 -3498 12940 -3122
rect 12882 -3510 12940 -3498
rect 13000 -3122 13058 -3110
rect 13000 -3498 13012 -3122
rect 13046 -3498 13058 -3122
rect 13000 -3510 13058 -3498
rect 13118 -3122 13176 -3110
rect 13118 -3498 13130 -3122
rect 13164 -3498 13176 -3122
rect 13118 -3510 13176 -3498
rect 13236 -3122 13294 -3110
rect 13236 -3498 13248 -3122
rect 13282 -3498 13294 -3122
rect 13236 -3510 13294 -3498
rect 13354 -3122 13412 -3110
rect 13354 -3498 13366 -3122
rect 13400 -3498 13412 -3122
rect 13354 -3510 13412 -3498
rect 13472 -3122 13530 -3110
rect 13472 -3498 13484 -3122
rect 13518 -3498 13530 -3122
rect 13472 -3510 13530 -3498
rect 13590 -3122 13648 -3110
rect 13590 -3498 13602 -3122
rect 13636 -3498 13648 -3122
rect 13590 -3510 13648 -3498
rect 13922 -3122 13980 -3110
rect 13922 -3498 13934 -3122
rect 13968 -3498 13980 -3122
rect 13922 -3510 13980 -3498
rect 14040 -3122 14098 -3110
rect 14040 -3498 14052 -3122
rect 14086 -3498 14098 -3122
rect 14040 -3510 14098 -3498
rect 14158 -3122 14216 -3110
rect 14158 -3498 14170 -3122
rect 14204 -3498 14216 -3122
rect 14158 -3510 14216 -3498
rect 14276 -3122 14334 -3110
rect 14276 -3498 14288 -3122
rect 14322 -3498 14334 -3122
rect 14276 -3510 14334 -3498
rect 14394 -3122 14452 -3110
rect 14394 -3498 14406 -3122
rect 14440 -3498 14452 -3122
rect 14394 -3510 14452 -3498
rect 14512 -3122 14570 -3110
rect 14512 -3498 14524 -3122
rect 14558 -3498 14570 -3122
rect 14512 -3510 14570 -3498
rect 14630 -3122 14688 -3110
rect 14630 -3498 14642 -3122
rect 14676 -3498 14688 -3122
rect 14630 -3510 14688 -3498
rect 14962 -3122 15020 -3110
rect 14962 -3498 14974 -3122
rect 15008 -3498 15020 -3122
rect 14962 -3510 15020 -3498
rect 15080 -3122 15138 -3110
rect 15080 -3498 15092 -3122
rect 15126 -3498 15138 -3122
rect 15080 -3510 15138 -3498
rect 15198 -3122 15256 -3110
rect 15198 -3498 15210 -3122
rect 15244 -3498 15256 -3122
rect 15198 -3510 15256 -3498
rect 15316 -3122 15374 -3110
rect 15316 -3498 15328 -3122
rect 15362 -3498 15374 -3122
rect 15316 -3510 15374 -3498
rect 15434 -3122 15492 -3110
rect 15434 -3498 15446 -3122
rect 15480 -3498 15492 -3122
rect 15434 -3510 15492 -3498
rect 15552 -3122 15610 -3110
rect 15552 -3498 15564 -3122
rect 15598 -3498 15610 -3122
rect 15552 -3510 15610 -3498
rect 15670 -3122 15728 -3110
rect 15670 -3498 15682 -3122
rect 15716 -3498 15728 -3122
rect 15670 -3510 15728 -3498
rect 16002 -3122 16060 -3110
rect 16002 -3498 16014 -3122
rect 16048 -3498 16060 -3122
rect 16002 -3510 16060 -3498
rect 16120 -3122 16178 -3110
rect 16120 -3498 16132 -3122
rect 16166 -3498 16178 -3122
rect 16120 -3510 16178 -3498
rect 16238 -3122 16296 -3110
rect 16238 -3498 16250 -3122
rect 16284 -3498 16296 -3122
rect 16238 -3510 16296 -3498
rect 16356 -3122 16414 -3110
rect 16356 -3498 16368 -3122
rect 16402 -3498 16414 -3122
rect 16356 -3510 16414 -3498
rect 16474 -3122 16532 -3110
rect 16474 -3498 16486 -3122
rect 16520 -3498 16532 -3122
rect 16474 -3510 16532 -3498
rect 16592 -3122 16650 -3110
rect 16592 -3498 16604 -3122
rect 16638 -3498 16650 -3122
rect 16592 -3510 16650 -3498
rect 16710 -3122 16768 -3110
rect 16710 -3498 16722 -3122
rect 16756 -3498 16768 -3122
rect 16710 -3510 16768 -3498
<< ndiffc >>
rect -1030 3222 -996 3598
rect -934 3222 -900 3598
rect -838 3222 -804 3598
rect -742 3222 -708 3598
rect -646 3222 -612 3598
rect -550 3222 -516 3598
rect -454 3222 -420 3598
rect -358 3222 -324 3598
rect -262 3222 -228 3598
rect -166 3222 -132 3598
rect -70 3222 -36 3598
rect 1770 3222 1804 3598
rect 1866 3222 1900 3598
rect 1962 3222 1996 3598
rect 2058 3222 2092 3598
rect 2154 3222 2188 3598
rect 2250 3222 2284 3598
rect 2346 3222 2380 3598
rect 2442 3222 2476 3598
rect 2538 3222 2572 3598
rect 2634 3222 2668 3598
rect 2730 3222 2764 3598
rect 4434 5076 4468 5452
rect 4530 5076 4564 5452
rect 4626 5076 4660 5452
rect 4722 5076 4756 5452
rect 4818 5076 4852 5452
rect 4914 5076 4948 5452
rect 5010 5076 5044 5452
rect 5106 5076 5140 5452
rect 5202 5076 5236 5452
rect 5298 5076 5332 5452
rect 5394 5076 5428 5452
rect 5490 5076 5524 5452
rect 5586 5076 5620 5452
rect 5682 5076 5716 5452
rect 5778 5076 5812 5452
rect 5874 5076 5908 5452
rect 5970 5076 6004 5452
rect 6066 5076 6100 5452
rect 6162 5076 6196 5452
rect 6258 5076 6292 5452
rect 6354 5076 6388 5452
rect 6450 5076 6484 5452
rect 6546 5076 6580 5452
rect 6642 5076 6676 5452
rect 6738 5076 6772 5452
rect 6834 5076 6868 5452
rect 6930 5076 6964 5452
rect 7026 5076 7060 5452
rect 7122 5076 7156 5452
rect 7218 5076 7252 5452
rect 7314 5076 7348 5452
rect 4434 4458 4468 4834
rect 4530 4458 4564 4834
rect 4626 4458 4660 4834
rect 4722 4458 4756 4834
rect 4818 4458 4852 4834
rect 4914 4458 4948 4834
rect 5010 4458 5044 4834
rect 5106 4458 5140 4834
rect 5202 4458 5236 4834
rect 5298 4458 5332 4834
rect 5394 4458 5428 4834
rect 5490 4458 5524 4834
rect 5586 4458 5620 4834
rect 5682 4458 5716 4834
rect 5778 4458 5812 4834
rect 5874 4458 5908 4834
rect 5970 4458 6004 4834
rect 6066 4458 6100 4834
rect 6162 4458 6196 4834
rect 6258 4458 6292 4834
rect 6354 4458 6388 4834
rect 6450 4458 6484 4834
rect 6546 4458 6580 4834
rect 6642 4458 6676 4834
rect 6738 4458 6772 4834
rect 6834 4458 6868 4834
rect 6930 4458 6964 4834
rect 7026 4458 7060 4834
rect 7122 4458 7156 4834
rect 7218 4458 7252 4834
rect 7314 4458 7348 4834
rect 4434 3840 4468 4216
rect 4530 3840 4564 4216
rect 4626 3840 4660 4216
rect 4722 3840 4756 4216
rect 4818 3840 4852 4216
rect 4914 3840 4948 4216
rect 5010 3840 5044 4216
rect 5106 3840 5140 4216
rect 5202 3840 5236 4216
rect 5298 3840 5332 4216
rect 5394 3840 5428 4216
rect 5490 3840 5524 4216
rect 5586 3840 5620 4216
rect 5682 3840 5716 4216
rect 5778 3840 5812 4216
rect 5874 3840 5908 4216
rect 5970 3840 6004 4216
rect 6066 3840 6100 4216
rect 6162 3840 6196 4216
rect 6258 3840 6292 4216
rect 6354 3840 6388 4216
rect 6450 3840 6484 4216
rect 6546 3840 6580 4216
rect 6642 3840 6676 4216
rect 6738 3840 6772 4216
rect 6834 3840 6868 4216
rect 6930 3840 6964 4216
rect 7026 3840 7060 4216
rect 7122 3840 7156 4216
rect 7218 3840 7252 4216
rect 7314 3840 7348 4216
rect 4434 3222 4468 3598
rect 4530 3222 4564 3598
rect 4626 3222 4660 3598
rect 4722 3222 4756 3598
rect 4818 3222 4852 3598
rect 4914 3222 4948 3598
rect 5010 3222 5044 3598
rect 5106 3222 5140 3598
rect 5202 3222 5236 3598
rect 5298 3222 5332 3598
rect 5394 3222 5428 3598
rect 5490 3222 5524 3598
rect 5586 3222 5620 3598
rect 5682 3222 5716 3598
rect 5778 3222 5812 3598
rect 5874 3222 5908 3598
rect 5970 3222 6004 3598
rect 6066 3222 6100 3598
rect 6162 3222 6196 3598
rect 6258 3222 6292 3598
rect 6354 3222 6388 3598
rect 6450 3222 6484 3598
rect 6546 3222 6580 3598
rect 6642 3222 6676 3598
rect 6738 3222 6772 3598
rect 6834 3222 6868 3598
rect 6930 3222 6964 3598
rect 7026 3222 7060 3598
rect 7122 3222 7156 3598
rect 7218 3222 7252 3598
rect 7314 3222 7348 3598
rect 8074 5076 8108 5452
rect 8170 5076 8204 5452
rect 8266 5076 8300 5452
rect 8362 5076 8396 5452
rect 8458 5076 8492 5452
rect 8554 5076 8588 5452
rect 8650 5076 8684 5452
rect 8746 5076 8780 5452
rect 8842 5076 8876 5452
rect 8938 5076 8972 5452
rect 9034 5076 9068 5452
rect 9130 5076 9164 5452
rect 9226 5076 9260 5452
rect 9322 5076 9356 5452
rect 9418 5076 9452 5452
rect 9514 5076 9548 5452
rect 9610 5076 9644 5452
rect 9706 5076 9740 5452
rect 9802 5076 9836 5452
rect 9898 5076 9932 5452
rect 9994 5076 10028 5452
rect 10090 5076 10124 5452
rect 10186 5076 10220 5452
rect 10282 5076 10316 5452
rect 10378 5076 10412 5452
rect 10474 5076 10508 5452
rect 10570 5076 10604 5452
rect 10666 5076 10700 5452
rect 10762 5076 10796 5452
rect 10858 5076 10892 5452
rect 10954 5076 10988 5452
rect 8074 4458 8108 4834
rect 8170 4458 8204 4834
rect 8266 4458 8300 4834
rect 8362 4458 8396 4834
rect 8458 4458 8492 4834
rect 8554 4458 8588 4834
rect 8650 4458 8684 4834
rect 8746 4458 8780 4834
rect 8842 4458 8876 4834
rect 8938 4458 8972 4834
rect 9034 4458 9068 4834
rect 9130 4458 9164 4834
rect 9226 4458 9260 4834
rect 9322 4458 9356 4834
rect 9418 4458 9452 4834
rect 9514 4458 9548 4834
rect 9610 4458 9644 4834
rect 9706 4458 9740 4834
rect 9802 4458 9836 4834
rect 9898 4458 9932 4834
rect 9994 4458 10028 4834
rect 10090 4458 10124 4834
rect 10186 4458 10220 4834
rect 10282 4458 10316 4834
rect 10378 4458 10412 4834
rect 10474 4458 10508 4834
rect 10570 4458 10604 4834
rect 10666 4458 10700 4834
rect 10762 4458 10796 4834
rect 10858 4458 10892 4834
rect 10954 4458 10988 4834
rect 8074 3840 8108 4216
rect 8170 3840 8204 4216
rect 8266 3840 8300 4216
rect 8362 3840 8396 4216
rect 8458 3840 8492 4216
rect 8554 3840 8588 4216
rect 8650 3840 8684 4216
rect 8746 3840 8780 4216
rect 8842 3840 8876 4216
rect 8938 3840 8972 4216
rect 9034 3840 9068 4216
rect 9130 3840 9164 4216
rect 9226 3840 9260 4216
rect 9322 3840 9356 4216
rect 9418 3840 9452 4216
rect 9514 3840 9548 4216
rect 9610 3840 9644 4216
rect 9706 3840 9740 4216
rect 9802 3840 9836 4216
rect 9898 3840 9932 4216
rect 9994 3840 10028 4216
rect 10090 3840 10124 4216
rect 10186 3840 10220 4216
rect 10282 3840 10316 4216
rect 10378 3840 10412 4216
rect 10474 3840 10508 4216
rect 10570 3840 10604 4216
rect 10666 3840 10700 4216
rect 10762 3840 10796 4216
rect 10858 3840 10892 4216
rect 10954 3840 10988 4216
rect 8074 3222 8108 3598
rect 8170 3222 8204 3598
rect 8266 3222 8300 3598
rect 8362 3222 8396 3598
rect 8458 3222 8492 3598
rect 8554 3222 8588 3598
rect 8650 3222 8684 3598
rect 8746 3222 8780 3598
rect 8842 3222 8876 3598
rect 8938 3222 8972 3598
rect 9034 3222 9068 3598
rect 9130 3222 9164 3598
rect 9226 3222 9260 3598
rect 9322 3222 9356 3598
rect 9418 3222 9452 3598
rect 9514 3222 9548 3598
rect 9610 3222 9644 3598
rect 9706 3222 9740 3598
rect 9802 3222 9836 3598
rect 9898 3222 9932 3598
rect 9994 3222 10028 3598
rect 10090 3222 10124 3598
rect 10186 3222 10220 3598
rect 10282 3222 10316 3598
rect 10378 3222 10412 3598
rect 10474 3222 10508 3598
rect 10570 3222 10604 3598
rect 10666 3222 10700 3598
rect 10762 3222 10796 3598
rect 10858 3222 10892 3598
rect 10954 3222 10988 3598
rect 12054 5076 12088 5452
rect 12150 5076 12184 5452
rect 12246 5076 12280 5452
rect 12342 5076 12376 5452
rect 12438 5076 12472 5452
rect 12534 5076 12568 5452
rect 12630 5076 12664 5452
rect 12726 5076 12760 5452
rect 12822 5076 12856 5452
rect 12918 5076 12952 5452
rect 13014 5076 13048 5452
rect 13110 5076 13144 5452
rect 13206 5076 13240 5452
rect 13302 5076 13336 5452
rect 13398 5076 13432 5452
rect 13494 5076 13528 5452
rect 13590 5076 13624 5452
rect 13686 5076 13720 5452
rect 13782 5076 13816 5452
rect 13878 5076 13912 5452
rect 13974 5076 14008 5452
rect 14070 5076 14104 5452
rect 14166 5076 14200 5452
rect 14262 5076 14296 5452
rect 14358 5076 14392 5452
rect 14454 5076 14488 5452
rect 14550 5076 14584 5452
rect 14646 5076 14680 5452
rect 14742 5076 14776 5452
rect 14838 5076 14872 5452
rect 14934 5076 14968 5452
rect 12054 4458 12088 4834
rect 12150 4458 12184 4834
rect 12246 4458 12280 4834
rect 12342 4458 12376 4834
rect 12438 4458 12472 4834
rect 12534 4458 12568 4834
rect 12630 4458 12664 4834
rect 12726 4458 12760 4834
rect 12822 4458 12856 4834
rect 12918 4458 12952 4834
rect 13014 4458 13048 4834
rect 13110 4458 13144 4834
rect 13206 4458 13240 4834
rect 13302 4458 13336 4834
rect 13398 4458 13432 4834
rect 13494 4458 13528 4834
rect 13590 4458 13624 4834
rect 13686 4458 13720 4834
rect 13782 4458 13816 4834
rect 13878 4458 13912 4834
rect 13974 4458 14008 4834
rect 14070 4458 14104 4834
rect 14166 4458 14200 4834
rect 14262 4458 14296 4834
rect 14358 4458 14392 4834
rect 14454 4458 14488 4834
rect 14550 4458 14584 4834
rect 14646 4458 14680 4834
rect 14742 4458 14776 4834
rect 14838 4458 14872 4834
rect 14934 4458 14968 4834
rect 12054 3840 12088 4216
rect 12150 3840 12184 4216
rect 12246 3840 12280 4216
rect 12342 3840 12376 4216
rect 12438 3840 12472 4216
rect 12534 3840 12568 4216
rect 12630 3840 12664 4216
rect 12726 3840 12760 4216
rect 12822 3840 12856 4216
rect 12918 3840 12952 4216
rect 13014 3840 13048 4216
rect 13110 3840 13144 4216
rect 13206 3840 13240 4216
rect 13302 3840 13336 4216
rect 13398 3840 13432 4216
rect 13494 3840 13528 4216
rect 13590 3840 13624 4216
rect 13686 3840 13720 4216
rect 13782 3840 13816 4216
rect 13878 3840 13912 4216
rect 13974 3840 14008 4216
rect 14070 3840 14104 4216
rect 14166 3840 14200 4216
rect 14262 3840 14296 4216
rect 14358 3840 14392 4216
rect 14454 3840 14488 4216
rect 14550 3840 14584 4216
rect 14646 3840 14680 4216
rect 14742 3840 14776 4216
rect 14838 3840 14872 4216
rect 14934 3840 14968 4216
rect 12054 3222 12088 3598
rect 12150 3222 12184 3598
rect 12246 3222 12280 3598
rect 12342 3222 12376 3598
rect 12438 3222 12472 3598
rect 12534 3222 12568 3598
rect 12630 3222 12664 3598
rect 12726 3222 12760 3598
rect 12822 3222 12856 3598
rect 12918 3222 12952 3598
rect 13014 3222 13048 3598
rect 13110 3222 13144 3598
rect 13206 3222 13240 3598
rect 13302 3222 13336 3598
rect 13398 3222 13432 3598
rect 13494 3222 13528 3598
rect 13590 3222 13624 3598
rect 13686 3222 13720 3598
rect 13782 3222 13816 3598
rect 13878 3222 13912 3598
rect 13974 3222 14008 3598
rect 14070 3222 14104 3598
rect 14166 3222 14200 3598
rect 14262 3222 14296 3598
rect 14358 3222 14392 3598
rect 14454 3222 14488 3598
rect 14550 3222 14584 3598
rect 14646 3222 14680 3598
rect 14742 3222 14776 3598
rect 14838 3222 14872 3598
rect 14934 3222 14968 3598
rect 15694 5076 15728 5452
rect 15790 5076 15824 5452
rect 15886 5076 15920 5452
rect 15982 5076 16016 5452
rect 16078 5076 16112 5452
rect 16174 5076 16208 5452
rect 16270 5076 16304 5452
rect 16366 5076 16400 5452
rect 16462 5076 16496 5452
rect 16558 5076 16592 5452
rect 16654 5076 16688 5452
rect 16750 5076 16784 5452
rect 16846 5076 16880 5452
rect 16942 5076 16976 5452
rect 17038 5076 17072 5452
rect 17134 5076 17168 5452
rect 17230 5076 17264 5452
rect 17326 5076 17360 5452
rect 17422 5076 17456 5452
rect 17518 5076 17552 5452
rect 17614 5076 17648 5452
rect 17710 5076 17744 5452
rect 17806 5076 17840 5452
rect 17902 5076 17936 5452
rect 17998 5076 18032 5452
rect 18094 5076 18128 5452
rect 18190 5076 18224 5452
rect 18286 5076 18320 5452
rect 18382 5076 18416 5452
rect 18478 5076 18512 5452
rect 18574 5076 18608 5452
rect 15694 4458 15728 4834
rect 15790 4458 15824 4834
rect 15886 4458 15920 4834
rect 15982 4458 16016 4834
rect 16078 4458 16112 4834
rect 16174 4458 16208 4834
rect 16270 4458 16304 4834
rect 16366 4458 16400 4834
rect 16462 4458 16496 4834
rect 16558 4458 16592 4834
rect 16654 4458 16688 4834
rect 16750 4458 16784 4834
rect 16846 4458 16880 4834
rect 16942 4458 16976 4834
rect 17038 4458 17072 4834
rect 17134 4458 17168 4834
rect 17230 4458 17264 4834
rect 17326 4458 17360 4834
rect 17422 4458 17456 4834
rect 17518 4458 17552 4834
rect 17614 4458 17648 4834
rect 17710 4458 17744 4834
rect 17806 4458 17840 4834
rect 17902 4458 17936 4834
rect 17998 4458 18032 4834
rect 18094 4458 18128 4834
rect 18190 4458 18224 4834
rect 18286 4458 18320 4834
rect 18382 4458 18416 4834
rect 18478 4458 18512 4834
rect 18574 4458 18608 4834
rect 15694 3840 15728 4216
rect 15790 3840 15824 4216
rect 15886 3840 15920 4216
rect 15982 3840 16016 4216
rect 16078 3840 16112 4216
rect 16174 3840 16208 4216
rect 16270 3840 16304 4216
rect 16366 3840 16400 4216
rect 16462 3840 16496 4216
rect 16558 3840 16592 4216
rect 16654 3840 16688 4216
rect 16750 3840 16784 4216
rect 16846 3840 16880 4216
rect 16942 3840 16976 4216
rect 17038 3840 17072 4216
rect 17134 3840 17168 4216
rect 17230 3840 17264 4216
rect 17326 3840 17360 4216
rect 17422 3840 17456 4216
rect 17518 3840 17552 4216
rect 17614 3840 17648 4216
rect 17710 3840 17744 4216
rect 17806 3840 17840 4216
rect 17902 3840 17936 4216
rect 17998 3840 18032 4216
rect 18094 3840 18128 4216
rect 18190 3840 18224 4216
rect 18286 3840 18320 4216
rect 18382 3840 18416 4216
rect 18478 3840 18512 4216
rect 18574 3840 18608 4216
rect 15694 3222 15728 3598
rect 15790 3222 15824 3598
rect 15886 3222 15920 3598
rect 15982 3222 16016 3598
rect 16078 3222 16112 3598
rect 16174 3222 16208 3598
rect 16270 3222 16304 3598
rect 16366 3222 16400 3598
rect 16462 3222 16496 3598
rect 16558 3222 16592 3598
rect 16654 3222 16688 3598
rect 16750 3222 16784 3598
rect 16846 3222 16880 3598
rect 16942 3222 16976 3598
rect 17038 3222 17072 3598
rect 17134 3222 17168 3598
rect 17230 3222 17264 3598
rect 17326 3222 17360 3598
rect 17422 3222 17456 3598
rect 17518 3222 17552 3598
rect 17614 3222 17648 3598
rect 17710 3222 17744 3598
rect 17806 3222 17840 3598
rect 17902 3222 17936 3598
rect 17998 3222 18032 3598
rect 18094 3222 18128 3598
rect 18190 3222 18224 3598
rect 18286 3222 18320 3598
rect 18382 3222 18416 3598
rect 18478 3222 18512 3598
rect 18574 3222 18608 3598
rect -1570 2244 -1536 2620
rect -1474 2244 -1440 2620
rect -1378 2244 -1344 2620
rect -1282 2244 -1248 2620
rect -1186 2244 -1152 2620
rect -1090 2244 -1056 2620
rect -994 2244 -960 2620
rect -1570 1626 -1536 2002
rect -1474 1626 -1440 2002
rect -1378 1626 -1344 2002
rect -1282 1626 -1248 2002
rect -1186 1626 -1152 2002
rect -1090 1626 -1056 2002
rect -994 1626 -960 2002
rect -530 2244 -496 2620
rect -434 2244 -400 2620
rect -338 2244 -304 2620
rect -242 2244 -208 2620
rect -146 2244 -112 2620
rect -50 2244 -16 2620
rect 46 2244 80 2620
rect -530 1626 -496 2002
rect -434 1626 -400 2002
rect -338 1626 -304 2002
rect -242 1626 -208 2002
rect -146 1626 -112 2002
rect -50 1626 -16 2002
rect 46 1626 80 2002
rect 510 2244 544 2620
rect 606 2244 640 2620
rect 702 2244 736 2620
rect 798 2244 832 2620
rect 894 2244 928 2620
rect 990 2244 1024 2620
rect 1086 2244 1120 2620
rect 510 1626 544 2002
rect 606 1626 640 2002
rect 702 1626 736 2002
rect 798 1626 832 2002
rect 894 1626 928 2002
rect 990 1626 1024 2002
rect 1086 1626 1120 2002
rect 1550 2244 1584 2620
rect 1646 2244 1680 2620
rect 1742 2244 1776 2620
rect 1838 2244 1872 2620
rect 1934 2244 1968 2620
rect 2030 2244 2064 2620
rect 2126 2244 2160 2620
rect 1550 1626 1584 2002
rect 1646 1626 1680 2002
rect 1742 1626 1776 2002
rect 1838 1626 1872 2002
rect 1934 1626 1968 2002
rect 2030 1626 2064 2002
rect 2126 1626 2160 2002
rect 2590 2244 2624 2620
rect 2686 2244 2720 2620
rect 2782 2244 2816 2620
rect 2878 2244 2912 2620
rect 2974 2244 3008 2620
rect 3070 2244 3104 2620
rect 3166 2244 3200 2620
rect 2590 1626 2624 2002
rect 2686 1626 2720 2002
rect 2782 1626 2816 2002
rect 2878 1626 2912 2002
rect 2974 1626 3008 2002
rect 3070 1626 3104 2002
rect 3166 1626 3200 2002
rect 4234 2404 4268 2780
rect 4330 2404 4364 2780
rect 4426 2404 4460 2780
rect 4522 2404 4556 2780
rect 4618 2404 4652 2780
rect 4714 2404 4748 2780
rect 4810 2404 4844 2780
rect 4234 1786 4268 2162
rect 4330 1786 4364 2162
rect 4426 1786 4460 2162
rect 4522 1786 4556 2162
rect 4618 1786 4652 2162
rect 4714 1786 4748 2162
rect 4810 1786 4844 2162
rect 5274 2404 5308 2780
rect 5370 2404 5404 2780
rect 5466 2404 5500 2780
rect 5562 2404 5596 2780
rect 5658 2404 5692 2780
rect 5754 2404 5788 2780
rect 5850 2404 5884 2780
rect 5274 1786 5308 2162
rect 5370 1786 5404 2162
rect 5466 1786 5500 2162
rect 5562 1786 5596 2162
rect 5658 1786 5692 2162
rect 5754 1786 5788 2162
rect 5850 1786 5884 2162
rect 6314 2404 6348 2780
rect 6410 2404 6444 2780
rect 6506 2404 6540 2780
rect 6602 2404 6636 2780
rect 6698 2404 6732 2780
rect 6794 2404 6828 2780
rect 6890 2404 6924 2780
rect 6314 1786 6348 2162
rect 6410 1786 6444 2162
rect 6506 1786 6540 2162
rect 6602 1786 6636 2162
rect 6698 1786 6732 2162
rect 6794 1786 6828 2162
rect 6890 1786 6924 2162
rect 7354 2404 7388 2780
rect 7450 2404 7484 2780
rect 7546 2404 7580 2780
rect 7642 2404 7676 2780
rect 7738 2404 7772 2780
rect 7834 2404 7868 2780
rect 7930 2404 7964 2780
rect 7354 1786 7388 2162
rect 7450 1786 7484 2162
rect 7546 1786 7580 2162
rect 7642 1786 7676 2162
rect 7738 1786 7772 2162
rect 7834 1786 7868 2162
rect 7930 1786 7964 2162
rect 8394 2404 8428 2780
rect 8490 2404 8524 2780
rect 8586 2404 8620 2780
rect 8682 2404 8716 2780
rect 8778 2404 8812 2780
rect 8874 2404 8908 2780
rect 8970 2404 9004 2780
rect 8394 1786 8428 2162
rect 8490 1786 8524 2162
rect 8586 1786 8620 2162
rect 8682 1786 8716 2162
rect 8778 1786 8812 2162
rect 8874 1786 8908 2162
rect 8970 1786 9004 2162
rect 9434 2404 9468 2780
rect 9530 2404 9564 2780
rect 9626 2404 9660 2780
rect 9722 2404 9756 2780
rect 9818 2404 9852 2780
rect 9914 2404 9948 2780
rect 10010 2404 10044 2780
rect 9434 1786 9468 2162
rect 9530 1786 9564 2162
rect 9626 1786 9660 2162
rect 9722 1786 9756 2162
rect 9818 1786 9852 2162
rect 9914 1786 9948 2162
rect 10010 1786 10044 2162
rect 10474 2404 10508 2780
rect 10570 2404 10604 2780
rect 10666 2404 10700 2780
rect 10762 2404 10796 2780
rect 10858 2404 10892 2780
rect 10954 2404 10988 2780
rect 11050 2404 11084 2780
rect 10474 1786 10508 2162
rect 10570 1786 10604 2162
rect 10666 1786 10700 2162
rect 10762 1786 10796 2162
rect 10858 1786 10892 2162
rect 10954 1786 10988 2162
rect 11050 1786 11084 2162
rect 11854 2404 11888 2780
rect 11950 2404 11984 2780
rect 12046 2404 12080 2780
rect 12142 2404 12176 2780
rect 12238 2404 12272 2780
rect 12334 2404 12368 2780
rect 12430 2404 12464 2780
rect 11854 1786 11888 2162
rect 11950 1786 11984 2162
rect 12046 1786 12080 2162
rect 12142 1786 12176 2162
rect 12238 1786 12272 2162
rect 12334 1786 12368 2162
rect 12430 1786 12464 2162
rect 12894 2404 12928 2780
rect 12990 2404 13024 2780
rect 13086 2404 13120 2780
rect 13182 2404 13216 2780
rect 13278 2404 13312 2780
rect 13374 2404 13408 2780
rect 13470 2404 13504 2780
rect 12894 1786 12928 2162
rect 12990 1786 13024 2162
rect 13086 1786 13120 2162
rect 13182 1786 13216 2162
rect 13278 1786 13312 2162
rect 13374 1786 13408 2162
rect 13470 1786 13504 2162
rect 13934 2404 13968 2780
rect 14030 2404 14064 2780
rect 14126 2404 14160 2780
rect 14222 2404 14256 2780
rect 14318 2404 14352 2780
rect 14414 2404 14448 2780
rect 14510 2404 14544 2780
rect 13934 1786 13968 2162
rect 14030 1786 14064 2162
rect 14126 1786 14160 2162
rect 14222 1786 14256 2162
rect 14318 1786 14352 2162
rect 14414 1786 14448 2162
rect 14510 1786 14544 2162
rect 14974 2404 15008 2780
rect 15070 2404 15104 2780
rect 15166 2404 15200 2780
rect 15262 2404 15296 2780
rect 15358 2404 15392 2780
rect 15454 2404 15488 2780
rect 15550 2404 15584 2780
rect 14974 1786 15008 2162
rect 15070 1786 15104 2162
rect 15166 1786 15200 2162
rect 15262 1786 15296 2162
rect 15358 1786 15392 2162
rect 15454 1786 15488 2162
rect 15550 1786 15584 2162
rect 16014 2404 16048 2780
rect 16110 2404 16144 2780
rect 16206 2404 16240 2780
rect 16302 2404 16336 2780
rect 16398 2404 16432 2780
rect 16494 2404 16528 2780
rect 16590 2404 16624 2780
rect 16014 1786 16048 2162
rect 16110 1786 16144 2162
rect 16206 1786 16240 2162
rect 16302 1786 16336 2162
rect 16398 1786 16432 2162
rect 16494 1786 16528 2162
rect 16590 1786 16624 2162
rect 17054 2404 17088 2780
rect 17150 2404 17184 2780
rect 17246 2404 17280 2780
rect 17342 2404 17376 2780
rect 17438 2404 17472 2780
rect 17534 2404 17568 2780
rect 17630 2404 17664 2780
rect 17054 1786 17088 2162
rect 17150 1786 17184 2162
rect 17246 1786 17280 2162
rect 17342 1786 17376 2162
rect 17438 1786 17472 2162
rect 17534 1786 17568 2162
rect 17630 1786 17664 2162
rect 18094 2404 18128 2780
rect 18190 2404 18224 2780
rect 18286 2404 18320 2780
rect 18382 2404 18416 2780
rect 18478 2404 18512 2780
rect 18574 2404 18608 2780
rect 18670 2404 18704 2780
rect 18094 1786 18128 2162
rect 18190 1786 18224 2162
rect 18286 1786 18320 2162
rect 18382 1786 18416 2162
rect 18478 1786 18512 2162
rect 18574 1786 18608 2162
rect 18670 1786 18704 2162
rect -1570 822 -1536 1198
rect -1452 822 -1418 1198
rect -1334 822 -1300 1198
rect -1216 822 -1182 1198
rect -1098 822 -1064 1198
rect -980 822 -946 1198
rect -862 822 -828 1198
rect -530 822 -496 1198
rect -412 822 -378 1198
rect -294 822 -260 1198
rect -176 822 -142 1198
rect -58 822 -24 1198
rect 60 822 94 1198
rect 178 822 212 1198
rect 510 822 544 1198
rect 628 822 662 1198
rect 746 822 780 1198
rect 864 822 898 1198
rect 982 822 1016 1198
rect 1100 822 1134 1198
rect 1218 822 1252 1198
rect 1550 822 1584 1198
rect 1668 822 1702 1198
rect 1786 822 1820 1198
rect 1904 822 1938 1198
rect 2022 822 2056 1198
rect 2140 822 2174 1198
rect 2258 822 2292 1198
rect 2590 822 2624 1198
rect 2708 822 2742 1198
rect 2826 822 2860 1198
rect 2944 822 2978 1198
rect 3062 822 3096 1198
rect 3180 822 3214 1198
rect 3298 822 3332 1198
rect 4234 982 4268 1358
rect 4352 982 4386 1358
rect 4470 982 4504 1358
rect 4588 982 4622 1358
rect 4706 982 4740 1358
rect 4824 982 4858 1358
rect 4942 982 4976 1358
rect 5274 982 5308 1358
rect 5392 982 5426 1358
rect 5510 982 5544 1358
rect 5628 982 5662 1358
rect 5746 982 5780 1358
rect 5864 982 5898 1358
rect 5982 982 6016 1358
rect 6314 982 6348 1358
rect 6432 982 6466 1358
rect 6550 982 6584 1358
rect 6668 982 6702 1358
rect 6786 982 6820 1358
rect 6904 982 6938 1358
rect 7022 982 7056 1358
rect 7354 982 7388 1358
rect 7472 982 7506 1358
rect 7590 982 7624 1358
rect 7708 982 7742 1358
rect 7826 982 7860 1358
rect 7944 982 7978 1358
rect 8062 982 8096 1358
rect 8394 982 8428 1358
rect 8512 982 8546 1358
rect 8630 982 8664 1358
rect 8748 982 8782 1358
rect 8866 982 8900 1358
rect 8984 982 9018 1358
rect 9102 982 9136 1358
rect 9434 982 9468 1358
rect 9552 982 9586 1358
rect 9670 982 9704 1358
rect 9788 982 9822 1358
rect 9906 982 9940 1358
rect 10024 982 10058 1358
rect 10142 982 10176 1358
rect 10474 982 10508 1358
rect 10592 982 10626 1358
rect 10710 982 10744 1358
rect 10828 982 10862 1358
rect 10946 982 10980 1358
rect 11064 982 11098 1358
rect 11182 982 11216 1358
rect 11854 982 11888 1358
rect 11972 982 12006 1358
rect 12090 982 12124 1358
rect 12208 982 12242 1358
rect 12326 982 12360 1358
rect 12444 982 12478 1358
rect 12562 982 12596 1358
rect 12894 982 12928 1358
rect 13012 982 13046 1358
rect 13130 982 13164 1358
rect 13248 982 13282 1358
rect 13366 982 13400 1358
rect 13484 982 13518 1358
rect 13602 982 13636 1358
rect 13934 982 13968 1358
rect 14052 982 14086 1358
rect 14170 982 14204 1358
rect 14288 982 14322 1358
rect 14406 982 14440 1358
rect 14524 982 14558 1358
rect 14642 982 14676 1358
rect 14974 982 15008 1358
rect 15092 982 15126 1358
rect 15210 982 15244 1358
rect 15328 982 15362 1358
rect 15446 982 15480 1358
rect 15564 982 15598 1358
rect 15682 982 15716 1358
rect 16014 982 16048 1358
rect 16132 982 16166 1358
rect 16250 982 16284 1358
rect 16368 982 16402 1358
rect 16486 982 16520 1358
rect 16604 982 16638 1358
rect 16722 982 16756 1358
rect 17054 982 17088 1358
rect 17172 982 17206 1358
rect 17290 982 17324 1358
rect 17408 982 17442 1358
rect 17526 982 17560 1358
rect 17644 982 17678 1358
rect 17762 982 17796 1358
rect 18094 982 18128 1358
rect 18212 982 18246 1358
rect 18330 982 18364 1358
rect 18448 982 18482 1358
rect 18566 982 18600 1358
rect 18684 982 18718 1358
rect 18802 982 18836 1358
rect -7400 -442 -7366 -66
rect -7304 -442 -7270 -66
rect -7208 -442 -7174 -66
rect -7112 -442 -7078 -66
rect -7016 -442 -6982 -66
rect -6920 -442 -6886 -66
rect -6824 -442 -6790 -66
rect -6728 -442 -6694 -66
rect -6632 -442 -6598 -66
rect -6536 -442 -6502 -66
rect -6440 -442 -6406 -66
rect -7400 -1060 -7366 -684
rect -7304 -1060 -7270 -684
rect -7208 -1060 -7174 -684
rect -7112 -1060 -7078 -684
rect -7016 -1060 -6982 -684
rect -6920 -1060 -6886 -684
rect -6824 -1060 -6790 -684
rect -6728 -1060 -6694 -684
rect -6632 -1060 -6598 -684
rect -6536 -1060 -6502 -684
rect -6440 -1060 -6406 -684
rect -7400 -2278 -7366 -1902
rect -7304 -2278 -7270 -1902
rect -7208 -2278 -7174 -1902
rect -7112 -2278 -7078 -1902
rect -7016 -2278 -6982 -1902
rect -6920 -2278 -6886 -1902
rect -6824 -2278 -6790 -1902
rect -7400 -2896 -7366 -2520
rect -7304 -2896 -7270 -2520
rect -7208 -2896 -7174 -2520
rect -7112 -2896 -7078 -2520
rect -7016 -2896 -6982 -2520
rect -6920 -2896 -6886 -2520
rect -6824 -2896 -6790 -2520
rect -5988 -42 -5812 -8
rect -5988 -1700 -5812 -1666
rect 4234 164 4268 540
rect 4330 164 4364 540
rect 4426 164 4460 540
rect 4522 164 4556 540
rect 4618 164 4652 540
rect 4714 164 4748 540
rect 4810 164 4844 540
rect 4234 -454 4268 -78
rect 4330 -454 4364 -78
rect 4426 -454 4460 -78
rect 4522 -454 4556 -78
rect 4618 -454 4652 -78
rect 4714 -454 4748 -78
rect 4810 -454 4844 -78
rect 5274 164 5308 540
rect 5370 164 5404 540
rect 5466 164 5500 540
rect 5562 164 5596 540
rect 5658 164 5692 540
rect 5754 164 5788 540
rect 5850 164 5884 540
rect 5274 -454 5308 -78
rect 5370 -454 5404 -78
rect 5466 -454 5500 -78
rect 5562 -454 5596 -78
rect 5658 -454 5692 -78
rect 5754 -454 5788 -78
rect 5850 -454 5884 -78
rect 6314 164 6348 540
rect 6410 164 6444 540
rect 6506 164 6540 540
rect 6602 164 6636 540
rect 6698 164 6732 540
rect 6794 164 6828 540
rect 6890 164 6924 540
rect 6314 -454 6348 -78
rect 6410 -454 6444 -78
rect 6506 -454 6540 -78
rect 6602 -454 6636 -78
rect 6698 -454 6732 -78
rect 6794 -454 6828 -78
rect 6890 -454 6924 -78
rect 7354 164 7388 540
rect 7450 164 7484 540
rect 7546 164 7580 540
rect 7642 164 7676 540
rect 7738 164 7772 540
rect 7834 164 7868 540
rect 7930 164 7964 540
rect 7354 -454 7388 -78
rect 7450 -454 7484 -78
rect 7546 -454 7580 -78
rect 7642 -454 7676 -78
rect 7738 -454 7772 -78
rect 7834 -454 7868 -78
rect 7930 -454 7964 -78
rect 8394 164 8428 540
rect 8490 164 8524 540
rect 8586 164 8620 540
rect 8682 164 8716 540
rect 8778 164 8812 540
rect 8874 164 8908 540
rect 8970 164 9004 540
rect 8394 -454 8428 -78
rect 8490 -454 8524 -78
rect 8586 -454 8620 -78
rect 8682 -454 8716 -78
rect 8778 -454 8812 -78
rect 8874 -454 8908 -78
rect 8970 -454 9004 -78
rect 9434 164 9468 540
rect 9530 164 9564 540
rect 9626 164 9660 540
rect 9722 164 9756 540
rect 9818 164 9852 540
rect 9914 164 9948 540
rect 10010 164 10044 540
rect 9434 -454 9468 -78
rect 9530 -454 9564 -78
rect 9626 -454 9660 -78
rect 9722 -454 9756 -78
rect 9818 -454 9852 -78
rect 9914 -454 9948 -78
rect 10010 -454 10044 -78
rect 10474 164 10508 540
rect 10570 164 10604 540
rect 10666 164 10700 540
rect 10762 164 10796 540
rect 10858 164 10892 540
rect 10954 164 10988 540
rect 11050 164 11084 540
rect 10474 -454 10508 -78
rect 10570 -454 10604 -78
rect 10666 -454 10700 -78
rect 10762 -454 10796 -78
rect 10858 -454 10892 -78
rect 10954 -454 10988 -78
rect 11050 -454 11084 -78
rect 11854 164 11888 540
rect 11950 164 11984 540
rect 12046 164 12080 540
rect 12142 164 12176 540
rect 12238 164 12272 540
rect 12334 164 12368 540
rect 12430 164 12464 540
rect 11854 -454 11888 -78
rect 11950 -454 11984 -78
rect 12046 -454 12080 -78
rect 12142 -454 12176 -78
rect 12238 -454 12272 -78
rect 12334 -454 12368 -78
rect 12430 -454 12464 -78
rect 12894 164 12928 540
rect 12990 164 13024 540
rect 13086 164 13120 540
rect 13182 164 13216 540
rect 13278 164 13312 540
rect 13374 164 13408 540
rect 13470 164 13504 540
rect 12894 -454 12928 -78
rect 12990 -454 13024 -78
rect 13086 -454 13120 -78
rect 13182 -454 13216 -78
rect 13278 -454 13312 -78
rect 13374 -454 13408 -78
rect 13470 -454 13504 -78
rect 13934 164 13968 540
rect 14030 164 14064 540
rect 14126 164 14160 540
rect 14222 164 14256 540
rect 14318 164 14352 540
rect 14414 164 14448 540
rect 14510 164 14544 540
rect 13934 -454 13968 -78
rect 14030 -454 14064 -78
rect 14126 -454 14160 -78
rect 14222 -454 14256 -78
rect 14318 -454 14352 -78
rect 14414 -454 14448 -78
rect 14510 -454 14544 -78
rect 14974 164 15008 540
rect 15070 164 15104 540
rect 15166 164 15200 540
rect 15262 164 15296 540
rect 15358 164 15392 540
rect 15454 164 15488 540
rect 15550 164 15584 540
rect 14974 -454 15008 -78
rect 15070 -454 15104 -78
rect 15166 -454 15200 -78
rect 15262 -454 15296 -78
rect 15358 -454 15392 -78
rect 15454 -454 15488 -78
rect 15550 -454 15584 -78
rect 16014 164 16048 540
rect 16110 164 16144 540
rect 16206 164 16240 540
rect 16302 164 16336 540
rect 16398 164 16432 540
rect 16494 164 16528 540
rect 16590 164 16624 540
rect 16014 -454 16048 -78
rect 16110 -454 16144 -78
rect 16206 -454 16240 -78
rect 16302 -454 16336 -78
rect 16398 -454 16432 -78
rect 16494 -454 16528 -78
rect 16590 -454 16624 -78
rect 17054 164 17088 540
rect 17150 164 17184 540
rect 17246 164 17280 540
rect 17342 164 17376 540
rect 17438 164 17472 540
rect 17534 164 17568 540
rect 17630 164 17664 540
rect 17054 -454 17088 -78
rect 17150 -454 17184 -78
rect 17246 -454 17280 -78
rect 17342 -454 17376 -78
rect 17438 -454 17472 -78
rect 17534 -454 17568 -78
rect 17630 -454 17664 -78
rect 18094 164 18128 540
rect 18190 164 18224 540
rect 18286 164 18320 540
rect 18382 164 18416 540
rect 18478 164 18512 540
rect 18574 164 18608 540
rect 18670 164 18704 540
rect 18094 -454 18128 -78
rect 18190 -454 18224 -78
rect 18286 -454 18320 -78
rect 18382 -454 18416 -78
rect 18478 -454 18512 -78
rect 18574 -454 18608 -78
rect 18670 -454 18704 -78
rect 4234 -1258 4268 -882
rect 4352 -1258 4386 -882
rect 4470 -1258 4504 -882
rect 4588 -1258 4622 -882
rect 4706 -1258 4740 -882
rect 4824 -1258 4858 -882
rect 4942 -1258 4976 -882
rect 5274 -1258 5308 -882
rect 5392 -1258 5426 -882
rect 5510 -1258 5544 -882
rect 5628 -1258 5662 -882
rect 5746 -1258 5780 -882
rect 5864 -1258 5898 -882
rect 5982 -1258 6016 -882
rect 6314 -1258 6348 -882
rect 6432 -1258 6466 -882
rect 6550 -1258 6584 -882
rect 6668 -1258 6702 -882
rect 6786 -1258 6820 -882
rect 6904 -1258 6938 -882
rect 7022 -1258 7056 -882
rect 7354 -1258 7388 -882
rect 7472 -1258 7506 -882
rect 7590 -1258 7624 -882
rect 7708 -1258 7742 -882
rect 7826 -1258 7860 -882
rect 7944 -1258 7978 -882
rect 8062 -1258 8096 -882
rect 8394 -1258 8428 -882
rect 8512 -1258 8546 -882
rect 8630 -1258 8664 -882
rect 8748 -1258 8782 -882
rect 8866 -1258 8900 -882
rect 8984 -1258 9018 -882
rect 9102 -1258 9136 -882
rect 9434 -1258 9468 -882
rect 9552 -1258 9586 -882
rect 9670 -1258 9704 -882
rect 9788 -1258 9822 -882
rect 9906 -1258 9940 -882
rect 10024 -1258 10058 -882
rect 10142 -1258 10176 -882
rect 10474 -1258 10508 -882
rect 10592 -1258 10626 -882
rect 10710 -1258 10744 -882
rect 10828 -1258 10862 -882
rect 10946 -1258 10980 -882
rect 11064 -1258 11098 -882
rect 11182 -1258 11216 -882
rect 11854 -1258 11888 -882
rect 11972 -1258 12006 -882
rect 12090 -1258 12124 -882
rect 12208 -1258 12242 -882
rect 12326 -1258 12360 -882
rect 12444 -1258 12478 -882
rect 12562 -1258 12596 -882
rect 12894 -1258 12928 -882
rect 13012 -1258 13046 -882
rect 13130 -1258 13164 -882
rect 13248 -1258 13282 -882
rect 13366 -1258 13400 -882
rect 13484 -1258 13518 -882
rect 13602 -1258 13636 -882
rect 13934 -1258 13968 -882
rect 14052 -1258 14086 -882
rect 14170 -1258 14204 -882
rect 14288 -1258 14322 -882
rect 14406 -1258 14440 -882
rect 14524 -1258 14558 -882
rect 14642 -1258 14676 -882
rect 14974 -1258 15008 -882
rect 15092 -1258 15126 -882
rect 15210 -1258 15244 -882
rect 15328 -1258 15362 -882
rect 15446 -1258 15480 -882
rect 15564 -1258 15598 -882
rect 15682 -1258 15716 -882
rect 16014 -1258 16048 -882
rect 16132 -1258 16166 -882
rect 16250 -1258 16284 -882
rect 16368 -1258 16402 -882
rect 16486 -1258 16520 -882
rect 16604 -1258 16638 -882
rect 16722 -1258 16756 -882
rect 17054 -1258 17088 -882
rect 17172 -1258 17206 -882
rect 17290 -1258 17324 -882
rect 17408 -1258 17442 -882
rect 17526 -1258 17560 -882
rect 17644 -1258 17678 -882
rect 17762 -1258 17796 -882
rect 18094 -1258 18128 -882
rect 18212 -1258 18246 -882
rect 18330 -1258 18364 -882
rect 18448 -1258 18482 -882
rect 18566 -1258 18600 -882
rect 18684 -1258 18718 -882
rect 18802 -1258 18836 -882
rect 4234 -2076 4268 -1700
rect 4330 -2076 4364 -1700
rect 4426 -2076 4460 -1700
rect 4522 -2076 4556 -1700
rect 4618 -2076 4652 -1700
rect 4714 -2076 4748 -1700
rect 4810 -2076 4844 -1700
rect 4234 -2694 4268 -2318
rect 4330 -2694 4364 -2318
rect 4426 -2694 4460 -2318
rect 4522 -2694 4556 -2318
rect 4618 -2694 4652 -2318
rect 4714 -2694 4748 -2318
rect 4810 -2694 4844 -2318
rect 5274 -2076 5308 -1700
rect 5370 -2076 5404 -1700
rect 5466 -2076 5500 -1700
rect 5562 -2076 5596 -1700
rect 5658 -2076 5692 -1700
rect 5754 -2076 5788 -1700
rect 5850 -2076 5884 -1700
rect 5274 -2694 5308 -2318
rect 5370 -2694 5404 -2318
rect 5466 -2694 5500 -2318
rect 5562 -2694 5596 -2318
rect 5658 -2694 5692 -2318
rect 5754 -2694 5788 -2318
rect 5850 -2694 5884 -2318
rect 6314 -2076 6348 -1700
rect 6410 -2076 6444 -1700
rect 6506 -2076 6540 -1700
rect 6602 -2076 6636 -1700
rect 6698 -2076 6732 -1700
rect 6794 -2076 6828 -1700
rect 6890 -2076 6924 -1700
rect 6314 -2694 6348 -2318
rect 6410 -2694 6444 -2318
rect 6506 -2694 6540 -2318
rect 6602 -2694 6636 -2318
rect 6698 -2694 6732 -2318
rect 6794 -2694 6828 -2318
rect 6890 -2694 6924 -2318
rect 7354 -2076 7388 -1700
rect 7450 -2076 7484 -1700
rect 7546 -2076 7580 -1700
rect 7642 -2076 7676 -1700
rect 7738 -2076 7772 -1700
rect 7834 -2076 7868 -1700
rect 7930 -2076 7964 -1700
rect 7354 -2694 7388 -2318
rect 7450 -2694 7484 -2318
rect 7546 -2694 7580 -2318
rect 7642 -2694 7676 -2318
rect 7738 -2694 7772 -2318
rect 7834 -2694 7868 -2318
rect 7930 -2694 7964 -2318
rect 8394 -2076 8428 -1700
rect 8490 -2076 8524 -1700
rect 8586 -2076 8620 -1700
rect 8682 -2076 8716 -1700
rect 8778 -2076 8812 -1700
rect 8874 -2076 8908 -1700
rect 8970 -2076 9004 -1700
rect 8394 -2694 8428 -2318
rect 8490 -2694 8524 -2318
rect 8586 -2694 8620 -2318
rect 8682 -2694 8716 -2318
rect 8778 -2694 8812 -2318
rect 8874 -2694 8908 -2318
rect 8970 -2694 9004 -2318
rect 11854 -2076 11888 -1700
rect 11950 -2076 11984 -1700
rect 12046 -2076 12080 -1700
rect 12142 -2076 12176 -1700
rect 12238 -2076 12272 -1700
rect 12334 -2076 12368 -1700
rect 12430 -2076 12464 -1700
rect 11854 -2694 11888 -2318
rect 11950 -2694 11984 -2318
rect 12046 -2694 12080 -2318
rect 12142 -2694 12176 -2318
rect 12238 -2694 12272 -2318
rect 12334 -2694 12368 -2318
rect 12430 -2694 12464 -2318
rect 12894 -2076 12928 -1700
rect 12990 -2076 13024 -1700
rect 13086 -2076 13120 -1700
rect 13182 -2076 13216 -1700
rect 13278 -2076 13312 -1700
rect 13374 -2076 13408 -1700
rect 13470 -2076 13504 -1700
rect 12894 -2694 12928 -2318
rect 12990 -2694 13024 -2318
rect 13086 -2694 13120 -2318
rect 13182 -2694 13216 -2318
rect 13278 -2694 13312 -2318
rect 13374 -2694 13408 -2318
rect 13470 -2694 13504 -2318
rect 13934 -2076 13968 -1700
rect 14030 -2076 14064 -1700
rect 14126 -2076 14160 -1700
rect 14222 -2076 14256 -1700
rect 14318 -2076 14352 -1700
rect 14414 -2076 14448 -1700
rect 14510 -2076 14544 -1700
rect 13934 -2694 13968 -2318
rect 14030 -2694 14064 -2318
rect 14126 -2694 14160 -2318
rect 14222 -2694 14256 -2318
rect 14318 -2694 14352 -2318
rect 14414 -2694 14448 -2318
rect 14510 -2694 14544 -2318
rect 14974 -2076 15008 -1700
rect 15070 -2076 15104 -1700
rect 15166 -2076 15200 -1700
rect 15262 -2076 15296 -1700
rect 15358 -2076 15392 -1700
rect 15454 -2076 15488 -1700
rect 15550 -2076 15584 -1700
rect 14974 -2694 15008 -2318
rect 15070 -2694 15104 -2318
rect 15166 -2694 15200 -2318
rect 15262 -2694 15296 -2318
rect 15358 -2694 15392 -2318
rect 15454 -2694 15488 -2318
rect 15550 -2694 15584 -2318
rect 16014 -2076 16048 -1700
rect 16110 -2076 16144 -1700
rect 16206 -2076 16240 -1700
rect 16302 -2076 16336 -1700
rect 16398 -2076 16432 -1700
rect 16494 -2076 16528 -1700
rect 16590 -2076 16624 -1700
rect 16014 -2694 16048 -2318
rect 16110 -2694 16144 -2318
rect 16206 -2694 16240 -2318
rect 16302 -2694 16336 -2318
rect 16398 -2694 16432 -2318
rect 16494 -2694 16528 -2318
rect 16590 -2694 16624 -2318
rect -7400 -3700 -7366 -3324
rect -7282 -3700 -7248 -3324
rect -7164 -3700 -7130 -3324
rect -7046 -3700 -7012 -3324
rect -6928 -3700 -6894 -3324
rect -6810 -3700 -6776 -3324
rect -6692 -3700 -6658 -3324
rect 4234 -3498 4268 -3122
rect 4352 -3498 4386 -3122
rect 4470 -3498 4504 -3122
rect 4588 -3498 4622 -3122
rect 4706 -3498 4740 -3122
rect 4824 -3498 4858 -3122
rect 4942 -3498 4976 -3122
rect 5274 -3498 5308 -3122
rect 5392 -3498 5426 -3122
rect 5510 -3498 5544 -3122
rect 5628 -3498 5662 -3122
rect 5746 -3498 5780 -3122
rect 5864 -3498 5898 -3122
rect 5982 -3498 6016 -3122
rect 6314 -3498 6348 -3122
rect 6432 -3498 6466 -3122
rect 6550 -3498 6584 -3122
rect 6668 -3498 6702 -3122
rect 6786 -3498 6820 -3122
rect 6904 -3498 6938 -3122
rect 7022 -3498 7056 -3122
rect 7354 -3498 7388 -3122
rect 7472 -3498 7506 -3122
rect 7590 -3498 7624 -3122
rect 7708 -3498 7742 -3122
rect 7826 -3498 7860 -3122
rect 7944 -3498 7978 -3122
rect 8062 -3498 8096 -3122
rect 8394 -3498 8428 -3122
rect 8512 -3498 8546 -3122
rect 8630 -3498 8664 -3122
rect 8748 -3498 8782 -3122
rect 8866 -3498 8900 -3122
rect 8984 -3498 9018 -3122
rect 9102 -3498 9136 -3122
rect 11854 -3498 11888 -3122
rect 11972 -3498 12006 -3122
rect 12090 -3498 12124 -3122
rect 12208 -3498 12242 -3122
rect 12326 -3498 12360 -3122
rect 12444 -3498 12478 -3122
rect 12562 -3498 12596 -3122
rect 12894 -3498 12928 -3122
rect 13012 -3498 13046 -3122
rect 13130 -3498 13164 -3122
rect 13248 -3498 13282 -3122
rect 13366 -3498 13400 -3122
rect 13484 -3498 13518 -3122
rect 13602 -3498 13636 -3122
rect 13934 -3498 13968 -3122
rect 14052 -3498 14086 -3122
rect 14170 -3498 14204 -3122
rect 14288 -3498 14322 -3122
rect 14406 -3498 14440 -3122
rect 14524 -3498 14558 -3122
rect 14642 -3498 14676 -3122
rect 14974 -3498 15008 -3122
rect 15092 -3498 15126 -3122
rect 15210 -3498 15244 -3122
rect 15328 -3498 15362 -3122
rect 15446 -3498 15480 -3122
rect 15564 -3498 15598 -3122
rect 15682 -3498 15716 -3122
rect 16014 -3498 16048 -3122
rect 16132 -3498 16166 -3122
rect 16250 -3498 16284 -3122
rect 16368 -3498 16402 -3122
rect 16486 -3498 16520 -3122
rect 16604 -3498 16638 -3122
rect 16722 -3498 16756 -3122
<< psubdiff >>
rect -1564 6698 -1468 6732
rect 394 6698 490 6732
rect -1564 6636 -1530 6698
rect 456 6636 490 6698
rect -1564 3874 -1530 3936
rect 456 3874 490 3936
rect -1564 3840 -1468 3874
rect 394 3840 490 3874
rect 1236 6698 1332 6732
rect 3194 6698 3290 6732
rect 1236 6636 1270 6698
rect 3256 6636 3290 6698
rect 1236 3874 1270 3936
rect 3256 3874 3290 3936
rect 1236 3840 1332 3874
rect 3194 3840 3290 3874
rect 4320 5604 4416 5638
rect 7366 5604 7462 5638
rect 4320 5542 4354 5604
rect -1144 3750 -1048 3784
rect -18 3750 78 3784
rect -1144 3688 -1110 3750
rect 44 3688 78 3750
rect -1144 3070 -1110 3132
rect 44 3070 78 3132
rect -1144 3036 -1048 3070
rect -18 3036 78 3070
rect 1656 3750 1752 3784
rect 2782 3750 2878 3784
rect 1656 3688 1690 3750
rect 2844 3688 2878 3750
rect 1656 3070 1690 3132
rect 2844 3070 2878 3132
rect 1656 3036 1752 3070
rect 2782 3036 2878 3070
rect 7428 5542 7462 5604
rect 4320 3070 4354 3132
rect 7428 3070 7462 3132
rect 4320 3036 4416 3070
rect 7366 3036 7462 3070
rect 7960 5604 8056 5638
rect 11006 5604 11102 5638
rect 7960 5542 7994 5604
rect 11068 5542 11102 5604
rect 7960 3070 7994 3132
rect 11068 3070 11102 3132
rect 7960 3036 8056 3070
rect 11006 3036 11102 3070
rect 11940 5604 12036 5638
rect 14986 5604 15082 5638
rect 11940 5542 11974 5604
rect 15048 5542 15082 5604
rect 11940 3070 11974 3132
rect 15048 3070 15082 3132
rect 11940 3036 12036 3070
rect 14986 3036 15082 3070
rect 15580 5604 15676 5638
rect 18626 5604 18722 5638
rect 15580 5542 15614 5604
rect 18688 5542 18722 5604
rect 15580 3070 15614 3132
rect 18688 3070 18722 3132
rect 15580 3036 15676 3070
rect 18626 3036 18722 3070
rect 4120 2932 4216 2966
rect 4862 2932 4958 2966
rect 4120 2870 4154 2932
rect -1684 2772 -1588 2806
rect -942 2772 -846 2806
rect -1684 2710 -1650 2772
rect -880 2710 -846 2772
rect -1684 1474 -1650 1536
rect -880 1474 -846 1536
rect -1684 1440 -1588 1474
rect -942 1440 -846 1474
rect -644 2772 -548 2806
rect 98 2772 194 2806
rect -644 2710 -610 2772
rect 160 2710 194 2772
rect -644 1474 -610 1536
rect 160 1474 194 1536
rect -644 1440 -548 1474
rect 98 1440 194 1474
rect 396 2772 492 2806
rect 1138 2772 1234 2806
rect 396 2710 430 2772
rect 1200 2710 1234 2772
rect 396 1474 430 1536
rect 1200 1474 1234 1536
rect 396 1440 492 1474
rect 1138 1440 1234 1474
rect 1436 2772 1532 2806
rect 2178 2772 2274 2806
rect 1436 2710 1470 2772
rect 2240 2710 2274 2772
rect 1436 1474 1470 1536
rect 2240 1474 2274 1536
rect 1436 1440 1532 1474
rect 2178 1440 2274 1474
rect 2476 2772 2572 2806
rect 3218 2772 3314 2806
rect 2476 2710 2510 2772
rect 3280 2710 3314 2772
rect 2476 1474 2510 1536
rect 4924 2870 4958 2932
rect 4120 1634 4154 1696
rect 4924 1634 4958 1696
rect 4120 1600 4216 1634
rect 4862 1600 4958 1634
rect 5160 2932 5256 2966
rect 5902 2932 5998 2966
rect 5160 2870 5194 2932
rect 5964 2870 5998 2932
rect 5160 1634 5194 1696
rect 5964 1634 5998 1696
rect 5160 1600 5256 1634
rect 5902 1600 5998 1634
rect 6200 2932 6296 2966
rect 6942 2932 7038 2966
rect 6200 2870 6234 2932
rect 7004 2870 7038 2932
rect 6200 1634 6234 1696
rect 7004 1634 7038 1696
rect 6200 1600 6296 1634
rect 6942 1600 7038 1634
rect 7240 2932 7336 2966
rect 7982 2932 8078 2966
rect 7240 2870 7274 2932
rect 8044 2870 8078 2932
rect 7240 1634 7274 1696
rect 8044 1634 8078 1696
rect 7240 1600 7336 1634
rect 7982 1600 8078 1634
rect 8280 2932 8376 2966
rect 9022 2932 9118 2966
rect 8280 2870 8314 2932
rect 9084 2870 9118 2932
rect 8280 1634 8314 1696
rect 9084 1634 9118 1696
rect 8280 1600 8376 1634
rect 9022 1600 9118 1634
rect 9320 2932 9416 2966
rect 10062 2932 10158 2966
rect 9320 2870 9354 2932
rect 10124 2870 10158 2932
rect 9320 1634 9354 1696
rect 10124 1634 10158 1696
rect 9320 1600 9416 1634
rect 10062 1600 10158 1634
rect 10360 2932 10456 2966
rect 11102 2932 11198 2966
rect 10360 2870 10394 2932
rect 11164 2870 11198 2932
rect 10360 1634 10394 1696
rect 11164 1634 11198 1696
rect 10360 1600 10456 1634
rect 11102 1600 11198 1634
rect 11740 2932 11836 2966
rect 12482 2932 12578 2966
rect 11740 2870 11774 2932
rect 12544 2870 12578 2932
rect 11740 1634 11774 1696
rect 12544 1634 12578 1696
rect 11740 1600 11836 1634
rect 12482 1600 12578 1634
rect 12780 2932 12876 2966
rect 13522 2932 13618 2966
rect 12780 2870 12814 2932
rect 13584 2870 13618 2932
rect 12780 1634 12814 1696
rect 13584 1634 13618 1696
rect 12780 1600 12876 1634
rect 13522 1600 13618 1634
rect 13820 2932 13916 2966
rect 14562 2932 14658 2966
rect 13820 2870 13854 2932
rect 14624 2870 14658 2932
rect 13820 1634 13854 1696
rect 14624 1634 14658 1696
rect 13820 1600 13916 1634
rect 14562 1600 14658 1634
rect 14860 2932 14956 2966
rect 15602 2932 15698 2966
rect 14860 2870 14894 2932
rect 15664 2870 15698 2932
rect 14860 1634 14894 1696
rect 15664 1634 15698 1696
rect 14860 1600 14956 1634
rect 15602 1600 15698 1634
rect 15900 2932 15996 2966
rect 16642 2932 16738 2966
rect 15900 2870 15934 2932
rect 16704 2870 16738 2932
rect 15900 1634 15934 1696
rect 16704 1634 16738 1696
rect 15900 1600 15996 1634
rect 16642 1600 16738 1634
rect 16940 2932 17036 2966
rect 17682 2932 17778 2966
rect 16940 2870 16974 2932
rect 17744 2870 17778 2932
rect 16940 1634 16974 1696
rect 17744 1634 17778 1696
rect 16940 1600 17036 1634
rect 17682 1600 17778 1634
rect 17980 2932 18076 2966
rect 18722 2932 18818 2966
rect 17980 2870 18014 2932
rect 18784 2870 18818 2932
rect 17980 1634 18014 1696
rect 18784 1634 18818 1696
rect 17980 1600 18076 1634
rect 18722 1600 18818 1634
rect 3280 1474 3314 1536
rect 2476 1440 2572 1474
rect 3218 1440 3314 1474
rect 4120 1510 4216 1544
rect 4994 1510 5090 1544
rect 4120 1448 4154 1510
rect -1684 1350 -1588 1384
rect -810 1350 -714 1384
rect -1684 1288 -1650 1350
rect -748 1288 -714 1350
rect -1684 670 -1650 732
rect -748 670 -714 732
rect -1684 636 -1588 670
rect -810 636 -714 670
rect -644 1350 -548 1384
rect 230 1350 326 1384
rect -644 1288 -610 1350
rect 292 1288 326 1350
rect -644 670 -610 732
rect 292 670 326 732
rect -644 636 -548 670
rect 230 636 326 670
rect 396 1350 492 1384
rect 1270 1350 1366 1384
rect 396 1288 430 1350
rect 1332 1288 1366 1350
rect 396 670 430 732
rect 1332 670 1366 732
rect 396 636 492 670
rect 1270 636 1366 670
rect 1436 1350 1532 1384
rect 2310 1350 2406 1384
rect 1436 1288 1470 1350
rect 2372 1288 2406 1350
rect 1436 670 1470 732
rect 2372 670 2406 732
rect 1436 636 1532 670
rect 2310 636 2406 670
rect 2476 1350 2572 1384
rect 3350 1350 3446 1384
rect 2476 1288 2510 1350
rect 3412 1288 3446 1350
rect 2476 670 2510 732
rect 5056 1448 5090 1510
rect 4120 830 4154 892
rect 5056 830 5090 892
rect 4120 796 4216 830
rect 4994 796 5090 830
rect 5160 1510 5256 1544
rect 6034 1510 6130 1544
rect 5160 1448 5194 1510
rect 6096 1448 6130 1510
rect 5160 830 5194 892
rect 6096 830 6130 892
rect 5160 796 5256 830
rect 6034 796 6130 830
rect 6200 1510 6296 1544
rect 7074 1510 7170 1544
rect 6200 1448 6234 1510
rect 7136 1448 7170 1510
rect 6200 830 6234 892
rect 7136 830 7170 892
rect 6200 796 6296 830
rect 7074 796 7170 830
rect 7240 1510 7336 1544
rect 8114 1510 8210 1544
rect 7240 1448 7274 1510
rect 8176 1448 8210 1510
rect 7240 830 7274 892
rect 8176 830 8210 892
rect 7240 796 7336 830
rect 8114 796 8210 830
rect 8280 1510 8376 1544
rect 9154 1510 9250 1544
rect 8280 1448 8314 1510
rect 9216 1448 9250 1510
rect 8280 830 8314 892
rect 9216 830 9250 892
rect 8280 796 8376 830
rect 9154 796 9250 830
rect 9320 1510 9416 1544
rect 10194 1510 10290 1544
rect 9320 1448 9354 1510
rect 10256 1448 10290 1510
rect 9320 830 9354 892
rect 10256 830 10290 892
rect 9320 796 9416 830
rect 10194 796 10290 830
rect 10360 1510 10456 1544
rect 11234 1510 11330 1544
rect 10360 1448 10394 1510
rect 11296 1448 11330 1510
rect 10360 830 10394 892
rect 11296 830 11330 892
rect 10360 796 10456 830
rect 11234 796 11330 830
rect 11740 1510 11836 1544
rect 12614 1510 12710 1544
rect 11740 1448 11774 1510
rect 12676 1448 12710 1510
rect 11740 830 11774 892
rect 12676 830 12710 892
rect 11740 796 11836 830
rect 12614 796 12710 830
rect 12780 1510 12876 1544
rect 13654 1510 13750 1544
rect 12780 1448 12814 1510
rect 13716 1448 13750 1510
rect 12780 830 12814 892
rect 13716 830 13750 892
rect 12780 796 12876 830
rect 13654 796 13750 830
rect 13820 1510 13916 1544
rect 14694 1510 14790 1544
rect 13820 1448 13854 1510
rect 14756 1448 14790 1510
rect 13820 830 13854 892
rect 14756 830 14790 892
rect 13820 796 13916 830
rect 14694 796 14790 830
rect 14860 1510 14956 1544
rect 15734 1510 15830 1544
rect 14860 1448 14894 1510
rect 15796 1448 15830 1510
rect 14860 830 14894 892
rect 15796 830 15830 892
rect 14860 796 14956 830
rect 15734 796 15830 830
rect 15900 1510 15996 1544
rect 16774 1510 16870 1544
rect 15900 1448 15934 1510
rect 16836 1448 16870 1510
rect 15900 830 15934 892
rect 16836 830 16870 892
rect 15900 796 15996 830
rect 16774 796 16870 830
rect 16940 1510 17036 1544
rect 17814 1510 17910 1544
rect 16940 1448 16974 1510
rect 17876 1448 17910 1510
rect 16940 830 16974 892
rect 17876 830 17910 892
rect 16940 796 17036 830
rect 17814 796 17910 830
rect 17980 1510 18076 1544
rect 18854 1510 18950 1544
rect 17980 1448 18014 1510
rect 18916 1448 18950 1510
rect 17980 830 18014 892
rect 18916 830 18950 892
rect 17980 796 18076 830
rect 18854 796 18950 830
rect 3412 670 3446 732
rect 2476 636 2572 670
rect 3350 636 3446 670
rect 4120 692 4216 726
rect 4862 692 4958 726
rect 4120 630 4154 692
rect -7514 86 -7418 120
rect -6388 86 -6292 120
rect -7514 24 -7480 86
rect -6326 24 -6292 86
rect -7514 -1212 -7480 -1150
rect -6326 -1212 -6292 -1150
rect -7514 -1246 -7418 -1212
rect -6388 -1246 -6292 -1212
rect -6174 72 -6078 106
rect -5722 72 -5626 106
rect -6174 10 -6140 72
rect -7514 -1750 -7418 -1716
rect -6772 -1750 -6676 -1716
rect -7514 -1812 -7480 -1750
rect -6710 -1812 -6676 -1750
rect -7514 -3048 -7480 -2986
rect -5660 10 -5626 72
rect -6174 -1780 -6140 -1718
rect 4924 630 4958 692
rect 4120 -606 4154 -544
rect 4924 -606 4958 -544
rect 4120 -640 4216 -606
rect 4862 -640 4958 -606
rect 5160 692 5256 726
rect 5902 692 5998 726
rect 5160 630 5194 692
rect 5964 630 5998 692
rect 5160 -606 5194 -544
rect 5964 -606 5998 -544
rect 5160 -640 5256 -606
rect 5902 -640 5998 -606
rect 6200 692 6296 726
rect 6942 692 7038 726
rect 6200 630 6234 692
rect 7004 630 7038 692
rect 6200 -606 6234 -544
rect 7004 -606 7038 -544
rect 6200 -640 6296 -606
rect 6942 -640 7038 -606
rect 7240 692 7336 726
rect 7982 692 8078 726
rect 7240 630 7274 692
rect 8044 630 8078 692
rect 7240 -606 7274 -544
rect 8044 -606 8078 -544
rect 7240 -640 7336 -606
rect 7982 -640 8078 -606
rect 8280 692 8376 726
rect 9022 692 9118 726
rect 8280 630 8314 692
rect 9084 630 9118 692
rect 8280 -606 8314 -544
rect 9084 -606 9118 -544
rect 8280 -640 8376 -606
rect 9022 -640 9118 -606
rect 9320 692 9416 726
rect 10062 692 10158 726
rect 9320 630 9354 692
rect 10124 630 10158 692
rect 9320 -606 9354 -544
rect 10124 -606 10158 -544
rect 9320 -640 9416 -606
rect 10062 -640 10158 -606
rect 10360 692 10456 726
rect 11102 692 11198 726
rect 10360 630 10394 692
rect 11164 630 11198 692
rect 10360 -606 10394 -544
rect 11164 -606 11198 -544
rect 10360 -640 10456 -606
rect 11102 -640 11198 -606
rect 11740 692 11836 726
rect 12482 692 12578 726
rect 11740 630 11774 692
rect 12544 630 12578 692
rect 11740 -606 11774 -544
rect 12544 -606 12578 -544
rect 11740 -640 11836 -606
rect 12482 -640 12578 -606
rect 12780 692 12876 726
rect 13522 692 13618 726
rect 12780 630 12814 692
rect 13584 630 13618 692
rect 12780 -606 12814 -544
rect 13584 -606 13618 -544
rect 12780 -640 12876 -606
rect 13522 -640 13618 -606
rect 13820 692 13916 726
rect 14562 692 14658 726
rect 13820 630 13854 692
rect 14624 630 14658 692
rect 13820 -606 13854 -544
rect 14624 -606 14658 -544
rect 13820 -640 13916 -606
rect 14562 -640 14658 -606
rect 14860 692 14956 726
rect 15602 692 15698 726
rect 14860 630 14894 692
rect 15664 630 15698 692
rect 14860 -606 14894 -544
rect 15664 -606 15698 -544
rect 14860 -640 14956 -606
rect 15602 -640 15698 -606
rect 15900 692 15996 726
rect 16642 692 16738 726
rect 15900 630 15934 692
rect 16704 630 16738 692
rect 15900 -606 15934 -544
rect 16704 -606 16738 -544
rect 15900 -640 15996 -606
rect 16642 -640 16738 -606
rect 16940 692 17036 726
rect 17682 692 17778 726
rect 16940 630 16974 692
rect 17744 630 17778 692
rect 16940 -606 16974 -544
rect 17744 -606 17778 -544
rect 16940 -640 17036 -606
rect 17682 -640 17778 -606
rect 17980 692 18076 726
rect 18722 692 18818 726
rect 17980 630 18014 692
rect 18784 630 18818 692
rect 17980 -606 18014 -544
rect 18784 -606 18818 -544
rect 17980 -640 18076 -606
rect 18722 -640 18818 -606
rect 4120 -730 4216 -696
rect 4994 -730 5090 -696
rect 4120 -792 4154 -730
rect 5056 -792 5090 -730
rect 4120 -1410 4154 -1348
rect 5056 -1410 5090 -1348
rect 4120 -1444 4216 -1410
rect 4994 -1444 5090 -1410
rect 5160 -730 5256 -696
rect 6034 -730 6130 -696
rect 5160 -792 5194 -730
rect 6096 -792 6130 -730
rect 5160 -1410 5194 -1348
rect 6096 -1410 6130 -1348
rect 5160 -1444 5256 -1410
rect 6034 -1444 6130 -1410
rect 6200 -730 6296 -696
rect 7074 -730 7170 -696
rect 6200 -792 6234 -730
rect 7136 -792 7170 -730
rect 6200 -1410 6234 -1348
rect 7136 -1410 7170 -1348
rect 6200 -1444 6296 -1410
rect 7074 -1444 7170 -1410
rect 7240 -730 7336 -696
rect 8114 -730 8210 -696
rect 7240 -792 7274 -730
rect 8176 -792 8210 -730
rect 7240 -1410 7274 -1348
rect 8176 -1410 8210 -1348
rect 7240 -1444 7336 -1410
rect 8114 -1444 8210 -1410
rect 8280 -730 8376 -696
rect 9154 -730 9250 -696
rect 8280 -792 8314 -730
rect 9216 -792 9250 -730
rect 8280 -1410 8314 -1348
rect 9216 -1410 9250 -1348
rect 8280 -1444 8376 -1410
rect 9154 -1444 9250 -1410
rect 9320 -730 9416 -696
rect 10194 -730 10290 -696
rect 9320 -792 9354 -730
rect 10256 -792 10290 -730
rect 9320 -1410 9354 -1348
rect 10256 -1410 10290 -1348
rect 9320 -1444 9416 -1410
rect 10194 -1444 10290 -1410
rect 10360 -730 10456 -696
rect 11234 -730 11330 -696
rect 10360 -792 10394 -730
rect 11296 -792 11330 -730
rect 10360 -1410 10394 -1348
rect 11296 -1410 11330 -1348
rect 10360 -1444 10456 -1410
rect 11234 -1444 11330 -1410
rect 11740 -730 11836 -696
rect 12614 -730 12710 -696
rect 11740 -792 11774 -730
rect 12676 -792 12710 -730
rect 11740 -1410 11774 -1348
rect 12676 -1410 12710 -1348
rect 11740 -1444 11836 -1410
rect 12614 -1444 12710 -1410
rect 12780 -730 12876 -696
rect 13654 -730 13750 -696
rect 12780 -792 12814 -730
rect 13716 -792 13750 -730
rect 12780 -1410 12814 -1348
rect 13716 -1410 13750 -1348
rect 12780 -1444 12876 -1410
rect 13654 -1444 13750 -1410
rect 13820 -730 13916 -696
rect 14694 -730 14790 -696
rect 13820 -792 13854 -730
rect 14756 -792 14790 -730
rect 13820 -1410 13854 -1348
rect 14756 -1410 14790 -1348
rect 13820 -1444 13916 -1410
rect 14694 -1444 14790 -1410
rect 14860 -730 14956 -696
rect 15734 -730 15830 -696
rect 14860 -792 14894 -730
rect 15796 -792 15830 -730
rect 14860 -1410 14894 -1348
rect 15796 -1410 15830 -1348
rect 14860 -1444 14956 -1410
rect 15734 -1444 15830 -1410
rect 15900 -730 15996 -696
rect 16774 -730 16870 -696
rect 15900 -792 15934 -730
rect 16836 -792 16870 -730
rect 15900 -1410 15934 -1348
rect 16836 -1410 16870 -1348
rect 15900 -1444 15996 -1410
rect 16774 -1444 16870 -1410
rect 16940 -730 17036 -696
rect 17814 -730 17910 -696
rect 16940 -792 16974 -730
rect 17876 -792 17910 -730
rect 16940 -1410 16974 -1348
rect 17876 -1410 17910 -1348
rect 16940 -1444 17036 -1410
rect 17814 -1444 17910 -1410
rect 17980 -730 18076 -696
rect 18854 -730 18950 -696
rect 17980 -792 18014 -730
rect 18916 -792 18950 -730
rect 17980 -1410 18014 -1348
rect 18916 -1410 18950 -1348
rect 17980 -1444 18076 -1410
rect 18854 -1444 18950 -1410
rect -5660 -1780 -5626 -1718
rect -6174 -1814 -6078 -1780
rect -5722 -1814 -5626 -1780
rect 4120 -1548 4216 -1514
rect 4862 -1548 4958 -1514
rect 4120 -1610 4154 -1548
rect 4924 -1610 4958 -1548
rect 4120 -2846 4154 -2784
rect 4924 -2846 4958 -2784
rect 4120 -2880 4216 -2846
rect 4862 -2880 4958 -2846
rect 5160 -1548 5256 -1514
rect 5902 -1548 5998 -1514
rect 5160 -1610 5194 -1548
rect 5964 -1610 5998 -1548
rect 5160 -2846 5194 -2784
rect 5964 -2846 5998 -2784
rect 5160 -2880 5256 -2846
rect 5902 -2880 5998 -2846
rect 6200 -1548 6296 -1514
rect 6942 -1548 7038 -1514
rect 6200 -1610 6234 -1548
rect 7004 -1610 7038 -1548
rect 6200 -2846 6234 -2784
rect 7004 -2846 7038 -2784
rect 6200 -2880 6296 -2846
rect 6942 -2880 7038 -2846
rect 7240 -1548 7336 -1514
rect 7982 -1548 8078 -1514
rect 7240 -1610 7274 -1548
rect 8044 -1610 8078 -1548
rect 7240 -2846 7274 -2784
rect 8044 -2846 8078 -2784
rect 7240 -2880 7336 -2846
rect 7982 -2880 8078 -2846
rect 8280 -1548 8376 -1514
rect 9022 -1548 9118 -1514
rect 8280 -1610 8314 -1548
rect 9084 -1610 9118 -1548
rect 8280 -2846 8314 -2784
rect 9084 -2846 9118 -2784
rect 8280 -2880 8376 -2846
rect 9022 -2880 9118 -2846
rect 11740 -1548 11836 -1514
rect 12482 -1548 12578 -1514
rect 11740 -1610 11774 -1548
rect 12544 -1610 12578 -1548
rect 11740 -2846 11774 -2784
rect 12544 -2846 12578 -2784
rect 11740 -2880 11836 -2846
rect 12482 -2880 12578 -2846
rect 12780 -1548 12876 -1514
rect 13522 -1548 13618 -1514
rect 12780 -1610 12814 -1548
rect 13584 -1610 13618 -1548
rect 12780 -2846 12814 -2784
rect 13584 -2846 13618 -2784
rect 12780 -2880 12876 -2846
rect 13522 -2880 13618 -2846
rect 13820 -1548 13916 -1514
rect 14562 -1548 14658 -1514
rect 13820 -1610 13854 -1548
rect 14624 -1610 14658 -1548
rect 13820 -2846 13854 -2784
rect 14624 -2846 14658 -2784
rect 13820 -2880 13916 -2846
rect 14562 -2880 14658 -2846
rect 14860 -1548 14956 -1514
rect 15602 -1548 15698 -1514
rect 14860 -1610 14894 -1548
rect 15664 -1610 15698 -1548
rect 14860 -2846 14894 -2784
rect 15664 -2846 15698 -2784
rect 14860 -2880 14956 -2846
rect 15602 -2880 15698 -2846
rect 15900 -1548 15996 -1514
rect 16642 -1548 16738 -1514
rect 15900 -1610 15934 -1548
rect 16704 -1610 16738 -1548
rect 15900 -2846 15934 -2784
rect 16704 -2846 16738 -2784
rect 15900 -2880 15996 -2846
rect 16642 -2880 16738 -2846
rect -6710 -3048 -6676 -2986
rect -7514 -3082 -7418 -3048
rect -6772 -3082 -6676 -3048
rect 4120 -2970 4216 -2936
rect 4994 -2970 5090 -2936
rect 4120 -3032 4154 -2970
rect -7514 -3172 -7418 -3138
rect -6640 -3172 -6544 -3138
rect -7514 -3234 -7480 -3172
rect -6578 -3234 -6544 -3172
rect -7514 -3852 -7480 -3790
rect 5056 -3032 5090 -2970
rect 4120 -3650 4154 -3588
rect 5056 -3650 5090 -3588
rect 4120 -3684 4216 -3650
rect 4994 -3684 5090 -3650
rect 5160 -2970 5256 -2936
rect 6034 -2970 6130 -2936
rect 5160 -3032 5194 -2970
rect 6096 -3032 6130 -2970
rect 5160 -3650 5194 -3588
rect 6096 -3650 6130 -3588
rect 5160 -3684 5256 -3650
rect 6034 -3684 6130 -3650
rect 6200 -2970 6296 -2936
rect 7074 -2970 7170 -2936
rect 6200 -3032 6234 -2970
rect 7136 -3032 7170 -2970
rect 6200 -3650 6234 -3588
rect 7136 -3650 7170 -3588
rect 6200 -3684 6296 -3650
rect 7074 -3684 7170 -3650
rect 7240 -2970 7336 -2936
rect 8114 -2970 8210 -2936
rect 7240 -3032 7274 -2970
rect 8176 -3032 8210 -2970
rect 7240 -3650 7274 -3588
rect 8176 -3650 8210 -3588
rect 7240 -3684 7336 -3650
rect 8114 -3684 8210 -3650
rect 8280 -2970 8376 -2936
rect 9154 -2970 9250 -2936
rect 8280 -3032 8314 -2970
rect 9216 -3032 9250 -2970
rect 8280 -3650 8314 -3588
rect 9216 -3650 9250 -3588
rect 8280 -3684 8376 -3650
rect 9154 -3684 9250 -3650
rect 11740 -2970 11836 -2936
rect 12614 -2970 12710 -2936
rect 11740 -3032 11774 -2970
rect 12676 -3032 12710 -2970
rect 11740 -3650 11774 -3588
rect 12676 -3650 12710 -3588
rect 11740 -3684 11836 -3650
rect 12614 -3684 12710 -3650
rect 12780 -2970 12876 -2936
rect 13654 -2970 13750 -2936
rect 12780 -3032 12814 -2970
rect 13716 -3032 13750 -2970
rect 12780 -3650 12814 -3588
rect 13716 -3650 13750 -3588
rect 12780 -3684 12876 -3650
rect 13654 -3684 13750 -3650
rect 13820 -2970 13916 -2936
rect 14694 -2970 14790 -2936
rect 13820 -3032 13854 -2970
rect 14756 -3032 14790 -2970
rect 13820 -3650 13854 -3588
rect 14756 -3650 14790 -3588
rect 13820 -3684 13916 -3650
rect 14694 -3684 14790 -3650
rect 14860 -2970 14956 -2936
rect 15734 -2970 15830 -2936
rect 14860 -3032 14894 -2970
rect 15796 -3032 15830 -2970
rect 14860 -3650 14894 -3588
rect 15796 -3650 15830 -3588
rect 14860 -3684 14956 -3650
rect 15734 -3684 15830 -3650
rect 15900 -2970 15996 -2936
rect 16774 -2970 16870 -2936
rect 15900 -3032 15934 -2970
rect 16836 -3032 16870 -2970
rect 15900 -3650 15934 -3588
rect 16836 -3650 16870 -3588
rect 15900 -3684 15996 -3650
rect 16774 -3684 16870 -3650
rect -6578 -3852 -6544 -3790
rect -7514 -3886 -7418 -3852
rect -6640 -3886 -6544 -3852
rect -7940 -6448 -7160 -5416
<< psubdiffcont >>
rect -1468 6698 394 6732
rect -1564 3936 -1530 6636
rect 456 3936 490 6636
rect -1468 3840 394 3874
rect 1332 6698 3194 6732
rect 1236 3936 1270 6636
rect 3256 3936 3290 6636
rect 1332 3840 3194 3874
rect 4416 5604 7366 5638
rect -1048 3750 -18 3784
rect -1144 3132 -1110 3688
rect 44 3132 78 3688
rect -1048 3036 -18 3070
rect 1752 3750 2782 3784
rect 1656 3132 1690 3688
rect 2844 3132 2878 3688
rect 1752 3036 2782 3070
rect 4320 3132 4354 5542
rect 7428 3132 7462 5542
rect 4416 3036 7366 3070
rect 8056 5604 11006 5638
rect 7960 3132 7994 5542
rect 11068 3132 11102 5542
rect 8056 3036 11006 3070
rect 12036 5604 14986 5638
rect 11940 3132 11974 5542
rect 15048 3132 15082 5542
rect 12036 3036 14986 3070
rect 15676 5604 18626 5638
rect 15580 3132 15614 5542
rect 18688 3132 18722 5542
rect 15676 3036 18626 3070
rect 4216 2932 4862 2966
rect -1588 2772 -942 2806
rect -1684 1536 -1650 2710
rect -880 1536 -846 2710
rect -1588 1440 -942 1474
rect -548 2772 98 2806
rect -644 1536 -610 2710
rect 160 1536 194 2710
rect -548 1440 98 1474
rect 492 2772 1138 2806
rect 396 1536 430 2710
rect 1200 1536 1234 2710
rect 492 1440 1138 1474
rect 1532 2772 2178 2806
rect 1436 1536 1470 2710
rect 2240 1536 2274 2710
rect 1532 1440 2178 1474
rect 2572 2772 3218 2806
rect 2476 1536 2510 2710
rect 3280 1536 3314 2710
rect 4120 1696 4154 2870
rect 4924 1696 4958 2870
rect 4216 1600 4862 1634
rect 5256 2932 5902 2966
rect 5160 1696 5194 2870
rect 5964 1696 5998 2870
rect 5256 1600 5902 1634
rect 6296 2932 6942 2966
rect 6200 1696 6234 2870
rect 7004 1696 7038 2870
rect 6296 1600 6942 1634
rect 7336 2932 7982 2966
rect 7240 1696 7274 2870
rect 8044 1696 8078 2870
rect 7336 1600 7982 1634
rect 8376 2932 9022 2966
rect 8280 1696 8314 2870
rect 9084 1696 9118 2870
rect 8376 1600 9022 1634
rect 9416 2932 10062 2966
rect 9320 1696 9354 2870
rect 10124 1696 10158 2870
rect 9416 1600 10062 1634
rect 10456 2932 11102 2966
rect 10360 1696 10394 2870
rect 11164 1696 11198 2870
rect 10456 1600 11102 1634
rect 11836 2932 12482 2966
rect 11740 1696 11774 2870
rect 12544 1696 12578 2870
rect 11836 1600 12482 1634
rect 12876 2932 13522 2966
rect 12780 1696 12814 2870
rect 13584 1696 13618 2870
rect 12876 1600 13522 1634
rect 13916 2932 14562 2966
rect 13820 1696 13854 2870
rect 14624 1696 14658 2870
rect 13916 1600 14562 1634
rect 14956 2932 15602 2966
rect 14860 1696 14894 2870
rect 15664 1696 15698 2870
rect 14956 1600 15602 1634
rect 15996 2932 16642 2966
rect 15900 1696 15934 2870
rect 16704 1696 16738 2870
rect 15996 1600 16642 1634
rect 17036 2932 17682 2966
rect 16940 1696 16974 2870
rect 17744 1696 17778 2870
rect 17036 1600 17682 1634
rect 18076 2932 18722 2966
rect 17980 1696 18014 2870
rect 18784 1696 18818 2870
rect 18076 1600 18722 1634
rect 2572 1440 3218 1474
rect 4216 1510 4994 1544
rect -1588 1350 -810 1384
rect -1684 732 -1650 1288
rect -748 732 -714 1288
rect -1588 636 -810 670
rect -548 1350 230 1384
rect -644 732 -610 1288
rect 292 732 326 1288
rect -548 636 230 670
rect 492 1350 1270 1384
rect 396 732 430 1288
rect 1332 732 1366 1288
rect 492 636 1270 670
rect 1532 1350 2310 1384
rect 1436 732 1470 1288
rect 2372 732 2406 1288
rect 1532 636 2310 670
rect 2572 1350 3350 1384
rect 2476 732 2510 1288
rect 3412 732 3446 1288
rect 4120 892 4154 1448
rect 5056 892 5090 1448
rect 4216 796 4994 830
rect 5256 1510 6034 1544
rect 5160 892 5194 1448
rect 6096 892 6130 1448
rect 5256 796 6034 830
rect 6296 1510 7074 1544
rect 6200 892 6234 1448
rect 7136 892 7170 1448
rect 6296 796 7074 830
rect 7336 1510 8114 1544
rect 7240 892 7274 1448
rect 8176 892 8210 1448
rect 7336 796 8114 830
rect 8376 1510 9154 1544
rect 8280 892 8314 1448
rect 9216 892 9250 1448
rect 8376 796 9154 830
rect 9416 1510 10194 1544
rect 9320 892 9354 1448
rect 10256 892 10290 1448
rect 9416 796 10194 830
rect 10456 1510 11234 1544
rect 10360 892 10394 1448
rect 11296 892 11330 1448
rect 10456 796 11234 830
rect 11836 1510 12614 1544
rect 11740 892 11774 1448
rect 12676 892 12710 1448
rect 11836 796 12614 830
rect 12876 1510 13654 1544
rect 12780 892 12814 1448
rect 13716 892 13750 1448
rect 12876 796 13654 830
rect 13916 1510 14694 1544
rect 13820 892 13854 1448
rect 14756 892 14790 1448
rect 13916 796 14694 830
rect 14956 1510 15734 1544
rect 14860 892 14894 1448
rect 15796 892 15830 1448
rect 14956 796 15734 830
rect 15996 1510 16774 1544
rect 15900 892 15934 1448
rect 16836 892 16870 1448
rect 15996 796 16774 830
rect 17036 1510 17814 1544
rect 16940 892 16974 1448
rect 17876 892 17910 1448
rect 17036 796 17814 830
rect 18076 1510 18854 1544
rect 17980 892 18014 1448
rect 18916 892 18950 1448
rect 18076 796 18854 830
rect 2572 636 3350 670
rect 4216 692 4862 726
rect -7418 86 -6388 120
rect -7514 -1150 -7480 24
rect -6326 -1150 -6292 24
rect -7418 -1246 -6388 -1212
rect -6078 72 -5722 106
rect -7418 -1750 -6772 -1716
rect -7514 -2986 -7480 -1812
rect -6710 -2986 -6676 -1812
rect -6174 -1718 -6140 10
rect -5660 -1718 -5626 10
rect 4120 -544 4154 630
rect 4924 -544 4958 630
rect 4216 -640 4862 -606
rect 5256 692 5902 726
rect 5160 -544 5194 630
rect 5964 -544 5998 630
rect 5256 -640 5902 -606
rect 6296 692 6942 726
rect 6200 -544 6234 630
rect 7004 -544 7038 630
rect 6296 -640 6942 -606
rect 7336 692 7982 726
rect 7240 -544 7274 630
rect 8044 -544 8078 630
rect 7336 -640 7982 -606
rect 8376 692 9022 726
rect 8280 -544 8314 630
rect 9084 -544 9118 630
rect 8376 -640 9022 -606
rect 9416 692 10062 726
rect 9320 -544 9354 630
rect 10124 -544 10158 630
rect 9416 -640 10062 -606
rect 10456 692 11102 726
rect 10360 -544 10394 630
rect 11164 -544 11198 630
rect 10456 -640 11102 -606
rect 11836 692 12482 726
rect 11740 -544 11774 630
rect 12544 -544 12578 630
rect 11836 -640 12482 -606
rect 12876 692 13522 726
rect 12780 -544 12814 630
rect 13584 -544 13618 630
rect 12876 -640 13522 -606
rect 13916 692 14562 726
rect 13820 -544 13854 630
rect 14624 -544 14658 630
rect 13916 -640 14562 -606
rect 14956 692 15602 726
rect 14860 -544 14894 630
rect 15664 -544 15698 630
rect 14956 -640 15602 -606
rect 15996 692 16642 726
rect 15900 -544 15934 630
rect 16704 -544 16738 630
rect 15996 -640 16642 -606
rect 17036 692 17682 726
rect 16940 -544 16974 630
rect 17744 -544 17778 630
rect 17036 -640 17682 -606
rect 18076 692 18722 726
rect 17980 -544 18014 630
rect 18784 -544 18818 630
rect 18076 -640 18722 -606
rect 4216 -730 4994 -696
rect 4120 -1348 4154 -792
rect 5056 -1348 5090 -792
rect 4216 -1444 4994 -1410
rect 5256 -730 6034 -696
rect 5160 -1348 5194 -792
rect 6096 -1348 6130 -792
rect 5256 -1444 6034 -1410
rect 6296 -730 7074 -696
rect 6200 -1348 6234 -792
rect 7136 -1348 7170 -792
rect 6296 -1444 7074 -1410
rect 7336 -730 8114 -696
rect 7240 -1348 7274 -792
rect 8176 -1348 8210 -792
rect 7336 -1444 8114 -1410
rect 8376 -730 9154 -696
rect 8280 -1348 8314 -792
rect 9216 -1348 9250 -792
rect 8376 -1444 9154 -1410
rect 9416 -730 10194 -696
rect 9320 -1348 9354 -792
rect 10256 -1348 10290 -792
rect 9416 -1444 10194 -1410
rect 10456 -730 11234 -696
rect 10360 -1348 10394 -792
rect 11296 -1348 11330 -792
rect 10456 -1444 11234 -1410
rect 11836 -730 12614 -696
rect 11740 -1348 11774 -792
rect 12676 -1348 12710 -792
rect 11836 -1444 12614 -1410
rect 12876 -730 13654 -696
rect 12780 -1348 12814 -792
rect 13716 -1348 13750 -792
rect 12876 -1444 13654 -1410
rect 13916 -730 14694 -696
rect 13820 -1348 13854 -792
rect 14756 -1348 14790 -792
rect 13916 -1444 14694 -1410
rect 14956 -730 15734 -696
rect 14860 -1348 14894 -792
rect 15796 -1348 15830 -792
rect 14956 -1444 15734 -1410
rect 15996 -730 16774 -696
rect 15900 -1348 15934 -792
rect 16836 -1348 16870 -792
rect 15996 -1444 16774 -1410
rect 17036 -730 17814 -696
rect 16940 -1348 16974 -792
rect 17876 -1348 17910 -792
rect 17036 -1444 17814 -1410
rect 18076 -730 18854 -696
rect 17980 -1348 18014 -792
rect 18916 -1348 18950 -792
rect 18076 -1444 18854 -1410
rect -6078 -1814 -5722 -1780
rect 4216 -1548 4862 -1514
rect 4120 -2784 4154 -1610
rect 4924 -2784 4958 -1610
rect 4216 -2880 4862 -2846
rect 5256 -1548 5902 -1514
rect 5160 -2784 5194 -1610
rect 5964 -2784 5998 -1610
rect 5256 -2880 5902 -2846
rect 6296 -1548 6942 -1514
rect 6200 -2784 6234 -1610
rect 7004 -2784 7038 -1610
rect 6296 -2880 6942 -2846
rect 7336 -1548 7982 -1514
rect 7240 -2784 7274 -1610
rect 8044 -2784 8078 -1610
rect 7336 -2880 7982 -2846
rect 8376 -1548 9022 -1514
rect 8280 -2784 8314 -1610
rect 9084 -2784 9118 -1610
rect 8376 -2880 9022 -2846
rect 11836 -1548 12482 -1514
rect 11740 -2784 11774 -1610
rect 12544 -2784 12578 -1610
rect 11836 -2880 12482 -2846
rect 12876 -1548 13522 -1514
rect 12780 -2784 12814 -1610
rect 13584 -2784 13618 -1610
rect 12876 -2880 13522 -2846
rect 13916 -1548 14562 -1514
rect 13820 -2784 13854 -1610
rect 14624 -2784 14658 -1610
rect 13916 -2880 14562 -2846
rect 14956 -1548 15602 -1514
rect 14860 -2784 14894 -1610
rect 15664 -2784 15698 -1610
rect 14956 -2880 15602 -2846
rect 15996 -1548 16642 -1514
rect 15900 -2784 15934 -1610
rect 16704 -2784 16738 -1610
rect 15996 -2880 16642 -2846
rect -7418 -3082 -6772 -3048
rect 4216 -2970 4994 -2936
rect -7418 -3172 -6640 -3138
rect -7514 -3790 -7480 -3234
rect -6578 -3790 -6544 -3234
rect 4120 -3588 4154 -3032
rect 5056 -3588 5090 -3032
rect 4216 -3684 4994 -3650
rect 5256 -2970 6034 -2936
rect 5160 -3588 5194 -3032
rect 6096 -3588 6130 -3032
rect 5256 -3684 6034 -3650
rect 6296 -2970 7074 -2936
rect 6200 -3588 6234 -3032
rect 7136 -3588 7170 -3032
rect 6296 -3684 7074 -3650
rect 7336 -2970 8114 -2936
rect 7240 -3588 7274 -3032
rect 8176 -3588 8210 -3032
rect 7336 -3684 8114 -3650
rect 8376 -2970 9154 -2936
rect 8280 -3588 8314 -3032
rect 9216 -3588 9250 -3032
rect 8376 -3684 9154 -3650
rect 11836 -2970 12614 -2936
rect 11740 -3588 11774 -3032
rect 12676 -3588 12710 -3032
rect 11836 -3684 12614 -3650
rect 12876 -2970 13654 -2936
rect 12780 -3588 12814 -3032
rect 13716 -3588 13750 -3032
rect 12876 -3684 13654 -3650
rect 13916 -2970 14694 -2936
rect 13820 -3588 13854 -3032
rect 14756 -3588 14790 -3032
rect 13916 -3684 14694 -3650
rect 14956 -2970 15734 -2936
rect 14860 -3588 14894 -3032
rect 15796 -3588 15830 -3032
rect 14956 -3684 15734 -3650
rect 15996 -2970 16774 -2936
rect 15900 -3588 15934 -3032
rect 16836 -3588 16870 -3032
rect 15996 -3684 16774 -3650
rect -7418 -3886 -6640 -3852
<< poly >>
rect -902 3682 -836 3698
rect -902 3648 -886 3682
rect -852 3648 -836 3682
rect -980 3610 -950 3636
rect -902 3632 -836 3648
rect -710 3682 -644 3698
rect -710 3648 -694 3682
rect -660 3648 -644 3682
rect -884 3610 -854 3632
rect -788 3610 -758 3636
rect -710 3632 -644 3648
rect -518 3682 -452 3698
rect -518 3648 -502 3682
rect -468 3648 -452 3682
rect -692 3610 -662 3632
rect -596 3610 -566 3636
rect -518 3632 -452 3648
rect -326 3682 -260 3698
rect -326 3648 -310 3682
rect -276 3648 -260 3682
rect -500 3610 -470 3632
rect -404 3610 -374 3636
rect -326 3632 -260 3648
rect -134 3682 -68 3698
rect -134 3648 -118 3682
rect -84 3648 -68 3682
rect -308 3610 -278 3632
rect -212 3610 -182 3636
rect -134 3632 -68 3648
rect -116 3610 -86 3632
rect -980 3188 -950 3210
rect -998 3172 -932 3188
rect -884 3184 -854 3210
rect -788 3188 -758 3210
rect -998 3138 -982 3172
rect -948 3138 -932 3172
rect -998 3122 -932 3138
rect -806 3172 -740 3188
rect -692 3184 -662 3210
rect -596 3188 -566 3210
rect -806 3138 -790 3172
rect -756 3138 -740 3172
rect -806 3122 -740 3138
rect -614 3172 -548 3188
rect -500 3184 -470 3210
rect -404 3188 -374 3210
rect -614 3138 -598 3172
rect -564 3138 -548 3172
rect -614 3122 -548 3138
rect -422 3172 -356 3188
rect -308 3184 -278 3210
rect -212 3188 -182 3210
rect -422 3138 -406 3172
rect -372 3138 -356 3172
rect -422 3122 -356 3138
rect -230 3172 -164 3188
rect -116 3184 -86 3210
rect -230 3138 -214 3172
rect -180 3138 -164 3172
rect -230 3122 -164 3138
rect 1898 3682 1964 3698
rect 1898 3648 1914 3682
rect 1948 3648 1964 3682
rect 1820 3610 1850 3636
rect 1898 3632 1964 3648
rect 2090 3682 2156 3698
rect 2090 3648 2106 3682
rect 2140 3648 2156 3682
rect 1916 3610 1946 3632
rect 2012 3610 2042 3636
rect 2090 3632 2156 3648
rect 2282 3682 2348 3698
rect 2282 3648 2298 3682
rect 2332 3648 2348 3682
rect 2108 3610 2138 3632
rect 2204 3610 2234 3636
rect 2282 3632 2348 3648
rect 2474 3682 2540 3698
rect 2474 3648 2490 3682
rect 2524 3648 2540 3682
rect 2300 3610 2330 3632
rect 2396 3610 2426 3636
rect 2474 3632 2540 3648
rect 2666 3682 2732 3698
rect 2666 3648 2682 3682
rect 2716 3648 2732 3682
rect 2492 3610 2522 3632
rect 2588 3610 2618 3636
rect 2666 3632 2732 3648
rect 2684 3610 2714 3632
rect 1820 3188 1850 3210
rect 1802 3172 1868 3188
rect 1916 3184 1946 3210
rect 2012 3188 2042 3210
rect 1802 3138 1818 3172
rect 1852 3138 1868 3172
rect 1802 3122 1868 3138
rect 1994 3172 2060 3188
rect 2108 3184 2138 3210
rect 2204 3188 2234 3210
rect 1994 3138 2010 3172
rect 2044 3138 2060 3172
rect 1994 3122 2060 3138
rect 2186 3172 2252 3188
rect 2300 3184 2330 3210
rect 2396 3188 2426 3210
rect 2186 3138 2202 3172
rect 2236 3138 2252 3172
rect 2186 3122 2252 3138
rect 2378 3172 2444 3188
rect 2492 3184 2522 3210
rect 2588 3188 2618 3210
rect 2378 3138 2394 3172
rect 2428 3138 2444 3172
rect 2378 3122 2444 3138
rect 2570 3172 2636 3188
rect 2684 3184 2714 3210
rect 2570 3138 2586 3172
rect 2620 3138 2636 3172
rect 2570 3122 2636 3138
rect 4466 5536 4532 5552
rect 4466 5502 4482 5536
rect 4516 5502 4532 5536
rect 4466 5486 4532 5502
rect 4658 5536 4724 5552
rect 4658 5502 4674 5536
rect 4708 5502 4724 5536
rect 4484 5464 4514 5486
rect 4580 5464 4610 5490
rect 4658 5486 4724 5502
rect 4850 5536 4916 5552
rect 4850 5502 4866 5536
rect 4900 5502 4916 5536
rect 4676 5464 4706 5486
rect 4772 5464 4802 5490
rect 4850 5486 4916 5502
rect 5042 5536 5108 5552
rect 5042 5502 5058 5536
rect 5092 5502 5108 5536
rect 4868 5464 4898 5486
rect 4964 5464 4994 5490
rect 5042 5486 5108 5502
rect 5234 5536 5300 5552
rect 5234 5502 5250 5536
rect 5284 5502 5300 5536
rect 5060 5464 5090 5486
rect 5156 5464 5186 5490
rect 5234 5486 5300 5502
rect 5426 5536 5492 5552
rect 5426 5502 5442 5536
rect 5476 5502 5492 5536
rect 5252 5464 5282 5486
rect 5348 5464 5378 5490
rect 5426 5486 5492 5502
rect 5618 5536 5684 5552
rect 5618 5502 5634 5536
rect 5668 5502 5684 5536
rect 5444 5464 5474 5486
rect 5540 5464 5570 5490
rect 5618 5486 5684 5502
rect 5810 5536 5876 5552
rect 5810 5502 5826 5536
rect 5860 5502 5876 5536
rect 5636 5464 5666 5486
rect 5732 5464 5762 5490
rect 5810 5486 5876 5502
rect 6002 5536 6068 5552
rect 6002 5502 6018 5536
rect 6052 5502 6068 5536
rect 5828 5464 5858 5486
rect 5924 5464 5954 5490
rect 6002 5486 6068 5502
rect 6194 5536 6260 5552
rect 6194 5502 6210 5536
rect 6244 5502 6260 5536
rect 6020 5464 6050 5486
rect 6116 5464 6146 5490
rect 6194 5486 6260 5502
rect 6386 5536 6452 5552
rect 6386 5502 6402 5536
rect 6436 5502 6452 5536
rect 6212 5464 6242 5486
rect 6308 5464 6338 5490
rect 6386 5486 6452 5502
rect 6578 5536 6644 5552
rect 6578 5502 6594 5536
rect 6628 5502 6644 5536
rect 6404 5464 6434 5486
rect 6500 5464 6530 5490
rect 6578 5486 6644 5502
rect 6770 5536 6836 5552
rect 6770 5502 6786 5536
rect 6820 5502 6836 5536
rect 6596 5464 6626 5486
rect 6692 5464 6722 5490
rect 6770 5486 6836 5502
rect 6962 5536 7028 5552
rect 6962 5502 6978 5536
rect 7012 5502 7028 5536
rect 6788 5464 6818 5486
rect 6884 5464 6914 5490
rect 6962 5486 7028 5502
rect 7154 5536 7220 5552
rect 7154 5502 7170 5536
rect 7204 5502 7220 5536
rect 6980 5464 7010 5486
rect 7076 5464 7106 5490
rect 7154 5486 7220 5502
rect 7172 5464 7202 5486
rect 7268 5464 7298 5490
rect 4484 5038 4514 5064
rect 4580 5042 4610 5064
rect 4562 5026 4628 5042
rect 4676 5038 4706 5064
rect 4772 5042 4802 5064
rect 4562 4992 4578 5026
rect 4612 4992 4628 5026
rect 4562 4976 4628 4992
rect 4754 5026 4820 5042
rect 4868 5038 4898 5064
rect 4964 5042 4994 5064
rect 4754 4992 4770 5026
rect 4804 4992 4820 5026
rect 4754 4976 4820 4992
rect 4946 5026 5012 5042
rect 5060 5038 5090 5064
rect 5156 5042 5186 5064
rect 4946 4992 4962 5026
rect 4996 4992 5012 5026
rect 4946 4976 5012 4992
rect 5138 5026 5204 5042
rect 5252 5038 5282 5064
rect 5348 5042 5378 5064
rect 5138 4992 5154 5026
rect 5188 4992 5204 5026
rect 5138 4976 5204 4992
rect 5330 5026 5396 5042
rect 5444 5038 5474 5064
rect 5540 5042 5570 5064
rect 5330 4992 5346 5026
rect 5380 4992 5396 5026
rect 5330 4976 5396 4992
rect 5522 5026 5588 5042
rect 5636 5038 5666 5064
rect 5732 5042 5762 5064
rect 5522 4992 5538 5026
rect 5572 4992 5588 5026
rect 5522 4976 5588 4992
rect 5714 5026 5780 5042
rect 5828 5038 5858 5064
rect 5924 5042 5954 5064
rect 5714 4992 5730 5026
rect 5764 4992 5780 5026
rect 5714 4976 5780 4992
rect 5906 5026 5972 5042
rect 6020 5038 6050 5064
rect 6116 5042 6146 5064
rect 5906 4992 5922 5026
rect 5956 4992 5972 5026
rect 5906 4976 5972 4992
rect 6098 5026 6164 5042
rect 6212 5038 6242 5064
rect 6308 5042 6338 5064
rect 6098 4992 6114 5026
rect 6148 4992 6164 5026
rect 6098 4976 6164 4992
rect 6290 5026 6356 5042
rect 6404 5038 6434 5064
rect 6500 5042 6530 5064
rect 6290 4992 6306 5026
rect 6340 4992 6356 5026
rect 6290 4976 6356 4992
rect 6482 5026 6548 5042
rect 6596 5038 6626 5064
rect 6692 5042 6722 5064
rect 6482 4992 6498 5026
rect 6532 4992 6548 5026
rect 6482 4976 6548 4992
rect 6674 5026 6740 5042
rect 6788 5038 6818 5064
rect 6884 5042 6914 5064
rect 6674 4992 6690 5026
rect 6724 4992 6740 5026
rect 6674 4976 6740 4992
rect 6866 5026 6932 5042
rect 6980 5038 7010 5064
rect 7076 5042 7106 5064
rect 6866 4992 6882 5026
rect 6916 4992 6932 5026
rect 6866 4976 6932 4992
rect 7058 5026 7124 5042
rect 7172 5038 7202 5064
rect 7268 5042 7298 5064
rect 7058 4992 7074 5026
rect 7108 4992 7124 5026
rect 7058 4976 7124 4992
rect 7250 5026 7316 5042
rect 7250 4992 7266 5026
rect 7300 4992 7316 5026
rect 7250 4976 7316 4992
rect 4562 4918 4628 4934
rect 4562 4884 4578 4918
rect 4612 4884 4628 4918
rect 4484 4846 4514 4872
rect 4562 4868 4628 4884
rect 4754 4918 4820 4934
rect 4754 4884 4770 4918
rect 4804 4884 4820 4918
rect 4580 4846 4610 4868
rect 4676 4846 4706 4872
rect 4754 4868 4820 4884
rect 4946 4918 5012 4934
rect 4946 4884 4962 4918
rect 4996 4884 5012 4918
rect 4772 4846 4802 4868
rect 4868 4846 4898 4872
rect 4946 4868 5012 4884
rect 5138 4918 5204 4934
rect 5138 4884 5154 4918
rect 5188 4884 5204 4918
rect 4964 4846 4994 4868
rect 5060 4846 5090 4872
rect 5138 4868 5204 4884
rect 5330 4918 5396 4934
rect 5330 4884 5346 4918
rect 5380 4884 5396 4918
rect 5156 4846 5186 4868
rect 5252 4846 5282 4872
rect 5330 4868 5396 4884
rect 5522 4918 5588 4934
rect 5522 4884 5538 4918
rect 5572 4884 5588 4918
rect 5348 4846 5378 4868
rect 5444 4846 5474 4872
rect 5522 4868 5588 4884
rect 5714 4918 5780 4934
rect 5714 4884 5730 4918
rect 5764 4884 5780 4918
rect 5540 4846 5570 4868
rect 5636 4846 5666 4872
rect 5714 4868 5780 4884
rect 5906 4918 5972 4934
rect 5906 4884 5922 4918
rect 5956 4884 5972 4918
rect 5732 4846 5762 4868
rect 5828 4846 5858 4872
rect 5906 4868 5972 4884
rect 6098 4918 6164 4934
rect 6098 4884 6114 4918
rect 6148 4884 6164 4918
rect 5924 4846 5954 4868
rect 6020 4846 6050 4872
rect 6098 4868 6164 4884
rect 6290 4918 6356 4934
rect 6290 4884 6306 4918
rect 6340 4884 6356 4918
rect 6116 4846 6146 4868
rect 6212 4846 6242 4872
rect 6290 4868 6356 4884
rect 6482 4918 6548 4934
rect 6482 4884 6498 4918
rect 6532 4884 6548 4918
rect 6308 4846 6338 4868
rect 6404 4846 6434 4872
rect 6482 4868 6548 4884
rect 6674 4918 6740 4934
rect 6674 4884 6690 4918
rect 6724 4884 6740 4918
rect 6500 4846 6530 4868
rect 6596 4846 6626 4872
rect 6674 4868 6740 4884
rect 6866 4918 6932 4934
rect 6866 4884 6882 4918
rect 6916 4884 6932 4918
rect 6692 4846 6722 4868
rect 6788 4846 6818 4872
rect 6866 4868 6932 4884
rect 7058 4918 7124 4934
rect 7058 4884 7074 4918
rect 7108 4884 7124 4918
rect 6884 4846 6914 4868
rect 6980 4846 7010 4872
rect 7058 4868 7124 4884
rect 7250 4918 7316 4934
rect 7250 4884 7266 4918
rect 7300 4884 7316 4918
rect 7076 4846 7106 4868
rect 7172 4846 7202 4872
rect 7250 4868 7316 4884
rect 7268 4846 7298 4868
rect 4484 4424 4514 4446
rect 4466 4408 4532 4424
rect 4580 4420 4610 4446
rect 4676 4424 4706 4446
rect 4466 4374 4482 4408
rect 4516 4374 4532 4408
rect 4466 4358 4532 4374
rect 4658 4408 4724 4424
rect 4772 4420 4802 4446
rect 4868 4424 4898 4446
rect 4658 4374 4674 4408
rect 4708 4374 4724 4408
rect 4658 4358 4724 4374
rect 4850 4408 4916 4424
rect 4964 4420 4994 4446
rect 5060 4424 5090 4446
rect 4850 4374 4866 4408
rect 4900 4374 4916 4408
rect 4850 4358 4916 4374
rect 5042 4408 5108 4424
rect 5156 4420 5186 4446
rect 5252 4424 5282 4446
rect 5042 4374 5058 4408
rect 5092 4374 5108 4408
rect 5042 4358 5108 4374
rect 5234 4408 5300 4424
rect 5348 4420 5378 4446
rect 5444 4424 5474 4446
rect 5234 4374 5250 4408
rect 5284 4374 5300 4408
rect 5234 4358 5300 4374
rect 5426 4408 5492 4424
rect 5540 4420 5570 4446
rect 5636 4424 5666 4446
rect 5426 4374 5442 4408
rect 5476 4374 5492 4408
rect 5426 4358 5492 4374
rect 5618 4408 5684 4424
rect 5732 4420 5762 4446
rect 5828 4424 5858 4446
rect 5618 4374 5634 4408
rect 5668 4374 5684 4408
rect 5618 4358 5684 4374
rect 5810 4408 5876 4424
rect 5924 4420 5954 4446
rect 6020 4424 6050 4446
rect 5810 4374 5826 4408
rect 5860 4374 5876 4408
rect 5810 4358 5876 4374
rect 6002 4408 6068 4424
rect 6116 4420 6146 4446
rect 6212 4424 6242 4446
rect 6002 4374 6018 4408
rect 6052 4374 6068 4408
rect 6002 4358 6068 4374
rect 6194 4408 6260 4424
rect 6308 4420 6338 4446
rect 6404 4424 6434 4446
rect 6194 4374 6210 4408
rect 6244 4374 6260 4408
rect 6194 4358 6260 4374
rect 6386 4408 6452 4424
rect 6500 4420 6530 4446
rect 6596 4424 6626 4446
rect 6386 4374 6402 4408
rect 6436 4374 6452 4408
rect 6386 4358 6452 4374
rect 6578 4408 6644 4424
rect 6692 4420 6722 4446
rect 6788 4424 6818 4446
rect 6578 4374 6594 4408
rect 6628 4374 6644 4408
rect 6578 4358 6644 4374
rect 6770 4408 6836 4424
rect 6884 4420 6914 4446
rect 6980 4424 7010 4446
rect 6770 4374 6786 4408
rect 6820 4374 6836 4408
rect 6770 4358 6836 4374
rect 6962 4408 7028 4424
rect 7076 4420 7106 4446
rect 7172 4424 7202 4446
rect 6962 4374 6978 4408
rect 7012 4374 7028 4408
rect 6962 4358 7028 4374
rect 7154 4408 7220 4424
rect 7268 4420 7298 4446
rect 7154 4374 7170 4408
rect 7204 4374 7220 4408
rect 7154 4358 7220 4374
rect 4466 4300 4532 4316
rect 4466 4266 4482 4300
rect 4516 4266 4532 4300
rect 4466 4250 4532 4266
rect 4658 4300 4724 4316
rect 4658 4266 4674 4300
rect 4708 4266 4724 4300
rect 4484 4228 4514 4250
rect 4580 4228 4610 4254
rect 4658 4250 4724 4266
rect 4850 4300 4916 4316
rect 4850 4266 4866 4300
rect 4900 4266 4916 4300
rect 4676 4228 4706 4250
rect 4772 4228 4802 4254
rect 4850 4250 4916 4266
rect 5042 4300 5108 4316
rect 5042 4266 5058 4300
rect 5092 4266 5108 4300
rect 4868 4228 4898 4250
rect 4964 4228 4994 4254
rect 5042 4250 5108 4266
rect 5234 4300 5300 4316
rect 5234 4266 5250 4300
rect 5284 4266 5300 4300
rect 5060 4228 5090 4250
rect 5156 4228 5186 4254
rect 5234 4250 5300 4266
rect 5426 4300 5492 4316
rect 5426 4266 5442 4300
rect 5476 4266 5492 4300
rect 5252 4228 5282 4250
rect 5348 4228 5378 4254
rect 5426 4250 5492 4266
rect 5618 4300 5684 4316
rect 5618 4266 5634 4300
rect 5668 4266 5684 4300
rect 5444 4228 5474 4250
rect 5540 4228 5570 4254
rect 5618 4250 5684 4266
rect 5810 4300 5876 4316
rect 5810 4266 5826 4300
rect 5860 4266 5876 4300
rect 5636 4228 5666 4250
rect 5732 4228 5762 4254
rect 5810 4250 5876 4266
rect 6002 4300 6068 4316
rect 6002 4266 6018 4300
rect 6052 4266 6068 4300
rect 5828 4228 5858 4250
rect 5924 4228 5954 4254
rect 6002 4250 6068 4266
rect 6194 4300 6260 4316
rect 6194 4266 6210 4300
rect 6244 4266 6260 4300
rect 6020 4228 6050 4250
rect 6116 4228 6146 4254
rect 6194 4250 6260 4266
rect 6386 4300 6452 4316
rect 6386 4266 6402 4300
rect 6436 4266 6452 4300
rect 6212 4228 6242 4250
rect 6308 4228 6338 4254
rect 6386 4250 6452 4266
rect 6578 4300 6644 4316
rect 6578 4266 6594 4300
rect 6628 4266 6644 4300
rect 6404 4228 6434 4250
rect 6500 4228 6530 4254
rect 6578 4250 6644 4266
rect 6770 4300 6836 4316
rect 6770 4266 6786 4300
rect 6820 4266 6836 4300
rect 6596 4228 6626 4250
rect 6692 4228 6722 4254
rect 6770 4250 6836 4266
rect 6962 4300 7028 4316
rect 6962 4266 6978 4300
rect 7012 4266 7028 4300
rect 6788 4228 6818 4250
rect 6884 4228 6914 4254
rect 6962 4250 7028 4266
rect 7154 4300 7220 4316
rect 7154 4266 7170 4300
rect 7204 4266 7220 4300
rect 6980 4228 7010 4250
rect 7076 4228 7106 4254
rect 7154 4250 7220 4266
rect 7172 4228 7202 4250
rect 7268 4228 7298 4254
rect 4484 3802 4514 3828
rect 4580 3806 4610 3828
rect 4562 3790 4628 3806
rect 4676 3802 4706 3828
rect 4772 3806 4802 3828
rect 4562 3756 4578 3790
rect 4612 3756 4628 3790
rect 4562 3740 4628 3756
rect 4754 3790 4820 3806
rect 4868 3802 4898 3828
rect 4964 3806 4994 3828
rect 4754 3756 4770 3790
rect 4804 3756 4820 3790
rect 4754 3740 4820 3756
rect 4946 3790 5012 3806
rect 5060 3802 5090 3828
rect 5156 3806 5186 3828
rect 4946 3756 4962 3790
rect 4996 3756 5012 3790
rect 4946 3740 5012 3756
rect 5138 3790 5204 3806
rect 5252 3802 5282 3828
rect 5348 3806 5378 3828
rect 5138 3756 5154 3790
rect 5188 3756 5204 3790
rect 5138 3740 5204 3756
rect 5330 3790 5396 3806
rect 5444 3802 5474 3828
rect 5540 3806 5570 3828
rect 5330 3756 5346 3790
rect 5380 3756 5396 3790
rect 5330 3740 5396 3756
rect 5522 3790 5588 3806
rect 5636 3802 5666 3828
rect 5732 3806 5762 3828
rect 5522 3756 5538 3790
rect 5572 3756 5588 3790
rect 5522 3740 5588 3756
rect 5714 3790 5780 3806
rect 5828 3802 5858 3828
rect 5924 3806 5954 3828
rect 5714 3756 5730 3790
rect 5764 3756 5780 3790
rect 5714 3740 5780 3756
rect 5906 3790 5972 3806
rect 6020 3802 6050 3828
rect 6116 3806 6146 3828
rect 5906 3756 5922 3790
rect 5956 3756 5972 3790
rect 5906 3740 5972 3756
rect 6098 3790 6164 3806
rect 6212 3802 6242 3828
rect 6308 3806 6338 3828
rect 6098 3756 6114 3790
rect 6148 3756 6164 3790
rect 6098 3740 6164 3756
rect 6290 3790 6356 3806
rect 6404 3802 6434 3828
rect 6500 3806 6530 3828
rect 6290 3756 6306 3790
rect 6340 3756 6356 3790
rect 6290 3740 6356 3756
rect 6482 3790 6548 3806
rect 6596 3802 6626 3828
rect 6692 3806 6722 3828
rect 6482 3756 6498 3790
rect 6532 3756 6548 3790
rect 6482 3740 6548 3756
rect 6674 3790 6740 3806
rect 6788 3802 6818 3828
rect 6884 3806 6914 3828
rect 6674 3756 6690 3790
rect 6724 3756 6740 3790
rect 6674 3740 6740 3756
rect 6866 3790 6932 3806
rect 6980 3802 7010 3828
rect 7076 3806 7106 3828
rect 6866 3756 6882 3790
rect 6916 3756 6932 3790
rect 6866 3740 6932 3756
rect 7058 3790 7124 3806
rect 7172 3802 7202 3828
rect 7268 3806 7298 3828
rect 7058 3756 7074 3790
rect 7108 3756 7124 3790
rect 7058 3740 7124 3756
rect 7250 3790 7316 3806
rect 7250 3756 7266 3790
rect 7300 3756 7316 3790
rect 7250 3740 7316 3756
rect 4562 3682 4628 3698
rect 4562 3648 4578 3682
rect 4612 3648 4628 3682
rect 4484 3610 4514 3636
rect 4562 3632 4628 3648
rect 4754 3682 4820 3698
rect 4754 3648 4770 3682
rect 4804 3648 4820 3682
rect 4580 3610 4610 3632
rect 4676 3610 4706 3636
rect 4754 3632 4820 3648
rect 4946 3682 5012 3698
rect 4946 3648 4962 3682
rect 4996 3648 5012 3682
rect 4772 3610 4802 3632
rect 4868 3610 4898 3636
rect 4946 3632 5012 3648
rect 5138 3682 5204 3698
rect 5138 3648 5154 3682
rect 5188 3648 5204 3682
rect 4964 3610 4994 3632
rect 5060 3610 5090 3636
rect 5138 3632 5204 3648
rect 5330 3682 5396 3698
rect 5330 3648 5346 3682
rect 5380 3648 5396 3682
rect 5156 3610 5186 3632
rect 5252 3610 5282 3636
rect 5330 3632 5396 3648
rect 5522 3682 5588 3698
rect 5522 3648 5538 3682
rect 5572 3648 5588 3682
rect 5348 3610 5378 3632
rect 5444 3610 5474 3636
rect 5522 3632 5588 3648
rect 5714 3682 5780 3698
rect 5714 3648 5730 3682
rect 5764 3648 5780 3682
rect 5540 3610 5570 3632
rect 5636 3610 5666 3636
rect 5714 3632 5780 3648
rect 5906 3682 5972 3698
rect 5906 3648 5922 3682
rect 5956 3648 5972 3682
rect 5732 3610 5762 3632
rect 5828 3610 5858 3636
rect 5906 3632 5972 3648
rect 6098 3682 6164 3698
rect 6098 3648 6114 3682
rect 6148 3648 6164 3682
rect 5924 3610 5954 3632
rect 6020 3610 6050 3636
rect 6098 3632 6164 3648
rect 6290 3682 6356 3698
rect 6290 3648 6306 3682
rect 6340 3648 6356 3682
rect 6116 3610 6146 3632
rect 6212 3610 6242 3636
rect 6290 3632 6356 3648
rect 6482 3682 6548 3698
rect 6482 3648 6498 3682
rect 6532 3648 6548 3682
rect 6308 3610 6338 3632
rect 6404 3610 6434 3636
rect 6482 3632 6548 3648
rect 6674 3682 6740 3698
rect 6674 3648 6690 3682
rect 6724 3648 6740 3682
rect 6500 3610 6530 3632
rect 6596 3610 6626 3636
rect 6674 3632 6740 3648
rect 6866 3682 6932 3698
rect 6866 3648 6882 3682
rect 6916 3648 6932 3682
rect 6692 3610 6722 3632
rect 6788 3610 6818 3636
rect 6866 3632 6932 3648
rect 7058 3682 7124 3698
rect 7058 3648 7074 3682
rect 7108 3648 7124 3682
rect 6884 3610 6914 3632
rect 6980 3610 7010 3636
rect 7058 3632 7124 3648
rect 7250 3682 7316 3698
rect 7250 3648 7266 3682
rect 7300 3648 7316 3682
rect 7076 3610 7106 3632
rect 7172 3610 7202 3636
rect 7250 3632 7316 3648
rect 7268 3610 7298 3632
rect 4484 3188 4514 3210
rect 4466 3172 4532 3188
rect 4580 3184 4610 3210
rect 4676 3188 4706 3210
rect 4466 3138 4482 3172
rect 4516 3138 4532 3172
rect 4466 3122 4532 3138
rect 4658 3172 4724 3188
rect 4772 3184 4802 3210
rect 4868 3188 4898 3210
rect 4658 3138 4674 3172
rect 4708 3138 4724 3172
rect 4658 3122 4724 3138
rect 4850 3172 4916 3188
rect 4964 3184 4994 3210
rect 5060 3188 5090 3210
rect 4850 3138 4866 3172
rect 4900 3138 4916 3172
rect 4850 3122 4916 3138
rect 5042 3172 5108 3188
rect 5156 3184 5186 3210
rect 5252 3188 5282 3210
rect 5042 3138 5058 3172
rect 5092 3138 5108 3172
rect 5042 3122 5108 3138
rect 5234 3172 5300 3188
rect 5348 3184 5378 3210
rect 5444 3188 5474 3210
rect 5234 3138 5250 3172
rect 5284 3138 5300 3172
rect 5234 3122 5300 3138
rect 5426 3172 5492 3188
rect 5540 3184 5570 3210
rect 5636 3188 5666 3210
rect 5426 3138 5442 3172
rect 5476 3138 5492 3172
rect 5426 3122 5492 3138
rect 5618 3172 5684 3188
rect 5732 3184 5762 3210
rect 5828 3188 5858 3210
rect 5618 3138 5634 3172
rect 5668 3138 5684 3172
rect 5618 3122 5684 3138
rect 5810 3172 5876 3188
rect 5924 3184 5954 3210
rect 6020 3188 6050 3210
rect 5810 3138 5826 3172
rect 5860 3138 5876 3172
rect 5810 3122 5876 3138
rect 6002 3172 6068 3188
rect 6116 3184 6146 3210
rect 6212 3188 6242 3210
rect 6002 3138 6018 3172
rect 6052 3138 6068 3172
rect 6002 3122 6068 3138
rect 6194 3172 6260 3188
rect 6308 3184 6338 3210
rect 6404 3188 6434 3210
rect 6194 3138 6210 3172
rect 6244 3138 6260 3172
rect 6194 3122 6260 3138
rect 6386 3172 6452 3188
rect 6500 3184 6530 3210
rect 6596 3188 6626 3210
rect 6386 3138 6402 3172
rect 6436 3138 6452 3172
rect 6386 3122 6452 3138
rect 6578 3172 6644 3188
rect 6692 3184 6722 3210
rect 6788 3188 6818 3210
rect 6578 3138 6594 3172
rect 6628 3138 6644 3172
rect 6578 3122 6644 3138
rect 6770 3172 6836 3188
rect 6884 3184 6914 3210
rect 6980 3188 7010 3210
rect 6770 3138 6786 3172
rect 6820 3138 6836 3172
rect 6770 3122 6836 3138
rect 6962 3172 7028 3188
rect 7076 3184 7106 3210
rect 7172 3188 7202 3210
rect 6962 3138 6978 3172
rect 7012 3138 7028 3172
rect 6962 3122 7028 3138
rect 7154 3172 7220 3188
rect 7268 3184 7298 3210
rect 7154 3138 7170 3172
rect 7204 3138 7220 3172
rect 7154 3122 7220 3138
rect 8106 5536 8172 5552
rect 8106 5502 8122 5536
rect 8156 5502 8172 5536
rect 8106 5486 8172 5502
rect 8298 5536 8364 5552
rect 8298 5502 8314 5536
rect 8348 5502 8364 5536
rect 8124 5464 8154 5486
rect 8220 5464 8250 5490
rect 8298 5486 8364 5502
rect 8490 5536 8556 5552
rect 8490 5502 8506 5536
rect 8540 5502 8556 5536
rect 8316 5464 8346 5486
rect 8412 5464 8442 5490
rect 8490 5486 8556 5502
rect 8682 5536 8748 5552
rect 8682 5502 8698 5536
rect 8732 5502 8748 5536
rect 8508 5464 8538 5486
rect 8604 5464 8634 5490
rect 8682 5486 8748 5502
rect 8874 5536 8940 5552
rect 8874 5502 8890 5536
rect 8924 5502 8940 5536
rect 8700 5464 8730 5486
rect 8796 5464 8826 5490
rect 8874 5486 8940 5502
rect 9066 5536 9132 5552
rect 9066 5502 9082 5536
rect 9116 5502 9132 5536
rect 8892 5464 8922 5486
rect 8988 5464 9018 5490
rect 9066 5486 9132 5502
rect 9258 5536 9324 5552
rect 9258 5502 9274 5536
rect 9308 5502 9324 5536
rect 9084 5464 9114 5486
rect 9180 5464 9210 5490
rect 9258 5486 9324 5502
rect 9450 5536 9516 5552
rect 9450 5502 9466 5536
rect 9500 5502 9516 5536
rect 9276 5464 9306 5486
rect 9372 5464 9402 5490
rect 9450 5486 9516 5502
rect 9642 5536 9708 5552
rect 9642 5502 9658 5536
rect 9692 5502 9708 5536
rect 9468 5464 9498 5486
rect 9564 5464 9594 5490
rect 9642 5486 9708 5502
rect 9834 5536 9900 5552
rect 9834 5502 9850 5536
rect 9884 5502 9900 5536
rect 9660 5464 9690 5486
rect 9756 5464 9786 5490
rect 9834 5486 9900 5502
rect 10026 5536 10092 5552
rect 10026 5502 10042 5536
rect 10076 5502 10092 5536
rect 9852 5464 9882 5486
rect 9948 5464 9978 5490
rect 10026 5486 10092 5502
rect 10218 5536 10284 5552
rect 10218 5502 10234 5536
rect 10268 5502 10284 5536
rect 10044 5464 10074 5486
rect 10140 5464 10170 5490
rect 10218 5486 10284 5502
rect 10410 5536 10476 5552
rect 10410 5502 10426 5536
rect 10460 5502 10476 5536
rect 10236 5464 10266 5486
rect 10332 5464 10362 5490
rect 10410 5486 10476 5502
rect 10602 5536 10668 5552
rect 10602 5502 10618 5536
rect 10652 5502 10668 5536
rect 10428 5464 10458 5486
rect 10524 5464 10554 5490
rect 10602 5486 10668 5502
rect 10794 5536 10860 5552
rect 10794 5502 10810 5536
rect 10844 5502 10860 5536
rect 10620 5464 10650 5486
rect 10716 5464 10746 5490
rect 10794 5486 10860 5502
rect 10812 5464 10842 5486
rect 10908 5464 10938 5490
rect 8124 5038 8154 5064
rect 8220 5042 8250 5064
rect 8202 5026 8268 5042
rect 8316 5038 8346 5064
rect 8412 5042 8442 5064
rect 8202 4992 8218 5026
rect 8252 4992 8268 5026
rect 8202 4976 8268 4992
rect 8394 5026 8460 5042
rect 8508 5038 8538 5064
rect 8604 5042 8634 5064
rect 8394 4992 8410 5026
rect 8444 4992 8460 5026
rect 8394 4976 8460 4992
rect 8586 5026 8652 5042
rect 8700 5038 8730 5064
rect 8796 5042 8826 5064
rect 8586 4992 8602 5026
rect 8636 4992 8652 5026
rect 8586 4976 8652 4992
rect 8778 5026 8844 5042
rect 8892 5038 8922 5064
rect 8988 5042 9018 5064
rect 8778 4992 8794 5026
rect 8828 4992 8844 5026
rect 8778 4976 8844 4992
rect 8970 5026 9036 5042
rect 9084 5038 9114 5064
rect 9180 5042 9210 5064
rect 8970 4992 8986 5026
rect 9020 4992 9036 5026
rect 8970 4976 9036 4992
rect 9162 5026 9228 5042
rect 9276 5038 9306 5064
rect 9372 5042 9402 5064
rect 9162 4992 9178 5026
rect 9212 4992 9228 5026
rect 9162 4976 9228 4992
rect 9354 5026 9420 5042
rect 9468 5038 9498 5064
rect 9564 5042 9594 5064
rect 9354 4992 9370 5026
rect 9404 4992 9420 5026
rect 9354 4976 9420 4992
rect 9546 5026 9612 5042
rect 9660 5038 9690 5064
rect 9756 5042 9786 5064
rect 9546 4992 9562 5026
rect 9596 4992 9612 5026
rect 9546 4976 9612 4992
rect 9738 5026 9804 5042
rect 9852 5038 9882 5064
rect 9948 5042 9978 5064
rect 9738 4992 9754 5026
rect 9788 4992 9804 5026
rect 9738 4976 9804 4992
rect 9930 5026 9996 5042
rect 10044 5038 10074 5064
rect 10140 5042 10170 5064
rect 9930 4992 9946 5026
rect 9980 4992 9996 5026
rect 9930 4976 9996 4992
rect 10122 5026 10188 5042
rect 10236 5038 10266 5064
rect 10332 5042 10362 5064
rect 10122 4992 10138 5026
rect 10172 4992 10188 5026
rect 10122 4976 10188 4992
rect 10314 5026 10380 5042
rect 10428 5038 10458 5064
rect 10524 5042 10554 5064
rect 10314 4992 10330 5026
rect 10364 4992 10380 5026
rect 10314 4976 10380 4992
rect 10506 5026 10572 5042
rect 10620 5038 10650 5064
rect 10716 5042 10746 5064
rect 10506 4992 10522 5026
rect 10556 4992 10572 5026
rect 10506 4976 10572 4992
rect 10698 5026 10764 5042
rect 10812 5038 10842 5064
rect 10908 5042 10938 5064
rect 10698 4992 10714 5026
rect 10748 4992 10764 5026
rect 10698 4976 10764 4992
rect 10890 5026 10956 5042
rect 10890 4992 10906 5026
rect 10940 4992 10956 5026
rect 10890 4976 10956 4992
rect 8202 4918 8268 4934
rect 8202 4884 8218 4918
rect 8252 4884 8268 4918
rect 8124 4846 8154 4872
rect 8202 4868 8268 4884
rect 8394 4918 8460 4934
rect 8394 4884 8410 4918
rect 8444 4884 8460 4918
rect 8220 4846 8250 4868
rect 8316 4846 8346 4872
rect 8394 4868 8460 4884
rect 8586 4918 8652 4934
rect 8586 4884 8602 4918
rect 8636 4884 8652 4918
rect 8412 4846 8442 4868
rect 8508 4846 8538 4872
rect 8586 4868 8652 4884
rect 8778 4918 8844 4934
rect 8778 4884 8794 4918
rect 8828 4884 8844 4918
rect 8604 4846 8634 4868
rect 8700 4846 8730 4872
rect 8778 4868 8844 4884
rect 8970 4918 9036 4934
rect 8970 4884 8986 4918
rect 9020 4884 9036 4918
rect 8796 4846 8826 4868
rect 8892 4846 8922 4872
rect 8970 4868 9036 4884
rect 9162 4918 9228 4934
rect 9162 4884 9178 4918
rect 9212 4884 9228 4918
rect 8988 4846 9018 4868
rect 9084 4846 9114 4872
rect 9162 4868 9228 4884
rect 9354 4918 9420 4934
rect 9354 4884 9370 4918
rect 9404 4884 9420 4918
rect 9180 4846 9210 4868
rect 9276 4846 9306 4872
rect 9354 4868 9420 4884
rect 9546 4918 9612 4934
rect 9546 4884 9562 4918
rect 9596 4884 9612 4918
rect 9372 4846 9402 4868
rect 9468 4846 9498 4872
rect 9546 4868 9612 4884
rect 9738 4918 9804 4934
rect 9738 4884 9754 4918
rect 9788 4884 9804 4918
rect 9564 4846 9594 4868
rect 9660 4846 9690 4872
rect 9738 4868 9804 4884
rect 9930 4918 9996 4934
rect 9930 4884 9946 4918
rect 9980 4884 9996 4918
rect 9756 4846 9786 4868
rect 9852 4846 9882 4872
rect 9930 4868 9996 4884
rect 10122 4918 10188 4934
rect 10122 4884 10138 4918
rect 10172 4884 10188 4918
rect 9948 4846 9978 4868
rect 10044 4846 10074 4872
rect 10122 4868 10188 4884
rect 10314 4918 10380 4934
rect 10314 4884 10330 4918
rect 10364 4884 10380 4918
rect 10140 4846 10170 4868
rect 10236 4846 10266 4872
rect 10314 4868 10380 4884
rect 10506 4918 10572 4934
rect 10506 4884 10522 4918
rect 10556 4884 10572 4918
rect 10332 4846 10362 4868
rect 10428 4846 10458 4872
rect 10506 4868 10572 4884
rect 10698 4918 10764 4934
rect 10698 4884 10714 4918
rect 10748 4884 10764 4918
rect 10524 4846 10554 4868
rect 10620 4846 10650 4872
rect 10698 4868 10764 4884
rect 10890 4918 10956 4934
rect 10890 4884 10906 4918
rect 10940 4884 10956 4918
rect 10716 4846 10746 4868
rect 10812 4846 10842 4872
rect 10890 4868 10956 4884
rect 10908 4846 10938 4868
rect 8124 4424 8154 4446
rect 8106 4408 8172 4424
rect 8220 4420 8250 4446
rect 8316 4424 8346 4446
rect 8106 4374 8122 4408
rect 8156 4374 8172 4408
rect 8106 4358 8172 4374
rect 8298 4408 8364 4424
rect 8412 4420 8442 4446
rect 8508 4424 8538 4446
rect 8298 4374 8314 4408
rect 8348 4374 8364 4408
rect 8298 4358 8364 4374
rect 8490 4408 8556 4424
rect 8604 4420 8634 4446
rect 8700 4424 8730 4446
rect 8490 4374 8506 4408
rect 8540 4374 8556 4408
rect 8490 4358 8556 4374
rect 8682 4408 8748 4424
rect 8796 4420 8826 4446
rect 8892 4424 8922 4446
rect 8682 4374 8698 4408
rect 8732 4374 8748 4408
rect 8682 4358 8748 4374
rect 8874 4408 8940 4424
rect 8988 4420 9018 4446
rect 9084 4424 9114 4446
rect 8874 4374 8890 4408
rect 8924 4374 8940 4408
rect 8874 4358 8940 4374
rect 9066 4408 9132 4424
rect 9180 4420 9210 4446
rect 9276 4424 9306 4446
rect 9066 4374 9082 4408
rect 9116 4374 9132 4408
rect 9066 4358 9132 4374
rect 9258 4408 9324 4424
rect 9372 4420 9402 4446
rect 9468 4424 9498 4446
rect 9258 4374 9274 4408
rect 9308 4374 9324 4408
rect 9258 4358 9324 4374
rect 9450 4408 9516 4424
rect 9564 4420 9594 4446
rect 9660 4424 9690 4446
rect 9450 4374 9466 4408
rect 9500 4374 9516 4408
rect 9450 4358 9516 4374
rect 9642 4408 9708 4424
rect 9756 4420 9786 4446
rect 9852 4424 9882 4446
rect 9642 4374 9658 4408
rect 9692 4374 9708 4408
rect 9642 4358 9708 4374
rect 9834 4408 9900 4424
rect 9948 4420 9978 4446
rect 10044 4424 10074 4446
rect 9834 4374 9850 4408
rect 9884 4374 9900 4408
rect 9834 4358 9900 4374
rect 10026 4408 10092 4424
rect 10140 4420 10170 4446
rect 10236 4424 10266 4446
rect 10026 4374 10042 4408
rect 10076 4374 10092 4408
rect 10026 4358 10092 4374
rect 10218 4408 10284 4424
rect 10332 4420 10362 4446
rect 10428 4424 10458 4446
rect 10218 4374 10234 4408
rect 10268 4374 10284 4408
rect 10218 4358 10284 4374
rect 10410 4408 10476 4424
rect 10524 4420 10554 4446
rect 10620 4424 10650 4446
rect 10410 4374 10426 4408
rect 10460 4374 10476 4408
rect 10410 4358 10476 4374
rect 10602 4408 10668 4424
rect 10716 4420 10746 4446
rect 10812 4424 10842 4446
rect 10602 4374 10618 4408
rect 10652 4374 10668 4408
rect 10602 4358 10668 4374
rect 10794 4408 10860 4424
rect 10908 4420 10938 4446
rect 10794 4374 10810 4408
rect 10844 4374 10860 4408
rect 10794 4358 10860 4374
rect 8106 4300 8172 4316
rect 8106 4266 8122 4300
rect 8156 4266 8172 4300
rect 8106 4250 8172 4266
rect 8298 4300 8364 4316
rect 8298 4266 8314 4300
rect 8348 4266 8364 4300
rect 8124 4228 8154 4250
rect 8220 4228 8250 4254
rect 8298 4250 8364 4266
rect 8490 4300 8556 4316
rect 8490 4266 8506 4300
rect 8540 4266 8556 4300
rect 8316 4228 8346 4250
rect 8412 4228 8442 4254
rect 8490 4250 8556 4266
rect 8682 4300 8748 4316
rect 8682 4266 8698 4300
rect 8732 4266 8748 4300
rect 8508 4228 8538 4250
rect 8604 4228 8634 4254
rect 8682 4250 8748 4266
rect 8874 4300 8940 4316
rect 8874 4266 8890 4300
rect 8924 4266 8940 4300
rect 8700 4228 8730 4250
rect 8796 4228 8826 4254
rect 8874 4250 8940 4266
rect 9066 4300 9132 4316
rect 9066 4266 9082 4300
rect 9116 4266 9132 4300
rect 8892 4228 8922 4250
rect 8988 4228 9018 4254
rect 9066 4250 9132 4266
rect 9258 4300 9324 4316
rect 9258 4266 9274 4300
rect 9308 4266 9324 4300
rect 9084 4228 9114 4250
rect 9180 4228 9210 4254
rect 9258 4250 9324 4266
rect 9450 4300 9516 4316
rect 9450 4266 9466 4300
rect 9500 4266 9516 4300
rect 9276 4228 9306 4250
rect 9372 4228 9402 4254
rect 9450 4250 9516 4266
rect 9642 4300 9708 4316
rect 9642 4266 9658 4300
rect 9692 4266 9708 4300
rect 9468 4228 9498 4250
rect 9564 4228 9594 4254
rect 9642 4250 9708 4266
rect 9834 4300 9900 4316
rect 9834 4266 9850 4300
rect 9884 4266 9900 4300
rect 9660 4228 9690 4250
rect 9756 4228 9786 4254
rect 9834 4250 9900 4266
rect 10026 4300 10092 4316
rect 10026 4266 10042 4300
rect 10076 4266 10092 4300
rect 9852 4228 9882 4250
rect 9948 4228 9978 4254
rect 10026 4250 10092 4266
rect 10218 4300 10284 4316
rect 10218 4266 10234 4300
rect 10268 4266 10284 4300
rect 10044 4228 10074 4250
rect 10140 4228 10170 4254
rect 10218 4250 10284 4266
rect 10410 4300 10476 4316
rect 10410 4266 10426 4300
rect 10460 4266 10476 4300
rect 10236 4228 10266 4250
rect 10332 4228 10362 4254
rect 10410 4250 10476 4266
rect 10602 4300 10668 4316
rect 10602 4266 10618 4300
rect 10652 4266 10668 4300
rect 10428 4228 10458 4250
rect 10524 4228 10554 4254
rect 10602 4250 10668 4266
rect 10794 4300 10860 4316
rect 10794 4266 10810 4300
rect 10844 4266 10860 4300
rect 10620 4228 10650 4250
rect 10716 4228 10746 4254
rect 10794 4250 10860 4266
rect 10812 4228 10842 4250
rect 10908 4228 10938 4254
rect 8124 3802 8154 3828
rect 8220 3806 8250 3828
rect 8202 3790 8268 3806
rect 8316 3802 8346 3828
rect 8412 3806 8442 3828
rect 8202 3756 8218 3790
rect 8252 3756 8268 3790
rect 8202 3740 8268 3756
rect 8394 3790 8460 3806
rect 8508 3802 8538 3828
rect 8604 3806 8634 3828
rect 8394 3756 8410 3790
rect 8444 3756 8460 3790
rect 8394 3740 8460 3756
rect 8586 3790 8652 3806
rect 8700 3802 8730 3828
rect 8796 3806 8826 3828
rect 8586 3756 8602 3790
rect 8636 3756 8652 3790
rect 8586 3740 8652 3756
rect 8778 3790 8844 3806
rect 8892 3802 8922 3828
rect 8988 3806 9018 3828
rect 8778 3756 8794 3790
rect 8828 3756 8844 3790
rect 8778 3740 8844 3756
rect 8970 3790 9036 3806
rect 9084 3802 9114 3828
rect 9180 3806 9210 3828
rect 8970 3756 8986 3790
rect 9020 3756 9036 3790
rect 8970 3740 9036 3756
rect 9162 3790 9228 3806
rect 9276 3802 9306 3828
rect 9372 3806 9402 3828
rect 9162 3756 9178 3790
rect 9212 3756 9228 3790
rect 9162 3740 9228 3756
rect 9354 3790 9420 3806
rect 9468 3802 9498 3828
rect 9564 3806 9594 3828
rect 9354 3756 9370 3790
rect 9404 3756 9420 3790
rect 9354 3740 9420 3756
rect 9546 3790 9612 3806
rect 9660 3802 9690 3828
rect 9756 3806 9786 3828
rect 9546 3756 9562 3790
rect 9596 3756 9612 3790
rect 9546 3740 9612 3756
rect 9738 3790 9804 3806
rect 9852 3802 9882 3828
rect 9948 3806 9978 3828
rect 9738 3756 9754 3790
rect 9788 3756 9804 3790
rect 9738 3740 9804 3756
rect 9930 3790 9996 3806
rect 10044 3802 10074 3828
rect 10140 3806 10170 3828
rect 9930 3756 9946 3790
rect 9980 3756 9996 3790
rect 9930 3740 9996 3756
rect 10122 3790 10188 3806
rect 10236 3802 10266 3828
rect 10332 3806 10362 3828
rect 10122 3756 10138 3790
rect 10172 3756 10188 3790
rect 10122 3740 10188 3756
rect 10314 3790 10380 3806
rect 10428 3802 10458 3828
rect 10524 3806 10554 3828
rect 10314 3756 10330 3790
rect 10364 3756 10380 3790
rect 10314 3740 10380 3756
rect 10506 3790 10572 3806
rect 10620 3802 10650 3828
rect 10716 3806 10746 3828
rect 10506 3756 10522 3790
rect 10556 3756 10572 3790
rect 10506 3740 10572 3756
rect 10698 3790 10764 3806
rect 10812 3802 10842 3828
rect 10908 3806 10938 3828
rect 10698 3756 10714 3790
rect 10748 3756 10764 3790
rect 10698 3740 10764 3756
rect 10890 3790 10956 3806
rect 10890 3756 10906 3790
rect 10940 3756 10956 3790
rect 10890 3740 10956 3756
rect 8202 3682 8268 3698
rect 8202 3648 8218 3682
rect 8252 3648 8268 3682
rect 8124 3610 8154 3636
rect 8202 3632 8268 3648
rect 8394 3682 8460 3698
rect 8394 3648 8410 3682
rect 8444 3648 8460 3682
rect 8220 3610 8250 3632
rect 8316 3610 8346 3636
rect 8394 3632 8460 3648
rect 8586 3682 8652 3698
rect 8586 3648 8602 3682
rect 8636 3648 8652 3682
rect 8412 3610 8442 3632
rect 8508 3610 8538 3636
rect 8586 3632 8652 3648
rect 8778 3682 8844 3698
rect 8778 3648 8794 3682
rect 8828 3648 8844 3682
rect 8604 3610 8634 3632
rect 8700 3610 8730 3636
rect 8778 3632 8844 3648
rect 8970 3682 9036 3698
rect 8970 3648 8986 3682
rect 9020 3648 9036 3682
rect 8796 3610 8826 3632
rect 8892 3610 8922 3636
rect 8970 3632 9036 3648
rect 9162 3682 9228 3698
rect 9162 3648 9178 3682
rect 9212 3648 9228 3682
rect 8988 3610 9018 3632
rect 9084 3610 9114 3636
rect 9162 3632 9228 3648
rect 9354 3682 9420 3698
rect 9354 3648 9370 3682
rect 9404 3648 9420 3682
rect 9180 3610 9210 3632
rect 9276 3610 9306 3636
rect 9354 3632 9420 3648
rect 9546 3682 9612 3698
rect 9546 3648 9562 3682
rect 9596 3648 9612 3682
rect 9372 3610 9402 3632
rect 9468 3610 9498 3636
rect 9546 3632 9612 3648
rect 9738 3682 9804 3698
rect 9738 3648 9754 3682
rect 9788 3648 9804 3682
rect 9564 3610 9594 3632
rect 9660 3610 9690 3636
rect 9738 3632 9804 3648
rect 9930 3682 9996 3698
rect 9930 3648 9946 3682
rect 9980 3648 9996 3682
rect 9756 3610 9786 3632
rect 9852 3610 9882 3636
rect 9930 3632 9996 3648
rect 10122 3682 10188 3698
rect 10122 3648 10138 3682
rect 10172 3648 10188 3682
rect 9948 3610 9978 3632
rect 10044 3610 10074 3636
rect 10122 3632 10188 3648
rect 10314 3682 10380 3698
rect 10314 3648 10330 3682
rect 10364 3648 10380 3682
rect 10140 3610 10170 3632
rect 10236 3610 10266 3636
rect 10314 3632 10380 3648
rect 10506 3682 10572 3698
rect 10506 3648 10522 3682
rect 10556 3648 10572 3682
rect 10332 3610 10362 3632
rect 10428 3610 10458 3636
rect 10506 3632 10572 3648
rect 10698 3682 10764 3698
rect 10698 3648 10714 3682
rect 10748 3648 10764 3682
rect 10524 3610 10554 3632
rect 10620 3610 10650 3636
rect 10698 3632 10764 3648
rect 10890 3682 10956 3698
rect 10890 3648 10906 3682
rect 10940 3648 10956 3682
rect 10716 3610 10746 3632
rect 10812 3610 10842 3636
rect 10890 3632 10956 3648
rect 10908 3610 10938 3632
rect 8124 3188 8154 3210
rect 8106 3172 8172 3188
rect 8220 3184 8250 3210
rect 8316 3188 8346 3210
rect 8106 3138 8122 3172
rect 8156 3138 8172 3172
rect 8106 3122 8172 3138
rect 8298 3172 8364 3188
rect 8412 3184 8442 3210
rect 8508 3188 8538 3210
rect 8298 3138 8314 3172
rect 8348 3138 8364 3172
rect 8298 3122 8364 3138
rect 8490 3172 8556 3188
rect 8604 3184 8634 3210
rect 8700 3188 8730 3210
rect 8490 3138 8506 3172
rect 8540 3138 8556 3172
rect 8490 3122 8556 3138
rect 8682 3172 8748 3188
rect 8796 3184 8826 3210
rect 8892 3188 8922 3210
rect 8682 3138 8698 3172
rect 8732 3138 8748 3172
rect 8682 3122 8748 3138
rect 8874 3172 8940 3188
rect 8988 3184 9018 3210
rect 9084 3188 9114 3210
rect 8874 3138 8890 3172
rect 8924 3138 8940 3172
rect 8874 3122 8940 3138
rect 9066 3172 9132 3188
rect 9180 3184 9210 3210
rect 9276 3188 9306 3210
rect 9066 3138 9082 3172
rect 9116 3138 9132 3172
rect 9066 3122 9132 3138
rect 9258 3172 9324 3188
rect 9372 3184 9402 3210
rect 9468 3188 9498 3210
rect 9258 3138 9274 3172
rect 9308 3138 9324 3172
rect 9258 3122 9324 3138
rect 9450 3172 9516 3188
rect 9564 3184 9594 3210
rect 9660 3188 9690 3210
rect 9450 3138 9466 3172
rect 9500 3138 9516 3172
rect 9450 3122 9516 3138
rect 9642 3172 9708 3188
rect 9756 3184 9786 3210
rect 9852 3188 9882 3210
rect 9642 3138 9658 3172
rect 9692 3138 9708 3172
rect 9642 3122 9708 3138
rect 9834 3172 9900 3188
rect 9948 3184 9978 3210
rect 10044 3188 10074 3210
rect 9834 3138 9850 3172
rect 9884 3138 9900 3172
rect 9834 3122 9900 3138
rect 10026 3172 10092 3188
rect 10140 3184 10170 3210
rect 10236 3188 10266 3210
rect 10026 3138 10042 3172
rect 10076 3138 10092 3172
rect 10026 3122 10092 3138
rect 10218 3172 10284 3188
rect 10332 3184 10362 3210
rect 10428 3188 10458 3210
rect 10218 3138 10234 3172
rect 10268 3138 10284 3172
rect 10218 3122 10284 3138
rect 10410 3172 10476 3188
rect 10524 3184 10554 3210
rect 10620 3188 10650 3210
rect 10410 3138 10426 3172
rect 10460 3138 10476 3172
rect 10410 3122 10476 3138
rect 10602 3172 10668 3188
rect 10716 3184 10746 3210
rect 10812 3188 10842 3210
rect 10602 3138 10618 3172
rect 10652 3138 10668 3172
rect 10602 3122 10668 3138
rect 10794 3172 10860 3188
rect 10908 3184 10938 3210
rect 10794 3138 10810 3172
rect 10844 3138 10860 3172
rect 10794 3122 10860 3138
rect 12086 5536 12152 5552
rect 12086 5502 12102 5536
rect 12136 5502 12152 5536
rect 12086 5486 12152 5502
rect 12278 5536 12344 5552
rect 12278 5502 12294 5536
rect 12328 5502 12344 5536
rect 12104 5464 12134 5486
rect 12200 5464 12230 5490
rect 12278 5486 12344 5502
rect 12470 5536 12536 5552
rect 12470 5502 12486 5536
rect 12520 5502 12536 5536
rect 12296 5464 12326 5486
rect 12392 5464 12422 5490
rect 12470 5486 12536 5502
rect 12662 5536 12728 5552
rect 12662 5502 12678 5536
rect 12712 5502 12728 5536
rect 12488 5464 12518 5486
rect 12584 5464 12614 5490
rect 12662 5486 12728 5502
rect 12854 5536 12920 5552
rect 12854 5502 12870 5536
rect 12904 5502 12920 5536
rect 12680 5464 12710 5486
rect 12776 5464 12806 5490
rect 12854 5486 12920 5502
rect 13046 5536 13112 5552
rect 13046 5502 13062 5536
rect 13096 5502 13112 5536
rect 12872 5464 12902 5486
rect 12968 5464 12998 5490
rect 13046 5486 13112 5502
rect 13238 5536 13304 5552
rect 13238 5502 13254 5536
rect 13288 5502 13304 5536
rect 13064 5464 13094 5486
rect 13160 5464 13190 5490
rect 13238 5486 13304 5502
rect 13430 5536 13496 5552
rect 13430 5502 13446 5536
rect 13480 5502 13496 5536
rect 13256 5464 13286 5486
rect 13352 5464 13382 5490
rect 13430 5486 13496 5502
rect 13622 5536 13688 5552
rect 13622 5502 13638 5536
rect 13672 5502 13688 5536
rect 13448 5464 13478 5486
rect 13544 5464 13574 5490
rect 13622 5486 13688 5502
rect 13814 5536 13880 5552
rect 13814 5502 13830 5536
rect 13864 5502 13880 5536
rect 13640 5464 13670 5486
rect 13736 5464 13766 5490
rect 13814 5486 13880 5502
rect 14006 5536 14072 5552
rect 14006 5502 14022 5536
rect 14056 5502 14072 5536
rect 13832 5464 13862 5486
rect 13928 5464 13958 5490
rect 14006 5486 14072 5502
rect 14198 5536 14264 5552
rect 14198 5502 14214 5536
rect 14248 5502 14264 5536
rect 14024 5464 14054 5486
rect 14120 5464 14150 5490
rect 14198 5486 14264 5502
rect 14390 5536 14456 5552
rect 14390 5502 14406 5536
rect 14440 5502 14456 5536
rect 14216 5464 14246 5486
rect 14312 5464 14342 5490
rect 14390 5486 14456 5502
rect 14582 5536 14648 5552
rect 14582 5502 14598 5536
rect 14632 5502 14648 5536
rect 14408 5464 14438 5486
rect 14504 5464 14534 5490
rect 14582 5486 14648 5502
rect 14774 5536 14840 5552
rect 14774 5502 14790 5536
rect 14824 5502 14840 5536
rect 14600 5464 14630 5486
rect 14696 5464 14726 5490
rect 14774 5486 14840 5502
rect 14792 5464 14822 5486
rect 14888 5464 14918 5490
rect 12104 5038 12134 5064
rect 12200 5042 12230 5064
rect 12182 5026 12248 5042
rect 12296 5038 12326 5064
rect 12392 5042 12422 5064
rect 12182 4992 12198 5026
rect 12232 4992 12248 5026
rect 12182 4976 12248 4992
rect 12374 5026 12440 5042
rect 12488 5038 12518 5064
rect 12584 5042 12614 5064
rect 12374 4992 12390 5026
rect 12424 4992 12440 5026
rect 12374 4976 12440 4992
rect 12566 5026 12632 5042
rect 12680 5038 12710 5064
rect 12776 5042 12806 5064
rect 12566 4992 12582 5026
rect 12616 4992 12632 5026
rect 12566 4976 12632 4992
rect 12758 5026 12824 5042
rect 12872 5038 12902 5064
rect 12968 5042 12998 5064
rect 12758 4992 12774 5026
rect 12808 4992 12824 5026
rect 12758 4976 12824 4992
rect 12950 5026 13016 5042
rect 13064 5038 13094 5064
rect 13160 5042 13190 5064
rect 12950 4992 12966 5026
rect 13000 4992 13016 5026
rect 12950 4976 13016 4992
rect 13142 5026 13208 5042
rect 13256 5038 13286 5064
rect 13352 5042 13382 5064
rect 13142 4992 13158 5026
rect 13192 4992 13208 5026
rect 13142 4976 13208 4992
rect 13334 5026 13400 5042
rect 13448 5038 13478 5064
rect 13544 5042 13574 5064
rect 13334 4992 13350 5026
rect 13384 4992 13400 5026
rect 13334 4976 13400 4992
rect 13526 5026 13592 5042
rect 13640 5038 13670 5064
rect 13736 5042 13766 5064
rect 13526 4992 13542 5026
rect 13576 4992 13592 5026
rect 13526 4976 13592 4992
rect 13718 5026 13784 5042
rect 13832 5038 13862 5064
rect 13928 5042 13958 5064
rect 13718 4992 13734 5026
rect 13768 4992 13784 5026
rect 13718 4976 13784 4992
rect 13910 5026 13976 5042
rect 14024 5038 14054 5064
rect 14120 5042 14150 5064
rect 13910 4992 13926 5026
rect 13960 4992 13976 5026
rect 13910 4976 13976 4992
rect 14102 5026 14168 5042
rect 14216 5038 14246 5064
rect 14312 5042 14342 5064
rect 14102 4992 14118 5026
rect 14152 4992 14168 5026
rect 14102 4976 14168 4992
rect 14294 5026 14360 5042
rect 14408 5038 14438 5064
rect 14504 5042 14534 5064
rect 14294 4992 14310 5026
rect 14344 4992 14360 5026
rect 14294 4976 14360 4992
rect 14486 5026 14552 5042
rect 14600 5038 14630 5064
rect 14696 5042 14726 5064
rect 14486 4992 14502 5026
rect 14536 4992 14552 5026
rect 14486 4976 14552 4992
rect 14678 5026 14744 5042
rect 14792 5038 14822 5064
rect 14888 5042 14918 5064
rect 14678 4992 14694 5026
rect 14728 4992 14744 5026
rect 14678 4976 14744 4992
rect 14870 5026 14936 5042
rect 14870 4992 14886 5026
rect 14920 4992 14936 5026
rect 14870 4976 14936 4992
rect 12182 4918 12248 4934
rect 12182 4884 12198 4918
rect 12232 4884 12248 4918
rect 12104 4846 12134 4872
rect 12182 4868 12248 4884
rect 12374 4918 12440 4934
rect 12374 4884 12390 4918
rect 12424 4884 12440 4918
rect 12200 4846 12230 4868
rect 12296 4846 12326 4872
rect 12374 4868 12440 4884
rect 12566 4918 12632 4934
rect 12566 4884 12582 4918
rect 12616 4884 12632 4918
rect 12392 4846 12422 4868
rect 12488 4846 12518 4872
rect 12566 4868 12632 4884
rect 12758 4918 12824 4934
rect 12758 4884 12774 4918
rect 12808 4884 12824 4918
rect 12584 4846 12614 4868
rect 12680 4846 12710 4872
rect 12758 4868 12824 4884
rect 12950 4918 13016 4934
rect 12950 4884 12966 4918
rect 13000 4884 13016 4918
rect 12776 4846 12806 4868
rect 12872 4846 12902 4872
rect 12950 4868 13016 4884
rect 13142 4918 13208 4934
rect 13142 4884 13158 4918
rect 13192 4884 13208 4918
rect 12968 4846 12998 4868
rect 13064 4846 13094 4872
rect 13142 4868 13208 4884
rect 13334 4918 13400 4934
rect 13334 4884 13350 4918
rect 13384 4884 13400 4918
rect 13160 4846 13190 4868
rect 13256 4846 13286 4872
rect 13334 4868 13400 4884
rect 13526 4918 13592 4934
rect 13526 4884 13542 4918
rect 13576 4884 13592 4918
rect 13352 4846 13382 4868
rect 13448 4846 13478 4872
rect 13526 4868 13592 4884
rect 13718 4918 13784 4934
rect 13718 4884 13734 4918
rect 13768 4884 13784 4918
rect 13544 4846 13574 4868
rect 13640 4846 13670 4872
rect 13718 4868 13784 4884
rect 13910 4918 13976 4934
rect 13910 4884 13926 4918
rect 13960 4884 13976 4918
rect 13736 4846 13766 4868
rect 13832 4846 13862 4872
rect 13910 4868 13976 4884
rect 14102 4918 14168 4934
rect 14102 4884 14118 4918
rect 14152 4884 14168 4918
rect 13928 4846 13958 4868
rect 14024 4846 14054 4872
rect 14102 4868 14168 4884
rect 14294 4918 14360 4934
rect 14294 4884 14310 4918
rect 14344 4884 14360 4918
rect 14120 4846 14150 4868
rect 14216 4846 14246 4872
rect 14294 4868 14360 4884
rect 14486 4918 14552 4934
rect 14486 4884 14502 4918
rect 14536 4884 14552 4918
rect 14312 4846 14342 4868
rect 14408 4846 14438 4872
rect 14486 4868 14552 4884
rect 14678 4918 14744 4934
rect 14678 4884 14694 4918
rect 14728 4884 14744 4918
rect 14504 4846 14534 4868
rect 14600 4846 14630 4872
rect 14678 4868 14744 4884
rect 14870 4918 14936 4934
rect 14870 4884 14886 4918
rect 14920 4884 14936 4918
rect 14696 4846 14726 4868
rect 14792 4846 14822 4872
rect 14870 4868 14936 4884
rect 14888 4846 14918 4868
rect 12104 4424 12134 4446
rect 12086 4408 12152 4424
rect 12200 4420 12230 4446
rect 12296 4424 12326 4446
rect 12086 4374 12102 4408
rect 12136 4374 12152 4408
rect 12086 4358 12152 4374
rect 12278 4408 12344 4424
rect 12392 4420 12422 4446
rect 12488 4424 12518 4446
rect 12278 4374 12294 4408
rect 12328 4374 12344 4408
rect 12278 4358 12344 4374
rect 12470 4408 12536 4424
rect 12584 4420 12614 4446
rect 12680 4424 12710 4446
rect 12470 4374 12486 4408
rect 12520 4374 12536 4408
rect 12470 4358 12536 4374
rect 12662 4408 12728 4424
rect 12776 4420 12806 4446
rect 12872 4424 12902 4446
rect 12662 4374 12678 4408
rect 12712 4374 12728 4408
rect 12662 4358 12728 4374
rect 12854 4408 12920 4424
rect 12968 4420 12998 4446
rect 13064 4424 13094 4446
rect 12854 4374 12870 4408
rect 12904 4374 12920 4408
rect 12854 4358 12920 4374
rect 13046 4408 13112 4424
rect 13160 4420 13190 4446
rect 13256 4424 13286 4446
rect 13046 4374 13062 4408
rect 13096 4374 13112 4408
rect 13046 4358 13112 4374
rect 13238 4408 13304 4424
rect 13352 4420 13382 4446
rect 13448 4424 13478 4446
rect 13238 4374 13254 4408
rect 13288 4374 13304 4408
rect 13238 4358 13304 4374
rect 13430 4408 13496 4424
rect 13544 4420 13574 4446
rect 13640 4424 13670 4446
rect 13430 4374 13446 4408
rect 13480 4374 13496 4408
rect 13430 4358 13496 4374
rect 13622 4408 13688 4424
rect 13736 4420 13766 4446
rect 13832 4424 13862 4446
rect 13622 4374 13638 4408
rect 13672 4374 13688 4408
rect 13622 4358 13688 4374
rect 13814 4408 13880 4424
rect 13928 4420 13958 4446
rect 14024 4424 14054 4446
rect 13814 4374 13830 4408
rect 13864 4374 13880 4408
rect 13814 4358 13880 4374
rect 14006 4408 14072 4424
rect 14120 4420 14150 4446
rect 14216 4424 14246 4446
rect 14006 4374 14022 4408
rect 14056 4374 14072 4408
rect 14006 4358 14072 4374
rect 14198 4408 14264 4424
rect 14312 4420 14342 4446
rect 14408 4424 14438 4446
rect 14198 4374 14214 4408
rect 14248 4374 14264 4408
rect 14198 4358 14264 4374
rect 14390 4408 14456 4424
rect 14504 4420 14534 4446
rect 14600 4424 14630 4446
rect 14390 4374 14406 4408
rect 14440 4374 14456 4408
rect 14390 4358 14456 4374
rect 14582 4408 14648 4424
rect 14696 4420 14726 4446
rect 14792 4424 14822 4446
rect 14582 4374 14598 4408
rect 14632 4374 14648 4408
rect 14582 4358 14648 4374
rect 14774 4408 14840 4424
rect 14888 4420 14918 4446
rect 14774 4374 14790 4408
rect 14824 4374 14840 4408
rect 14774 4358 14840 4374
rect 12086 4300 12152 4316
rect 12086 4266 12102 4300
rect 12136 4266 12152 4300
rect 12086 4250 12152 4266
rect 12278 4300 12344 4316
rect 12278 4266 12294 4300
rect 12328 4266 12344 4300
rect 12104 4228 12134 4250
rect 12200 4228 12230 4254
rect 12278 4250 12344 4266
rect 12470 4300 12536 4316
rect 12470 4266 12486 4300
rect 12520 4266 12536 4300
rect 12296 4228 12326 4250
rect 12392 4228 12422 4254
rect 12470 4250 12536 4266
rect 12662 4300 12728 4316
rect 12662 4266 12678 4300
rect 12712 4266 12728 4300
rect 12488 4228 12518 4250
rect 12584 4228 12614 4254
rect 12662 4250 12728 4266
rect 12854 4300 12920 4316
rect 12854 4266 12870 4300
rect 12904 4266 12920 4300
rect 12680 4228 12710 4250
rect 12776 4228 12806 4254
rect 12854 4250 12920 4266
rect 13046 4300 13112 4316
rect 13046 4266 13062 4300
rect 13096 4266 13112 4300
rect 12872 4228 12902 4250
rect 12968 4228 12998 4254
rect 13046 4250 13112 4266
rect 13238 4300 13304 4316
rect 13238 4266 13254 4300
rect 13288 4266 13304 4300
rect 13064 4228 13094 4250
rect 13160 4228 13190 4254
rect 13238 4250 13304 4266
rect 13430 4300 13496 4316
rect 13430 4266 13446 4300
rect 13480 4266 13496 4300
rect 13256 4228 13286 4250
rect 13352 4228 13382 4254
rect 13430 4250 13496 4266
rect 13622 4300 13688 4316
rect 13622 4266 13638 4300
rect 13672 4266 13688 4300
rect 13448 4228 13478 4250
rect 13544 4228 13574 4254
rect 13622 4250 13688 4266
rect 13814 4300 13880 4316
rect 13814 4266 13830 4300
rect 13864 4266 13880 4300
rect 13640 4228 13670 4250
rect 13736 4228 13766 4254
rect 13814 4250 13880 4266
rect 14006 4300 14072 4316
rect 14006 4266 14022 4300
rect 14056 4266 14072 4300
rect 13832 4228 13862 4250
rect 13928 4228 13958 4254
rect 14006 4250 14072 4266
rect 14198 4300 14264 4316
rect 14198 4266 14214 4300
rect 14248 4266 14264 4300
rect 14024 4228 14054 4250
rect 14120 4228 14150 4254
rect 14198 4250 14264 4266
rect 14390 4300 14456 4316
rect 14390 4266 14406 4300
rect 14440 4266 14456 4300
rect 14216 4228 14246 4250
rect 14312 4228 14342 4254
rect 14390 4250 14456 4266
rect 14582 4300 14648 4316
rect 14582 4266 14598 4300
rect 14632 4266 14648 4300
rect 14408 4228 14438 4250
rect 14504 4228 14534 4254
rect 14582 4250 14648 4266
rect 14774 4300 14840 4316
rect 14774 4266 14790 4300
rect 14824 4266 14840 4300
rect 14600 4228 14630 4250
rect 14696 4228 14726 4254
rect 14774 4250 14840 4266
rect 14792 4228 14822 4250
rect 14888 4228 14918 4254
rect 12104 3802 12134 3828
rect 12200 3806 12230 3828
rect 12182 3790 12248 3806
rect 12296 3802 12326 3828
rect 12392 3806 12422 3828
rect 12182 3756 12198 3790
rect 12232 3756 12248 3790
rect 12182 3740 12248 3756
rect 12374 3790 12440 3806
rect 12488 3802 12518 3828
rect 12584 3806 12614 3828
rect 12374 3756 12390 3790
rect 12424 3756 12440 3790
rect 12374 3740 12440 3756
rect 12566 3790 12632 3806
rect 12680 3802 12710 3828
rect 12776 3806 12806 3828
rect 12566 3756 12582 3790
rect 12616 3756 12632 3790
rect 12566 3740 12632 3756
rect 12758 3790 12824 3806
rect 12872 3802 12902 3828
rect 12968 3806 12998 3828
rect 12758 3756 12774 3790
rect 12808 3756 12824 3790
rect 12758 3740 12824 3756
rect 12950 3790 13016 3806
rect 13064 3802 13094 3828
rect 13160 3806 13190 3828
rect 12950 3756 12966 3790
rect 13000 3756 13016 3790
rect 12950 3740 13016 3756
rect 13142 3790 13208 3806
rect 13256 3802 13286 3828
rect 13352 3806 13382 3828
rect 13142 3756 13158 3790
rect 13192 3756 13208 3790
rect 13142 3740 13208 3756
rect 13334 3790 13400 3806
rect 13448 3802 13478 3828
rect 13544 3806 13574 3828
rect 13334 3756 13350 3790
rect 13384 3756 13400 3790
rect 13334 3740 13400 3756
rect 13526 3790 13592 3806
rect 13640 3802 13670 3828
rect 13736 3806 13766 3828
rect 13526 3756 13542 3790
rect 13576 3756 13592 3790
rect 13526 3740 13592 3756
rect 13718 3790 13784 3806
rect 13832 3802 13862 3828
rect 13928 3806 13958 3828
rect 13718 3756 13734 3790
rect 13768 3756 13784 3790
rect 13718 3740 13784 3756
rect 13910 3790 13976 3806
rect 14024 3802 14054 3828
rect 14120 3806 14150 3828
rect 13910 3756 13926 3790
rect 13960 3756 13976 3790
rect 13910 3740 13976 3756
rect 14102 3790 14168 3806
rect 14216 3802 14246 3828
rect 14312 3806 14342 3828
rect 14102 3756 14118 3790
rect 14152 3756 14168 3790
rect 14102 3740 14168 3756
rect 14294 3790 14360 3806
rect 14408 3802 14438 3828
rect 14504 3806 14534 3828
rect 14294 3756 14310 3790
rect 14344 3756 14360 3790
rect 14294 3740 14360 3756
rect 14486 3790 14552 3806
rect 14600 3802 14630 3828
rect 14696 3806 14726 3828
rect 14486 3756 14502 3790
rect 14536 3756 14552 3790
rect 14486 3740 14552 3756
rect 14678 3790 14744 3806
rect 14792 3802 14822 3828
rect 14888 3806 14918 3828
rect 14678 3756 14694 3790
rect 14728 3756 14744 3790
rect 14678 3740 14744 3756
rect 14870 3790 14936 3806
rect 14870 3756 14886 3790
rect 14920 3756 14936 3790
rect 14870 3740 14936 3756
rect 12182 3682 12248 3698
rect 12182 3648 12198 3682
rect 12232 3648 12248 3682
rect 12104 3610 12134 3636
rect 12182 3632 12248 3648
rect 12374 3682 12440 3698
rect 12374 3648 12390 3682
rect 12424 3648 12440 3682
rect 12200 3610 12230 3632
rect 12296 3610 12326 3636
rect 12374 3632 12440 3648
rect 12566 3682 12632 3698
rect 12566 3648 12582 3682
rect 12616 3648 12632 3682
rect 12392 3610 12422 3632
rect 12488 3610 12518 3636
rect 12566 3632 12632 3648
rect 12758 3682 12824 3698
rect 12758 3648 12774 3682
rect 12808 3648 12824 3682
rect 12584 3610 12614 3632
rect 12680 3610 12710 3636
rect 12758 3632 12824 3648
rect 12950 3682 13016 3698
rect 12950 3648 12966 3682
rect 13000 3648 13016 3682
rect 12776 3610 12806 3632
rect 12872 3610 12902 3636
rect 12950 3632 13016 3648
rect 13142 3682 13208 3698
rect 13142 3648 13158 3682
rect 13192 3648 13208 3682
rect 12968 3610 12998 3632
rect 13064 3610 13094 3636
rect 13142 3632 13208 3648
rect 13334 3682 13400 3698
rect 13334 3648 13350 3682
rect 13384 3648 13400 3682
rect 13160 3610 13190 3632
rect 13256 3610 13286 3636
rect 13334 3632 13400 3648
rect 13526 3682 13592 3698
rect 13526 3648 13542 3682
rect 13576 3648 13592 3682
rect 13352 3610 13382 3632
rect 13448 3610 13478 3636
rect 13526 3632 13592 3648
rect 13718 3682 13784 3698
rect 13718 3648 13734 3682
rect 13768 3648 13784 3682
rect 13544 3610 13574 3632
rect 13640 3610 13670 3636
rect 13718 3632 13784 3648
rect 13910 3682 13976 3698
rect 13910 3648 13926 3682
rect 13960 3648 13976 3682
rect 13736 3610 13766 3632
rect 13832 3610 13862 3636
rect 13910 3632 13976 3648
rect 14102 3682 14168 3698
rect 14102 3648 14118 3682
rect 14152 3648 14168 3682
rect 13928 3610 13958 3632
rect 14024 3610 14054 3636
rect 14102 3632 14168 3648
rect 14294 3682 14360 3698
rect 14294 3648 14310 3682
rect 14344 3648 14360 3682
rect 14120 3610 14150 3632
rect 14216 3610 14246 3636
rect 14294 3632 14360 3648
rect 14486 3682 14552 3698
rect 14486 3648 14502 3682
rect 14536 3648 14552 3682
rect 14312 3610 14342 3632
rect 14408 3610 14438 3636
rect 14486 3632 14552 3648
rect 14678 3682 14744 3698
rect 14678 3648 14694 3682
rect 14728 3648 14744 3682
rect 14504 3610 14534 3632
rect 14600 3610 14630 3636
rect 14678 3632 14744 3648
rect 14870 3682 14936 3698
rect 14870 3648 14886 3682
rect 14920 3648 14936 3682
rect 14696 3610 14726 3632
rect 14792 3610 14822 3636
rect 14870 3632 14936 3648
rect 14888 3610 14918 3632
rect 12104 3188 12134 3210
rect 12086 3172 12152 3188
rect 12200 3184 12230 3210
rect 12296 3188 12326 3210
rect 12086 3138 12102 3172
rect 12136 3138 12152 3172
rect 12086 3122 12152 3138
rect 12278 3172 12344 3188
rect 12392 3184 12422 3210
rect 12488 3188 12518 3210
rect 12278 3138 12294 3172
rect 12328 3138 12344 3172
rect 12278 3122 12344 3138
rect 12470 3172 12536 3188
rect 12584 3184 12614 3210
rect 12680 3188 12710 3210
rect 12470 3138 12486 3172
rect 12520 3138 12536 3172
rect 12470 3122 12536 3138
rect 12662 3172 12728 3188
rect 12776 3184 12806 3210
rect 12872 3188 12902 3210
rect 12662 3138 12678 3172
rect 12712 3138 12728 3172
rect 12662 3122 12728 3138
rect 12854 3172 12920 3188
rect 12968 3184 12998 3210
rect 13064 3188 13094 3210
rect 12854 3138 12870 3172
rect 12904 3138 12920 3172
rect 12854 3122 12920 3138
rect 13046 3172 13112 3188
rect 13160 3184 13190 3210
rect 13256 3188 13286 3210
rect 13046 3138 13062 3172
rect 13096 3138 13112 3172
rect 13046 3122 13112 3138
rect 13238 3172 13304 3188
rect 13352 3184 13382 3210
rect 13448 3188 13478 3210
rect 13238 3138 13254 3172
rect 13288 3138 13304 3172
rect 13238 3122 13304 3138
rect 13430 3172 13496 3188
rect 13544 3184 13574 3210
rect 13640 3188 13670 3210
rect 13430 3138 13446 3172
rect 13480 3138 13496 3172
rect 13430 3122 13496 3138
rect 13622 3172 13688 3188
rect 13736 3184 13766 3210
rect 13832 3188 13862 3210
rect 13622 3138 13638 3172
rect 13672 3138 13688 3172
rect 13622 3122 13688 3138
rect 13814 3172 13880 3188
rect 13928 3184 13958 3210
rect 14024 3188 14054 3210
rect 13814 3138 13830 3172
rect 13864 3138 13880 3172
rect 13814 3122 13880 3138
rect 14006 3172 14072 3188
rect 14120 3184 14150 3210
rect 14216 3188 14246 3210
rect 14006 3138 14022 3172
rect 14056 3138 14072 3172
rect 14006 3122 14072 3138
rect 14198 3172 14264 3188
rect 14312 3184 14342 3210
rect 14408 3188 14438 3210
rect 14198 3138 14214 3172
rect 14248 3138 14264 3172
rect 14198 3122 14264 3138
rect 14390 3172 14456 3188
rect 14504 3184 14534 3210
rect 14600 3188 14630 3210
rect 14390 3138 14406 3172
rect 14440 3138 14456 3172
rect 14390 3122 14456 3138
rect 14582 3172 14648 3188
rect 14696 3184 14726 3210
rect 14792 3188 14822 3210
rect 14582 3138 14598 3172
rect 14632 3138 14648 3172
rect 14582 3122 14648 3138
rect 14774 3172 14840 3188
rect 14888 3184 14918 3210
rect 14774 3138 14790 3172
rect 14824 3138 14840 3172
rect 14774 3122 14840 3138
rect 15726 5536 15792 5552
rect 15726 5502 15742 5536
rect 15776 5502 15792 5536
rect 15726 5486 15792 5502
rect 15918 5536 15984 5552
rect 15918 5502 15934 5536
rect 15968 5502 15984 5536
rect 15744 5464 15774 5486
rect 15840 5464 15870 5490
rect 15918 5486 15984 5502
rect 16110 5536 16176 5552
rect 16110 5502 16126 5536
rect 16160 5502 16176 5536
rect 15936 5464 15966 5486
rect 16032 5464 16062 5490
rect 16110 5486 16176 5502
rect 16302 5536 16368 5552
rect 16302 5502 16318 5536
rect 16352 5502 16368 5536
rect 16128 5464 16158 5486
rect 16224 5464 16254 5490
rect 16302 5486 16368 5502
rect 16494 5536 16560 5552
rect 16494 5502 16510 5536
rect 16544 5502 16560 5536
rect 16320 5464 16350 5486
rect 16416 5464 16446 5490
rect 16494 5486 16560 5502
rect 16686 5536 16752 5552
rect 16686 5502 16702 5536
rect 16736 5502 16752 5536
rect 16512 5464 16542 5486
rect 16608 5464 16638 5490
rect 16686 5486 16752 5502
rect 16878 5536 16944 5552
rect 16878 5502 16894 5536
rect 16928 5502 16944 5536
rect 16704 5464 16734 5486
rect 16800 5464 16830 5490
rect 16878 5486 16944 5502
rect 17070 5536 17136 5552
rect 17070 5502 17086 5536
rect 17120 5502 17136 5536
rect 16896 5464 16926 5486
rect 16992 5464 17022 5490
rect 17070 5486 17136 5502
rect 17262 5536 17328 5552
rect 17262 5502 17278 5536
rect 17312 5502 17328 5536
rect 17088 5464 17118 5486
rect 17184 5464 17214 5490
rect 17262 5486 17328 5502
rect 17454 5536 17520 5552
rect 17454 5502 17470 5536
rect 17504 5502 17520 5536
rect 17280 5464 17310 5486
rect 17376 5464 17406 5490
rect 17454 5486 17520 5502
rect 17646 5536 17712 5552
rect 17646 5502 17662 5536
rect 17696 5502 17712 5536
rect 17472 5464 17502 5486
rect 17568 5464 17598 5490
rect 17646 5486 17712 5502
rect 17838 5536 17904 5552
rect 17838 5502 17854 5536
rect 17888 5502 17904 5536
rect 17664 5464 17694 5486
rect 17760 5464 17790 5490
rect 17838 5486 17904 5502
rect 18030 5536 18096 5552
rect 18030 5502 18046 5536
rect 18080 5502 18096 5536
rect 17856 5464 17886 5486
rect 17952 5464 17982 5490
rect 18030 5486 18096 5502
rect 18222 5536 18288 5552
rect 18222 5502 18238 5536
rect 18272 5502 18288 5536
rect 18048 5464 18078 5486
rect 18144 5464 18174 5490
rect 18222 5486 18288 5502
rect 18414 5536 18480 5552
rect 18414 5502 18430 5536
rect 18464 5502 18480 5536
rect 18240 5464 18270 5486
rect 18336 5464 18366 5490
rect 18414 5486 18480 5502
rect 18432 5464 18462 5486
rect 18528 5464 18558 5490
rect 15744 5038 15774 5064
rect 15840 5042 15870 5064
rect 15822 5026 15888 5042
rect 15936 5038 15966 5064
rect 16032 5042 16062 5064
rect 15822 4992 15838 5026
rect 15872 4992 15888 5026
rect 15822 4976 15888 4992
rect 16014 5026 16080 5042
rect 16128 5038 16158 5064
rect 16224 5042 16254 5064
rect 16014 4992 16030 5026
rect 16064 4992 16080 5026
rect 16014 4976 16080 4992
rect 16206 5026 16272 5042
rect 16320 5038 16350 5064
rect 16416 5042 16446 5064
rect 16206 4992 16222 5026
rect 16256 4992 16272 5026
rect 16206 4976 16272 4992
rect 16398 5026 16464 5042
rect 16512 5038 16542 5064
rect 16608 5042 16638 5064
rect 16398 4992 16414 5026
rect 16448 4992 16464 5026
rect 16398 4976 16464 4992
rect 16590 5026 16656 5042
rect 16704 5038 16734 5064
rect 16800 5042 16830 5064
rect 16590 4992 16606 5026
rect 16640 4992 16656 5026
rect 16590 4976 16656 4992
rect 16782 5026 16848 5042
rect 16896 5038 16926 5064
rect 16992 5042 17022 5064
rect 16782 4992 16798 5026
rect 16832 4992 16848 5026
rect 16782 4976 16848 4992
rect 16974 5026 17040 5042
rect 17088 5038 17118 5064
rect 17184 5042 17214 5064
rect 16974 4992 16990 5026
rect 17024 4992 17040 5026
rect 16974 4976 17040 4992
rect 17166 5026 17232 5042
rect 17280 5038 17310 5064
rect 17376 5042 17406 5064
rect 17166 4992 17182 5026
rect 17216 4992 17232 5026
rect 17166 4976 17232 4992
rect 17358 5026 17424 5042
rect 17472 5038 17502 5064
rect 17568 5042 17598 5064
rect 17358 4992 17374 5026
rect 17408 4992 17424 5026
rect 17358 4976 17424 4992
rect 17550 5026 17616 5042
rect 17664 5038 17694 5064
rect 17760 5042 17790 5064
rect 17550 4992 17566 5026
rect 17600 4992 17616 5026
rect 17550 4976 17616 4992
rect 17742 5026 17808 5042
rect 17856 5038 17886 5064
rect 17952 5042 17982 5064
rect 17742 4992 17758 5026
rect 17792 4992 17808 5026
rect 17742 4976 17808 4992
rect 17934 5026 18000 5042
rect 18048 5038 18078 5064
rect 18144 5042 18174 5064
rect 17934 4992 17950 5026
rect 17984 4992 18000 5026
rect 17934 4976 18000 4992
rect 18126 5026 18192 5042
rect 18240 5038 18270 5064
rect 18336 5042 18366 5064
rect 18126 4992 18142 5026
rect 18176 4992 18192 5026
rect 18126 4976 18192 4992
rect 18318 5026 18384 5042
rect 18432 5038 18462 5064
rect 18528 5042 18558 5064
rect 18318 4992 18334 5026
rect 18368 4992 18384 5026
rect 18318 4976 18384 4992
rect 18510 5026 18576 5042
rect 18510 4992 18526 5026
rect 18560 4992 18576 5026
rect 18510 4976 18576 4992
rect 15822 4918 15888 4934
rect 15822 4884 15838 4918
rect 15872 4884 15888 4918
rect 15744 4846 15774 4872
rect 15822 4868 15888 4884
rect 16014 4918 16080 4934
rect 16014 4884 16030 4918
rect 16064 4884 16080 4918
rect 15840 4846 15870 4868
rect 15936 4846 15966 4872
rect 16014 4868 16080 4884
rect 16206 4918 16272 4934
rect 16206 4884 16222 4918
rect 16256 4884 16272 4918
rect 16032 4846 16062 4868
rect 16128 4846 16158 4872
rect 16206 4868 16272 4884
rect 16398 4918 16464 4934
rect 16398 4884 16414 4918
rect 16448 4884 16464 4918
rect 16224 4846 16254 4868
rect 16320 4846 16350 4872
rect 16398 4868 16464 4884
rect 16590 4918 16656 4934
rect 16590 4884 16606 4918
rect 16640 4884 16656 4918
rect 16416 4846 16446 4868
rect 16512 4846 16542 4872
rect 16590 4868 16656 4884
rect 16782 4918 16848 4934
rect 16782 4884 16798 4918
rect 16832 4884 16848 4918
rect 16608 4846 16638 4868
rect 16704 4846 16734 4872
rect 16782 4868 16848 4884
rect 16974 4918 17040 4934
rect 16974 4884 16990 4918
rect 17024 4884 17040 4918
rect 16800 4846 16830 4868
rect 16896 4846 16926 4872
rect 16974 4868 17040 4884
rect 17166 4918 17232 4934
rect 17166 4884 17182 4918
rect 17216 4884 17232 4918
rect 16992 4846 17022 4868
rect 17088 4846 17118 4872
rect 17166 4868 17232 4884
rect 17358 4918 17424 4934
rect 17358 4884 17374 4918
rect 17408 4884 17424 4918
rect 17184 4846 17214 4868
rect 17280 4846 17310 4872
rect 17358 4868 17424 4884
rect 17550 4918 17616 4934
rect 17550 4884 17566 4918
rect 17600 4884 17616 4918
rect 17376 4846 17406 4868
rect 17472 4846 17502 4872
rect 17550 4868 17616 4884
rect 17742 4918 17808 4934
rect 17742 4884 17758 4918
rect 17792 4884 17808 4918
rect 17568 4846 17598 4868
rect 17664 4846 17694 4872
rect 17742 4868 17808 4884
rect 17934 4918 18000 4934
rect 17934 4884 17950 4918
rect 17984 4884 18000 4918
rect 17760 4846 17790 4868
rect 17856 4846 17886 4872
rect 17934 4868 18000 4884
rect 18126 4918 18192 4934
rect 18126 4884 18142 4918
rect 18176 4884 18192 4918
rect 17952 4846 17982 4868
rect 18048 4846 18078 4872
rect 18126 4868 18192 4884
rect 18318 4918 18384 4934
rect 18318 4884 18334 4918
rect 18368 4884 18384 4918
rect 18144 4846 18174 4868
rect 18240 4846 18270 4872
rect 18318 4868 18384 4884
rect 18510 4918 18576 4934
rect 18510 4884 18526 4918
rect 18560 4884 18576 4918
rect 18336 4846 18366 4868
rect 18432 4846 18462 4872
rect 18510 4868 18576 4884
rect 18528 4846 18558 4868
rect 15744 4424 15774 4446
rect 15726 4408 15792 4424
rect 15840 4420 15870 4446
rect 15936 4424 15966 4446
rect 15726 4374 15742 4408
rect 15776 4374 15792 4408
rect 15726 4358 15792 4374
rect 15918 4408 15984 4424
rect 16032 4420 16062 4446
rect 16128 4424 16158 4446
rect 15918 4374 15934 4408
rect 15968 4374 15984 4408
rect 15918 4358 15984 4374
rect 16110 4408 16176 4424
rect 16224 4420 16254 4446
rect 16320 4424 16350 4446
rect 16110 4374 16126 4408
rect 16160 4374 16176 4408
rect 16110 4358 16176 4374
rect 16302 4408 16368 4424
rect 16416 4420 16446 4446
rect 16512 4424 16542 4446
rect 16302 4374 16318 4408
rect 16352 4374 16368 4408
rect 16302 4358 16368 4374
rect 16494 4408 16560 4424
rect 16608 4420 16638 4446
rect 16704 4424 16734 4446
rect 16494 4374 16510 4408
rect 16544 4374 16560 4408
rect 16494 4358 16560 4374
rect 16686 4408 16752 4424
rect 16800 4420 16830 4446
rect 16896 4424 16926 4446
rect 16686 4374 16702 4408
rect 16736 4374 16752 4408
rect 16686 4358 16752 4374
rect 16878 4408 16944 4424
rect 16992 4420 17022 4446
rect 17088 4424 17118 4446
rect 16878 4374 16894 4408
rect 16928 4374 16944 4408
rect 16878 4358 16944 4374
rect 17070 4408 17136 4424
rect 17184 4420 17214 4446
rect 17280 4424 17310 4446
rect 17070 4374 17086 4408
rect 17120 4374 17136 4408
rect 17070 4358 17136 4374
rect 17262 4408 17328 4424
rect 17376 4420 17406 4446
rect 17472 4424 17502 4446
rect 17262 4374 17278 4408
rect 17312 4374 17328 4408
rect 17262 4358 17328 4374
rect 17454 4408 17520 4424
rect 17568 4420 17598 4446
rect 17664 4424 17694 4446
rect 17454 4374 17470 4408
rect 17504 4374 17520 4408
rect 17454 4358 17520 4374
rect 17646 4408 17712 4424
rect 17760 4420 17790 4446
rect 17856 4424 17886 4446
rect 17646 4374 17662 4408
rect 17696 4374 17712 4408
rect 17646 4358 17712 4374
rect 17838 4408 17904 4424
rect 17952 4420 17982 4446
rect 18048 4424 18078 4446
rect 17838 4374 17854 4408
rect 17888 4374 17904 4408
rect 17838 4358 17904 4374
rect 18030 4408 18096 4424
rect 18144 4420 18174 4446
rect 18240 4424 18270 4446
rect 18030 4374 18046 4408
rect 18080 4374 18096 4408
rect 18030 4358 18096 4374
rect 18222 4408 18288 4424
rect 18336 4420 18366 4446
rect 18432 4424 18462 4446
rect 18222 4374 18238 4408
rect 18272 4374 18288 4408
rect 18222 4358 18288 4374
rect 18414 4408 18480 4424
rect 18528 4420 18558 4446
rect 18414 4374 18430 4408
rect 18464 4374 18480 4408
rect 18414 4358 18480 4374
rect 15726 4300 15792 4316
rect 15726 4266 15742 4300
rect 15776 4266 15792 4300
rect 15726 4250 15792 4266
rect 15918 4300 15984 4316
rect 15918 4266 15934 4300
rect 15968 4266 15984 4300
rect 15744 4228 15774 4250
rect 15840 4228 15870 4254
rect 15918 4250 15984 4266
rect 16110 4300 16176 4316
rect 16110 4266 16126 4300
rect 16160 4266 16176 4300
rect 15936 4228 15966 4250
rect 16032 4228 16062 4254
rect 16110 4250 16176 4266
rect 16302 4300 16368 4316
rect 16302 4266 16318 4300
rect 16352 4266 16368 4300
rect 16128 4228 16158 4250
rect 16224 4228 16254 4254
rect 16302 4250 16368 4266
rect 16494 4300 16560 4316
rect 16494 4266 16510 4300
rect 16544 4266 16560 4300
rect 16320 4228 16350 4250
rect 16416 4228 16446 4254
rect 16494 4250 16560 4266
rect 16686 4300 16752 4316
rect 16686 4266 16702 4300
rect 16736 4266 16752 4300
rect 16512 4228 16542 4250
rect 16608 4228 16638 4254
rect 16686 4250 16752 4266
rect 16878 4300 16944 4316
rect 16878 4266 16894 4300
rect 16928 4266 16944 4300
rect 16704 4228 16734 4250
rect 16800 4228 16830 4254
rect 16878 4250 16944 4266
rect 17070 4300 17136 4316
rect 17070 4266 17086 4300
rect 17120 4266 17136 4300
rect 16896 4228 16926 4250
rect 16992 4228 17022 4254
rect 17070 4250 17136 4266
rect 17262 4300 17328 4316
rect 17262 4266 17278 4300
rect 17312 4266 17328 4300
rect 17088 4228 17118 4250
rect 17184 4228 17214 4254
rect 17262 4250 17328 4266
rect 17454 4300 17520 4316
rect 17454 4266 17470 4300
rect 17504 4266 17520 4300
rect 17280 4228 17310 4250
rect 17376 4228 17406 4254
rect 17454 4250 17520 4266
rect 17646 4300 17712 4316
rect 17646 4266 17662 4300
rect 17696 4266 17712 4300
rect 17472 4228 17502 4250
rect 17568 4228 17598 4254
rect 17646 4250 17712 4266
rect 17838 4300 17904 4316
rect 17838 4266 17854 4300
rect 17888 4266 17904 4300
rect 17664 4228 17694 4250
rect 17760 4228 17790 4254
rect 17838 4250 17904 4266
rect 18030 4300 18096 4316
rect 18030 4266 18046 4300
rect 18080 4266 18096 4300
rect 17856 4228 17886 4250
rect 17952 4228 17982 4254
rect 18030 4250 18096 4266
rect 18222 4300 18288 4316
rect 18222 4266 18238 4300
rect 18272 4266 18288 4300
rect 18048 4228 18078 4250
rect 18144 4228 18174 4254
rect 18222 4250 18288 4266
rect 18414 4300 18480 4316
rect 18414 4266 18430 4300
rect 18464 4266 18480 4300
rect 18240 4228 18270 4250
rect 18336 4228 18366 4254
rect 18414 4250 18480 4266
rect 18432 4228 18462 4250
rect 18528 4228 18558 4254
rect 15744 3802 15774 3828
rect 15840 3806 15870 3828
rect 15822 3790 15888 3806
rect 15936 3802 15966 3828
rect 16032 3806 16062 3828
rect 15822 3756 15838 3790
rect 15872 3756 15888 3790
rect 15822 3740 15888 3756
rect 16014 3790 16080 3806
rect 16128 3802 16158 3828
rect 16224 3806 16254 3828
rect 16014 3756 16030 3790
rect 16064 3756 16080 3790
rect 16014 3740 16080 3756
rect 16206 3790 16272 3806
rect 16320 3802 16350 3828
rect 16416 3806 16446 3828
rect 16206 3756 16222 3790
rect 16256 3756 16272 3790
rect 16206 3740 16272 3756
rect 16398 3790 16464 3806
rect 16512 3802 16542 3828
rect 16608 3806 16638 3828
rect 16398 3756 16414 3790
rect 16448 3756 16464 3790
rect 16398 3740 16464 3756
rect 16590 3790 16656 3806
rect 16704 3802 16734 3828
rect 16800 3806 16830 3828
rect 16590 3756 16606 3790
rect 16640 3756 16656 3790
rect 16590 3740 16656 3756
rect 16782 3790 16848 3806
rect 16896 3802 16926 3828
rect 16992 3806 17022 3828
rect 16782 3756 16798 3790
rect 16832 3756 16848 3790
rect 16782 3740 16848 3756
rect 16974 3790 17040 3806
rect 17088 3802 17118 3828
rect 17184 3806 17214 3828
rect 16974 3756 16990 3790
rect 17024 3756 17040 3790
rect 16974 3740 17040 3756
rect 17166 3790 17232 3806
rect 17280 3802 17310 3828
rect 17376 3806 17406 3828
rect 17166 3756 17182 3790
rect 17216 3756 17232 3790
rect 17166 3740 17232 3756
rect 17358 3790 17424 3806
rect 17472 3802 17502 3828
rect 17568 3806 17598 3828
rect 17358 3756 17374 3790
rect 17408 3756 17424 3790
rect 17358 3740 17424 3756
rect 17550 3790 17616 3806
rect 17664 3802 17694 3828
rect 17760 3806 17790 3828
rect 17550 3756 17566 3790
rect 17600 3756 17616 3790
rect 17550 3740 17616 3756
rect 17742 3790 17808 3806
rect 17856 3802 17886 3828
rect 17952 3806 17982 3828
rect 17742 3756 17758 3790
rect 17792 3756 17808 3790
rect 17742 3740 17808 3756
rect 17934 3790 18000 3806
rect 18048 3802 18078 3828
rect 18144 3806 18174 3828
rect 17934 3756 17950 3790
rect 17984 3756 18000 3790
rect 17934 3740 18000 3756
rect 18126 3790 18192 3806
rect 18240 3802 18270 3828
rect 18336 3806 18366 3828
rect 18126 3756 18142 3790
rect 18176 3756 18192 3790
rect 18126 3740 18192 3756
rect 18318 3790 18384 3806
rect 18432 3802 18462 3828
rect 18528 3806 18558 3828
rect 18318 3756 18334 3790
rect 18368 3756 18384 3790
rect 18318 3740 18384 3756
rect 18510 3790 18576 3806
rect 18510 3756 18526 3790
rect 18560 3756 18576 3790
rect 18510 3740 18576 3756
rect 15822 3682 15888 3698
rect 15822 3648 15838 3682
rect 15872 3648 15888 3682
rect 15744 3610 15774 3636
rect 15822 3632 15888 3648
rect 16014 3682 16080 3698
rect 16014 3648 16030 3682
rect 16064 3648 16080 3682
rect 15840 3610 15870 3632
rect 15936 3610 15966 3636
rect 16014 3632 16080 3648
rect 16206 3682 16272 3698
rect 16206 3648 16222 3682
rect 16256 3648 16272 3682
rect 16032 3610 16062 3632
rect 16128 3610 16158 3636
rect 16206 3632 16272 3648
rect 16398 3682 16464 3698
rect 16398 3648 16414 3682
rect 16448 3648 16464 3682
rect 16224 3610 16254 3632
rect 16320 3610 16350 3636
rect 16398 3632 16464 3648
rect 16590 3682 16656 3698
rect 16590 3648 16606 3682
rect 16640 3648 16656 3682
rect 16416 3610 16446 3632
rect 16512 3610 16542 3636
rect 16590 3632 16656 3648
rect 16782 3682 16848 3698
rect 16782 3648 16798 3682
rect 16832 3648 16848 3682
rect 16608 3610 16638 3632
rect 16704 3610 16734 3636
rect 16782 3632 16848 3648
rect 16974 3682 17040 3698
rect 16974 3648 16990 3682
rect 17024 3648 17040 3682
rect 16800 3610 16830 3632
rect 16896 3610 16926 3636
rect 16974 3632 17040 3648
rect 17166 3682 17232 3698
rect 17166 3648 17182 3682
rect 17216 3648 17232 3682
rect 16992 3610 17022 3632
rect 17088 3610 17118 3636
rect 17166 3632 17232 3648
rect 17358 3682 17424 3698
rect 17358 3648 17374 3682
rect 17408 3648 17424 3682
rect 17184 3610 17214 3632
rect 17280 3610 17310 3636
rect 17358 3632 17424 3648
rect 17550 3682 17616 3698
rect 17550 3648 17566 3682
rect 17600 3648 17616 3682
rect 17376 3610 17406 3632
rect 17472 3610 17502 3636
rect 17550 3632 17616 3648
rect 17742 3682 17808 3698
rect 17742 3648 17758 3682
rect 17792 3648 17808 3682
rect 17568 3610 17598 3632
rect 17664 3610 17694 3636
rect 17742 3632 17808 3648
rect 17934 3682 18000 3698
rect 17934 3648 17950 3682
rect 17984 3648 18000 3682
rect 17760 3610 17790 3632
rect 17856 3610 17886 3636
rect 17934 3632 18000 3648
rect 18126 3682 18192 3698
rect 18126 3648 18142 3682
rect 18176 3648 18192 3682
rect 17952 3610 17982 3632
rect 18048 3610 18078 3636
rect 18126 3632 18192 3648
rect 18318 3682 18384 3698
rect 18318 3648 18334 3682
rect 18368 3648 18384 3682
rect 18144 3610 18174 3632
rect 18240 3610 18270 3636
rect 18318 3632 18384 3648
rect 18510 3682 18576 3698
rect 18510 3648 18526 3682
rect 18560 3648 18576 3682
rect 18336 3610 18366 3632
rect 18432 3610 18462 3636
rect 18510 3632 18576 3648
rect 18528 3610 18558 3632
rect 15744 3188 15774 3210
rect 15726 3172 15792 3188
rect 15840 3184 15870 3210
rect 15936 3188 15966 3210
rect 15726 3138 15742 3172
rect 15776 3138 15792 3172
rect 15726 3122 15792 3138
rect 15918 3172 15984 3188
rect 16032 3184 16062 3210
rect 16128 3188 16158 3210
rect 15918 3138 15934 3172
rect 15968 3138 15984 3172
rect 15918 3122 15984 3138
rect 16110 3172 16176 3188
rect 16224 3184 16254 3210
rect 16320 3188 16350 3210
rect 16110 3138 16126 3172
rect 16160 3138 16176 3172
rect 16110 3122 16176 3138
rect 16302 3172 16368 3188
rect 16416 3184 16446 3210
rect 16512 3188 16542 3210
rect 16302 3138 16318 3172
rect 16352 3138 16368 3172
rect 16302 3122 16368 3138
rect 16494 3172 16560 3188
rect 16608 3184 16638 3210
rect 16704 3188 16734 3210
rect 16494 3138 16510 3172
rect 16544 3138 16560 3172
rect 16494 3122 16560 3138
rect 16686 3172 16752 3188
rect 16800 3184 16830 3210
rect 16896 3188 16926 3210
rect 16686 3138 16702 3172
rect 16736 3138 16752 3172
rect 16686 3122 16752 3138
rect 16878 3172 16944 3188
rect 16992 3184 17022 3210
rect 17088 3188 17118 3210
rect 16878 3138 16894 3172
rect 16928 3138 16944 3172
rect 16878 3122 16944 3138
rect 17070 3172 17136 3188
rect 17184 3184 17214 3210
rect 17280 3188 17310 3210
rect 17070 3138 17086 3172
rect 17120 3138 17136 3172
rect 17070 3122 17136 3138
rect 17262 3172 17328 3188
rect 17376 3184 17406 3210
rect 17472 3188 17502 3210
rect 17262 3138 17278 3172
rect 17312 3138 17328 3172
rect 17262 3122 17328 3138
rect 17454 3172 17520 3188
rect 17568 3184 17598 3210
rect 17664 3188 17694 3210
rect 17454 3138 17470 3172
rect 17504 3138 17520 3172
rect 17454 3122 17520 3138
rect 17646 3172 17712 3188
rect 17760 3184 17790 3210
rect 17856 3188 17886 3210
rect 17646 3138 17662 3172
rect 17696 3138 17712 3172
rect 17646 3122 17712 3138
rect 17838 3172 17904 3188
rect 17952 3184 17982 3210
rect 18048 3188 18078 3210
rect 17838 3138 17854 3172
rect 17888 3138 17904 3172
rect 17838 3122 17904 3138
rect 18030 3172 18096 3188
rect 18144 3184 18174 3210
rect 18240 3188 18270 3210
rect 18030 3138 18046 3172
rect 18080 3138 18096 3172
rect 18030 3122 18096 3138
rect 18222 3172 18288 3188
rect 18336 3184 18366 3210
rect 18432 3188 18462 3210
rect 18222 3138 18238 3172
rect 18272 3138 18288 3172
rect 18222 3122 18288 3138
rect 18414 3172 18480 3188
rect 18528 3184 18558 3210
rect 18414 3138 18430 3172
rect 18464 3138 18480 3172
rect 18414 3122 18480 3138
rect -1538 2704 -1472 2720
rect -1538 2670 -1522 2704
rect -1488 2670 -1472 2704
rect -1538 2654 -1472 2670
rect -1346 2704 -1280 2720
rect -1346 2670 -1330 2704
rect -1296 2670 -1280 2704
rect -1520 2632 -1490 2654
rect -1424 2632 -1394 2658
rect -1346 2654 -1280 2670
rect -1154 2704 -1088 2720
rect -1154 2670 -1138 2704
rect -1104 2670 -1088 2704
rect -1328 2632 -1298 2654
rect -1232 2632 -1202 2658
rect -1154 2654 -1088 2670
rect -1136 2632 -1106 2654
rect -1040 2632 -1010 2658
rect -1520 2206 -1490 2232
rect -1424 2210 -1394 2232
rect -1442 2194 -1376 2210
rect -1328 2206 -1298 2232
rect -1232 2210 -1202 2232
rect -1442 2160 -1426 2194
rect -1392 2160 -1376 2194
rect -1442 2144 -1376 2160
rect -1250 2194 -1184 2210
rect -1136 2206 -1106 2232
rect -1040 2210 -1010 2232
rect -1250 2160 -1234 2194
rect -1200 2160 -1184 2194
rect -1250 2144 -1184 2160
rect -1058 2194 -992 2210
rect -1058 2160 -1042 2194
rect -1008 2160 -992 2194
rect -1058 2144 -992 2160
rect -1442 2086 -1376 2102
rect -1442 2052 -1426 2086
rect -1392 2052 -1376 2086
rect -1520 2014 -1490 2040
rect -1442 2036 -1376 2052
rect -1250 2086 -1184 2102
rect -1250 2052 -1234 2086
rect -1200 2052 -1184 2086
rect -1424 2014 -1394 2036
rect -1328 2014 -1298 2040
rect -1250 2036 -1184 2052
rect -1058 2086 -992 2102
rect -1058 2052 -1042 2086
rect -1008 2052 -992 2086
rect -1232 2014 -1202 2036
rect -1136 2014 -1106 2040
rect -1058 2036 -992 2052
rect -1040 2014 -1010 2036
rect -1520 1592 -1490 1614
rect -1538 1576 -1472 1592
rect -1424 1588 -1394 1614
rect -1328 1592 -1298 1614
rect -1538 1542 -1522 1576
rect -1488 1542 -1472 1576
rect -1538 1526 -1472 1542
rect -1346 1576 -1280 1592
rect -1232 1588 -1202 1614
rect -1136 1592 -1106 1614
rect -1346 1542 -1330 1576
rect -1296 1542 -1280 1576
rect -1346 1526 -1280 1542
rect -1154 1576 -1088 1592
rect -1040 1588 -1010 1614
rect -1154 1542 -1138 1576
rect -1104 1542 -1088 1576
rect -1154 1526 -1088 1542
rect -498 2704 -432 2720
rect -498 2670 -482 2704
rect -448 2670 -432 2704
rect -498 2654 -432 2670
rect -306 2704 -240 2720
rect -306 2670 -290 2704
rect -256 2670 -240 2704
rect -480 2632 -450 2654
rect -384 2632 -354 2658
rect -306 2654 -240 2670
rect -114 2704 -48 2720
rect -114 2670 -98 2704
rect -64 2670 -48 2704
rect -288 2632 -258 2654
rect -192 2632 -162 2658
rect -114 2654 -48 2670
rect -96 2632 -66 2654
rect 0 2632 30 2658
rect -480 2206 -450 2232
rect -384 2210 -354 2232
rect -402 2194 -336 2210
rect -288 2206 -258 2232
rect -192 2210 -162 2232
rect -402 2160 -386 2194
rect -352 2160 -336 2194
rect -402 2144 -336 2160
rect -210 2194 -144 2210
rect -96 2206 -66 2232
rect 0 2210 30 2232
rect -210 2160 -194 2194
rect -160 2160 -144 2194
rect -210 2144 -144 2160
rect -18 2194 48 2210
rect -18 2160 -2 2194
rect 32 2160 48 2194
rect -18 2144 48 2160
rect -402 2086 -336 2102
rect -402 2052 -386 2086
rect -352 2052 -336 2086
rect -480 2014 -450 2040
rect -402 2036 -336 2052
rect -210 2086 -144 2102
rect -210 2052 -194 2086
rect -160 2052 -144 2086
rect -384 2014 -354 2036
rect -288 2014 -258 2040
rect -210 2036 -144 2052
rect -18 2086 48 2102
rect -18 2052 -2 2086
rect 32 2052 48 2086
rect -192 2014 -162 2036
rect -96 2014 -66 2040
rect -18 2036 48 2052
rect 0 2014 30 2036
rect -480 1592 -450 1614
rect -498 1576 -432 1592
rect -384 1588 -354 1614
rect -288 1592 -258 1614
rect -498 1542 -482 1576
rect -448 1542 -432 1576
rect -498 1526 -432 1542
rect -306 1576 -240 1592
rect -192 1588 -162 1614
rect -96 1592 -66 1614
rect -306 1542 -290 1576
rect -256 1542 -240 1576
rect -306 1526 -240 1542
rect -114 1576 -48 1592
rect 0 1588 30 1614
rect -114 1542 -98 1576
rect -64 1542 -48 1576
rect -114 1526 -48 1542
rect 542 2704 608 2720
rect 542 2670 558 2704
rect 592 2670 608 2704
rect 542 2654 608 2670
rect 734 2704 800 2720
rect 734 2670 750 2704
rect 784 2670 800 2704
rect 560 2632 590 2654
rect 656 2632 686 2658
rect 734 2654 800 2670
rect 926 2704 992 2720
rect 926 2670 942 2704
rect 976 2670 992 2704
rect 752 2632 782 2654
rect 848 2632 878 2658
rect 926 2654 992 2670
rect 944 2632 974 2654
rect 1040 2632 1070 2658
rect 560 2206 590 2232
rect 656 2210 686 2232
rect 638 2194 704 2210
rect 752 2206 782 2232
rect 848 2210 878 2232
rect 638 2160 654 2194
rect 688 2160 704 2194
rect 638 2144 704 2160
rect 830 2194 896 2210
rect 944 2206 974 2232
rect 1040 2210 1070 2232
rect 830 2160 846 2194
rect 880 2160 896 2194
rect 830 2144 896 2160
rect 1022 2194 1088 2210
rect 1022 2160 1038 2194
rect 1072 2160 1088 2194
rect 1022 2144 1088 2160
rect 638 2086 704 2102
rect 638 2052 654 2086
rect 688 2052 704 2086
rect 560 2014 590 2040
rect 638 2036 704 2052
rect 830 2086 896 2102
rect 830 2052 846 2086
rect 880 2052 896 2086
rect 656 2014 686 2036
rect 752 2014 782 2040
rect 830 2036 896 2052
rect 1022 2086 1088 2102
rect 1022 2052 1038 2086
rect 1072 2052 1088 2086
rect 848 2014 878 2036
rect 944 2014 974 2040
rect 1022 2036 1088 2052
rect 1040 2014 1070 2036
rect 560 1592 590 1614
rect 542 1576 608 1592
rect 656 1588 686 1614
rect 752 1592 782 1614
rect 542 1542 558 1576
rect 592 1542 608 1576
rect 542 1526 608 1542
rect 734 1576 800 1592
rect 848 1588 878 1614
rect 944 1592 974 1614
rect 734 1542 750 1576
rect 784 1542 800 1576
rect 734 1526 800 1542
rect 926 1576 992 1592
rect 1040 1588 1070 1614
rect 926 1542 942 1576
rect 976 1542 992 1576
rect 926 1526 992 1542
rect 1582 2704 1648 2720
rect 1582 2670 1598 2704
rect 1632 2670 1648 2704
rect 1582 2654 1648 2670
rect 1774 2704 1840 2720
rect 1774 2670 1790 2704
rect 1824 2670 1840 2704
rect 1600 2632 1630 2654
rect 1696 2632 1726 2658
rect 1774 2654 1840 2670
rect 1966 2704 2032 2720
rect 1966 2670 1982 2704
rect 2016 2670 2032 2704
rect 1792 2632 1822 2654
rect 1888 2632 1918 2658
rect 1966 2654 2032 2670
rect 1984 2632 2014 2654
rect 2080 2632 2110 2658
rect 1600 2206 1630 2232
rect 1696 2210 1726 2232
rect 1678 2194 1744 2210
rect 1792 2206 1822 2232
rect 1888 2210 1918 2232
rect 1678 2160 1694 2194
rect 1728 2160 1744 2194
rect 1678 2144 1744 2160
rect 1870 2194 1936 2210
rect 1984 2206 2014 2232
rect 2080 2210 2110 2232
rect 1870 2160 1886 2194
rect 1920 2160 1936 2194
rect 1870 2144 1936 2160
rect 2062 2194 2128 2210
rect 2062 2160 2078 2194
rect 2112 2160 2128 2194
rect 2062 2144 2128 2160
rect 1678 2086 1744 2102
rect 1678 2052 1694 2086
rect 1728 2052 1744 2086
rect 1600 2014 1630 2040
rect 1678 2036 1744 2052
rect 1870 2086 1936 2102
rect 1870 2052 1886 2086
rect 1920 2052 1936 2086
rect 1696 2014 1726 2036
rect 1792 2014 1822 2040
rect 1870 2036 1936 2052
rect 2062 2086 2128 2102
rect 2062 2052 2078 2086
rect 2112 2052 2128 2086
rect 1888 2014 1918 2036
rect 1984 2014 2014 2040
rect 2062 2036 2128 2052
rect 2080 2014 2110 2036
rect 1600 1592 1630 1614
rect 1582 1576 1648 1592
rect 1696 1588 1726 1614
rect 1792 1592 1822 1614
rect 1582 1542 1598 1576
rect 1632 1542 1648 1576
rect 1582 1526 1648 1542
rect 1774 1576 1840 1592
rect 1888 1588 1918 1614
rect 1984 1592 2014 1614
rect 1774 1542 1790 1576
rect 1824 1542 1840 1576
rect 1774 1526 1840 1542
rect 1966 1576 2032 1592
rect 2080 1588 2110 1614
rect 1966 1542 1982 1576
rect 2016 1542 2032 1576
rect 1966 1526 2032 1542
rect 2622 2704 2688 2720
rect 2622 2670 2638 2704
rect 2672 2670 2688 2704
rect 2622 2654 2688 2670
rect 2814 2704 2880 2720
rect 2814 2670 2830 2704
rect 2864 2670 2880 2704
rect 2640 2632 2670 2654
rect 2736 2632 2766 2658
rect 2814 2654 2880 2670
rect 3006 2704 3072 2720
rect 3006 2670 3022 2704
rect 3056 2670 3072 2704
rect 2832 2632 2862 2654
rect 2928 2632 2958 2658
rect 3006 2654 3072 2670
rect 3024 2632 3054 2654
rect 3120 2632 3150 2658
rect 2640 2206 2670 2232
rect 2736 2210 2766 2232
rect 2718 2194 2784 2210
rect 2832 2206 2862 2232
rect 2928 2210 2958 2232
rect 2718 2160 2734 2194
rect 2768 2160 2784 2194
rect 2718 2144 2784 2160
rect 2910 2194 2976 2210
rect 3024 2206 3054 2232
rect 3120 2210 3150 2232
rect 2910 2160 2926 2194
rect 2960 2160 2976 2194
rect 2910 2144 2976 2160
rect 3102 2194 3168 2210
rect 3102 2160 3118 2194
rect 3152 2160 3168 2194
rect 3102 2144 3168 2160
rect 2718 2086 2784 2102
rect 2718 2052 2734 2086
rect 2768 2052 2784 2086
rect 2640 2014 2670 2040
rect 2718 2036 2784 2052
rect 2910 2086 2976 2102
rect 2910 2052 2926 2086
rect 2960 2052 2976 2086
rect 2736 2014 2766 2036
rect 2832 2014 2862 2040
rect 2910 2036 2976 2052
rect 3102 2086 3168 2102
rect 3102 2052 3118 2086
rect 3152 2052 3168 2086
rect 2928 2014 2958 2036
rect 3024 2014 3054 2040
rect 3102 2036 3168 2052
rect 3120 2014 3150 2036
rect 2640 1592 2670 1614
rect 2622 1576 2688 1592
rect 2736 1588 2766 1614
rect 2832 1592 2862 1614
rect 2622 1542 2638 1576
rect 2672 1542 2688 1576
rect 2622 1526 2688 1542
rect 2814 1576 2880 1592
rect 2928 1588 2958 1614
rect 3024 1592 3054 1614
rect 2814 1542 2830 1576
rect 2864 1542 2880 1576
rect 2814 1526 2880 1542
rect 3006 1576 3072 1592
rect 3120 1588 3150 1614
rect 3006 1542 3022 1576
rect 3056 1542 3072 1576
rect 3006 1526 3072 1542
rect 4266 2864 4332 2880
rect 4266 2830 4282 2864
rect 4316 2830 4332 2864
rect 4266 2814 4332 2830
rect 4458 2864 4524 2880
rect 4458 2830 4474 2864
rect 4508 2830 4524 2864
rect 4284 2792 4314 2814
rect 4380 2792 4410 2818
rect 4458 2814 4524 2830
rect 4650 2864 4716 2880
rect 4650 2830 4666 2864
rect 4700 2830 4716 2864
rect 4476 2792 4506 2814
rect 4572 2792 4602 2818
rect 4650 2814 4716 2830
rect 4668 2792 4698 2814
rect 4764 2792 4794 2818
rect 4284 2366 4314 2392
rect 4380 2370 4410 2392
rect 4362 2354 4428 2370
rect 4476 2366 4506 2392
rect 4572 2370 4602 2392
rect 4362 2320 4378 2354
rect 4412 2320 4428 2354
rect 4362 2304 4428 2320
rect 4554 2354 4620 2370
rect 4668 2366 4698 2392
rect 4764 2370 4794 2392
rect 4554 2320 4570 2354
rect 4604 2320 4620 2354
rect 4554 2304 4620 2320
rect 4746 2354 4812 2370
rect 4746 2320 4762 2354
rect 4796 2320 4812 2354
rect 4746 2304 4812 2320
rect 4362 2246 4428 2262
rect 4362 2212 4378 2246
rect 4412 2212 4428 2246
rect 4284 2174 4314 2200
rect 4362 2196 4428 2212
rect 4554 2246 4620 2262
rect 4554 2212 4570 2246
rect 4604 2212 4620 2246
rect 4380 2174 4410 2196
rect 4476 2174 4506 2200
rect 4554 2196 4620 2212
rect 4746 2246 4812 2262
rect 4746 2212 4762 2246
rect 4796 2212 4812 2246
rect 4572 2174 4602 2196
rect 4668 2174 4698 2200
rect 4746 2196 4812 2212
rect 4764 2174 4794 2196
rect 4284 1752 4314 1774
rect 4266 1736 4332 1752
rect 4380 1748 4410 1774
rect 4476 1752 4506 1774
rect 4266 1702 4282 1736
rect 4316 1702 4332 1736
rect 4266 1686 4332 1702
rect 4458 1736 4524 1752
rect 4572 1748 4602 1774
rect 4668 1752 4698 1774
rect 4458 1702 4474 1736
rect 4508 1702 4524 1736
rect 4458 1686 4524 1702
rect 4650 1736 4716 1752
rect 4764 1748 4794 1774
rect 4650 1702 4666 1736
rect 4700 1702 4716 1736
rect 4650 1686 4716 1702
rect 5306 2864 5372 2880
rect 5306 2830 5322 2864
rect 5356 2830 5372 2864
rect 5306 2814 5372 2830
rect 5498 2864 5564 2880
rect 5498 2830 5514 2864
rect 5548 2830 5564 2864
rect 5324 2792 5354 2814
rect 5420 2792 5450 2818
rect 5498 2814 5564 2830
rect 5690 2864 5756 2880
rect 5690 2830 5706 2864
rect 5740 2830 5756 2864
rect 5516 2792 5546 2814
rect 5612 2792 5642 2818
rect 5690 2814 5756 2830
rect 5708 2792 5738 2814
rect 5804 2792 5834 2818
rect 5324 2366 5354 2392
rect 5420 2370 5450 2392
rect 5402 2354 5468 2370
rect 5516 2366 5546 2392
rect 5612 2370 5642 2392
rect 5402 2320 5418 2354
rect 5452 2320 5468 2354
rect 5402 2304 5468 2320
rect 5594 2354 5660 2370
rect 5708 2366 5738 2392
rect 5804 2370 5834 2392
rect 5594 2320 5610 2354
rect 5644 2320 5660 2354
rect 5594 2304 5660 2320
rect 5786 2354 5852 2370
rect 5786 2320 5802 2354
rect 5836 2320 5852 2354
rect 5786 2304 5852 2320
rect 5402 2246 5468 2262
rect 5402 2212 5418 2246
rect 5452 2212 5468 2246
rect 5324 2174 5354 2200
rect 5402 2196 5468 2212
rect 5594 2246 5660 2262
rect 5594 2212 5610 2246
rect 5644 2212 5660 2246
rect 5420 2174 5450 2196
rect 5516 2174 5546 2200
rect 5594 2196 5660 2212
rect 5786 2246 5852 2262
rect 5786 2212 5802 2246
rect 5836 2212 5852 2246
rect 5612 2174 5642 2196
rect 5708 2174 5738 2200
rect 5786 2196 5852 2212
rect 5804 2174 5834 2196
rect 5324 1752 5354 1774
rect 5306 1736 5372 1752
rect 5420 1748 5450 1774
rect 5516 1752 5546 1774
rect 5306 1702 5322 1736
rect 5356 1702 5372 1736
rect 5306 1686 5372 1702
rect 5498 1736 5564 1752
rect 5612 1748 5642 1774
rect 5708 1752 5738 1774
rect 5498 1702 5514 1736
rect 5548 1702 5564 1736
rect 5498 1686 5564 1702
rect 5690 1736 5756 1752
rect 5804 1748 5834 1774
rect 5690 1702 5706 1736
rect 5740 1702 5756 1736
rect 5690 1686 5756 1702
rect 6346 2864 6412 2880
rect 6346 2830 6362 2864
rect 6396 2830 6412 2864
rect 6346 2814 6412 2830
rect 6538 2864 6604 2880
rect 6538 2830 6554 2864
rect 6588 2830 6604 2864
rect 6364 2792 6394 2814
rect 6460 2792 6490 2818
rect 6538 2814 6604 2830
rect 6730 2864 6796 2880
rect 6730 2830 6746 2864
rect 6780 2830 6796 2864
rect 6556 2792 6586 2814
rect 6652 2792 6682 2818
rect 6730 2814 6796 2830
rect 6748 2792 6778 2814
rect 6844 2792 6874 2818
rect 6364 2366 6394 2392
rect 6460 2370 6490 2392
rect 6442 2354 6508 2370
rect 6556 2366 6586 2392
rect 6652 2370 6682 2392
rect 6442 2320 6458 2354
rect 6492 2320 6508 2354
rect 6442 2304 6508 2320
rect 6634 2354 6700 2370
rect 6748 2366 6778 2392
rect 6844 2370 6874 2392
rect 6634 2320 6650 2354
rect 6684 2320 6700 2354
rect 6634 2304 6700 2320
rect 6826 2354 6892 2370
rect 6826 2320 6842 2354
rect 6876 2320 6892 2354
rect 6826 2304 6892 2320
rect 6442 2246 6508 2262
rect 6442 2212 6458 2246
rect 6492 2212 6508 2246
rect 6364 2174 6394 2200
rect 6442 2196 6508 2212
rect 6634 2246 6700 2262
rect 6634 2212 6650 2246
rect 6684 2212 6700 2246
rect 6460 2174 6490 2196
rect 6556 2174 6586 2200
rect 6634 2196 6700 2212
rect 6826 2246 6892 2262
rect 6826 2212 6842 2246
rect 6876 2212 6892 2246
rect 6652 2174 6682 2196
rect 6748 2174 6778 2200
rect 6826 2196 6892 2212
rect 6844 2174 6874 2196
rect 6364 1752 6394 1774
rect 6346 1736 6412 1752
rect 6460 1748 6490 1774
rect 6556 1752 6586 1774
rect 6346 1702 6362 1736
rect 6396 1702 6412 1736
rect 6346 1686 6412 1702
rect 6538 1736 6604 1752
rect 6652 1748 6682 1774
rect 6748 1752 6778 1774
rect 6538 1702 6554 1736
rect 6588 1702 6604 1736
rect 6538 1686 6604 1702
rect 6730 1736 6796 1752
rect 6844 1748 6874 1774
rect 6730 1702 6746 1736
rect 6780 1702 6796 1736
rect 6730 1686 6796 1702
rect 7386 2864 7452 2880
rect 7386 2830 7402 2864
rect 7436 2830 7452 2864
rect 7386 2814 7452 2830
rect 7578 2864 7644 2880
rect 7578 2830 7594 2864
rect 7628 2830 7644 2864
rect 7404 2792 7434 2814
rect 7500 2792 7530 2818
rect 7578 2814 7644 2830
rect 7770 2864 7836 2880
rect 7770 2830 7786 2864
rect 7820 2830 7836 2864
rect 7596 2792 7626 2814
rect 7692 2792 7722 2818
rect 7770 2814 7836 2830
rect 7788 2792 7818 2814
rect 7884 2792 7914 2818
rect 7404 2366 7434 2392
rect 7500 2370 7530 2392
rect 7482 2354 7548 2370
rect 7596 2366 7626 2392
rect 7692 2370 7722 2392
rect 7482 2320 7498 2354
rect 7532 2320 7548 2354
rect 7482 2304 7548 2320
rect 7674 2354 7740 2370
rect 7788 2366 7818 2392
rect 7884 2370 7914 2392
rect 7674 2320 7690 2354
rect 7724 2320 7740 2354
rect 7674 2304 7740 2320
rect 7866 2354 7932 2370
rect 7866 2320 7882 2354
rect 7916 2320 7932 2354
rect 7866 2304 7932 2320
rect 7482 2246 7548 2262
rect 7482 2212 7498 2246
rect 7532 2212 7548 2246
rect 7404 2174 7434 2200
rect 7482 2196 7548 2212
rect 7674 2246 7740 2262
rect 7674 2212 7690 2246
rect 7724 2212 7740 2246
rect 7500 2174 7530 2196
rect 7596 2174 7626 2200
rect 7674 2196 7740 2212
rect 7866 2246 7932 2262
rect 7866 2212 7882 2246
rect 7916 2212 7932 2246
rect 7692 2174 7722 2196
rect 7788 2174 7818 2200
rect 7866 2196 7932 2212
rect 7884 2174 7914 2196
rect 7404 1752 7434 1774
rect 7386 1736 7452 1752
rect 7500 1748 7530 1774
rect 7596 1752 7626 1774
rect 7386 1702 7402 1736
rect 7436 1702 7452 1736
rect 7386 1686 7452 1702
rect 7578 1736 7644 1752
rect 7692 1748 7722 1774
rect 7788 1752 7818 1774
rect 7578 1702 7594 1736
rect 7628 1702 7644 1736
rect 7578 1686 7644 1702
rect 7770 1736 7836 1752
rect 7884 1748 7914 1774
rect 7770 1702 7786 1736
rect 7820 1702 7836 1736
rect 7770 1686 7836 1702
rect 8426 2864 8492 2880
rect 8426 2830 8442 2864
rect 8476 2830 8492 2864
rect 8426 2814 8492 2830
rect 8618 2864 8684 2880
rect 8618 2830 8634 2864
rect 8668 2830 8684 2864
rect 8444 2792 8474 2814
rect 8540 2792 8570 2818
rect 8618 2814 8684 2830
rect 8810 2864 8876 2880
rect 8810 2830 8826 2864
rect 8860 2830 8876 2864
rect 8636 2792 8666 2814
rect 8732 2792 8762 2818
rect 8810 2814 8876 2830
rect 8828 2792 8858 2814
rect 8924 2792 8954 2818
rect 8444 2366 8474 2392
rect 8540 2370 8570 2392
rect 8522 2354 8588 2370
rect 8636 2366 8666 2392
rect 8732 2370 8762 2392
rect 8522 2320 8538 2354
rect 8572 2320 8588 2354
rect 8522 2304 8588 2320
rect 8714 2354 8780 2370
rect 8828 2366 8858 2392
rect 8924 2370 8954 2392
rect 8714 2320 8730 2354
rect 8764 2320 8780 2354
rect 8714 2304 8780 2320
rect 8906 2354 8972 2370
rect 8906 2320 8922 2354
rect 8956 2320 8972 2354
rect 8906 2304 8972 2320
rect 8522 2246 8588 2262
rect 8522 2212 8538 2246
rect 8572 2212 8588 2246
rect 8444 2174 8474 2200
rect 8522 2196 8588 2212
rect 8714 2246 8780 2262
rect 8714 2212 8730 2246
rect 8764 2212 8780 2246
rect 8540 2174 8570 2196
rect 8636 2174 8666 2200
rect 8714 2196 8780 2212
rect 8906 2246 8972 2262
rect 8906 2212 8922 2246
rect 8956 2212 8972 2246
rect 8732 2174 8762 2196
rect 8828 2174 8858 2200
rect 8906 2196 8972 2212
rect 8924 2174 8954 2196
rect 8444 1752 8474 1774
rect 8426 1736 8492 1752
rect 8540 1748 8570 1774
rect 8636 1752 8666 1774
rect 8426 1702 8442 1736
rect 8476 1702 8492 1736
rect 8426 1686 8492 1702
rect 8618 1736 8684 1752
rect 8732 1748 8762 1774
rect 8828 1752 8858 1774
rect 8618 1702 8634 1736
rect 8668 1702 8684 1736
rect 8618 1686 8684 1702
rect 8810 1736 8876 1752
rect 8924 1748 8954 1774
rect 8810 1702 8826 1736
rect 8860 1702 8876 1736
rect 8810 1686 8876 1702
rect 9466 2864 9532 2880
rect 9466 2830 9482 2864
rect 9516 2830 9532 2864
rect 9466 2814 9532 2830
rect 9658 2864 9724 2880
rect 9658 2830 9674 2864
rect 9708 2830 9724 2864
rect 9484 2792 9514 2814
rect 9580 2792 9610 2818
rect 9658 2814 9724 2830
rect 9850 2864 9916 2880
rect 9850 2830 9866 2864
rect 9900 2830 9916 2864
rect 9676 2792 9706 2814
rect 9772 2792 9802 2818
rect 9850 2814 9916 2830
rect 9868 2792 9898 2814
rect 9964 2792 9994 2818
rect 9484 2366 9514 2392
rect 9580 2370 9610 2392
rect 9562 2354 9628 2370
rect 9676 2366 9706 2392
rect 9772 2370 9802 2392
rect 9562 2320 9578 2354
rect 9612 2320 9628 2354
rect 9562 2304 9628 2320
rect 9754 2354 9820 2370
rect 9868 2366 9898 2392
rect 9964 2370 9994 2392
rect 9754 2320 9770 2354
rect 9804 2320 9820 2354
rect 9754 2304 9820 2320
rect 9946 2354 10012 2370
rect 9946 2320 9962 2354
rect 9996 2320 10012 2354
rect 9946 2304 10012 2320
rect 9562 2246 9628 2262
rect 9562 2212 9578 2246
rect 9612 2212 9628 2246
rect 9484 2174 9514 2200
rect 9562 2196 9628 2212
rect 9754 2246 9820 2262
rect 9754 2212 9770 2246
rect 9804 2212 9820 2246
rect 9580 2174 9610 2196
rect 9676 2174 9706 2200
rect 9754 2196 9820 2212
rect 9946 2246 10012 2262
rect 9946 2212 9962 2246
rect 9996 2212 10012 2246
rect 9772 2174 9802 2196
rect 9868 2174 9898 2200
rect 9946 2196 10012 2212
rect 9964 2174 9994 2196
rect 9484 1752 9514 1774
rect 9466 1736 9532 1752
rect 9580 1748 9610 1774
rect 9676 1752 9706 1774
rect 9466 1702 9482 1736
rect 9516 1702 9532 1736
rect 9466 1686 9532 1702
rect 9658 1736 9724 1752
rect 9772 1748 9802 1774
rect 9868 1752 9898 1774
rect 9658 1702 9674 1736
rect 9708 1702 9724 1736
rect 9658 1686 9724 1702
rect 9850 1736 9916 1752
rect 9964 1748 9994 1774
rect 9850 1702 9866 1736
rect 9900 1702 9916 1736
rect 9850 1686 9916 1702
rect 10506 2864 10572 2880
rect 10506 2830 10522 2864
rect 10556 2830 10572 2864
rect 10506 2814 10572 2830
rect 10698 2864 10764 2880
rect 10698 2830 10714 2864
rect 10748 2830 10764 2864
rect 10524 2792 10554 2814
rect 10620 2792 10650 2818
rect 10698 2814 10764 2830
rect 10890 2864 10956 2880
rect 10890 2830 10906 2864
rect 10940 2830 10956 2864
rect 10716 2792 10746 2814
rect 10812 2792 10842 2818
rect 10890 2814 10956 2830
rect 10908 2792 10938 2814
rect 11004 2792 11034 2818
rect 10524 2366 10554 2392
rect 10620 2370 10650 2392
rect 10602 2354 10668 2370
rect 10716 2366 10746 2392
rect 10812 2370 10842 2392
rect 10602 2320 10618 2354
rect 10652 2320 10668 2354
rect 10602 2304 10668 2320
rect 10794 2354 10860 2370
rect 10908 2366 10938 2392
rect 11004 2370 11034 2392
rect 10794 2320 10810 2354
rect 10844 2320 10860 2354
rect 10794 2304 10860 2320
rect 10986 2354 11052 2370
rect 10986 2320 11002 2354
rect 11036 2320 11052 2354
rect 10986 2304 11052 2320
rect 10602 2246 10668 2262
rect 10602 2212 10618 2246
rect 10652 2212 10668 2246
rect 10524 2174 10554 2200
rect 10602 2196 10668 2212
rect 10794 2246 10860 2262
rect 10794 2212 10810 2246
rect 10844 2212 10860 2246
rect 10620 2174 10650 2196
rect 10716 2174 10746 2200
rect 10794 2196 10860 2212
rect 10986 2246 11052 2262
rect 10986 2212 11002 2246
rect 11036 2212 11052 2246
rect 10812 2174 10842 2196
rect 10908 2174 10938 2200
rect 10986 2196 11052 2212
rect 11004 2174 11034 2196
rect 10524 1752 10554 1774
rect 10506 1736 10572 1752
rect 10620 1748 10650 1774
rect 10716 1752 10746 1774
rect 10506 1702 10522 1736
rect 10556 1702 10572 1736
rect 10506 1686 10572 1702
rect 10698 1736 10764 1752
rect 10812 1748 10842 1774
rect 10908 1752 10938 1774
rect 10698 1702 10714 1736
rect 10748 1702 10764 1736
rect 10698 1686 10764 1702
rect 10890 1736 10956 1752
rect 11004 1748 11034 1774
rect 10890 1702 10906 1736
rect 10940 1702 10956 1736
rect 10890 1686 10956 1702
rect 11886 2864 11952 2880
rect 11886 2830 11902 2864
rect 11936 2830 11952 2864
rect 11886 2814 11952 2830
rect 12078 2864 12144 2880
rect 12078 2830 12094 2864
rect 12128 2830 12144 2864
rect 11904 2792 11934 2814
rect 12000 2792 12030 2818
rect 12078 2814 12144 2830
rect 12270 2864 12336 2880
rect 12270 2830 12286 2864
rect 12320 2830 12336 2864
rect 12096 2792 12126 2814
rect 12192 2792 12222 2818
rect 12270 2814 12336 2830
rect 12288 2792 12318 2814
rect 12384 2792 12414 2818
rect 11904 2366 11934 2392
rect 12000 2370 12030 2392
rect 11982 2354 12048 2370
rect 12096 2366 12126 2392
rect 12192 2370 12222 2392
rect 11982 2320 11998 2354
rect 12032 2320 12048 2354
rect 11982 2304 12048 2320
rect 12174 2354 12240 2370
rect 12288 2366 12318 2392
rect 12384 2370 12414 2392
rect 12174 2320 12190 2354
rect 12224 2320 12240 2354
rect 12174 2304 12240 2320
rect 12366 2354 12432 2370
rect 12366 2320 12382 2354
rect 12416 2320 12432 2354
rect 12366 2304 12432 2320
rect 11982 2246 12048 2262
rect 11982 2212 11998 2246
rect 12032 2212 12048 2246
rect 11904 2174 11934 2200
rect 11982 2196 12048 2212
rect 12174 2246 12240 2262
rect 12174 2212 12190 2246
rect 12224 2212 12240 2246
rect 12000 2174 12030 2196
rect 12096 2174 12126 2200
rect 12174 2196 12240 2212
rect 12366 2246 12432 2262
rect 12366 2212 12382 2246
rect 12416 2212 12432 2246
rect 12192 2174 12222 2196
rect 12288 2174 12318 2200
rect 12366 2196 12432 2212
rect 12384 2174 12414 2196
rect 11904 1752 11934 1774
rect 11886 1736 11952 1752
rect 12000 1748 12030 1774
rect 12096 1752 12126 1774
rect 11886 1702 11902 1736
rect 11936 1702 11952 1736
rect 11886 1686 11952 1702
rect 12078 1736 12144 1752
rect 12192 1748 12222 1774
rect 12288 1752 12318 1774
rect 12078 1702 12094 1736
rect 12128 1702 12144 1736
rect 12078 1686 12144 1702
rect 12270 1736 12336 1752
rect 12384 1748 12414 1774
rect 12270 1702 12286 1736
rect 12320 1702 12336 1736
rect 12270 1686 12336 1702
rect 12926 2864 12992 2880
rect 12926 2830 12942 2864
rect 12976 2830 12992 2864
rect 12926 2814 12992 2830
rect 13118 2864 13184 2880
rect 13118 2830 13134 2864
rect 13168 2830 13184 2864
rect 12944 2792 12974 2814
rect 13040 2792 13070 2818
rect 13118 2814 13184 2830
rect 13310 2864 13376 2880
rect 13310 2830 13326 2864
rect 13360 2830 13376 2864
rect 13136 2792 13166 2814
rect 13232 2792 13262 2818
rect 13310 2814 13376 2830
rect 13328 2792 13358 2814
rect 13424 2792 13454 2818
rect 12944 2366 12974 2392
rect 13040 2370 13070 2392
rect 13022 2354 13088 2370
rect 13136 2366 13166 2392
rect 13232 2370 13262 2392
rect 13022 2320 13038 2354
rect 13072 2320 13088 2354
rect 13022 2304 13088 2320
rect 13214 2354 13280 2370
rect 13328 2366 13358 2392
rect 13424 2370 13454 2392
rect 13214 2320 13230 2354
rect 13264 2320 13280 2354
rect 13214 2304 13280 2320
rect 13406 2354 13472 2370
rect 13406 2320 13422 2354
rect 13456 2320 13472 2354
rect 13406 2304 13472 2320
rect 13022 2246 13088 2262
rect 13022 2212 13038 2246
rect 13072 2212 13088 2246
rect 12944 2174 12974 2200
rect 13022 2196 13088 2212
rect 13214 2246 13280 2262
rect 13214 2212 13230 2246
rect 13264 2212 13280 2246
rect 13040 2174 13070 2196
rect 13136 2174 13166 2200
rect 13214 2196 13280 2212
rect 13406 2246 13472 2262
rect 13406 2212 13422 2246
rect 13456 2212 13472 2246
rect 13232 2174 13262 2196
rect 13328 2174 13358 2200
rect 13406 2196 13472 2212
rect 13424 2174 13454 2196
rect 12944 1752 12974 1774
rect 12926 1736 12992 1752
rect 13040 1748 13070 1774
rect 13136 1752 13166 1774
rect 12926 1702 12942 1736
rect 12976 1702 12992 1736
rect 12926 1686 12992 1702
rect 13118 1736 13184 1752
rect 13232 1748 13262 1774
rect 13328 1752 13358 1774
rect 13118 1702 13134 1736
rect 13168 1702 13184 1736
rect 13118 1686 13184 1702
rect 13310 1736 13376 1752
rect 13424 1748 13454 1774
rect 13310 1702 13326 1736
rect 13360 1702 13376 1736
rect 13310 1686 13376 1702
rect 13966 2864 14032 2880
rect 13966 2830 13982 2864
rect 14016 2830 14032 2864
rect 13966 2814 14032 2830
rect 14158 2864 14224 2880
rect 14158 2830 14174 2864
rect 14208 2830 14224 2864
rect 13984 2792 14014 2814
rect 14080 2792 14110 2818
rect 14158 2814 14224 2830
rect 14350 2864 14416 2880
rect 14350 2830 14366 2864
rect 14400 2830 14416 2864
rect 14176 2792 14206 2814
rect 14272 2792 14302 2818
rect 14350 2814 14416 2830
rect 14368 2792 14398 2814
rect 14464 2792 14494 2818
rect 13984 2366 14014 2392
rect 14080 2370 14110 2392
rect 14062 2354 14128 2370
rect 14176 2366 14206 2392
rect 14272 2370 14302 2392
rect 14062 2320 14078 2354
rect 14112 2320 14128 2354
rect 14062 2304 14128 2320
rect 14254 2354 14320 2370
rect 14368 2366 14398 2392
rect 14464 2370 14494 2392
rect 14254 2320 14270 2354
rect 14304 2320 14320 2354
rect 14254 2304 14320 2320
rect 14446 2354 14512 2370
rect 14446 2320 14462 2354
rect 14496 2320 14512 2354
rect 14446 2304 14512 2320
rect 14062 2246 14128 2262
rect 14062 2212 14078 2246
rect 14112 2212 14128 2246
rect 13984 2174 14014 2200
rect 14062 2196 14128 2212
rect 14254 2246 14320 2262
rect 14254 2212 14270 2246
rect 14304 2212 14320 2246
rect 14080 2174 14110 2196
rect 14176 2174 14206 2200
rect 14254 2196 14320 2212
rect 14446 2246 14512 2262
rect 14446 2212 14462 2246
rect 14496 2212 14512 2246
rect 14272 2174 14302 2196
rect 14368 2174 14398 2200
rect 14446 2196 14512 2212
rect 14464 2174 14494 2196
rect 13984 1752 14014 1774
rect 13966 1736 14032 1752
rect 14080 1748 14110 1774
rect 14176 1752 14206 1774
rect 13966 1702 13982 1736
rect 14016 1702 14032 1736
rect 13966 1686 14032 1702
rect 14158 1736 14224 1752
rect 14272 1748 14302 1774
rect 14368 1752 14398 1774
rect 14158 1702 14174 1736
rect 14208 1702 14224 1736
rect 14158 1686 14224 1702
rect 14350 1736 14416 1752
rect 14464 1748 14494 1774
rect 14350 1702 14366 1736
rect 14400 1702 14416 1736
rect 14350 1686 14416 1702
rect 15006 2864 15072 2880
rect 15006 2830 15022 2864
rect 15056 2830 15072 2864
rect 15006 2814 15072 2830
rect 15198 2864 15264 2880
rect 15198 2830 15214 2864
rect 15248 2830 15264 2864
rect 15024 2792 15054 2814
rect 15120 2792 15150 2818
rect 15198 2814 15264 2830
rect 15390 2864 15456 2880
rect 15390 2830 15406 2864
rect 15440 2830 15456 2864
rect 15216 2792 15246 2814
rect 15312 2792 15342 2818
rect 15390 2814 15456 2830
rect 15408 2792 15438 2814
rect 15504 2792 15534 2818
rect 15024 2366 15054 2392
rect 15120 2370 15150 2392
rect 15102 2354 15168 2370
rect 15216 2366 15246 2392
rect 15312 2370 15342 2392
rect 15102 2320 15118 2354
rect 15152 2320 15168 2354
rect 15102 2304 15168 2320
rect 15294 2354 15360 2370
rect 15408 2366 15438 2392
rect 15504 2370 15534 2392
rect 15294 2320 15310 2354
rect 15344 2320 15360 2354
rect 15294 2304 15360 2320
rect 15486 2354 15552 2370
rect 15486 2320 15502 2354
rect 15536 2320 15552 2354
rect 15486 2304 15552 2320
rect 15102 2246 15168 2262
rect 15102 2212 15118 2246
rect 15152 2212 15168 2246
rect 15024 2174 15054 2200
rect 15102 2196 15168 2212
rect 15294 2246 15360 2262
rect 15294 2212 15310 2246
rect 15344 2212 15360 2246
rect 15120 2174 15150 2196
rect 15216 2174 15246 2200
rect 15294 2196 15360 2212
rect 15486 2246 15552 2262
rect 15486 2212 15502 2246
rect 15536 2212 15552 2246
rect 15312 2174 15342 2196
rect 15408 2174 15438 2200
rect 15486 2196 15552 2212
rect 15504 2174 15534 2196
rect 15024 1752 15054 1774
rect 15006 1736 15072 1752
rect 15120 1748 15150 1774
rect 15216 1752 15246 1774
rect 15006 1702 15022 1736
rect 15056 1702 15072 1736
rect 15006 1686 15072 1702
rect 15198 1736 15264 1752
rect 15312 1748 15342 1774
rect 15408 1752 15438 1774
rect 15198 1702 15214 1736
rect 15248 1702 15264 1736
rect 15198 1686 15264 1702
rect 15390 1736 15456 1752
rect 15504 1748 15534 1774
rect 15390 1702 15406 1736
rect 15440 1702 15456 1736
rect 15390 1686 15456 1702
rect 16046 2864 16112 2880
rect 16046 2830 16062 2864
rect 16096 2830 16112 2864
rect 16046 2814 16112 2830
rect 16238 2864 16304 2880
rect 16238 2830 16254 2864
rect 16288 2830 16304 2864
rect 16064 2792 16094 2814
rect 16160 2792 16190 2818
rect 16238 2814 16304 2830
rect 16430 2864 16496 2880
rect 16430 2830 16446 2864
rect 16480 2830 16496 2864
rect 16256 2792 16286 2814
rect 16352 2792 16382 2818
rect 16430 2814 16496 2830
rect 16448 2792 16478 2814
rect 16544 2792 16574 2818
rect 16064 2366 16094 2392
rect 16160 2370 16190 2392
rect 16142 2354 16208 2370
rect 16256 2366 16286 2392
rect 16352 2370 16382 2392
rect 16142 2320 16158 2354
rect 16192 2320 16208 2354
rect 16142 2304 16208 2320
rect 16334 2354 16400 2370
rect 16448 2366 16478 2392
rect 16544 2370 16574 2392
rect 16334 2320 16350 2354
rect 16384 2320 16400 2354
rect 16334 2304 16400 2320
rect 16526 2354 16592 2370
rect 16526 2320 16542 2354
rect 16576 2320 16592 2354
rect 16526 2304 16592 2320
rect 16142 2246 16208 2262
rect 16142 2212 16158 2246
rect 16192 2212 16208 2246
rect 16064 2174 16094 2200
rect 16142 2196 16208 2212
rect 16334 2246 16400 2262
rect 16334 2212 16350 2246
rect 16384 2212 16400 2246
rect 16160 2174 16190 2196
rect 16256 2174 16286 2200
rect 16334 2196 16400 2212
rect 16526 2246 16592 2262
rect 16526 2212 16542 2246
rect 16576 2212 16592 2246
rect 16352 2174 16382 2196
rect 16448 2174 16478 2200
rect 16526 2196 16592 2212
rect 16544 2174 16574 2196
rect 16064 1752 16094 1774
rect 16046 1736 16112 1752
rect 16160 1748 16190 1774
rect 16256 1752 16286 1774
rect 16046 1702 16062 1736
rect 16096 1702 16112 1736
rect 16046 1686 16112 1702
rect 16238 1736 16304 1752
rect 16352 1748 16382 1774
rect 16448 1752 16478 1774
rect 16238 1702 16254 1736
rect 16288 1702 16304 1736
rect 16238 1686 16304 1702
rect 16430 1736 16496 1752
rect 16544 1748 16574 1774
rect 16430 1702 16446 1736
rect 16480 1702 16496 1736
rect 16430 1686 16496 1702
rect 17086 2864 17152 2880
rect 17086 2830 17102 2864
rect 17136 2830 17152 2864
rect 17086 2814 17152 2830
rect 17278 2864 17344 2880
rect 17278 2830 17294 2864
rect 17328 2830 17344 2864
rect 17104 2792 17134 2814
rect 17200 2792 17230 2818
rect 17278 2814 17344 2830
rect 17470 2864 17536 2880
rect 17470 2830 17486 2864
rect 17520 2830 17536 2864
rect 17296 2792 17326 2814
rect 17392 2792 17422 2818
rect 17470 2814 17536 2830
rect 17488 2792 17518 2814
rect 17584 2792 17614 2818
rect 17104 2366 17134 2392
rect 17200 2370 17230 2392
rect 17182 2354 17248 2370
rect 17296 2366 17326 2392
rect 17392 2370 17422 2392
rect 17182 2320 17198 2354
rect 17232 2320 17248 2354
rect 17182 2304 17248 2320
rect 17374 2354 17440 2370
rect 17488 2366 17518 2392
rect 17584 2370 17614 2392
rect 17374 2320 17390 2354
rect 17424 2320 17440 2354
rect 17374 2304 17440 2320
rect 17566 2354 17632 2370
rect 17566 2320 17582 2354
rect 17616 2320 17632 2354
rect 17566 2304 17632 2320
rect 17182 2246 17248 2262
rect 17182 2212 17198 2246
rect 17232 2212 17248 2246
rect 17104 2174 17134 2200
rect 17182 2196 17248 2212
rect 17374 2246 17440 2262
rect 17374 2212 17390 2246
rect 17424 2212 17440 2246
rect 17200 2174 17230 2196
rect 17296 2174 17326 2200
rect 17374 2196 17440 2212
rect 17566 2246 17632 2262
rect 17566 2212 17582 2246
rect 17616 2212 17632 2246
rect 17392 2174 17422 2196
rect 17488 2174 17518 2200
rect 17566 2196 17632 2212
rect 17584 2174 17614 2196
rect 17104 1752 17134 1774
rect 17086 1736 17152 1752
rect 17200 1748 17230 1774
rect 17296 1752 17326 1774
rect 17086 1702 17102 1736
rect 17136 1702 17152 1736
rect 17086 1686 17152 1702
rect 17278 1736 17344 1752
rect 17392 1748 17422 1774
rect 17488 1752 17518 1774
rect 17278 1702 17294 1736
rect 17328 1702 17344 1736
rect 17278 1686 17344 1702
rect 17470 1736 17536 1752
rect 17584 1748 17614 1774
rect 17470 1702 17486 1736
rect 17520 1702 17536 1736
rect 17470 1686 17536 1702
rect 18126 2864 18192 2880
rect 18126 2830 18142 2864
rect 18176 2830 18192 2864
rect 18126 2814 18192 2830
rect 18318 2864 18384 2880
rect 18318 2830 18334 2864
rect 18368 2830 18384 2864
rect 18144 2792 18174 2814
rect 18240 2792 18270 2818
rect 18318 2814 18384 2830
rect 18510 2864 18576 2880
rect 18510 2830 18526 2864
rect 18560 2830 18576 2864
rect 18336 2792 18366 2814
rect 18432 2792 18462 2818
rect 18510 2814 18576 2830
rect 18528 2792 18558 2814
rect 18624 2792 18654 2818
rect 18144 2366 18174 2392
rect 18240 2370 18270 2392
rect 18222 2354 18288 2370
rect 18336 2366 18366 2392
rect 18432 2370 18462 2392
rect 18222 2320 18238 2354
rect 18272 2320 18288 2354
rect 18222 2304 18288 2320
rect 18414 2354 18480 2370
rect 18528 2366 18558 2392
rect 18624 2370 18654 2392
rect 18414 2320 18430 2354
rect 18464 2320 18480 2354
rect 18414 2304 18480 2320
rect 18606 2354 18672 2370
rect 18606 2320 18622 2354
rect 18656 2320 18672 2354
rect 18606 2304 18672 2320
rect 18222 2246 18288 2262
rect 18222 2212 18238 2246
rect 18272 2212 18288 2246
rect 18144 2174 18174 2200
rect 18222 2196 18288 2212
rect 18414 2246 18480 2262
rect 18414 2212 18430 2246
rect 18464 2212 18480 2246
rect 18240 2174 18270 2196
rect 18336 2174 18366 2200
rect 18414 2196 18480 2212
rect 18606 2246 18672 2262
rect 18606 2212 18622 2246
rect 18656 2212 18672 2246
rect 18432 2174 18462 2196
rect 18528 2174 18558 2200
rect 18606 2196 18672 2212
rect 18624 2174 18654 2196
rect 18144 1752 18174 1774
rect 18126 1736 18192 1752
rect 18240 1748 18270 1774
rect 18336 1752 18366 1774
rect 18126 1702 18142 1736
rect 18176 1702 18192 1736
rect 18126 1686 18192 1702
rect 18318 1736 18384 1752
rect 18432 1748 18462 1774
rect 18528 1752 18558 1774
rect 18318 1702 18334 1736
rect 18368 1702 18384 1736
rect 18318 1686 18384 1702
rect 18510 1736 18576 1752
rect 18624 1748 18654 1774
rect 18510 1702 18526 1736
rect 18560 1702 18576 1736
rect 18510 1686 18576 1702
rect -1527 1282 -1461 1298
rect -1527 1248 -1511 1282
rect -1477 1248 -1461 1282
rect -1527 1232 -1461 1248
rect -1409 1282 -1343 1298
rect -1409 1248 -1393 1282
rect -1359 1248 -1343 1282
rect -1409 1232 -1343 1248
rect -1291 1282 -1225 1298
rect -1291 1248 -1275 1282
rect -1241 1248 -1225 1282
rect -1291 1232 -1225 1248
rect -1173 1282 -1107 1298
rect -1173 1248 -1157 1282
rect -1123 1248 -1107 1282
rect -1173 1232 -1107 1248
rect -1055 1282 -989 1298
rect -1055 1248 -1039 1282
rect -1005 1248 -989 1282
rect -1055 1232 -989 1248
rect -937 1282 -871 1298
rect -937 1248 -921 1282
rect -887 1248 -871 1282
rect -937 1232 -871 1248
rect -1524 1210 -1464 1232
rect -1406 1210 -1346 1232
rect -1288 1210 -1228 1232
rect -1170 1210 -1110 1232
rect -1052 1210 -992 1232
rect -934 1210 -874 1232
rect -1524 788 -1464 810
rect -1406 788 -1346 810
rect -1288 788 -1228 810
rect -1170 788 -1110 810
rect -1052 788 -992 810
rect -934 788 -874 810
rect -1527 772 -1461 788
rect -1527 738 -1511 772
rect -1477 738 -1461 772
rect -1527 722 -1461 738
rect -1409 772 -1343 788
rect -1409 738 -1393 772
rect -1359 738 -1343 772
rect -1409 722 -1343 738
rect -1291 772 -1225 788
rect -1291 738 -1275 772
rect -1241 738 -1225 772
rect -1291 722 -1225 738
rect -1173 772 -1107 788
rect -1173 738 -1157 772
rect -1123 738 -1107 772
rect -1173 722 -1107 738
rect -1055 772 -989 788
rect -1055 738 -1039 772
rect -1005 738 -989 772
rect -1055 722 -989 738
rect -937 772 -871 788
rect -937 738 -921 772
rect -887 738 -871 772
rect -937 722 -871 738
rect -487 1282 -421 1298
rect -487 1248 -471 1282
rect -437 1248 -421 1282
rect -487 1232 -421 1248
rect -369 1282 -303 1298
rect -369 1248 -353 1282
rect -319 1248 -303 1282
rect -369 1232 -303 1248
rect -251 1282 -185 1298
rect -251 1248 -235 1282
rect -201 1248 -185 1282
rect -251 1232 -185 1248
rect -133 1282 -67 1298
rect -133 1248 -117 1282
rect -83 1248 -67 1282
rect -133 1232 -67 1248
rect -15 1282 51 1298
rect -15 1248 1 1282
rect 35 1248 51 1282
rect -15 1232 51 1248
rect 103 1282 169 1298
rect 103 1248 119 1282
rect 153 1248 169 1282
rect 103 1232 169 1248
rect -484 1210 -424 1232
rect -366 1210 -306 1232
rect -248 1210 -188 1232
rect -130 1210 -70 1232
rect -12 1210 48 1232
rect 106 1210 166 1232
rect -484 788 -424 810
rect -366 788 -306 810
rect -248 788 -188 810
rect -130 788 -70 810
rect -12 788 48 810
rect 106 788 166 810
rect -487 772 -421 788
rect -487 738 -471 772
rect -437 738 -421 772
rect -487 722 -421 738
rect -369 772 -303 788
rect -369 738 -353 772
rect -319 738 -303 772
rect -369 722 -303 738
rect -251 772 -185 788
rect -251 738 -235 772
rect -201 738 -185 772
rect -251 722 -185 738
rect -133 772 -67 788
rect -133 738 -117 772
rect -83 738 -67 772
rect -133 722 -67 738
rect -15 772 51 788
rect -15 738 1 772
rect 35 738 51 772
rect -15 722 51 738
rect 103 772 169 788
rect 103 738 119 772
rect 153 738 169 772
rect 103 722 169 738
rect 553 1282 619 1298
rect 553 1248 569 1282
rect 603 1248 619 1282
rect 553 1232 619 1248
rect 671 1282 737 1298
rect 671 1248 687 1282
rect 721 1248 737 1282
rect 671 1232 737 1248
rect 789 1282 855 1298
rect 789 1248 805 1282
rect 839 1248 855 1282
rect 789 1232 855 1248
rect 907 1282 973 1298
rect 907 1248 923 1282
rect 957 1248 973 1282
rect 907 1232 973 1248
rect 1025 1282 1091 1298
rect 1025 1248 1041 1282
rect 1075 1248 1091 1282
rect 1025 1232 1091 1248
rect 1143 1282 1209 1298
rect 1143 1248 1159 1282
rect 1193 1248 1209 1282
rect 1143 1232 1209 1248
rect 556 1210 616 1232
rect 674 1210 734 1232
rect 792 1210 852 1232
rect 910 1210 970 1232
rect 1028 1210 1088 1232
rect 1146 1210 1206 1232
rect 556 788 616 810
rect 674 788 734 810
rect 792 788 852 810
rect 910 788 970 810
rect 1028 788 1088 810
rect 1146 788 1206 810
rect 553 772 619 788
rect 553 738 569 772
rect 603 738 619 772
rect 553 722 619 738
rect 671 772 737 788
rect 671 738 687 772
rect 721 738 737 772
rect 671 722 737 738
rect 789 772 855 788
rect 789 738 805 772
rect 839 738 855 772
rect 789 722 855 738
rect 907 772 973 788
rect 907 738 923 772
rect 957 738 973 772
rect 907 722 973 738
rect 1025 772 1091 788
rect 1025 738 1041 772
rect 1075 738 1091 772
rect 1025 722 1091 738
rect 1143 772 1209 788
rect 1143 738 1159 772
rect 1193 738 1209 772
rect 1143 722 1209 738
rect 1593 1282 1659 1298
rect 1593 1248 1609 1282
rect 1643 1248 1659 1282
rect 1593 1232 1659 1248
rect 1711 1282 1777 1298
rect 1711 1248 1727 1282
rect 1761 1248 1777 1282
rect 1711 1232 1777 1248
rect 1829 1282 1895 1298
rect 1829 1248 1845 1282
rect 1879 1248 1895 1282
rect 1829 1232 1895 1248
rect 1947 1282 2013 1298
rect 1947 1248 1963 1282
rect 1997 1248 2013 1282
rect 1947 1232 2013 1248
rect 2065 1282 2131 1298
rect 2065 1248 2081 1282
rect 2115 1248 2131 1282
rect 2065 1232 2131 1248
rect 2183 1282 2249 1298
rect 2183 1248 2199 1282
rect 2233 1248 2249 1282
rect 2183 1232 2249 1248
rect 1596 1210 1656 1232
rect 1714 1210 1774 1232
rect 1832 1210 1892 1232
rect 1950 1210 2010 1232
rect 2068 1210 2128 1232
rect 2186 1210 2246 1232
rect 1596 788 1656 810
rect 1714 788 1774 810
rect 1832 788 1892 810
rect 1950 788 2010 810
rect 2068 788 2128 810
rect 2186 788 2246 810
rect 1593 772 1659 788
rect 1593 738 1609 772
rect 1643 738 1659 772
rect 1593 722 1659 738
rect 1711 772 1777 788
rect 1711 738 1727 772
rect 1761 738 1777 772
rect 1711 722 1777 738
rect 1829 772 1895 788
rect 1829 738 1845 772
rect 1879 738 1895 772
rect 1829 722 1895 738
rect 1947 772 2013 788
rect 1947 738 1963 772
rect 1997 738 2013 772
rect 1947 722 2013 738
rect 2065 772 2131 788
rect 2065 738 2081 772
rect 2115 738 2131 772
rect 2065 722 2131 738
rect 2183 772 2249 788
rect 2183 738 2199 772
rect 2233 738 2249 772
rect 2183 722 2249 738
rect 2633 1282 2699 1298
rect 2633 1248 2649 1282
rect 2683 1248 2699 1282
rect 2633 1232 2699 1248
rect 2751 1282 2817 1298
rect 2751 1248 2767 1282
rect 2801 1248 2817 1282
rect 2751 1232 2817 1248
rect 2869 1282 2935 1298
rect 2869 1248 2885 1282
rect 2919 1248 2935 1282
rect 2869 1232 2935 1248
rect 2987 1282 3053 1298
rect 2987 1248 3003 1282
rect 3037 1248 3053 1282
rect 2987 1232 3053 1248
rect 3105 1282 3171 1298
rect 3105 1248 3121 1282
rect 3155 1248 3171 1282
rect 3105 1232 3171 1248
rect 3223 1282 3289 1298
rect 3223 1248 3239 1282
rect 3273 1248 3289 1282
rect 3223 1232 3289 1248
rect 2636 1210 2696 1232
rect 2754 1210 2814 1232
rect 2872 1210 2932 1232
rect 2990 1210 3050 1232
rect 3108 1210 3168 1232
rect 3226 1210 3286 1232
rect 2636 788 2696 810
rect 2754 788 2814 810
rect 2872 788 2932 810
rect 2990 788 3050 810
rect 3108 788 3168 810
rect 3226 788 3286 810
rect 2633 772 2699 788
rect 2633 738 2649 772
rect 2683 738 2699 772
rect 2633 722 2699 738
rect 2751 772 2817 788
rect 2751 738 2767 772
rect 2801 738 2817 772
rect 2751 722 2817 738
rect 2869 772 2935 788
rect 2869 738 2885 772
rect 2919 738 2935 772
rect 2869 722 2935 738
rect 2987 772 3053 788
rect 2987 738 3003 772
rect 3037 738 3053 772
rect 2987 722 3053 738
rect 3105 772 3171 788
rect 3105 738 3121 772
rect 3155 738 3171 772
rect 3105 722 3171 738
rect 3223 772 3289 788
rect 3223 738 3239 772
rect 3273 738 3289 772
rect 3223 722 3289 738
rect 4277 1442 4343 1458
rect 4277 1408 4293 1442
rect 4327 1408 4343 1442
rect 4277 1392 4343 1408
rect 4395 1442 4461 1458
rect 4395 1408 4411 1442
rect 4445 1408 4461 1442
rect 4395 1392 4461 1408
rect 4513 1442 4579 1458
rect 4513 1408 4529 1442
rect 4563 1408 4579 1442
rect 4513 1392 4579 1408
rect 4631 1442 4697 1458
rect 4631 1408 4647 1442
rect 4681 1408 4697 1442
rect 4631 1392 4697 1408
rect 4749 1442 4815 1458
rect 4749 1408 4765 1442
rect 4799 1408 4815 1442
rect 4749 1392 4815 1408
rect 4867 1442 4933 1458
rect 4867 1408 4883 1442
rect 4917 1408 4933 1442
rect 4867 1392 4933 1408
rect 4280 1370 4340 1392
rect 4398 1370 4458 1392
rect 4516 1370 4576 1392
rect 4634 1370 4694 1392
rect 4752 1370 4812 1392
rect 4870 1370 4930 1392
rect 4280 948 4340 970
rect 4398 948 4458 970
rect 4516 948 4576 970
rect 4634 948 4694 970
rect 4752 948 4812 970
rect 4870 948 4930 970
rect 4277 932 4343 948
rect 4277 898 4293 932
rect 4327 898 4343 932
rect 4277 882 4343 898
rect 4395 932 4461 948
rect 4395 898 4411 932
rect 4445 898 4461 932
rect 4395 882 4461 898
rect 4513 932 4579 948
rect 4513 898 4529 932
rect 4563 898 4579 932
rect 4513 882 4579 898
rect 4631 932 4697 948
rect 4631 898 4647 932
rect 4681 898 4697 932
rect 4631 882 4697 898
rect 4749 932 4815 948
rect 4749 898 4765 932
rect 4799 898 4815 932
rect 4749 882 4815 898
rect 4867 932 4933 948
rect 4867 898 4883 932
rect 4917 898 4933 932
rect 4867 882 4933 898
rect 5317 1442 5383 1458
rect 5317 1408 5333 1442
rect 5367 1408 5383 1442
rect 5317 1392 5383 1408
rect 5435 1442 5501 1458
rect 5435 1408 5451 1442
rect 5485 1408 5501 1442
rect 5435 1392 5501 1408
rect 5553 1442 5619 1458
rect 5553 1408 5569 1442
rect 5603 1408 5619 1442
rect 5553 1392 5619 1408
rect 5671 1442 5737 1458
rect 5671 1408 5687 1442
rect 5721 1408 5737 1442
rect 5671 1392 5737 1408
rect 5789 1442 5855 1458
rect 5789 1408 5805 1442
rect 5839 1408 5855 1442
rect 5789 1392 5855 1408
rect 5907 1442 5973 1458
rect 5907 1408 5923 1442
rect 5957 1408 5973 1442
rect 5907 1392 5973 1408
rect 5320 1370 5380 1392
rect 5438 1370 5498 1392
rect 5556 1370 5616 1392
rect 5674 1370 5734 1392
rect 5792 1370 5852 1392
rect 5910 1370 5970 1392
rect 5320 948 5380 970
rect 5438 948 5498 970
rect 5556 948 5616 970
rect 5674 948 5734 970
rect 5792 948 5852 970
rect 5910 948 5970 970
rect 5317 932 5383 948
rect 5317 898 5333 932
rect 5367 898 5383 932
rect 5317 882 5383 898
rect 5435 932 5501 948
rect 5435 898 5451 932
rect 5485 898 5501 932
rect 5435 882 5501 898
rect 5553 932 5619 948
rect 5553 898 5569 932
rect 5603 898 5619 932
rect 5553 882 5619 898
rect 5671 932 5737 948
rect 5671 898 5687 932
rect 5721 898 5737 932
rect 5671 882 5737 898
rect 5789 932 5855 948
rect 5789 898 5805 932
rect 5839 898 5855 932
rect 5789 882 5855 898
rect 5907 932 5973 948
rect 5907 898 5923 932
rect 5957 898 5973 932
rect 5907 882 5973 898
rect 6357 1442 6423 1458
rect 6357 1408 6373 1442
rect 6407 1408 6423 1442
rect 6357 1392 6423 1408
rect 6475 1442 6541 1458
rect 6475 1408 6491 1442
rect 6525 1408 6541 1442
rect 6475 1392 6541 1408
rect 6593 1442 6659 1458
rect 6593 1408 6609 1442
rect 6643 1408 6659 1442
rect 6593 1392 6659 1408
rect 6711 1442 6777 1458
rect 6711 1408 6727 1442
rect 6761 1408 6777 1442
rect 6711 1392 6777 1408
rect 6829 1442 6895 1458
rect 6829 1408 6845 1442
rect 6879 1408 6895 1442
rect 6829 1392 6895 1408
rect 6947 1442 7013 1458
rect 6947 1408 6963 1442
rect 6997 1408 7013 1442
rect 6947 1392 7013 1408
rect 6360 1370 6420 1392
rect 6478 1370 6538 1392
rect 6596 1370 6656 1392
rect 6714 1370 6774 1392
rect 6832 1370 6892 1392
rect 6950 1370 7010 1392
rect 6360 948 6420 970
rect 6478 948 6538 970
rect 6596 948 6656 970
rect 6714 948 6774 970
rect 6832 948 6892 970
rect 6950 948 7010 970
rect 6357 932 6423 948
rect 6357 898 6373 932
rect 6407 898 6423 932
rect 6357 882 6423 898
rect 6475 932 6541 948
rect 6475 898 6491 932
rect 6525 898 6541 932
rect 6475 882 6541 898
rect 6593 932 6659 948
rect 6593 898 6609 932
rect 6643 898 6659 932
rect 6593 882 6659 898
rect 6711 932 6777 948
rect 6711 898 6727 932
rect 6761 898 6777 932
rect 6711 882 6777 898
rect 6829 932 6895 948
rect 6829 898 6845 932
rect 6879 898 6895 932
rect 6829 882 6895 898
rect 6947 932 7013 948
rect 6947 898 6963 932
rect 6997 898 7013 932
rect 6947 882 7013 898
rect 7397 1442 7463 1458
rect 7397 1408 7413 1442
rect 7447 1408 7463 1442
rect 7397 1392 7463 1408
rect 7515 1442 7581 1458
rect 7515 1408 7531 1442
rect 7565 1408 7581 1442
rect 7515 1392 7581 1408
rect 7633 1442 7699 1458
rect 7633 1408 7649 1442
rect 7683 1408 7699 1442
rect 7633 1392 7699 1408
rect 7751 1442 7817 1458
rect 7751 1408 7767 1442
rect 7801 1408 7817 1442
rect 7751 1392 7817 1408
rect 7869 1442 7935 1458
rect 7869 1408 7885 1442
rect 7919 1408 7935 1442
rect 7869 1392 7935 1408
rect 7987 1442 8053 1458
rect 7987 1408 8003 1442
rect 8037 1408 8053 1442
rect 7987 1392 8053 1408
rect 7400 1370 7460 1392
rect 7518 1370 7578 1392
rect 7636 1370 7696 1392
rect 7754 1370 7814 1392
rect 7872 1370 7932 1392
rect 7990 1370 8050 1392
rect 7400 948 7460 970
rect 7518 948 7578 970
rect 7636 948 7696 970
rect 7754 948 7814 970
rect 7872 948 7932 970
rect 7990 948 8050 970
rect 7397 932 7463 948
rect 7397 898 7413 932
rect 7447 898 7463 932
rect 7397 882 7463 898
rect 7515 932 7581 948
rect 7515 898 7531 932
rect 7565 898 7581 932
rect 7515 882 7581 898
rect 7633 932 7699 948
rect 7633 898 7649 932
rect 7683 898 7699 932
rect 7633 882 7699 898
rect 7751 932 7817 948
rect 7751 898 7767 932
rect 7801 898 7817 932
rect 7751 882 7817 898
rect 7869 932 7935 948
rect 7869 898 7885 932
rect 7919 898 7935 932
rect 7869 882 7935 898
rect 7987 932 8053 948
rect 7987 898 8003 932
rect 8037 898 8053 932
rect 7987 882 8053 898
rect 8437 1442 8503 1458
rect 8437 1408 8453 1442
rect 8487 1408 8503 1442
rect 8437 1392 8503 1408
rect 8555 1442 8621 1458
rect 8555 1408 8571 1442
rect 8605 1408 8621 1442
rect 8555 1392 8621 1408
rect 8673 1442 8739 1458
rect 8673 1408 8689 1442
rect 8723 1408 8739 1442
rect 8673 1392 8739 1408
rect 8791 1442 8857 1458
rect 8791 1408 8807 1442
rect 8841 1408 8857 1442
rect 8791 1392 8857 1408
rect 8909 1442 8975 1458
rect 8909 1408 8925 1442
rect 8959 1408 8975 1442
rect 8909 1392 8975 1408
rect 9027 1442 9093 1458
rect 9027 1408 9043 1442
rect 9077 1408 9093 1442
rect 9027 1392 9093 1408
rect 8440 1370 8500 1392
rect 8558 1370 8618 1392
rect 8676 1370 8736 1392
rect 8794 1370 8854 1392
rect 8912 1370 8972 1392
rect 9030 1370 9090 1392
rect 8440 948 8500 970
rect 8558 948 8618 970
rect 8676 948 8736 970
rect 8794 948 8854 970
rect 8912 948 8972 970
rect 9030 948 9090 970
rect 8437 932 8503 948
rect 8437 898 8453 932
rect 8487 898 8503 932
rect 8437 882 8503 898
rect 8555 932 8621 948
rect 8555 898 8571 932
rect 8605 898 8621 932
rect 8555 882 8621 898
rect 8673 932 8739 948
rect 8673 898 8689 932
rect 8723 898 8739 932
rect 8673 882 8739 898
rect 8791 932 8857 948
rect 8791 898 8807 932
rect 8841 898 8857 932
rect 8791 882 8857 898
rect 8909 932 8975 948
rect 8909 898 8925 932
rect 8959 898 8975 932
rect 8909 882 8975 898
rect 9027 932 9093 948
rect 9027 898 9043 932
rect 9077 898 9093 932
rect 9027 882 9093 898
rect 9477 1442 9543 1458
rect 9477 1408 9493 1442
rect 9527 1408 9543 1442
rect 9477 1392 9543 1408
rect 9595 1442 9661 1458
rect 9595 1408 9611 1442
rect 9645 1408 9661 1442
rect 9595 1392 9661 1408
rect 9713 1442 9779 1458
rect 9713 1408 9729 1442
rect 9763 1408 9779 1442
rect 9713 1392 9779 1408
rect 9831 1442 9897 1458
rect 9831 1408 9847 1442
rect 9881 1408 9897 1442
rect 9831 1392 9897 1408
rect 9949 1442 10015 1458
rect 9949 1408 9965 1442
rect 9999 1408 10015 1442
rect 9949 1392 10015 1408
rect 10067 1442 10133 1458
rect 10067 1408 10083 1442
rect 10117 1408 10133 1442
rect 10067 1392 10133 1408
rect 9480 1370 9540 1392
rect 9598 1370 9658 1392
rect 9716 1370 9776 1392
rect 9834 1370 9894 1392
rect 9952 1370 10012 1392
rect 10070 1370 10130 1392
rect 9480 948 9540 970
rect 9598 948 9658 970
rect 9716 948 9776 970
rect 9834 948 9894 970
rect 9952 948 10012 970
rect 10070 948 10130 970
rect 9477 932 9543 948
rect 9477 898 9493 932
rect 9527 898 9543 932
rect 9477 882 9543 898
rect 9595 932 9661 948
rect 9595 898 9611 932
rect 9645 898 9661 932
rect 9595 882 9661 898
rect 9713 932 9779 948
rect 9713 898 9729 932
rect 9763 898 9779 932
rect 9713 882 9779 898
rect 9831 932 9897 948
rect 9831 898 9847 932
rect 9881 898 9897 932
rect 9831 882 9897 898
rect 9949 932 10015 948
rect 9949 898 9965 932
rect 9999 898 10015 932
rect 9949 882 10015 898
rect 10067 932 10133 948
rect 10067 898 10083 932
rect 10117 898 10133 932
rect 10067 882 10133 898
rect 10517 1442 10583 1458
rect 10517 1408 10533 1442
rect 10567 1408 10583 1442
rect 10517 1392 10583 1408
rect 10635 1442 10701 1458
rect 10635 1408 10651 1442
rect 10685 1408 10701 1442
rect 10635 1392 10701 1408
rect 10753 1442 10819 1458
rect 10753 1408 10769 1442
rect 10803 1408 10819 1442
rect 10753 1392 10819 1408
rect 10871 1442 10937 1458
rect 10871 1408 10887 1442
rect 10921 1408 10937 1442
rect 10871 1392 10937 1408
rect 10989 1442 11055 1458
rect 10989 1408 11005 1442
rect 11039 1408 11055 1442
rect 10989 1392 11055 1408
rect 11107 1442 11173 1458
rect 11107 1408 11123 1442
rect 11157 1408 11173 1442
rect 11107 1392 11173 1408
rect 10520 1370 10580 1392
rect 10638 1370 10698 1392
rect 10756 1370 10816 1392
rect 10874 1370 10934 1392
rect 10992 1370 11052 1392
rect 11110 1370 11170 1392
rect 10520 948 10580 970
rect 10638 948 10698 970
rect 10756 948 10816 970
rect 10874 948 10934 970
rect 10992 948 11052 970
rect 11110 948 11170 970
rect 10517 932 10583 948
rect 10517 898 10533 932
rect 10567 898 10583 932
rect 10517 882 10583 898
rect 10635 932 10701 948
rect 10635 898 10651 932
rect 10685 898 10701 932
rect 10635 882 10701 898
rect 10753 932 10819 948
rect 10753 898 10769 932
rect 10803 898 10819 932
rect 10753 882 10819 898
rect 10871 932 10937 948
rect 10871 898 10887 932
rect 10921 898 10937 932
rect 10871 882 10937 898
rect 10989 932 11055 948
rect 10989 898 11005 932
rect 11039 898 11055 932
rect 10989 882 11055 898
rect 11107 932 11173 948
rect 11107 898 11123 932
rect 11157 898 11173 932
rect 11107 882 11173 898
rect 11897 1442 11963 1458
rect 11897 1408 11913 1442
rect 11947 1408 11963 1442
rect 11897 1392 11963 1408
rect 12015 1442 12081 1458
rect 12015 1408 12031 1442
rect 12065 1408 12081 1442
rect 12015 1392 12081 1408
rect 12133 1442 12199 1458
rect 12133 1408 12149 1442
rect 12183 1408 12199 1442
rect 12133 1392 12199 1408
rect 12251 1442 12317 1458
rect 12251 1408 12267 1442
rect 12301 1408 12317 1442
rect 12251 1392 12317 1408
rect 12369 1442 12435 1458
rect 12369 1408 12385 1442
rect 12419 1408 12435 1442
rect 12369 1392 12435 1408
rect 12487 1442 12553 1458
rect 12487 1408 12503 1442
rect 12537 1408 12553 1442
rect 12487 1392 12553 1408
rect 11900 1370 11960 1392
rect 12018 1370 12078 1392
rect 12136 1370 12196 1392
rect 12254 1370 12314 1392
rect 12372 1370 12432 1392
rect 12490 1370 12550 1392
rect 11900 948 11960 970
rect 12018 948 12078 970
rect 12136 948 12196 970
rect 12254 948 12314 970
rect 12372 948 12432 970
rect 12490 948 12550 970
rect 11897 932 11963 948
rect 11897 898 11913 932
rect 11947 898 11963 932
rect 11897 882 11963 898
rect 12015 932 12081 948
rect 12015 898 12031 932
rect 12065 898 12081 932
rect 12015 882 12081 898
rect 12133 932 12199 948
rect 12133 898 12149 932
rect 12183 898 12199 932
rect 12133 882 12199 898
rect 12251 932 12317 948
rect 12251 898 12267 932
rect 12301 898 12317 932
rect 12251 882 12317 898
rect 12369 932 12435 948
rect 12369 898 12385 932
rect 12419 898 12435 932
rect 12369 882 12435 898
rect 12487 932 12553 948
rect 12487 898 12503 932
rect 12537 898 12553 932
rect 12487 882 12553 898
rect 12937 1442 13003 1458
rect 12937 1408 12953 1442
rect 12987 1408 13003 1442
rect 12937 1392 13003 1408
rect 13055 1442 13121 1458
rect 13055 1408 13071 1442
rect 13105 1408 13121 1442
rect 13055 1392 13121 1408
rect 13173 1442 13239 1458
rect 13173 1408 13189 1442
rect 13223 1408 13239 1442
rect 13173 1392 13239 1408
rect 13291 1442 13357 1458
rect 13291 1408 13307 1442
rect 13341 1408 13357 1442
rect 13291 1392 13357 1408
rect 13409 1442 13475 1458
rect 13409 1408 13425 1442
rect 13459 1408 13475 1442
rect 13409 1392 13475 1408
rect 13527 1442 13593 1458
rect 13527 1408 13543 1442
rect 13577 1408 13593 1442
rect 13527 1392 13593 1408
rect 12940 1370 13000 1392
rect 13058 1370 13118 1392
rect 13176 1370 13236 1392
rect 13294 1370 13354 1392
rect 13412 1370 13472 1392
rect 13530 1370 13590 1392
rect 12940 948 13000 970
rect 13058 948 13118 970
rect 13176 948 13236 970
rect 13294 948 13354 970
rect 13412 948 13472 970
rect 13530 948 13590 970
rect 12937 932 13003 948
rect 12937 898 12953 932
rect 12987 898 13003 932
rect 12937 882 13003 898
rect 13055 932 13121 948
rect 13055 898 13071 932
rect 13105 898 13121 932
rect 13055 882 13121 898
rect 13173 932 13239 948
rect 13173 898 13189 932
rect 13223 898 13239 932
rect 13173 882 13239 898
rect 13291 932 13357 948
rect 13291 898 13307 932
rect 13341 898 13357 932
rect 13291 882 13357 898
rect 13409 932 13475 948
rect 13409 898 13425 932
rect 13459 898 13475 932
rect 13409 882 13475 898
rect 13527 932 13593 948
rect 13527 898 13543 932
rect 13577 898 13593 932
rect 13527 882 13593 898
rect 13977 1442 14043 1458
rect 13977 1408 13993 1442
rect 14027 1408 14043 1442
rect 13977 1392 14043 1408
rect 14095 1442 14161 1458
rect 14095 1408 14111 1442
rect 14145 1408 14161 1442
rect 14095 1392 14161 1408
rect 14213 1442 14279 1458
rect 14213 1408 14229 1442
rect 14263 1408 14279 1442
rect 14213 1392 14279 1408
rect 14331 1442 14397 1458
rect 14331 1408 14347 1442
rect 14381 1408 14397 1442
rect 14331 1392 14397 1408
rect 14449 1442 14515 1458
rect 14449 1408 14465 1442
rect 14499 1408 14515 1442
rect 14449 1392 14515 1408
rect 14567 1442 14633 1458
rect 14567 1408 14583 1442
rect 14617 1408 14633 1442
rect 14567 1392 14633 1408
rect 13980 1370 14040 1392
rect 14098 1370 14158 1392
rect 14216 1370 14276 1392
rect 14334 1370 14394 1392
rect 14452 1370 14512 1392
rect 14570 1370 14630 1392
rect 13980 948 14040 970
rect 14098 948 14158 970
rect 14216 948 14276 970
rect 14334 948 14394 970
rect 14452 948 14512 970
rect 14570 948 14630 970
rect 13977 932 14043 948
rect 13977 898 13993 932
rect 14027 898 14043 932
rect 13977 882 14043 898
rect 14095 932 14161 948
rect 14095 898 14111 932
rect 14145 898 14161 932
rect 14095 882 14161 898
rect 14213 932 14279 948
rect 14213 898 14229 932
rect 14263 898 14279 932
rect 14213 882 14279 898
rect 14331 932 14397 948
rect 14331 898 14347 932
rect 14381 898 14397 932
rect 14331 882 14397 898
rect 14449 932 14515 948
rect 14449 898 14465 932
rect 14499 898 14515 932
rect 14449 882 14515 898
rect 14567 932 14633 948
rect 14567 898 14583 932
rect 14617 898 14633 932
rect 14567 882 14633 898
rect 15017 1442 15083 1458
rect 15017 1408 15033 1442
rect 15067 1408 15083 1442
rect 15017 1392 15083 1408
rect 15135 1442 15201 1458
rect 15135 1408 15151 1442
rect 15185 1408 15201 1442
rect 15135 1392 15201 1408
rect 15253 1442 15319 1458
rect 15253 1408 15269 1442
rect 15303 1408 15319 1442
rect 15253 1392 15319 1408
rect 15371 1442 15437 1458
rect 15371 1408 15387 1442
rect 15421 1408 15437 1442
rect 15371 1392 15437 1408
rect 15489 1442 15555 1458
rect 15489 1408 15505 1442
rect 15539 1408 15555 1442
rect 15489 1392 15555 1408
rect 15607 1442 15673 1458
rect 15607 1408 15623 1442
rect 15657 1408 15673 1442
rect 15607 1392 15673 1408
rect 15020 1370 15080 1392
rect 15138 1370 15198 1392
rect 15256 1370 15316 1392
rect 15374 1370 15434 1392
rect 15492 1370 15552 1392
rect 15610 1370 15670 1392
rect 15020 948 15080 970
rect 15138 948 15198 970
rect 15256 948 15316 970
rect 15374 948 15434 970
rect 15492 948 15552 970
rect 15610 948 15670 970
rect 15017 932 15083 948
rect 15017 898 15033 932
rect 15067 898 15083 932
rect 15017 882 15083 898
rect 15135 932 15201 948
rect 15135 898 15151 932
rect 15185 898 15201 932
rect 15135 882 15201 898
rect 15253 932 15319 948
rect 15253 898 15269 932
rect 15303 898 15319 932
rect 15253 882 15319 898
rect 15371 932 15437 948
rect 15371 898 15387 932
rect 15421 898 15437 932
rect 15371 882 15437 898
rect 15489 932 15555 948
rect 15489 898 15505 932
rect 15539 898 15555 932
rect 15489 882 15555 898
rect 15607 932 15673 948
rect 15607 898 15623 932
rect 15657 898 15673 932
rect 15607 882 15673 898
rect 16057 1442 16123 1458
rect 16057 1408 16073 1442
rect 16107 1408 16123 1442
rect 16057 1392 16123 1408
rect 16175 1442 16241 1458
rect 16175 1408 16191 1442
rect 16225 1408 16241 1442
rect 16175 1392 16241 1408
rect 16293 1442 16359 1458
rect 16293 1408 16309 1442
rect 16343 1408 16359 1442
rect 16293 1392 16359 1408
rect 16411 1442 16477 1458
rect 16411 1408 16427 1442
rect 16461 1408 16477 1442
rect 16411 1392 16477 1408
rect 16529 1442 16595 1458
rect 16529 1408 16545 1442
rect 16579 1408 16595 1442
rect 16529 1392 16595 1408
rect 16647 1442 16713 1458
rect 16647 1408 16663 1442
rect 16697 1408 16713 1442
rect 16647 1392 16713 1408
rect 16060 1370 16120 1392
rect 16178 1370 16238 1392
rect 16296 1370 16356 1392
rect 16414 1370 16474 1392
rect 16532 1370 16592 1392
rect 16650 1370 16710 1392
rect 16060 948 16120 970
rect 16178 948 16238 970
rect 16296 948 16356 970
rect 16414 948 16474 970
rect 16532 948 16592 970
rect 16650 948 16710 970
rect 16057 932 16123 948
rect 16057 898 16073 932
rect 16107 898 16123 932
rect 16057 882 16123 898
rect 16175 932 16241 948
rect 16175 898 16191 932
rect 16225 898 16241 932
rect 16175 882 16241 898
rect 16293 932 16359 948
rect 16293 898 16309 932
rect 16343 898 16359 932
rect 16293 882 16359 898
rect 16411 932 16477 948
rect 16411 898 16427 932
rect 16461 898 16477 932
rect 16411 882 16477 898
rect 16529 932 16595 948
rect 16529 898 16545 932
rect 16579 898 16595 932
rect 16529 882 16595 898
rect 16647 932 16713 948
rect 16647 898 16663 932
rect 16697 898 16713 932
rect 16647 882 16713 898
rect 17097 1442 17163 1458
rect 17097 1408 17113 1442
rect 17147 1408 17163 1442
rect 17097 1392 17163 1408
rect 17215 1442 17281 1458
rect 17215 1408 17231 1442
rect 17265 1408 17281 1442
rect 17215 1392 17281 1408
rect 17333 1442 17399 1458
rect 17333 1408 17349 1442
rect 17383 1408 17399 1442
rect 17333 1392 17399 1408
rect 17451 1442 17517 1458
rect 17451 1408 17467 1442
rect 17501 1408 17517 1442
rect 17451 1392 17517 1408
rect 17569 1442 17635 1458
rect 17569 1408 17585 1442
rect 17619 1408 17635 1442
rect 17569 1392 17635 1408
rect 17687 1442 17753 1458
rect 17687 1408 17703 1442
rect 17737 1408 17753 1442
rect 17687 1392 17753 1408
rect 17100 1370 17160 1392
rect 17218 1370 17278 1392
rect 17336 1370 17396 1392
rect 17454 1370 17514 1392
rect 17572 1370 17632 1392
rect 17690 1370 17750 1392
rect 17100 948 17160 970
rect 17218 948 17278 970
rect 17336 948 17396 970
rect 17454 948 17514 970
rect 17572 948 17632 970
rect 17690 948 17750 970
rect 17097 932 17163 948
rect 17097 898 17113 932
rect 17147 898 17163 932
rect 17097 882 17163 898
rect 17215 932 17281 948
rect 17215 898 17231 932
rect 17265 898 17281 932
rect 17215 882 17281 898
rect 17333 932 17399 948
rect 17333 898 17349 932
rect 17383 898 17399 932
rect 17333 882 17399 898
rect 17451 932 17517 948
rect 17451 898 17467 932
rect 17501 898 17517 932
rect 17451 882 17517 898
rect 17569 932 17635 948
rect 17569 898 17585 932
rect 17619 898 17635 932
rect 17569 882 17635 898
rect 17687 932 17753 948
rect 17687 898 17703 932
rect 17737 898 17753 932
rect 17687 882 17753 898
rect 18137 1442 18203 1458
rect 18137 1408 18153 1442
rect 18187 1408 18203 1442
rect 18137 1392 18203 1408
rect 18255 1442 18321 1458
rect 18255 1408 18271 1442
rect 18305 1408 18321 1442
rect 18255 1392 18321 1408
rect 18373 1442 18439 1458
rect 18373 1408 18389 1442
rect 18423 1408 18439 1442
rect 18373 1392 18439 1408
rect 18491 1442 18557 1458
rect 18491 1408 18507 1442
rect 18541 1408 18557 1442
rect 18491 1392 18557 1408
rect 18609 1442 18675 1458
rect 18609 1408 18625 1442
rect 18659 1408 18675 1442
rect 18609 1392 18675 1408
rect 18727 1442 18793 1458
rect 18727 1408 18743 1442
rect 18777 1408 18793 1442
rect 18727 1392 18793 1408
rect 18140 1370 18200 1392
rect 18258 1370 18318 1392
rect 18376 1370 18436 1392
rect 18494 1370 18554 1392
rect 18612 1370 18672 1392
rect 18730 1370 18790 1392
rect 18140 948 18200 970
rect 18258 948 18318 970
rect 18376 948 18436 970
rect 18494 948 18554 970
rect 18612 948 18672 970
rect 18730 948 18790 970
rect 18137 932 18203 948
rect 18137 898 18153 932
rect 18187 898 18203 932
rect 18137 882 18203 898
rect 18255 932 18321 948
rect 18255 898 18271 932
rect 18305 898 18321 932
rect 18255 882 18321 898
rect 18373 932 18439 948
rect 18373 898 18389 932
rect 18423 898 18439 932
rect 18373 882 18439 898
rect 18491 932 18557 948
rect 18491 898 18507 932
rect 18541 898 18557 932
rect 18491 882 18557 898
rect 18609 932 18675 948
rect 18609 898 18625 932
rect 18659 898 18675 932
rect 18609 882 18675 898
rect 18727 932 18793 948
rect 18727 898 18743 932
rect 18777 898 18793 932
rect 18727 882 18793 898
rect -7368 18 -7302 34
rect -7368 -16 -7352 18
rect -7318 -16 -7302 18
rect -7368 -32 -7302 -16
rect -7176 18 -7110 34
rect -7176 -16 -7160 18
rect -7126 -16 -7110 18
rect -7350 -54 -7320 -32
rect -7254 -54 -7224 -28
rect -7176 -32 -7110 -16
rect -6984 18 -6918 34
rect -6984 -16 -6968 18
rect -6934 -16 -6918 18
rect -7158 -54 -7128 -32
rect -7062 -54 -7032 -28
rect -6984 -32 -6918 -16
rect -6792 18 -6726 34
rect -6792 -16 -6776 18
rect -6742 -16 -6726 18
rect -6966 -54 -6936 -32
rect -6870 -54 -6840 -28
rect -6792 -32 -6726 -16
rect -6600 18 -6534 34
rect -6600 -16 -6584 18
rect -6550 -16 -6534 18
rect -6774 -54 -6744 -32
rect -6678 -54 -6648 -28
rect -6600 -32 -6534 -16
rect -6582 -54 -6552 -32
rect -6486 -54 -6456 -28
rect -7350 -480 -7320 -454
rect -7254 -476 -7224 -454
rect -7272 -492 -7206 -476
rect -7158 -480 -7128 -454
rect -7062 -476 -7032 -454
rect -7272 -526 -7256 -492
rect -7222 -526 -7206 -492
rect -7272 -542 -7206 -526
rect -7080 -492 -7014 -476
rect -6966 -480 -6936 -454
rect -6870 -476 -6840 -454
rect -7080 -526 -7064 -492
rect -7030 -526 -7014 -492
rect -7080 -542 -7014 -526
rect -6888 -492 -6822 -476
rect -6774 -480 -6744 -454
rect -6678 -476 -6648 -454
rect -6888 -526 -6872 -492
rect -6838 -526 -6822 -492
rect -6888 -542 -6822 -526
rect -6696 -492 -6630 -476
rect -6582 -480 -6552 -454
rect -6486 -476 -6456 -454
rect -6696 -526 -6680 -492
rect -6646 -526 -6630 -492
rect -6696 -542 -6630 -526
rect -6504 -492 -6438 -476
rect -6504 -526 -6488 -492
rect -6454 -526 -6438 -492
rect -6504 -542 -6438 -526
rect -7272 -600 -7206 -584
rect -7272 -634 -7256 -600
rect -7222 -634 -7206 -600
rect -7350 -672 -7320 -646
rect -7272 -650 -7206 -634
rect -7080 -600 -7014 -584
rect -7080 -634 -7064 -600
rect -7030 -634 -7014 -600
rect -7254 -672 -7224 -650
rect -7158 -672 -7128 -646
rect -7080 -650 -7014 -634
rect -6888 -600 -6822 -584
rect -6888 -634 -6872 -600
rect -6838 -634 -6822 -600
rect -7062 -672 -7032 -650
rect -6966 -672 -6936 -646
rect -6888 -650 -6822 -634
rect -6696 -600 -6630 -584
rect -6696 -634 -6680 -600
rect -6646 -634 -6630 -600
rect -6870 -672 -6840 -650
rect -6774 -672 -6744 -646
rect -6696 -650 -6630 -634
rect -6504 -600 -6438 -584
rect -6504 -634 -6488 -600
rect -6454 -634 -6438 -600
rect -6678 -672 -6648 -650
rect -6582 -672 -6552 -646
rect -6504 -650 -6438 -634
rect -6486 -672 -6456 -650
rect -7350 -1094 -7320 -1072
rect -7368 -1110 -7302 -1094
rect -7254 -1098 -7224 -1072
rect -7158 -1094 -7128 -1072
rect -7368 -1144 -7352 -1110
rect -7318 -1144 -7302 -1110
rect -7368 -1160 -7302 -1144
rect -7176 -1110 -7110 -1094
rect -7062 -1098 -7032 -1072
rect -6966 -1094 -6936 -1072
rect -7176 -1144 -7160 -1110
rect -7126 -1144 -7110 -1110
rect -7176 -1160 -7110 -1144
rect -6984 -1110 -6918 -1094
rect -6870 -1098 -6840 -1072
rect -6774 -1094 -6744 -1072
rect -6984 -1144 -6968 -1110
rect -6934 -1144 -6918 -1110
rect -6984 -1160 -6918 -1144
rect -6792 -1110 -6726 -1094
rect -6678 -1098 -6648 -1072
rect -6582 -1094 -6552 -1072
rect -6792 -1144 -6776 -1110
rect -6742 -1144 -6726 -1110
rect -6792 -1160 -6726 -1144
rect -6600 -1110 -6534 -1094
rect -6486 -1098 -6456 -1072
rect -6600 -1144 -6584 -1110
rect -6550 -1144 -6534 -1110
rect -6600 -1160 -6534 -1144
rect -7368 -1818 -7302 -1802
rect -7368 -1852 -7352 -1818
rect -7318 -1852 -7302 -1818
rect -7368 -1868 -7302 -1852
rect -7176 -1818 -7110 -1802
rect -7176 -1852 -7160 -1818
rect -7126 -1852 -7110 -1818
rect -7350 -1890 -7320 -1868
rect -7254 -1890 -7224 -1864
rect -7176 -1868 -7110 -1852
rect -6984 -1818 -6918 -1802
rect -6984 -1852 -6968 -1818
rect -6934 -1852 -6918 -1818
rect -7158 -1890 -7128 -1868
rect -7062 -1890 -7032 -1864
rect -6984 -1868 -6918 -1852
rect -6966 -1890 -6936 -1868
rect -6870 -1890 -6840 -1864
rect -7350 -2316 -7320 -2290
rect -7254 -2312 -7224 -2290
rect -7272 -2328 -7206 -2312
rect -7158 -2316 -7128 -2290
rect -7062 -2312 -7032 -2290
rect -7272 -2362 -7256 -2328
rect -7222 -2362 -7206 -2328
rect -7272 -2378 -7206 -2362
rect -7080 -2328 -7014 -2312
rect -6966 -2316 -6936 -2290
rect -6870 -2312 -6840 -2290
rect -7080 -2362 -7064 -2328
rect -7030 -2362 -7014 -2328
rect -7080 -2378 -7014 -2362
rect -6888 -2328 -6822 -2312
rect -6888 -2362 -6872 -2328
rect -6838 -2362 -6822 -2328
rect -6888 -2378 -6822 -2362
rect -7272 -2436 -7206 -2420
rect -7272 -2470 -7256 -2436
rect -7222 -2470 -7206 -2436
rect -7350 -2508 -7320 -2482
rect -7272 -2486 -7206 -2470
rect -7080 -2436 -7014 -2420
rect -7080 -2470 -7064 -2436
rect -7030 -2470 -7014 -2436
rect -7254 -2508 -7224 -2486
rect -7158 -2508 -7128 -2482
rect -7080 -2486 -7014 -2470
rect -6888 -2436 -6822 -2420
rect -6888 -2470 -6872 -2436
rect -6838 -2470 -6822 -2436
rect -7062 -2508 -7032 -2486
rect -6966 -2508 -6936 -2482
rect -6888 -2486 -6822 -2470
rect -6870 -2508 -6840 -2486
rect -7350 -2930 -7320 -2908
rect -7368 -2946 -7302 -2930
rect -7254 -2934 -7224 -2908
rect -7158 -2930 -7128 -2908
rect -7368 -2980 -7352 -2946
rect -7318 -2980 -7302 -2946
rect -7368 -2996 -7302 -2980
rect -7176 -2946 -7110 -2930
rect -7062 -2934 -7032 -2908
rect -6966 -2930 -6936 -2908
rect -7176 -2980 -7160 -2946
rect -7126 -2980 -7110 -2946
rect -7176 -2996 -7110 -2980
rect -6984 -2946 -6918 -2930
rect -6870 -2934 -6840 -2908
rect -6984 -2980 -6968 -2946
rect -6934 -2980 -6918 -2946
rect -6984 -2996 -6918 -2980
rect -6088 -70 -6000 -54
rect -6088 -1638 -6072 -70
rect -6038 -1638 -6000 -70
rect -6088 -1654 -6000 -1638
rect -5800 -70 -5712 -54
rect -5800 -1638 -5762 -70
rect -5728 -1638 -5712 -70
rect -5800 -1654 -5712 -1638
rect 4266 624 4332 640
rect 4266 590 4282 624
rect 4316 590 4332 624
rect 4266 574 4332 590
rect 4458 624 4524 640
rect 4458 590 4474 624
rect 4508 590 4524 624
rect 4284 552 4314 574
rect 4380 552 4410 578
rect 4458 574 4524 590
rect 4650 624 4716 640
rect 4650 590 4666 624
rect 4700 590 4716 624
rect 4476 552 4506 574
rect 4572 552 4602 578
rect 4650 574 4716 590
rect 4668 552 4698 574
rect 4764 552 4794 578
rect 4284 126 4314 152
rect 4380 130 4410 152
rect 4362 114 4428 130
rect 4476 126 4506 152
rect 4572 130 4602 152
rect 4362 80 4378 114
rect 4412 80 4428 114
rect 4362 64 4428 80
rect 4554 114 4620 130
rect 4668 126 4698 152
rect 4764 130 4794 152
rect 4554 80 4570 114
rect 4604 80 4620 114
rect 4554 64 4620 80
rect 4746 114 4812 130
rect 4746 80 4762 114
rect 4796 80 4812 114
rect 4746 64 4812 80
rect 4362 6 4428 22
rect 4362 -28 4378 6
rect 4412 -28 4428 6
rect 4284 -66 4314 -40
rect 4362 -44 4428 -28
rect 4554 6 4620 22
rect 4554 -28 4570 6
rect 4604 -28 4620 6
rect 4380 -66 4410 -44
rect 4476 -66 4506 -40
rect 4554 -44 4620 -28
rect 4746 6 4812 22
rect 4746 -28 4762 6
rect 4796 -28 4812 6
rect 4572 -66 4602 -44
rect 4668 -66 4698 -40
rect 4746 -44 4812 -28
rect 4764 -66 4794 -44
rect 4284 -488 4314 -466
rect 4266 -504 4332 -488
rect 4380 -492 4410 -466
rect 4476 -488 4506 -466
rect 4266 -538 4282 -504
rect 4316 -538 4332 -504
rect 4266 -554 4332 -538
rect 4458 -504 4524 -488
rect 4572 -492 4602 -466
rect 4668 -488 4698 -466
rect 4458 -538 4474 -504
rect 4508 -538 4524 -504
rect 4458 -554 4524 -538
rect 4650 -504 4716 -488
rect 4764 -492 4794 -466
rect 4650 -538 4666 -504
rect 4700 -538 4716 -504
rect 4650 -554 4716 -538
rect 5306 624 5372 640
rect 5306 590 5322 624
rect 5356 590 5372 624
rect 5306 574 5372 590
rect 5498 624 5564 640
rect 5498 590 5514 624
rect 5548 590 5564 624
rect 5324 552 5354 574
rect 5420 552 5450 578
rect 5498 574 5564 590
rect 5690 624 5756 640
rect 5690 590 5706 624
rect 5740 590 5756 624
rect 5516 552 5546 574
rect 5612 552 5642 578
rect 5690 574 5756 590
rect 5708 552 5738 574
rect 5804 552 5834 578
rect 5324 126 5354 152
rect 5420 130 5450 152
rect 5402 114 5468 130
rect 5516 126 5546 152
rect 5612 130 5642 152
rect 5402 80 5418 114
rect 5452 80 5468 114
rect 5402 64 5468 80
rect 5594 114 5660 130
rect 5708 126 5738 152
rect 5804 130 5834 152
rect 5594 80 5610 114
rect 5644 80 5660 114
rect 5594 64 5660 80
rect 5786 114 5852 130
rect 5786 80 5802 114
rect 5836 80 5852 114
rect 5786 64 5852 80
rect 5402 6 5468 22
rect 5402 -28 5418 6
rect 5452 -28 5468 6
rect 5324 -66 5354 -40
rect 5402 -44 5468 -28
rect 5594 6 5660 22
rect 5594 -28 5610 6
rect 5644 -28 5660 6
rect 5420 -66 5450 -44
rect 5516 -66 5546 -40
rect 5594 -44 5660 -28
rect 5786 6 5852 22
rect 5786 -28 5802 6
rect 5836 -28 5852 6
rect 5612 -66 5642 -44
rect 5708 -66 5738 -40
rect 5786 -44 5852 -28
rect 5804 -66 5834 -44
rect 5324 -488 5354 -466
rect 5306 -504 5372 -488
rect 5420 -492 5450 -466
rect 5516 -488 5546 -466
rect 5306 -538 5322 -504
rect 5356 -538 5372 -504
rect 5306 -554 5372 -538
rect 5498 -504 5564 -488
rect 5612 -492 5642 -466
rect 5708 -488 5738 -466
rect 5498 -538 5514 -504
rect 5548 -538 5564 -504
rect 5498 -554 5564 -538
rect 5690 -504 5756 -488
rect 5804 -492 5834 -466
rect 5690 -538 5706 -504
rect 5740 -538 5756 -504
rect 5690 -554 5756 -538
rect 6346 624 6412 640
rect 6346 590 6362 624
rect 6396 590 6412 624
rect 6346 574 6412 590
rect 6538 624 6604 640
rect 6538 590 6554 624
rect 6588 590 6604 624
rect 6364 552 6394 574
rect 6460 552 6490 578
rect 6538 574 6604 590
rect 6730 624 6796 640
rect 6730 590 6746 624
rect 6780 590 6796 624
rect 6556 552 6586 574
rect 6652 552 6682 578
rect 6730 574 6796 590
rect 6748 552 6778 574
rect 6844 552 6874 578
rect 6364 126 6394 152
rect 6460 130 6490 152
rect 6442 114 6508 130
rect 6556 126 6586 152
rect 6652 130 6682 152
rect 6442 80 6458 114
rect 6492 80 6508 114
rect 6442 64 6508 80
rect 6634 114 6700 130
rect 6748 126 6778 152
rect 6844 130 6874 152
rect 6634 80 6650 114
rect 6684 80 6700 114
rect 6634 64 6700 80
rect 6826 114 6892 130
rect 6826 80 6842 114
rect 6876 80 6892 114
rect 6826 64 6892 80
rect 6442 6 6508 22
rect 6442 -28 6458 6
rect 6492 -28 6508 6
rect 6364 -66 6394 -40
rect 6442 -44 6508 -28
rect 6634 6 6700 22
rect 6634 -28 6650 6
rect 6684 -28 6700 6
rect 6460 -66 6490 -44
rect 6556 -66 6586 -40
rect 6634 -44 6700 -28
rect 6826 6 6892 22
rect 6826 -28 6842 6
rect 6876 -28 6892 6
rect 6652 -66 6682 -44
rect 6748 -66 6778 -40
rect 6826 -44 6892 -28
rect 6844 -66 6874 -44
rect 6364 -488 6394 -466
rect 6346 -504 6412 -488
rect 6460 -492 6490 -466
rect 6556 -488 6586 -466
rect 6346 -538 6362 -504
rect 6396 -538 6412 -504
rect 6346 -554 6412 -538
rect 6538 -504 6604 -488
rect 6652 -492 6682 -466
rect 6748 -488 6778 -466
rect 6538 -538 6554 -504
rect 6588 -538 6604 -504
rect 6538 -554 6604 -538
rect 6730 -504 6796 -488
rect 6844 -492 6874 -466
rect 6730 -538 6746 -504
rect 6780 -538 6796 -504
rect 6730 -554 6796 -538
rect 7386 624 7452 640
rect 7386 590 7402 624
rect 7436 590 7452 624
rect 7386 574 7452 590
rect 7578 624 7644 640
rect 7578 590 7594 624
rect 7628 590 7644 624
rect 7404 552 7434 574
rect 7500 552 7530 578
rect 7578 574 7644 590
rect 7770 624 7836 640
rect 7770 590 7786 624
rect 7820 590 7836 624
rect 7596 552 7626 574
rect 7692 552 7722 578
rect 7770 574 7836 590
rect 7788 552 7818 574
rect 7884 552 7914 578
rect 7404 126 7434 152
rect 7500 130 7530 152
rect 7482 114 7548 130
rect 7596 126 7626 152
rect 7692 130 7722 152
rect 7482 80 7498 114
rect 7532 80 7548 114
rect 7482 64 7548 80
rect 7674 114 7740 130
rect 7788 126 7818 152
rect 7884 130 7914 152
rect 7674 80 7690 114
rect 7724 80 7740 114
rect 7674 64 7740 80
rect 7866 114 7932 130
rect 7866 80 7882 114
rect 7916 80 7932 114
rect 7866 64 7932 80
rect 7482 6 7548 22
rect 7482 -28 7498 6
rect 7532 -28 7548 6
rect 7404 -66 7434 -40
rect 7482 -44 7548 -28
rect 7674 6 7740 22
rect 7674 -28 7690 6
rect 7724 -28 7740 6
rect 7500 -66 7530 -44
rect 7596 -66 7626 -40
rect 7674 -44 7740 -28
rect 7866 6 7932 22
rect 7866 -28 7882 6
rect 7916 -28 7932 6
rect 7692 -66 7722 -44
rect 7788 -66 7818 -40
rect 7866 -44 7932 -28
rect 7884 -66 7914 -44
rect 7404 -488 7434 -466
rect 7386 -504 7452 -488
rect 7500 -492 7530 -466
rect 7596 -488 7626 -466
rect 7386 -538 7402 -504
rect 7436 -538 7452 -504
rect 7386 -554 7452 -538
rect 7578 -504 7644 -488
rect 7692 -492 7722 -466
rect 7788 -488 7818 -466
rect 7578 -538 7594 -504
rect 7628 -538 7644 -504
rect 7578 -554 7644 -538
rect 7770 -504 7836 -488
rect 7884 -492 7914 -466
rect 7770 -538 7786 -504
rect 7820 -538 7836 -504
rect 7770 -554 7836 -538
rect 8426 624 8492 640
rect 8426 590 8442 624
rect 8476 590 8492 624
rect 8426 574 8492 590
rect 8618 624 8684 640
rect 8618 590 8634 624
rect 8668 590 8684 624
rect 8444 552 8474 574
rect 8540 552 8570 578
rect 8618 574 8684 590
rect 8810 624 8876 640
rect 8810 590 8826 624
rect 8860 590 8876 624
rect 8636 552 8666 574
rect 8732 552 8762 578
rect 8810 574 8876 590
rect 8828 552 8858 574
rect 8924 552 8954 578
rect 8444 126 8474 152
rect 8540 130 8570 152
rect 8522 114 8588 130
rect 8636 126 8666 152
rect 8732 130 8762 152
rect 8522 80 8538 114
rect 8572 80 8588 114
rect 8522 64 8588 80
rect 8714 114 8780 130
rect 8828 126 8858 152
rect 8924 130 8954 152
rect 8714 80 8730 114
rect 8764 80 8780 114
rect 8714 64 8780 80
rect 8906 114 8972 130
rect 8906 80 8922 114
rect 8956 80 8972 114
rect 8906 64 8972 80
rect 8522 6 8588 22
rect 8522 -28 8538 6
rect 8572 -28 8588 6
rect 8444 -66 8474 -40
rect 8522 -44 8588 -28
rect 8714 6 8780 22
rect 8714 -28 8730 6
rect 8764 -28 8780 6
rect 8540 -66 8570 -44
rect 8636 -66 8666 -40
rect 8714 -44 8780 -28
rect 8906 6 8972 22
rect 8906 -28 8922 6
rect 8956 -28 8972 6
rect 8732 -66 8762 -44
rect 8828 -66 8858 -40
rect 8906 -44 8972 -28
rect 8924 -66 8954 -44
rect 8444 -488 8474 -466
rect 8426 -504 8492 -488
rect 8540 -492 8570 -466
rect 8636 -488 8666 -466
rect 8426 -538 8442 -504
rect 8476 -538 8492 -504
rect 8426 -554 8492 -538
rect 8618 -504 8684 -488
rect 8732 -492 8762 -466
rect 8828 -488 8858 -466
rect 8618 -538 8634 -504
rect 8668 -538 8684 -504
rect 8618 -554 8684 -538
rect 8810 -504 8876 -488
rect 8924 -492 8954 -466
rect 8810 -538 8826 -504
rect 8860 -538 8876 -504
rect 8810 -554 8876 -538
rect 9466 624 9532 640
rect 9466 590 9482 624
rect 9516 590 9532 624
rect 9466 574 9532 590
rect 9658 624 9724 640
rect 9658 590 9674 624
rect 9708 590 9724 624
rect 9484 552 9514 574
rect 9580 552 9610 578
rect 9658 574 9724 590
rect 9850 624 9916 640
rect 9850 590 9866 624
rect 9900 590 9916 624
rect 9676 552 9706 574
rect 9772 552 9802 578
rect 9850 574 9916 590
rect 9868 552 9898 574
rect 9964 552 9994 578
rect 9484 126 9514 152
rect 9580 130 9610 152
rect 9562 114 9628 130
rect 9676 126 9706 152
rect 9772 130 9802 152
rect 9562 80 9578 114
rect 9612 80 9628 114
rect 9562 64 9628 80
rect 9754 114 9820 130
rect 9868 126 9898 152
rect 9964 130 9994 152
rect 9754 80 9770 114
rect 9804 80 9820 114
rect 9754 64 9820 80
rect 9946 114 10012 130
rect 9946 80 9962 114
rect 9996 80 10012 114
rect 9946 64 10012 80
rect 9562 6 9628 22
rect 9562 -28 9578 6
rect 9612 -28 9628 6
rect 9484 -66 9514 -40
rect 9562 -44 9628 -28
rect 9754 6 9820 22
rect 9754 -28 9770 6
rect 9804 -28 9820 6
rect 9580 -66 9610 -44
rect 9676 -66 9706 -40
rect 9754 -44 9820 -28
rect 9946 6 10012 22
rect 9946 -28 9962 6
rect 9996 -28 10012 6
rect 9772 -66 9802 -44
rect 9868 -66 9898 -40
rect 9946 -44 10012 -28
rect 9964 -66 9994 -44
rect 9484 -488 9514 -466
rect 9466 -504 9532 -488
rect 9580 -492 9610 -466
rect 9676 -488 9706 -466
rect 9466 -538 9482 -504
rect 9516 -538 9532 -504
rect 9466 -554 9532 -538
rect 9658 -504 9724 -488
rect 9772 -492 9802 -466
rect 9868 -488 9898 -466
rect 9658 -538 9674 -504
rect 9708 -538 9724 -504
rect 9658 -554 9724 -538
rect 9850 -504 9916 -488
rect 9964 -492 9994 -466
rect 9850 -538 9866 -504
rect 9900 -538 9916 -504
rect 9850 -554 9916 -538
rect 10506 624 10572 640
rect 10506 590 10522 624
rect 10556 590 10572 624
rect 10506 574 10572 590
rect 10698 624 10764 640
rect 10698 590 10714 624
rect 10748 590 10764 624
rect 10524 552 10554 574
rect 10620 552 10650 578
rect 10698 574 10764 590
rect 10890 624 10956 640
rect 10890 590 10906 624
rect 10940 590 10956 624
rect 10716 552 10746 574
rect 10812 552 10842 578
rect 10890 574 10956 590
rect 10908 552 10938 574
rect 11004 552 11034 578
rect 10524 126 10554 152
rect 10620 130 10650 152
rect 10602 114 10668 130
rect 10716 126 10746 152
rect 10812 130 10842 152
rect 10602 80 10618 114
rect 10652 80 10668 114
rect 10602 64 10668 80
rect 10794 114 10860 130
rect 10908 126 10938 152
rect 11004 130 11034 152
rect 10794 80 10810 114
rect 10844 80 10860 114
rect 10794 64 10860 80
rect 10986 114 11052 130
rect 10986 80 11002 114
rect 11036 80 11052 114
rect 10986 64 11052 80
rect 10602 6 10668 22
rect 10602 -28 10618 6
rect 10652 -28 10668 6
rect 10524 -66 10554 -40
rect 10602 -44 10668 -28
rect 10794 6 10860 22
rect 10794 -28 10810 6
rect 10844 -28 10860 6
rect 10620 -66 10650 -44
rect 10716 -66 10746 -40
rect 10794 -44 10860 -28
rect 10986 6 11052 22
rect 10986 -28 11002 6
rect 11036 -28 11052 6
rect 10812 -66 10842 -44
rect 10908 -66 10938 -40
rect 10986 -44 11052 -28
rect 11004 -66 11034 -44
rect 10524 -488 10554 -466
rect 10506 -504 10572 -488
rect 10620 -492 10650 -466
rect 10716 -488 10746 -466
rect 10506 -538 10522 -504
rect 10556 -538 10572 -504
rect 10506 -554 10572 -538
rect 10698 -504 10764 -488
rect 10812 -492 10842 -466
rect 10908 -488 10938 -466
rect 10698 -538 10714 -504
rect 10748 -538 10764 -504
rect 10698 -554 10764 -538
rect 10890 -504 10956 -488
rect 11004 -492 11034 -466
rect 10890 -538 10906 -504
rect 10940 -538 10956 -504
rect 10890 -554 10956 -538
rect 11886 624 11952 640
rect 11886 590 11902 624
rect 11936 590 11952 624
rect 11886 574 11952 590
rect 12078 624 12144 640
rect 12078 590 12094 624
rect 12128 590 12144 624
rect 11904 552 11934 574
rect 12000 552 12030 578
rect 12078 574 12144 590
rect 12270 624 12336 640
rect 12270 590 12286 624
rect 12320 590 12336 624
rect 12096 552 12126 574
rect 12192 552 12222 578
rect 12270 574 12336 590
rect 12288 552 12318 574
rect 12384 552 12414 578
rect 11904 126 11934 152
rect 12000 130 12030 152
rect 11982 114 12048 130
rect 12096 126 12126 152
rect 12192 130 12222 152
rect 11982 80 11998 114
rect 12032 80 12048 114
rect 11982 64 12048 80
rect 12174 114 12240 130
rect 12288 126 12318 152
rect 12384 130 12414 152
rect 12174 80 12190 114
rect 12224 80 12240 114
rect 12174 64 12240 80
rect 12366 114 12432 130
rect 12366 80 12382 114
rect 12416 80 12432 114
rect 12366 64 12432 80
rect 11982 6 12048 22
rect 11982 -28 11998 6
rect 12032 -28 12048 6
rect 11904 -66 11934 -40
rect 11982 -44 12048 -28
rect 12174 6 12240 22
rect 12174 -28 12190 6
rect 12224 -28 12240 6
rect 12000 -66 12030 -44
rect 12096 -66 12126 -40
rect 12174 -44 12240 -28
rect 12366 6 12432 22
rect 12366 -28 12382 6
rect 12416 -28 12432 6
rect 12192 -66 12222 -44
rect 12288 -66 12318 -40
rect 12366 -44 12432 -28
rect 12384 -66 12414 -44
rect 11904 -488 11934 -466
rect 11886 -504 11952 -488
rect 12000 -492 12030 -466
rect 12096 -488 12126 -466
rect 11886 -538 11902 -504
rect 11936 -538 11952 -504
rect 11886 -554 11952 -538
rect 12078 -504 12144 -488
rect 12192 -492 12222 -466
rect 12288 -488 12318 -466
rect 12078 -538 12094 -504
rect 12128 -538 12144 -504
rect 12078 -554 12144 -538
rect 12270 -504 12336 -488
rect 12384 -492 12414 -466
rect 12270 -538 12286 -504
rect 12320 -538 12336 -504
rect 12270 -554 12336 -538
rect 12926 624 12992 640
rect 12926 590 12942 624
rect 12976 590 12992 624
rect 12926 574 12992 590
rect 13118 624 13184 640
rect 13118 590 13134 624
rect 13168 590 13184 624
rect 12944 552 12974 574
rect 13040 552 13070 578
rect 13118 574 13184 590
rect 13310 624 13376 640
rect 13310 590 13326 624
rect 13360 590 13376 624
rect 13136 552 13166 574
rect 13232 552 13262 578
rect 13310 574 13376 590
rect 13328 552 13358 574
rect 13424 552 13454 578
rect 12944 126 12974 152
rect 13040 130 13070 152
rect 13022 114 13088 130
rect 13136 126 13166 152
rect 13232 130 13262 152
rect 13022 80 13038 114
rect 13072 80 13088 114
rect 13022 64 13088 80
rect 13214 114 13280 130
rect 13328 126 13358 152
rect 13424 130 13454 152
rect 13214 80 13230 114
rect 13264 80 13280 114
rect 13214 64 13280 80
rect 13406 114 13472 130
rect 13406 80 13422 114
rect 13456 80 13472 114
rect 13406 64 13472 80
rect 13022 6 13088 22
rect 13022 -28 13038 6
rect 13072 -28 13088 6
rect 12944 -66 12974 -40
rect 13022 -44 13088 -28
rect 13214 6 13280 22
rect 13214 -28 13230 6
rect 13264 -28 13280 6
rect 13040 -66 13070 -44
rect 13136 -66 13166 -40
rect 13214 -44 13280 -28
rect 13406 6 13472 22
rect 13406 -28 13422 6
rect 13456 -28 13472 6
rect 13232 -66 13262 -44
rect 13328 -66 13358 -40
rect 13406 -44 13472 -28
rect 13424 -66 13454 -44
rect 12944 -488 12974 -466
rect 12926 -504 12992 -488
rect 13040 -492 13070 -466
rect 13136 -488 13166 -466
rect 12926 -538 12942 -504
rect 12976 -538 12992 -504
rect 12926 -554 12992 -538
rect 13118 -504 13184 -488
rect 13232 -492 13262 -466
rect 13328 -488 13358 -466
rect 13118 -538 13134 -504
rect 13168 -538 13184 -504
rect 13118 -554 13184 -538
rect 13310 -504 13376 -488
rect 13424 -492 13454 -466
rect 13310 -538 13326 -504
rect 13360 -538 13376 -504
rect 13310 -554 13376 -538
rect 13966 624 14032 640
rect 13966 590 13982 624
rect 14016 590 14032 624
rect 13966 574 14032 590
rect 14158 624 14224 640
rect 14158 590 14174 624
rect 14208 590 14224 624
rect 13984 552 14014 574
rect 14080 552 14110 578
rect 14158 574 14224 590
rect 14350 624 14416 640
rect 14350 590 14366 624
rect 14400 590 14416 624
rect 14176 552 14206 574
rect 14272 552 14302 578
rect 14350 574 14416 590
rect 14368 552 14398 574
rect 14464 552 14494 578
rect 13984 126 14014 152
rect 14080 130 14110 152
rect 14062 114 14128 130
rect 14176 126 14206 152
rect 14272 130 14302 152
rect 14062 80 14078 114
rect 14112 80 14128 114
rect 14062 64 14128 80
rect 14254 114 14320 130
rect 14368 126 14398 152
rect 14464 130 14494 152
rect 14254 80 14270 114
rect 14304 80 14320 114
rect 14254 64 14320 80
rect 14446 114 14512 130
rect 14446 80 14462 114
rect 14496 80 14512 114
rect 14446 64 14512 80
rect 14062 6 14128 22
rect 14062 -28 14078 6
rect 14112 -28 14128 6
rect 13984 -66 14014 -40
rect 14062 -44 14128 -28
rect 14254 6 14320 22
rect 14254 -28 14270 6
rect 14304 -28 14320 6
rect 14080 -66 14110 -44
rect 14176 -66 14206 -40
rect 14254 -44 14320 -28
rect 14446 6 14512 22
rect 14446 -28 14462 6
rect 14496 -28 14512 6
rect 14272 -66 14302 -44
rect 14368 -66 14398 -40
rect 14446 -44 14512 -28
rect 14464 -66 14494 -44
rect 13984 -488 14014 -466
rect 13966 -504 14032 -488
rect 14080 -492 14110 -466
rect 14176 -488 14206 -466
rect 13966 -538 13982 -504
rect 14016 -538 14032 -504
rect 13966 -554 14032 -538
rect 14158 -504 14224 -488
rect 14272 -492 14302 -466
rect 14368 -488 14398 -466
rect 14158 -538 14174 -504
rect 14208 -538 14224 -504
rect 14158 -554 14224 -538
rect 14350 -504 14416 -488
rect 14464 -492 14494 -466
rect 14350 -538 14366 -504
rect 14400 -538 14416 -504
rect 14350 -554 14416 -538
rect 15006 624 15072 640
rect 15006 590 15022 624
rect 15056 590 15072 624
rect 15006 574 15072 590
rect 15198 624 15264 640
rect 15198 590 15214 624
rect 15248 590 15264 624
rect 15024 552 15054 574
rect 15120 552 15150 578
rect 15198 574 15264 590
rect 15390 624 15456 640
rect 15390 590 15406 624
rect 15440 590 15456 624
rect 15216 552 15246 574
rect 15312 552 15342 578
rect 15390 574 15456 590
rect 15408 552 15438 574
rect 15504 552 15534 578
rect 15024 126 15054 152
rect 15120 130 15150 152
rect 15102 114 15168 130
rect 15216 126 15246 152
rect 15312 130 15342 152
rect 15102 80 15118 114
rect 15152 80 15168 114
rect 15102 64 15168 80
rect 15294 114 15360 130
rect 15408 126 15438 152
rect 15504 130 15534 152
rect 15294 80 15310 114
rect 15344 80 15360 114
rect 15294 64 15360 80
rect 15486 114 15552 130
rect 15486 80 15502 114
rect 15536 80 15552 114
rect 15486 64 15552 80
rect 15102 6 15168 22
rect 15102 -28 15118 6
rect 15152 -28 15168 6
rect 15024 -66 15054 -40
rect 15102 -44 15168 -28
rect 15294 6 15360 22
rect 15294 -28 15310 6
rect 15344 -28 15360 6
rect 15120 -66 15150 -44
rect 15216 -66 15246 -40
rect 15294 -44 15360 -28
rect 15486 6 15552 22
rect 15486 -28 15502 6
rect 15536 -28 15552 6
rect 15312 -66 15342 -44
rect 15408 -66 15438 -40
rect 15486 -44 15552 -28
rect 15504 -66 15534 -44
rect 15024 -488 15054 -466
rect 15006 -504 15072 -488
rect 15120 -492 15150 -466
rect 15216 -488 15246 -466
rect 15006 -538 15022 -504
rect 15056 -538 15072 -504
rect 15006 -554 15072 -538
rect 15198 -504 15264 -488
rect 15312 -492 15342 -466
rect 15408 -488 15438 -466
rect 15198 -538 15214 -504
rect 15248 -538 15264 -504
rect 15198 -554 15264 -538
rect 15390 -504 15456 -488
rect 15504 -492 15534 -466
rect 15390 -538 15406 -504
rect 15440 -538 15456 -504
rect 15390 -554 15456 -538
rect 16046 624 16112 640
rect 16046 590 16062 624
rect 16096 590 16112 624
rect 16046 574 16112 590
rect 16238 624 16304 640
rect 16238 590 16254 624
rect 16288 590 16304 624
rect 16064 552 16094 574
rect 16160 552 16190 578
rect 16238 574 16304 590
rect 16430 624 16496 640
rect 16430 590 16446 624
rect 16480 590 16496 624
rect 16256 552 16286 574
rect 16352 552 16382 578
rect 16430 574 16496 590
rect 16448 552 16478 574
rect 16544 552 16574 578
rect 16064 126 16094 152
rect 16160 130 16190 152
rect 16142 114 16208 130
rect 16256 126 16286 152
rect 16352 130 16382 152
rect 16142 80 16158 114
rect 16192 80 16208 114
rect 16142 64 16208 80
rect 16334 114 16400 130
rect 16448 126 16478 152
rect 16544 130 16574 152
rect 16334 80 16350 114
rect 16384 80 16400 114
rect 16334 64 16400 80
rect 16526 114 16592 130
rect 16526 80 16542 114
rect 16576 80 16592 114
rect 16526 64 16592 80
rect 16142 6 16208 22
rect 16142 -28 16158 6
rect 16192 -28 16208 6
rect 16064 -66 16094 -40
rect 16142 -44 16208 -28
rect 16334 6 16400 22
rect 16334 -28 16350 6
rect 16384 -28 16400 6
rect 16160 -66 16190 -44
rect 16256 -66 16286 -40
rect 16334 -44 16400 -28
rect 16526 6 16592 22
rect 16526 -28 16542 6
rect 16576 -28 16592 6
rect 16352 -66 16382 -44
rect 16448 -66 16478 -40
rect 16526 -44 16592 -28
rect 16544 -66 16574 -44
rect 16064 -488 16094 -466
rect 16046 -504 16112 -488
rect 16160 -492 16190 -466
rect 16256 -488 16286 -466
rect 16046 -538 16062 -504
rect 16096 -538 16112 -504
rect 16046 -554 16112 -538
rect 16238 -504 16304 -488
rect 16352 -492 16382 -466
rect 16448 -488 16478 -466
rect 16238 -538 16254 -504
rect 16288 -538 16304 -504
rect 16238 -554 16304 -538
rect 16430 -504 16496 -488
rect 16544 -492 16574 -466
rect 16430 -538 16446 -504
rect 16480 -538 16496 -504
rect 16430 -554 16496 -538
rect 17086 624 17152 640
rect 17086 590 17102 624
rect 17136 590 17152 624
rect 17086 574 17152 590
rect 17278 624 17344 640
rect 17278 590 17294 624
rect 17328 590 17344 624
rect 17104 552 17134 574
rect 17200 552 17230 578
rect 17278 574 17344 590
rect 17470 624 17536 640
rect 17470 590 17486 624
rect 17520 590 17536 624
rect 17296 552 17326 574
rect 17392 552 17422 578
rect 17470 574 17536 590
rect 17488 552 17518 574
rect 17584 552 17614 578
rect 17104 126 17134 152
rect 17200 130 17230 152
rect 17182 114 17248 130
rect 17296 126 17326 152
rect 17392 130 17422 152
rect 17182 80 17198 114
rect 17232 80 17248 114
rect 17182 64 17248 80
rect 17374 114 17440 130
rect 17488 126 17518 152
rect 17584 130 17614 152
rect 17374 80 17390 114
rect 17424 80 17440 114
rect 17374 64 17440 80
rect 17566 114 17632 130
rect 17566 80 17582 114
rect 17616 80 17632 114
rect 17566 64 17632 80
rect 17182 6 17248 22
rect 17182 -28 17198 6
rect 17232 -28 17248 6
rect 17104 -66 17134 -40
rect 17182 -44 17248 -28
rect 17374 6 17440 22
rect 17374 -28 17390 6
rect 17424 -28 17440 6
rect 17200 -66 17230 -44
rect 17296 -66 17326 -40
rect 17374 -44 17440 -28
rect 17566 6 17632 22
rect 17566 -28 17582 6
rect 17616 -28 17632 6
rect 17392 -66 17422 -44
rect 17488 -66 17518 -40
rect 17566 -44 17632 -28
rect 17584 -66 17614 -44
rect 17104 -488 17134 -466
rect 17086 -504 17152 -488
rect 17200 -492 17230 -466
rect 17296 -488 17326 -466
rect 17086 -538 17102 -504
rect 17136 -538 17152 -504
rect 17086 -554 17152 -538
rect 17278 -504 17344 -488
rect 17392 -492 17422 -466
rect 17488 -488 17518 -466
rect 17278 -538 17294 -504
rect 17328 -538 17344 -504
rect 17278 -554 17344 -538
rect 17470 -504 17536 -488
rect 17584 -492 17614 -466
rect 17470 -538 17486 -504
rect 17520 -538 17536 -504
rect 17470 -554 17536 -538
rect 18126 624 18192 640
rect 18126 590 18142 624
rect 18176 590 18192 624
rect 18126 574 18192 590
rect 18318 624 18384 640
rect 18318 590 18334 624
rect 18368 590 18384 624
rect 18144 552 18174 574
rect 18240 552 18270 578
rect 18318 574 18384 590
rect 18510 624 18576 640
rect 18510 590 18526 624
rect 18560 590 18576 624
rect 18336 552 18366 574
rect 18432 552 18462 578
rect 18510 574 18576 590
rect 18528 552 18558 574
rect 18624 552 18654 578
rect 18144 126 18174 152
rect 18240 130 18270 152
rect 18222 114 18288 130
rect 18336 126 18366 152
rect 18432 130 18462 152
rect 18222 80 18238 114
rect 18272 80 18288 114
rect 18222 64 18288 80
rect 18414 114 18480 130
rect 18528 126 18558 152
rect 18624 130 18654 152
rect 18414 80 18430 114
rect 18464 80 18480 114
rect 18414 64 18480 80
rect 18606 114 18672 130
rect 18606 80 18622 114
rect 18656 80 18672 114
rect 18606 64 18672 80
rect 18222 6 18288 22
rect 18222 -28 18238 6
rect 18272 -28 18288 6
rect 18144 -66 18174 -40
rect 18222 -44 18288 -28
rect 18414 6 18480 22
rect 18414 -28 18430 6
rect 18464 -28 18480 6
rect 18240 -66 18270 -44
rect 18336 -66 18366 -40
rect 18414 -44 18480 -28
rect 18606 6 18672 22
rect 18606 -28 18622 6
rect 18656 -28 18672 6
rect 18432 -66 18462 -44
rect 18528 -66 18558 -40
rect 18606 -44 18672 -28
rect 18624 -66 18654 -44
rect 18144 -488 18174 -466
rect 18126 -504 18192 -488
rect 18240 -492 18270 -466
rect 18336 -488 18366 -466
rect 18126 -538 18142 -504
rect 18176 -538 18192 -504
rect 18126 -554 18192 -538
rect 18318 -504 18384 -488
rect 18432 -492 18462 -466
rect 18528 -488 18558 -466
rect 18318 -538 18334 -504
rect 18368 -538 18384 -504
rect 18318 -554 18384 -538
rect 18510 -504 18576 -488
rect 18624 -492 18654 -466
rect 18510 -538 18526 -504
rect 18560 -538 18576 -504
rect 18510 -554 18576 -538
rect 4277 -798 4343 -782
rect 4277 -832 4293 -798
rect 4327 -832 4343 -798
rect 4277 -848 4343 -832
rect 4395 -798 4461 -782
rect 4395 -832 4411 -798
rect 4445 -832 4461 -798
rect 4395 -848 4461 -832
rect 4513 -798 4579 -782
rect 4513 -832 4529 -798
rect 4563 -832 4579 -798
rect 4513 -848 4579 -832
rect 4631 -798 4697 -782
rect 4631 -832 4647 -798
rect 4681 -832 4697 -798
rect 4631 -848 4697 -832
rect 4749 -798 4815 -782
rect 4749 -832 4765 -798
rect 4799 -832 4815 -798
rect 4749 -848 4815 -832
rect 4867 -798 4933 -782
rect 4867 -832 4883 -798
rect 4917 -832 4933 -798
rect 4867 -848 4933 -832
rect 4280 -870 4340 -848
rect 4398 -870 4458 -848
rect 4516 -870 4576 -848
rect 4634 -870 4694 -848
rect 4752 -870 4812 -848
rect 4870 -870 4930 -848
rect 4280 -1292 4340 -1270
rect 4398 -1292 4458 -1270
rect 4516 -1292 4576 -1270
rect 4634 -1292 4694 -1270
rect 4752 -1292 4812 -1270
rect 4870 -1292 4930 -1270
rect 4277 -1308 4343 -1292
rect 4277 -1342 4293 -1308
rect 4327 -1342 4343 -1308
rect 4277 -1358 4343 -1342
rect 4395 -1308 4461 -1292
rect 4395 -1342 4411 -1308
rect 4445 -1342 4461 -1308
rect 4395 -1358 4461 -1342
rect 4513 -1308 4579 -1292
rect 4513 -1342 4529 -1308
rect 4563 -1342 4579 -1308
rect 4513 -1358 4579 -1342
rect 4631 -1308 4697 -1292
rect 4631 -1342 4647 -1308
rect 4681 -1342 4697 -1308
rect 4631 -1358 4697 -1342
rect 4749 -1308 4815 -1292
rect 4749 -1342 4765 -1308
rect 4799 -1342 4815 -1308
rect 4749 -1358 4815 -1342
rect 4867 -1308 4933 -1292
rect 4867 -1342 4883 -1308
rect 4917 -1342 4933 -1308
rect 4867 -1358 4933 -1342
rect 5317 -798 5383 -782
rect 5317 -832 5333 -798
rect 5367 -832 5383 -798
rect 5317 -848 5383 -832
rect 5435 -798 5501 -782
rect 5435 -832 5451 -798
rect 5485 -832 5501 -798
rect 5435 -848 5501 -832
rect 5553 -798 5619 -782
rect 5553 -832 5569 -798
rect 5603 -832 5619 -798
rect 5553 -848 5619 -832
rect 5671 -798 5737 -782
rect 5671 -832 5687 -798
rect 5721 -832 5737 -798
rect 5671 -848 5737 -832
rect 5789 -798 5855 -782
rect 5789 -832 5805 -798
rect 5839 -832 5855 -798
rect 5789 -848 5855 -832
rect 5907 -798 5973 -782
rect 5907 -832 5923 -798
rect 5957 -832 5973 -798
rect 5907 -848 5973 -832
rect 5320 -870 5380 -848
rect 5438 -870 5498 -848
rect 5556 -870 5616 -848
rect 5674 -870 5734 -848
rect 5792 -870 5852 -848
rect 5910 -870 5970 -848
rect 5320 -1292 5380 -1270
rect 5438 -1292 5498 -1270
rect 5556 -1292 5616 -1270
rect 5674 -1292 5734 -1270
rect 5792 -1292 5852 -1270
rect 5910 -1292 5970 -1270
rect 5317 -1308 5383 -1292
rect 5317 -1342 5333 -1308
rect 5367 -1342 5383 -1308
rect 5317 -1358 5383 -1342
rect 5435 -1308 5501 -1292
rect 5435 -1342 5451 -1308
rect 5485 -1342 5501 -1308
rect 5435 -1358 5501 -1342
rect 5553 -1308 5619 -1292
rect 5553 -1342 5569 -1308
rect 5603 -1342 5619 -1308
rect 5553 -1358 5619 -1342
rect 5671 -1308 5737 -1292
rect 5671 -1342 5687 -1308
rect 5721 -1342 5737 -1308
rect 5671 -1358 5737 -1342
rect 5789 -1308 5855 -1292
rect 5789 -1342 5805 -1308
rect 5839 -1342 5855 -1308
rect 5789 -1358 5855 -1342
rect 5907 -1308 5973 -1292
rect 5907 -1342 5923 -1308
rect 5957 -1342 5973 -1308
rect 5907 -1358 5973 -1342
rect 6357 -798 6423 -782
rect 6357 -832 6373 -798
rect 6407 -832 6423 -798
rect 6357 -848 6423 -832
rect 6475 -798 6541 -782
rect 6475 -832 6491 -798
rect 6525 -832 6541 -798
rect 6475 -848 6541 -832
rect 6593 -798 6659 -782
rect 6593 -832 6609 -798
rect 6643 -832 6659 -798
rect 6593 -848 6659 -832
rect 6711 -798 6777 -782
rect 6711 -832 6727 -798
rect 6761 -832 6777 -798
rect 6711 -848 6777 -832
rect 6829 -798 6895 -782
rect 6829 -832 6845 -798
rect 6879 -832 6895 -798
rect 6829 -848 6895 -832
rect 6947 -798 7013 -782
rect 6947 -832 6963 -798
rect 6997 -832 7013 -798
rect 6947 -848 7013 -832
rect 6360 -870 6420 -848
rect 6478 -870 6538 -848
rect 6596 -870 6656 -848
rect 6714 -870 6774 -848
rect 6832 -870 6892 -848
rect 6950 -870 7010 -848
rect 6360 -1292 6420 -1270
rect 6478 -1292 6538 -1270
rect 6596 -1292 6656 -1270
rect 6714 -1292 6774 -1270
rect 6832 -1292 6892 -1270
rect 6950 -1292 7010 -1270
rect 6357 -1308 6423 -1292
rect 6357 -1342 6373 -1308
rect 6407 -1342 6423 -1308
rect 6357 -1358 6423 -1342
rect 6475 -1308 6541 -1292
rect 6475 -1342 6491 -1308
rect 6525 -1342 6541 -1308
rect 6475 -1358 6541 -1342
rect 6593 -1308 6659 -1292
rect 6593 -1342 6609 -1308
rect 6643 -1342 6659 -1308
rect 6593 -1358 6659 -1342
rect 6711 -1308 6777 -1292
rect 6711 -1342 6727 -1308
rect 6761 -1342 6777 -1308
rect 6711 -1358 6777 -1342
rect 6829 -1308 6895 -1292
rect 6829 -1342 6845 -1308
rect 6879 -1342 6895 -1308
rect 6829 -1358 6895 -1342
rect 6947 -1308 7013 -1292
rect 6947 -1342 6963 -1308
rect 6997 -1342 7013 -1308
rect 6947 -1358 7013 -1342
rect 7397 -798 7463 -782
rect 7397 -832 7413 -798
rect 7447 -832 7463 -798
rect 7397 -848 7463 -832
rect 7515 -798 7581 -782
rect 7515 -832 7531 -798
rect 7565 -832 7581 -798
rect 7515 -848 7581 -832
rect 7633 -798 7699 -782
rect 7633 -832 7649 -798
rect 7683 -832 7699 -798
rect 7633 -848 7699 -832
rect 7751 -798 7817 -782
rect 7751 -832 7767 -798
rect 7801 -832 7817 -798
rect 7751 -848 7817 -832
rect 7869 -798 7935 -782
rect 7869 -832 7885 -798
rect 7919 -832 7935 -798
rect 7869 -848 7935 -832
rect 7987 -798 8053 -782
rect 7987 -832 8003 -798
rect 8037 -832 8053 -798
rect 7987 -848 8053 -832
rect 7400 -870 7460 -848
rect 7518 -870 7578 -848
rect 7636 -870 7696 -848
rect 7754 -870 7814 -848
rect 7872 -870 7932 -848
rect 7990 -870 8050 -848
rect 7400 -1292 7460 -1270
rect 7518 -1292 7578 -1270
rect 7636 -1292 7696 -1270
rect 7754 -1292 7814 -1270
rect 7872 -1292 7932 -1270
rect 7990 -1292 8050 -1270
rect 7397 -1308 7463 -1292
rect 7397 -1342 7413 -1308
rect 7447 -1342 7463 -1308
rect 7397 -1358 7463 -1342
rect 7515 -1308 7581 -1292
rect 7515 -1342 7531 -1308
rect 7565 -1342 7581 -1308
rect 7515 -1358 7581 -1342
rect 7633 -1308 7699 -1292
rect 7633 -1342 7649 -1308
rect 7683 -1342 7699 -1308
rect 7633 -1358 7699 -1342
rect 7751 -1308 7817 -1292
rect 7751 -1342 7767 -1308
rect 7801 -1342 7817 -1308
rect 7751 -1358 7817 -1342
rect 7869 -1308 7935 -1292
rect 7869 -1342 7885 -1308
rect 7919 -1342 7935 -1308
rect 7869 -1358 7935 -1342
rect 7987 -1308 8053 -1292
rect 7987 -1342 8003 -1308
rect 8037 -1342 8053 -1308
rect 7987 -1358 8053 -1342
rect 8437 -798 8503 -782
rect 8437 -832 8453 -798
rect 8487 -832 8503 -798
rect 8437 -848 8503 -832
rect 8555 -798 8621 -782
rect 8555 -832 8571 -798
rect 8605 -832 8621 -798
rect 8555 -848 8621 -832
rect 8673 -798 8739 -782
rect 8673 -832 8689 -798
rect 8723 -832 8739 -798
rect 8673 -848 8739 -832
rect 8791 -798 8857 -782
rect 8791 -832 8807 -798
rect 8841 -832 8857 -798
rect 8791 -848 8857 -832
rect 8909 -798 8975 -782
rect 8909 -832 8925 -798
rect 8959 -832 8975 -798
rect 8909 -848 8975 -832
rect 9027 -798 9093 -782
rect 9027 -832 9043 -798
rect 9077 -832 9093 -798
rect 9027 -848 9093 -832
rect 8440 -870 8500 -848
rect 8558 -870 8618 -848
rect 8676 -870 8736 -848
rect 8794 -870 8854 -848
rect 8912 -870 8972 -848
rect 9030 -870 9090 -848
rect 8440 -1292 8500 -1270
rect 8558 -1292 8618 -1270
rect 8676 -1292 8736 -1270
rect 8794 -1292 8854 -1270
rect 8912 -1292 8972 -1270
rect 9030 -1292 9090 -1270
rect 8437 -1308 8503 -1292
rect 8437 -1342 8453 -1308
rect 8487 -1342 8503 -1308
rect 8437 -1358 8503 -1342
rect 8555 -1308 8621 -1292
rect 8555 -1342 8571 -1308
rect 8605 -1342 8621 -1308
rect 8555 -1358 8621 -1342
rect 8673 -1308 8739 -1292
rect 8673 -1342 8689 -1308
rect 8723 -1342 8739 -1308
rect 8673 -1358 8739 -1342
rect 8791 -1308 8857 -1292
rect 8791 -1342 8807 -1308
rect 8841 -1342 8857 -1308
rect 8791 -1358 8857 -1342
rect 8909 -1308 8975 -1292
rect 8909 -1342 8925 -1308
rect 8959 -1342 8975 -1308
rect 8909 -1358 8975 -1342
rect 9027 -1308 9093 -1292
rect 9027 -1342 9043 -1308
rect 9077 -1342 9093 -1308
rect 9027 -1358 9093 -1342
rect 9477 -798 9543 -782
rect 9477 -832 9493 -798
rect 9527 -832 9543 -798
rect 9477 -848 9543 -832
rect 9595 -798 9661 -782
rect 9595 -832 9611 -798
rect 9645 -832 9661 -798
rect 9595 -848 9661 -832
rect 9713 -798 9779 -782
rect 9713 -832 9729 -798
rect 9763 -832 9779 -798
rect 9713 -848 9779 -832
rect 9831 -798 9897 -782
rect 9831 -832 9847 -798
rect 9881 -832 9897 -798
rect 9831 -848 9897 -832
rect 9949 -798 10015 -782
rect 9949 -832 9965 -798
rect 9999 -832 10015 -798
rect 9949 -848 10015 -832
rect 10067 -798 10133 -782
rect 10067 -832 10083 -798
rect 10117 -832 10133 -798
rect 10067 -848 10133 -832
rect 9480 -870 9540 -848
rect 9598 -870 9658 -848
rect 9716 -870 9776 -848
rect 9834 -870 9894 -848
rect 9952 -870 10012 -848
rect 10070 -870 10130 -848
rect 9480 -1292 9540 -1270
rect 9598 -1292 9658 -1270
rect 9716 -1292 9776 -1270
rect 9834 -1292 9894 -1270
rect 9952 -1292 10012 -1270
rect 10070 -1292 10130 -1270
rect 9477 -1308 9543 -1292
rect 9477 -1342 9493 -1308
rect 9527 -1342 9543 -1308
rect 9477 -1358 9543 -1342
rect 9595 -1308 9661 -1292
rect 9595 -1342 9611 -1308
rect 9645 -1342 9661 -1308
rect 9595 -1358 9661 -1342
rect 9713 -1308 9779 -1292
rect 9713 -1342 9729 -1308
rect 9763 -1342 9779 -1308
rect 9713 -1358 9779 -1342
rect 9831 -1308 9897 -1292
rect 9831 -1342 9847 -1308
rect 9881 -1342 9897 -1308
rect 9831 -1358 9897 -1342
rect 9949 -1308 10015 -1292
rect 9949 -1342 9965 -1308
rect 9999 -1342 10015 -1308
rect 9949 -1358 10015 -1342
rect 10067 -1308 10133 -1292
rect 10067 -1342 10083 -1308
rect 10117 -1342 10133 -1308
rect 10067 -1358 10133 -1342
rect 10517 -798 10583 -782
rect 10517 -832 10533 -798
rect 10567 -832 10583 -798
rect 10517 -848 10583 -832
rect 10635 -798 10701 -782
rect 10635 -832 10651 -798
rect 10685 -832 10701 -798
rect 10635 -848 10701 -832
rect 10753 -798 10819 -782
rect 10753 -832 10769 -798
rect 10803 -832 10819 -798
rect 10753 -848 10819 -832
rect 10871 -798 10937 -782
rect 10871 -832 10887 -798
rect 10921 -832 10937 -798
rect 10871 -848 10937 -832
rect 10989 -798 11055 -782
rect 10989 -832 11005 -798
rect 11039 -832 11055 -798
rect 10989 -848 11055 -832
rect 11107 -798 11173 -782
rect 11107 -832 11123 -798
rect 11157 -832 11173 -798
rect 11107 -848 11173 -832
rect 10520 -870 10580 -848
rect 10638 -870 10698 -848
rect 10756 -870 10816 -848
rect 10874 -870 10934 -848
rect 10992 -870 11052 -848
rect 11110 -870 11170 -848
rect 10520 -1292 10580 -1270
rect 10638 -1292 10698 -1270
rect 10756 -1292 10816 -1270
rect 10874 -1292 10934 -1270
rect 10992 -1292 11052 -1270
rect 11110 -1292 11170 -1270
rect 10517 -1308 10583 -1292
rect 10517 -1342 10533 -1308
rect 10567 -1342 10583 -1308
rect 10517 -1358 10583 -1342
rect 10635 -1308 10701 -1292
rect 10635 -1342 10651 -1308
rect 10685 -1342 10701 -1308
rect 10635 -1358 10701 -1342
rect 10753 -1308 10819 -1292
rect 10753 -1342 10769 -1308
rect 10803 -1342 10819 -1308
rect 10753 -1358 10819 -1342
rect 10871 -1308 10937 -1292
rect 10871 -1342 10887 -1308
rect 10921 -1342 10937 -1308
rect 10871 -1358 10937 -1342
rect 10989 -1308 11055 -1292
rect 10989 -1342 11005 -1308
rect 11039 -1342 11055 -1308
rect 10989 -1358 11055 -1342
rect 11107 -1308 11173 -1292
rect 11107 -1342 11123 -1308
rect 11157 -1342 11173 -1308
rect 11107 -1358 11173 -1342
rect 11897 -798 11963 -782
rect 11897 -832 11913 -798
rect 11947 -832 11963 -798
rect 11897 -848 11963 -832
rect 12015 -798 12081 -782
rect 12015 -832 12031 -798
rect 12065 -832 12081 -798
rect 12015 -848 12081 -832
rect 12133 -798 12199 -782
rect 12133 -832 12149 -798
rect 12183 -832 12199 -798
rect 12133 -848 12199 -832
rect 12251 -798 12317 -782
rect 12251 -832 12267 -798
rect 12301 -832 12317 -798
rect 12251 -848 12317 -832
rect 12369 -798 12435 -782
rect 12369 -832 12385 -798
rect 12419 -832 12435 -798
rect 12369 -848 12435 -832
rect 12487 -798 12553 -782
rect 12487 -832 12503 -798
rect 12537 -832 12553 -798
rect 12487 -848 12553 -832
rect 11900 -870 11960 -848
rect 12018 -870 12078 -848
rect 12136 -870 12196 -848
rect 12254 -870 12314 -848
rect 12372 -870 12432 -848
rect 12490 -870 12550 -848
rect 11900 -1292 11960 -1270
rect 12018 -1292 12078 -1270
rect 12136 -1292 12196 -1270
rect 12254 -1292 12314 -1270
rect 12372 -1292 12432 -1270
rect 12490 -1292 12550 -1270
rect 11897 -1308 11963 -1292
rect 11897 -1342 11913 -1308
rect 11947 -1342 11963 -1308
rect 11897 -1358 11963 -1342
rect 12015 -1308 12081 -1292
rect 12015 -1342 12031 -1308
rect 12065 -1342 12081 -1308
rect 12015 -1358 12081 -1342
rect 12133 -1308 12199 -1292
rect 12133 -1342 12149 -1308
rect 12183 -1342 12199 -1308
rect 12133 -1358 12199 -1342
rect 12251 -1308 12317 -1292
rect 12251 -1342 12267 -1308
rect 12301 -1342 12317 -1308
rect 12251 -1358 12317 -1342
rect 12369 -1308 12435 -1292
rect 12369 -1342 12385 -1308
rect 12419 -1342 12435 -1308
rect 12369 -1358 12435 -1342
rect 12487 -1308 12553 -1292
rect 12487 -1342 12503 -1308
rect 12537 -1342 12553 -1308
rect 12487 -1358 12553 -1342
rect 12937 -798 13003 -782
rect 12937 -832 12953 -798
rect 12987 -832 13003 -798
rect 12937 -848 13003 -832
rect 13055 -798 13121 -782
rect 13055 -832 13071 -798
rect 13105 -832 13121 -798
rect 13055 -848 13121 -832
rect 13173 -798 13239 -782
rect 13173 -832 13189 -798
rect 13223 -832 13239 -798
rect 13173 -848 13239 -832
rect 13291 -798 13357 -782
rect 13291 -832 13307 -798
rect 13341 -832 13357 -798
rect 13291 -848 13357 -832
rect 13409 -798 13475 -782
rect 13409 -832 13425 -798
rect 13459 -832 13475 -798
rect 13409 -848 13475 -832
rect 13527 -798 13593 -782
rect 13527 -832 13543 -798
rect 13577 -832 13593 -798
rect 13527 -848 13593 -832
rect 12940 -870 13000 -848
rect 13058 -870 13118 -848
rect 13176 -870 13236 -848
rect 13294 -870 13354 -848
rect 13412 -870 13472 -848
rect 13530 -870 13590 -848
rect 12940 -1292 13000 -1270
rect 13058 -1292 13118 -1270
rect 13176 -1292 13236 -1270
rect 13294 -1292 13354 -1270
rect 13412 -1292 13472 -1270
rect 13530 -1292 13590 -1270
rect 12937 -1308 13003 -1292
rect 12937 -1342 12953 -1308
rect 12987 -1342 13003 -1308
rect 12937 -1358 13003 -1342
rect 13055 -1308 13121 -1292
rect 13055 -1342 13071 -1308
rect 13105 -1342 13121 -1308
rect 13055 -1358 13121 -1342
rect 13173 -1308 13239 -1292
rect 13173 -1342 13189 -1308
rect 13223 -1342 13239 -1308
rect 13173 -1358 13239 -1342
rect 13291 -1308 13357 -1292
rect 13291 -1342 13307 -1308
rect 13341 -1342 13357 -1308
rect 13291 -1358 13357 -1342
rect 13409 -1308 13475 -1292
rect 13409 -1342 13425 -1308
rect 13459 -1342 13475 -1308
rect 13409 -1358 13475 -1342
rect 13527 -1308 13593 -1292
rect 13527 -1342 13543 -1308
rect 13577 -1342 13593 -1308
rect 13527 -1358 13593 -1342
rect 13977 -798 14043 -782
rect 13977 -832 13993 -798
rect 14027 -832 14043 -798
rect 13977 -848 14043 -832
rect 14095 -798 14161 -782
rect 14095 -832 14111 -798
rect 14145 -832 14161 -798
rect 14095 -848 14161 -832
rect 14213 -798 14279 -782
rect 14213 -832 14229 -798
rect 14263 -832 14279 -798
rect 14213 -848 14279 -832
rect 14331 -798 14397 -782
rect 14331 -832 14347 -798
rect 14381 -832 14397 -798
rect 14331 -848 14397 -832
rect 14449 -798 14515 -782
rect 14449 -832 14465 -798
rect 14499 -832 14515 -798
rect 14449 -848 14515 -832
rect 14567 -798 14633 -782
rect 14567 -832 14583 -798
rect 14617 -832 14633 -798
rect 14567 -848 14633 -832
rect 13980 -870 14040 -848
rect 14098 -870 14158 -848
rect 14216 -870 14276 -848
rect 14334 -870 14394 -848
rect 14452 -870 14512 -848
rect 14570 -870 14630 -848
rect 13980 -1292 14040 -1270
rect 14098 -1292 14158 -1270
rect 14216 -1292 14276 -1270
rect 14334 -1292 14394 -1270
rect 14452 -1292 14512 -1270
rect 14570 -1292 14630 -1270
rect 13977 -1308 14043 -1292
rect 13977 -1342 13993 -1308
rect 14027 -1342 14043 -1308
rect 13977 -1358 14043 -1342
rect 14095 -1308 14161 -1292
rect 14095 -1342 14111 -1308
rect 14145 -1342 14161 -1308
rect 14095 -1358 14161 -1342
rect 14213 -1308 14279 -1292
rect 14213 -1342 14229 -1308
rect 14263 -1342 14279 -1308
rect 14213 -1358 14279 -1342
rect 14331 -1308 14397 -1292
rect 14331 -1342 14347 -1308
rect 14381 -1342 14397 -1308
rect 14331 -1358 14397 -1342
rect 14449 -1308 14515 -1292
rect 14449 -1342 14465 -1308
rect 14499 -1342 14515 -1308
rect 14449 -1358 14515 -1342
rect 14567 -1308 14633 -1292
rect 14567 -1342 14583 -1308
rect 14617 -1342 14633 -1308
rect 14567 -1358 14633 -1342
rect 15017 -798 15083 -782
rect 15017 -832 15033 -798
rect 15067 -832 15083 -798
rect 15017 -848 15083 -832
rect 15135 -798 15201 -782
rect 15135 -832 15151 -798
rect 15185 -832 15201 -798
rect 15135 -848 15201 -832
rect 15253 -798 15319 -782
rect 15253 -832 15269 -798
rect 15303 -832 15319 -798
rect 15253 -848 15319 -832
rect 15371 -798 15437 -782
rect 15371 -832 15387 -798
rect 15421 -832 15437 -798
rect 15371 -848 15437 -832
rect 15489 -798 15555 -782
rect 15489 -832 15505 -798
rect 15539 -832 15555 -798
rect 15489 -848 15555 -832
rect 15607 -798 15673 -782
rect 15607 -832 15623 -798
rect 15657 -832 15673 -798
rect 15607 -848 15673 -832
rect 15020 -870 15080 -848
rect 15138 -870 15198 -848
rect 15256 -870 15316 -848
rect 15374 -870 15434 -848
rect 15492 -870 15552 -848
rect 15610 -870 15670 -848
rect 15020 -1292 15080 -1270
rect 15138 -1292 15198 -1270
rect 15256 -1292 15316 -1270
rect 15374 -1292 15434 -1270
rect 15492 -1292 15552 -1270
rect 15610 -1292 15670 -1270
rect 15017 -1308 15083 -1292
rect 15017 -1342 15033 -1308
rect 15067 -1342 15083 -1308
rect 15017 -1358 15083 -1342
rect 15135 -1308 15201 -1292
rect 15135 -1342 15151 -1308
rect 15185 -1342 15201 -1308
rect 15135 -1358 15201 -1342
rect 15253 -1308 15319 -1292
rect 15253 -1342 15269 -1308
rect 15303 -1342 15319 -1308
rect 15253 -1358 15319 -1342
rect 15371 -1308 15437 -1292
rect 15371 -1342 15387 -1308
rect 15421 -1342 15437 -1308
rect 15371 -1358 15437 -1342
rect 15489 -1308 15555 -1292
rect 15489 -1342 15505 -1308
rect 15539 -1342 15555 -1308
rect 15489 -1358 15555 -1342
rect 15607 -1308 15673 -1292
rect 15607 -1342 15623 -1308
rect 15657 -1342 15673 -1308
rect 15607 -1358 15673 -1342
rect 16057 -798 16123 -782
rect 16057 -832 16073 -798
rect 16107 -832 16123 -798
rect 16057 -848 16123 -832
rect 16175 -798 16241 -782
rect 16175 -832 16191 -798
rect 16225 -832 16241 -798
rect 16175 -848 16241 -832
rect 16293 -798 16359 -782
rect 16293 -832 16309 -798
rect 16343 -832 16359 -798
rect 16293 -848 16359 -832
rect 16411 -798 16477 -782
rect 16411 -832 16427 -798
rect 16461 -832 16477 -798
rect 16411 -848 16477 -832
rect 16529 -798 16595 -782
rect 16529 -832 16545 -798
rect 16579 -832 16595 -798
rect 16529 -848 16595 -832
rect 16647 -798 16713 -782
rect 16647 -832 16663 -798
rect 16697 -832 16713 -798
rect 16647 -848 16713 -832
rect 16060 -870 16120 -848
rect 16178 -870 16238 -848
rect 16296 -870 16356 -848
rect 16414 -870 16474 -848
rect 16532 -870 16592 -848
rect 16650 -870 16710 -848
rect 16060 -1292 16120 -1270
rect 16178 -1292 16238 -1270
rect 16296 -1292 16356 -1270
rect 16414 -1292 16474 -1270
rect 16532 -1292 16592 -1270
rect 16650 -1292 16710 -1270
rect 16057 -1308 16123 -1292
rect 16057 -1342 16073 -1308
rect 16107 -1342 16123 -1308
rect 16057 -1358 16123 -1342
rect 16175 -1308 16241 -1292
rect 16175 -1342 16191 -1308
rect 16225 -1342 16241 -1308
rect 16175 -1358 16241 -1342
rect 16293 -1308 16359 -1292
rect 16293 -1342 16309 -1308
rect 16343 -1342 16359 -1308
rect 16293 -1358 16359 -1342
rect 16411 -1308 16477 -1292
rect 16411 -1342 16427 -1308
rect 16461 -1342 16477 -1308
rect 16411 -1358 16477 -1342
rect 16529 -1308 16595 -1292
rect 16529 -1342 16545 -1308
rect 16579 -1342 16595 -1308
rect 16529 -1358 16595 -1342
rect 16647 -1308 16713 -1292
rect 16647 -1342 16663 -1308
rect 16697 -1342 16713 -1308
rect 16647 -1358 16713 -1342
rect 17097 -798 17163 -782
rect 17097 -832 17113 -798
rect 17147 -832 17163 -798
rect 17097 -848 17163 -832
rect 17215 -798 17281 -782
rect 17215 -832 17231 -798
rect 17265 -832 17281 -798
rect 17215 -848 17281 -832
rect 17333 -798 17399 -782
rect 17333 -832 17349 -798
rect 17383 -832 17399 -798
rect 17333 -848 17399 -832
rect 17451 -798 17517 -782
rect 17451 -832 17467 -798
rect 17501 -832 17517 -798
rect 17451 -848 17517 -832
rect 17569 -798 17635 -782
rect 17569 -832 17585 -798
rect 17619 -832 17635 -798
rect 17569 -848 17635 -832
rect 17687 -798 17753 -782
rect 17687 -832 17703 -798
rect 17737 -832 17753 -798
rect 17687 -848 17753 -832
rect 17100 -870 17160 -848
rect 17218 -870 17278 -848
rect 17336 -870 17396 -848
rect 17454 -870 17514 -848
rect 17572 -870 17632 -848
rect 17690 -870 17750 -848
rect 17100 -1292 17160 -1270
rect 17218 -1292 17278 -1270
rect 17336 -1292 17396 -1270
rect 17454 -1292 17514 -1270
rect 17572 -1292 17632 -1270
rect 17690 -1292 17750 -1270
rect 17097 -1308 17163 -1292
rect 17097 -1342 17113 -1308
rect 17147 -1342 17163 -1308
rect 17097 -1358 17163 -1342
rect 17215 -1308 17281 -1292
rect 17215 -1342 17231 -1308
rect 17265 -1342 17281 -1308
rect 17215 -1358 17281 -1342
rect 17333 -1308 17399 -1292
rect 17333 -1342 17349 -1308
rect 17383 -1342 17399 -1308
rect 17333 -1358 17399 -1342
rect 17451 -1308 17517 -1292
rect 17451 -1342 17467 -1308
rect 17501 -1342 17517 -1308
rect 17451 -1358 17517 -1342
rect 17569 -1308 17635 -1292
rect 17569 -1342 17585 -1308
rect 17619 -1342 17635 -1308
rect 17569 -1358 17635 -1342
rect 17687 -1308 17753 -1292
rect 17687 -1342 17703 -1308
rect 17737 -1342 17753 -1308
rect 17687 -1358 17753 -1342
rect 18137 -798 18203 -782
rect 18137 -832 18153 -798
rect 18187 -832 18203 -798
rect 18137 -848 18203 -832
rect 18255 -798 18321 -782
rect 18255 -832 18271 -798
rect 18305 -832 18321 -798
rect 18255 -848 18321 -832
rect 18373 -798 18439 -782
rect 18373 -832 18389 -798
rect 18423 -832 18439 -798
rect 18373 -848 18439 -832
rect 18491 -798 18557 -782
rect 18491 -832 18507 -798
rect 18541 -832 18557 -798
rect 18491 -848 18557 -832
rect 18609 -798 18675 -782
rect 18609 -832 18625 -798
rect 18659 -832 18675 -798
rect 18609 -848 18675 -832
rect 18727 -798 18793 -782
rect 18727 -832 18743 -798
rect 18777 -832 18793 -798
rect 18727 -848 18793 -832
rect 18140 -870 18200 -848
rect 18258 -870 18318 -848
rect 18376 -870 18436 -848
rect 18494 -870 18554 -848
rect 18612 -870 18672 -848
rect 18730 -870 18790 -848
rect 18140 -1292 18200 -1270
rect 18258 -1292 18318 -1270
rect 18376 -1292 18436 -1270
rect 18494 -1292 18554 -1270
rect 18612 -1292 18672 -1270
rect 18730 -1292 18790 -1270
rect 18137 -1308 18203 -1292
rect 18137 -1342 18153 -1308
rect 18187 -1342 18203 -1308
rect 18137 -1358 18203 -1342
rect 18255 -1308 18321 -1292
rect 18255 -1342 18271 -1308
rect 18305 -1342 18321 -1308
rect 18255 -1358 18321 -1342
rect 18373 -1308 18439 -1292
rect 18373 -1342 18389 -1308
rect 18423 -1342 18439 -1308
rect 18373 -1358 18439 -1342
rect 18491 -1308 18557 -1292
rect 18491 -1342 18507 -1308
rect 18541 -1342 18557 -1308
rect 18491 -1358 18557 -1342
rect 18609 -1308 18675 -1292
rect 18609 -1342 18625 -1308
rect 18659 -1342 18675 -1308
rect 18609 -1358 18675 -1342
rect 18727 -1308 18793 -1292
rect 18727 -1342 18743 -1308
rect 18777 -1342 18793 -1308
rect 18727 -1358 18793 -1342
rect 4266 -1616 4332 -1600
rect 4266 -1650 4282 -1616
rect 4316 -1650 4332 -1616
rect 4266 -1666 4332 -1650
rect 4458 -1616 4524 -1600
rect 4458 -1650 4474 -1616
rect 4508 -1650 4524 -1616
rect 4284 -1688 4314 -1666
rect 4380 -1688 4410 -1662
rect 4458 -1666 4524 -1650
rect 4650 -1616 4716 -1600
rect 4650 -1650 4666 -1616
rect 4700 -1650 4716 -1616
rect 4476 -1688 4506 -1666
rect 4572 -1688 4602 -1662
rect 4650 -1666 4716 -1650
rect 4668 -1688 4698 -1666
rect 4764 -1688 4794 -1662
rect 4284 -2114 4314 -2088
rect 4380 -2110 4410 -2088
rect 4362 -2126 4428 -2110
rect 4476 -2114 4506 -2088
rect 4572 -2110 4602 -2088
rect 4362 -2160 4378 -2126
rect 4412 -2160 4428 -2126
rect 4362 -2176 4428 -2160
rect 4554 -2126 4620 -2110
rect 4668 -2114 4698 -2088
rect 4764 -2110 4794 -2088
rect 4554 -2160 4570 -2126
rect 4604 -2160 4620 -2126
rect 4554 -2176 4620 -2160
rect 4746 -2126 4812 -2110
rect 4746 -2160 4762 -2126
rect 4796 -2160 4812 -2126
rect 4746 -2176 4812 -2160
rect 4362 -2234 4428 -2218
rect 4362 -2268 4378 -2234
rect 4412 -2268 4428 -2234
rect 4284 -2306 4314 -2280
rect 4362 -2284 4428 -2268
rect 4554 -2234 4620 -2218
rect 4554 -2268 4570 -2234
rect 4604 -2268 4620 -2234
rect 4380 -2306 4410 -2284
rect 4476 -2306 4506 -2280
rect 4554 -2284 4620 -2268
rect 4746 -2234 4812 -2218
rect 4746 -2268 4762 -2234
rect 4796 -2268 4812 -2234
rect 4572 -2306 4602 -2284
rect 4668 -2306 4698 -2280
rect 4746 -2284 4812 -2268
rect 4764 -2306 4794 -2284
rect 4284 -2728 4314 -2706
rect 4266 -2744 4332 -2728
rect 4380 -2732 4410 -2706
rect 4476 -2728 4506 -2706
rect 4266 -2778 4282 -2744
rect 4316 -2778 4332 -2744
rect 4266 -2794 4332 -2778
rect 4458 -2744 4524 -2728
rect 4572 -2732 4602 -2706
rect 4668 -2728 4698 -2706
rect 4458 -2778 4474 -2744
rect 4508 -2778 4524 -2744
rect 4458 -2794 4524 -2778
rect 4650 -2744 4716 -2728
rect 4764 -2732 4794 -2706
rect 4650 -2778 4666 -2744
rect 4700 -2778 4716 -2744
rect 4650 -2794 4716 -2778
rect 5306 -1616 5372 -1600
rect 5306 -1650 5322 -1616
rect 5356 -1650 5372 -1616
rect 5306 -1666 5372 -1650
rect 5498 -1616 5564 -1600
rect 5498 -1650 5514 -1616
rect 5548 -1650 5564 -1616
rect 5324 -1688 5354 -1666
rect 5420 -1688 5450 -1662
rect 5498 -1666 5564 -1650
rect 5690 -1616 5756 -1600
rect 5690 -1650 5706 -1616
rect 5740 -1650 5756 -1616
rect 5516 -1688 5546 -1666
rect 5612 -1688 5642 -1662
rect 5690 -1666 5756 -1650
rect 5708 -1688 5738 -1666
rect 5804 -1688 5834 -1662
rect 5324 -2114 5354 -2088
rect 5420 -2110 5450 -2088
rect 5402 -2126 5468 -2110
rect 5516 -2114 5546 -2088
rect 5612 -2110 5642 -2088
rect 5402 -2160 5418 -2126
rect 5452 -2160 5468 -2126
rect 5402 -2176 5468 -2160
rect 5594 -2126 5660 -2110
rect 5708 -2114 5738 -2088
rect 5804 -2110 5834 -2088
rect 5594 -2160 5610 -2126
rect 5644 -2160 5660 -2126
rect 5594 -2176 5660 -2160
rect 5786 -2126 5852 -2110
rect 5786 -2160 5802 -2126
rect 5836 -2160 5852 -2126
rect 5786 -2176 5852 -2160
rect 5402 -2234 5468 -2218
rect 5402 -2268 5418 -2234
rect 5452 -2268 5468 -2234
rect 5324 -2306 5354 -2280
rect 5402 -2284 5468 -2268
rect 5594 -2234 5660 -2218
rect 5594 -2268 5610 -2234
rect 5644 -2268 5660 -2234
rect 5420 -2306 5450 -2284
rect 5516 -2306 5546 -2280
rect 5594 -2284 5660 -2268
rect 5786 -2234 5852 -2218
rect 5786 -2268 5802 -2234
rect 5836 -2268 5852 -2234
rect 5612 -2306 5642 -2284
rect 5708 -2306 5738 -2280
rect 5786 -2284 5852 -2268
rect 5804 -2306 5834 -2284
rect 5324 -2728 5354 -2706
rect 5306 -2744 5372 -2728
rect 5420 -2732 5450 -2706
rect 5516 -2728 5546 -2706
rect 5306 -2778 5322 -2744
rect 5356 -2778 5372 -2744
rect 5306 -2794 5372 -2778
rect 5498 -2744 5564 -2728
rect 5612 -2732 5642 -2706
rect 5708 -2728 5738 -2706
rect 5498 -2778 5514 -2744
rect 5548 -2778 5564 -2744
rect 5498 -2794 5564 -2778
rect 5690 -2744 5756 -2728
rect 5804 -2732 5834 -2706
rect 5690 -2778 5706 -2744
rect 5740 -2778 5756 -2744
rect 5690 -2794 5756 -2778
rect 6346 -1616 6412 -1600
rect 6346 -1650 6362 -1616
rect 6396 -1650 6412 -1616
rect 6346 -1666 6412 -1650
rect 6538 -1616 6604 -1600
rect 6538 -1650 6554 -1616
rect 6588 -1650 6604 -1616
rect 6364 -1688 6394 -1666
rect 6460 -1688 6490 -1662
rect 6538 -1666 6604 -1650
rect 6730 -1616 6796 -1600
rect 6730 -1650 6746 -1616
rect 6780 -1650 6796 -1616
rect 6556 -1688 6586 -1666
rect 6652 -1688 6682 -1662
rect 6730 -1666 6796 -1650
rect 6748 -1688 6778 -1666
rect 6844 -1688 6874 -1662
rect 6364 -2114 6394 -2088
rect 6460 -2110 6490 -2088
rect 6442 -2126 6508 -2110
rect 6556 -2114 6586 -2088
rect 6652 -2110 6682 -2088
rect 6442 -2160 6458 -2126
rect 6492 -2160 6508 -2126
rect 6442 -2176 6508 -2160
rect 6634 -2126 6700 -2110
rect 6748 -2114 6778 -2088
rect 6844 -2110 6874 -2088
rect 6634 -2160 6650 -2126
rect 6684 -2160 6700 -2126
rect 6634 -2176 6700 -2160
rect 6826 -2126 6892 -2110
rect 6826 -2160 6842 -2126
rect 6876 -2160 6892 -2126
rect 6826 -2176 6892 -2160
rect 6442 -2234 6508 -2218
rect 6442 -2268 6458 -2234
rect 6492 -2268 6508 -2234
rect 6364 -2306 6394 -2280
rect 6442 -2284 6508 -2268
rect 6634 -2234 6700 -2218
rect 6634 -2268 6650 -2234
rect 6684 -2268 6700 -2234
rect 6460 -2306 6490 -2284
rect 6556 -2306 6586 -2280
rect 6634 -2284 6700 -2268
rect 6826 -2234 6892 -2218
rect 6826 -2268 6842 -2234
rect 6876 -2268 6892 -2234
rect 6652 -2306 6682 -2284
rect 6748 -2306 6778 -2280
rect 6826 -2284 6892 -2268
rect 6844 -2306 6874 -2284
rect 6364 -2728 6394 -2706
rect 6346 -2744 6412 -2728
rect 6460 -2732 6490 -2706
rect 6556 -2728 6586 -2706
rect 6346 -2778 6362 -2744
rect 6396 -2778 6412 -2744
rect 6346 -2794 6412 -2778
rect 6538 -2744 6604 -2728
rect 6652 -2732 6682 -2706
rect 6748 -2728 6778 -2706
rect 6538 -2778 6554 -2744
rect 6588 -2778 6604 -2744
rect 6538 -2794 6604 -2778
rect 6730 -2744 6796 -2728
rect 6844 -2732 6874 -2706
rect 6730 -2778 6746 -2744
rect 6780 -2778 6796 -2744
rect 6730 -2794 6796 -2778
rect 7386 -1616 7452 -1600
rect 7386 -1650 7402 -1616
rect 7436 -1650 7452 -1616
rect 7386 -1666 7452 -1650
rect 7578 -1616 7644 -1600
rect 7578 -1650 7594 -1616
rect 7628 -1650 7644 -1616
rect 7404 -1688 7434 -1666
rect 7500 -1688 7530 -1662
rect 7578 -1666 7644 -1650
rect 7770 -1616 7836 -1600
rect 7770 -1650 7786 -1616
rect 7820 -1650 7836 -1616
rect 7596 -1688 7626 -1666
rect 7692 -1688 7722 -1662
rect 7770 -1666 7836 -1650
rect 7788 -1688 7818 -1666
rect 7884 -1688 7914 -1662
rect 7404 -2114 7434 -2088
rect 7500 -2110 7530 -2088
rect 7482 -2126 7548 -2110
rect 7596 -2114 7626 -2088
rect 7692 -2110 7722 -2088
rect 7482 -2160 7498 -2126
rect 7532 -2160 7548 -2126
rect 7482 -2176 7548 -2160
rect 7674 -2126 7740 -2110
rect 7788 -2114 7818 -2088
rect 7884 -2110 7914 -2088
rect 7674 -2160 7690 -2126
rect 7724 -2160 7740 -2126
rect 7674 -2176 7740 -2160
rect 7866 -2126 7932 -2110
rect 7866 -2160 7882 -2126
rect 7916 -2160 7932 -2126
rect 7866 -2176 7932 -2160
rect 7482 -2234 7548 -2218
rect 7482 -2268 7498 -2234
rect 7532 -2268 7548 -2234
rect 7404 -2306 7434 -2280
rect 7482 -2284 7548 -2268
rect 7674 -2234 7740 -2218
rect 7674 -2268 7690 -2234
rect 7724 -2268 7740 -2234
rect 7500 -2306 7530 -2284
rect 7596 -2306 7626 -2280
rect 7674 -2284 7740 -2268
rect 7866 -2234 7932 -2218
rect 7866 -2268 7882 -2234
rect 7916 -2268 7932 -2234
rect 7692 -2306 7722 -2284
rect 7788 -2306 7818 -2280
rect 7866 -2284 7932 -2268
rect 7884 -2306 7914 -2284
rect 7404 -2728 7434 -2706
rect 7386 -2744 7452 -2728
rect 7500 -2732 7530 -2706
rect 7596 -2728 7626 -2706
rect 7386 -2778 7402 -2744
rect 7436 -2778 7452 -2744
rect 7386 -2794 7452 -2778
rect 7578 -2744 7644 -2728
rect 7692 -2732 7722 -2706
rect 7788 -2728 7818 -2706
rect 7578 -2778 7594 -2744
rect 7628 -2778 7644 -2744
rect 7578 -2794 7644 -2778
rect 7770 -2744 7836 -2728
rect 7884 -2732 7914 -2706
rect 7770 -2778 7786 -2744
rect 7820 -2778 7836 -2744
rect 7770 -2794 7836 -2778
rect 8426 -1616 8492 -1600
rect 8426 -1650 8442 -1616
rect 8476 -1650 8492 -1616
rect 8426 -1666 8492 -1650
rect 8618 -1616 8684 -1600
rect 8618 -1650 8634 -1616
rect 8668 -1650 8684 -1616
rect 8444 -1688 8474 -1666
rect 8540 -1688 8570 -1662
rect 8618 -1666 8684 -1650
rect 8810 -1616 8876 -1600
rect 8810 -1650 8826 -1616
rect 8860 -1650 8876 -1616
rect 8636 -1688 8666 -1666
rect 8732 -1688 8762 -1662
rect 8810 -1666 8876 -1650
rect 8828 -1688 8858 -1666
rect 8924 -1688 8954 -1662
rect 8444 -2114 8474 -2088
rect 8540 -2110 8570 -2088
rect 8522 -2126 8588 -2110
rect 8636 -2114 8666 -2088
rect 8732 -2110 8762 -2088
rect 8522 -2160 8538 -2126
rect 8572 -2160 8588 -2126
rect 8522 -2176 8588 -2160
rect 8714 -2126 8780 -2110
rect 8828 -2114 8858 -2088
rect 8924 -2110 8954 -2088
rect 8714 -2160 8730 -2126
rect 8764 -2160 8780 -2126
rect 8714 -2176 8780 -2160
rect 8906 -2126 8972 -2110
rect 8906 -2160 8922 -2126
rect 8956 -2160 8972 -2126
rect 8906 -2176 8972 -2160
rect 8522 -2234 8588 -2218
rect 8522 -2268 8538 -2234
rect 8572 -2268 8588 -2234
rect 8444 -2306 8474 -2280
rect 8522 -2284 8588 -2268
rect 8714 -2234 8780 -2218
rect 8714 -2268 8730 -2234
rect 8764 -2268 8780 -2234
rect 8540 -2306 8570 -2284
rect 8636 -2306 8666 -2280
rect 8714 -2284 8780 -2268
rect 8906 -2234 8972 -2218
rect 8906 -2268 8922 -2234
rect 8956 -2268 8972 -2234
rect 8732 -2306 8762 -2284
rect 8828 -2306 8858 -2280
rect 8906 -2284 8972 -2268
rect 8924 -2306 8954 -2284
rect 8444 -2728 8474 -2706
rect 8426 -2744 8492 -2728
rect 8540 -2732 8570 -2706
rect 8636 -2728 8666 -2706
rect 8426 -2778 8442 -2744
rect 8476 -2778 8492 -2744
rect 8426 -2794 8492 -2778
rect 8618 -2744 8684 -2728
rect 8732 -2732 8762 -2706
rect 8828 -2728 8858 -2706
rect 8618 -2778 8634 -2744
rect 8668 -2778 8684 -2744
rect 8618 -2794 8684 -2778
rect 8810 -2744 8876 -2728
rect 8924 -2732 8954 -2706
rect 8810 -2778 8826 -2744
rect 8860 -2778 8876 -2744
rect 8810 -2794 8876 -2778
rect 11886 -1616 11952 -1600
rect 11886 -1650 11902 -1616
rect 11936 -1650 11952 -1616
rect 11886 -1666 11952 -1650
rect 12078 -1616 12144 -1600
rect 12078 -1650 12094 -1616
rect 12128 -1650 12144 -1616
rect 11904 -1688 11934 -1666
rect 12000 -1688 12030 -1662
rect 12078 -1666 12144 -1650
rect 12270 -1616 12336 -1600
rect 12270 -1650 12286 -1616
rect 12320 -1650 12336 -1616
rect 12096 -1688 12126 -1666
rect 12192 -1688 12222 -1662
rect 12270 -1666 12336 -1650
rect 12288 -1688 12318 -1666
rect 12384 -1688 12414 -1662
rect 11904 -2114 11934 -2088
rect 12000 -2110 12030 -2088
rect 11982 -2126 12048 -2110
rect 12096 -2114 12126 -2088
rect 12192 -2110 12222 -2088
rect 11982 -2160 11998 -2126
rect 12032 -2160 12048 -2126
rect 11982 -2176 12048 -2160
rect 12174 -2126 12240 -2110
rect 12288 -2114 12318 -2088
rect 12384 -2110 12414 -2088
rect 12174 -2160 12190 -2126
rect 12224 -2160 12240 -2126
rect 12174 -2176 12240 -2160
rect 12366 -2126 12432 -2110
rect 12366 -2160 12382 -2126
rect 12416 -2160 12432 -2126
rect 12366 -2176 12432 -2160
rect 11982 -2234 12048 -2218
rect 11982 -2268 11998 -2234
rect 12032 -2268 12048 -2234
rect 11904 -2306 11934 -2280
rect 11982 -2284 12048 -2268
rect 12174 -2234 12240 -2218
rect 12174 -2268 12190 -2234
rect 12224 -2268 12240 -2234
rect 12000 -2306 12030 -2284
rect 12096 -2306 12126 -2280
rect 12174 -2284 12240 -2268
rect 12366 -2234 12432 -2218
rect 12366 -2268 12382 -2234
rect 12416 -2268 12432 -2234
rect 12192 -2306 12222 -2284
rect 12288 -2306 12318 -2280
rect 12366 -2284 12432 -2268
rect 12384 -2306 12414 -2284
rect 11904 -2728 11934 -2706
rect 11886 -2744 11952 -2728
rect 12000 -2732 12030 -2706
rect 12096 -2728 12126 -2706
rect 11886 -2778 11902 -2744
rect 11936 -2778 11952 -2744
rect 11886 -2794 11952 -2778
rect 12078 -2744 12144 -2728
rect 12192 -2732 12222 -2706
rect 12288 -2728 12318 -2706
rect 12078 -2778 12094 -2744
rect 12128 -2778 12144 -2744
rect 12078 -2794 12144 -2778
rect 12270 -2744 12336 -2728
rect 12384 -2732 12414 -2706
rect 12270 -2778 12286 -2744
rect 12320 -2778 12336 -2744
rect 12270 -2794 12336 -2778
rect 12926 -1616 12992 -1600
rect 12926 -1650 12942 -1616
rect 12976 -1650 12992 -1616
rect 12926 -1666 12992 -1650
rect 13118 -1616 13184 -1600
rect 13118 -1650 13134 -1616
rect 13168 -1650 13184 -1616
rect 12944 -1688 12974 -1666
rect 13040 -1688 13070 -1662
rect 13118 -1666 13184 -1650
rect 13310 -1616 13376 -1600
rect 13310 -1650 13326 -1616
rect 13360 -1650 13376 -1616
rect 13136 -1688 13166 -1666
rect 13232 -1688 13262 -1662
rect 13310 -1666 13376 -1650
rect 13328 -1688 13358 -1666
rect 13424 -1688 13454 -1662
rect 12944 -2114 12974 -2088
rect 13040 -2110 13070 -2088
rect 13022 -2126 13088 -2110
rect 13136 -2114 13166 -2088
rect 13232 -2110 13262 -2088
rect 13022 -2160 13038 -2126
rect 13072 -2160 13088 -2126
rect 13022 -2176 13088 -2160
rect 13214 -2126 13280 -2110
rect 13328 -2114 13358 -2088
rect 13424 -2110 13454 -2088
rect 13214 -2160 13230 -2126
rect 13264 -2160 13280 -2126
rect 13214 -2176 13280 -2160
rect 13406 -2126 13472 -2110
rect 13406 -2160 13422 -2126
rect 13456 -2160 13472 -2126
rect 13406 -2176 13472 -2160
rect 13022 -2234 13088 -2218
rect 13022 -2268 13038 -2234
rect 13072 -2268 13088 -2234
rect 12944 -2306 12974 -2280
rect 13022 -2284 13088 -2268
rect 13214 -2234 13280 -2218
rect 13214 -2268 13230 -2234
rect 13264 -2268 13280 -2234
rect 13040 -2306 13070 -2284
rect 13136 -2306 13166 -2280
rect 13214 -2284 13280 -2268
rect 13406 -2234 13472 -2218
rect 13406 -2268 13422 -2234
rect 13456 -2268 13472 -2234
rect 13232 -2306 13262 -2284
rect 13328 -2306 13358 -2280
rect 13406 -2284 13472 -2268
rect 13424 -2306 13454 -2284
rect 12944 -2728 12974 -2706
rect 12926 -2744 12992 -2728
rect 13040 -2732 13070 -2706
rect 13136 -2728 13166 -2706
rect 12926 -2778 12942 -2744
rect 12976 -2778 12992 -2744
rect 12926 -2794 12992 -2778
rect 13118 -2744 13184 -2728
rect 13232 -2732 13262 -2706
rect 13328 -2728 13358 -2706
rect 13118 -2778 13134 -2744
rect 13168 -2778 13184 -2744
rect 13118 -2794 13184 -2778
rect 13310 -2744 13376 -2728
rect 13424 -2732 13454 -2706
rect 13310 -2778 13326 -2744
rect 13360 -2778 13376 -2744
rect 13310 -2794 13376 -2778
rect 13966 -1616 14032 -1600
rect 13966 -1650 13982 -1616
rect 14016 -1650 14032 -1616
rect 13966 -1666 14032 -1650
rect 14158 -1616 14224 -1600
rect 14158 -1650 14174 -1616
rect 14208 -1650 14224 -1616
rect 13984 -1688 14014 -1666
rect 14080 -1688 14110 -1662
rect 14158 -1666 14224 -1650
rect 14350 -1616 14416 -1600
rect 14350 -1650 14366 -1616
rect 14400 -1650 14416 -1616
rect 14176 -1688 14206 -1666
rect 14272 -1688 14302 -1662
rect 14350 -1666 14416 -1650
rect 14368 -1688 14398 -1666
rect 14464 -1688 14494 -1662
rect 13984 -2114 14014 -2088
rect 14080 -2110 14110 -2088
rect 14062 -2126 14128 -2110
rect 14176 -2114 14206 -2088
rect 14272 -2110 14302 -2088
rect 14062 -2160 14078 -2126
rect 14112 -2160 14128 -2126
rect 14062 -2176 14128 -2160
rect 14254 -2126 14320 -2110
rect 14368 -2114 14398 -2088
rect 14464 -2110 14494 -2088
rect 14254 -2160 14270 -2126
rect 14304 -2160 14320 -2126
rect 14254 -2176 14320 -2160
rect 14446 -2126 14512 -2110
rect 14446 -2160 14462 -2126
rect 14496 -2160 14512 -2126
rect 14446 -2176 14512 -2160
rect 14062 -2234 14128 -2218
rect 14062 -2268 14078 -2234
rect 14112 -2268 14128 -2234
rect 13984 -2306 14014 -2280
rect 14062 -2284 14128 -2268
rect 14254 -2234 14320 -2218
rect 14254 -2268 14270 -2234
rect 14304 -2268 14320 -2234
rect 14080 -2306 14110 -2284
rect 14176 -2306 14206 -2280
rect 14254 -2284 14320 -2268
rect 14446 -2234 14512 -2218
rect 14446 -2268 14462 -2234
rect 14496 -2268 14512 -2234
rect 14272 -2306 14302 -2284
rect 14368 -2306 14398 -2280
rect 14446 -2284 14512 -2268
rect 14464 -2306 14494 -2284
rect 13984 -2728 14014 -2706
rect 13966 -2744 14032 -2728
rect 14080 -2732 14110 -2706
rect 14176 -2728 14206 -2706
rect 13966 -2778 13982 -2744
rect 14016 -2778 14032 -2744
rect 13966 -2794 14032 -2778
rect 14158 -2744 14224 -2728
rect 14272 -2732 14302 -2706
rect 14368 -2728 14398 -2706
rect 14158 -2778 14174 -2744
rect 14208 -2778 14224 -2744
rect 14158 -2794 14224 -2778
rect 14350 -2744 14416 -2728
rect 14464 -2732 14494 -2706
rect 14350 -2778 14366 -2744
rect 14400 -2778 14416 -2744
rect 14350 -2794 14416 -2778
rect 15006 -1616 15072 -1600
rect 15006 -1650 15022 -1616
rect 15056 -1650 15072 -1616
rect 15006 -1666 15072 -1650
rect 15198 -1616 15264 -1600
rect 15198 -1650 15214 -1616
rect 15248 -1650 15264 -1616
rect 15024 -1688 15054 -1666
rect 15120 -1688 15150 -1662
rect 15198 -1666 15264 -1650
rect 15390 -1616 15456 -1600
rect 15390 -1650 15406 -1616
rect 15440 -1650 15456 -1616
rect 15216 -1688 15246 -1666
rect 15312 -1688 15342 -1662
rect 15390 -1666 15456 -1650
rect 15408 -1688 15438 -1666
rect 15504 -1688 15534 -1662
rect 15024 -2114 15054 -2088
rect 15120 -2110 15150 -2088
rect 15102 -2126 15168 -2110
rect 15216 -2114 15246 -2088
rect 15312 -2110 15342 -2088
rect 15102 -2160 15118 -2126
rect 15152 -2160 15168 -2126
rect 15102 -2176 15168 -2160
rect 15294 -2126 15360 -2110
rect 15408 -2114 15438 -2088
rect 15504 -2110 15534 -2088
rect 15294 -2160 15310 -2126
rect 15344 -2160 15360 -2126
rect 15294 -2176 15360 -2160
rect 15486 -2126 15552 -2110
rect 15486 -2160 15502 -2126
rect 15536 -2160 15552 -2126
rect 15486 -2176 15552 -2160
rect 15102 -2234 15168 -2218
rect 15102 -2268 15118 -2234
rect 15152 -2268 15168 -2234
rect 15024 -2306 15054 -2280
rect 15102 -2284 15168 -2268
rect 15294 -2234 15360 -2218
rect 15294 -2268 15310 -2234
rect 15344 -2268 15360 -2234
rect 15120 -2306 15150 -2284
rect 15216 -2306 15246 -2280
rect 15294 -2284 15360 -2268
rect 15486 -2234 15552 -2218
rect 15486 -2268 15502 -2234
rect 15536 -2268 15552 -2234
rect 15312 -2306 15342 -2284
rect 15408 -2306 15438 -2280
rect 15486 -2284 15552 -2268
rect 15504 -2306 15534 -2284
rect 15024 -2728 15054 -2706
rect 15006 -2744 15072 -2728
rect 15120 -2732 15150 -2706
rect 15216 -2728 15246 -2706
rect 15006 -2778 15022 -2744
rect 15056 -2778 15072 -2744
rect 15006 -2794 15072 -2778
rect 15198 -2744 15264 -2728
rect 15312 -2732 15342 -2706
rect 15408 -2728 15438 -2706
rect 15198 -2778 15214 -2744
rect 15248 -2778 15264 -2744
rect 15198 -2794 15264 -2778
rect 15390 -2744 15456 -2728
rect 15504 -2732 15534 -2706
rect 15390 -2778 15406 -2744
rect 15440 -2778 15456 -2744
rect 15390 -2794 15456 -2778
rect 16046 -1616 16112 -1600
rect 16046 -1650 16062 -1616
rect 16096 -1650 16112 -1616
rect 16046 -1666 16112 -1650
rect 16238 -1616 16304 -1600
rect 16238 -1650 16254 -1616
rect 16288 -1650 16304 -1616
rect 16064 -1688 16094 -1666
rect 16160 -1688 16190 -1662
rect 16238 -1666 16304 -1650
rect 16430 -1616 16496 -1600
rect 16430 -1650 16446 -1616
rect 16480 -1650 16496 -1616
rect 16256 -1688 16286 -1666
rect 16352 -1688 16382 -1662
rect 16430 -1666 16496 -1650
rect 16448 -1688 16478 -1666
rect 16544 -1688 16574 -1662
rect 16064 -2114 16094 -2088
rect 16160 -2110 16190 -2088
rect 16142 -2126 16208 -2110
rect 16256 -2114 16286 -2088
rect 16352 -2110 16382 -2088
rect 16142 -2160 16158 -2126
rect 16192 -2160 16208 -2126
rect 16142 -2176 16208 -2160
rect 16334 -2126 16400 -2110
rect 16448 -2114 16478 -2088
rect 16544 -2110 16574 -2088
rect 16334 -2160 16350 -2126
rect 16384 -2160 16400 -2126
rect 16334 -2176 16400 -2160
rect 16526 -2126 16592 -2110
rect 16526 -2160 16542 -2126
rect 16576 -2160 16592 -2126
rect 16526 -2176 16592 -2160
rect 16142 -2234 16208 -2218
rect 16142 -2268 16158 -2234
rect 16192 -2268 16208 -2234
rect 16064 -2306 16094 -2280
rect 16142 -2284 16208 -2268
rect 16334 -2234 16400 -2218
rect 16334 -2268 16350 -2234
rect 16384 -2268 16400 -2234
rect 16160 -2306 16190 -2284
rect 16256 -2306 16286 -2280
rect 16334 -2284 16400 -2268
rect 16526 -2234 16592 -2218
rect 16526 -2268 16542 -2234
rect 16576 -2268 16592 -2234
rect 16352 -2306 16382 -2284
rect 16448 -2306 16478 -2280
rect 16526 -2284 16592 -2268
rect 16544 -2306 16574 -2284
rect 16064 -2728 16094 -2706
rect 16046 -2744 16112 -2728
rect 16160 -2732 16190 -2706
rect 16256 -2728 16286 -2706
rect 16046 -2778 16062 -2744
rect 16096 -2778 16112 -2744
rect 16046 -2794 16112 -2778
rect 16238 -2744 16304 -2728
rect 16352 -2732 16382 -2706
rect 16448 -2728 16478 -2706
rect 16238 -2778 16254 -2744
rect 16288 -2778 16304 -2744
rect 16238 -2794 16304 -2778
rect 16430 -2744 16496 -2728
rect 16544 -2732 16574 -2706
rect 16430 -2778 16446 -2744
rect 16480 -2778 16496 -2744
rect 16430 -2794 16496 -2778
rect -7357 -3240 -7291 -3224
rect -7357 -3274 -7341 -3240
rect -7307 -3274 -7291 -3240
rect -7357 -3290 -7291 -3274
rect -7239 -3240 -7173 -3224
rect -7239 -3274 -7223 -3240
rect -7189 -3274 -7173 -3240
rect -7239 -3290 -7173 -3274
rect -7121 -3240 -7055 -3224
rect -7121 -3274 -7105 -3240
rect -7071 -3274 -7055 -3240
rect -7121 -3290 -7055 -3274
rect -7003 -3240 -6937 -3224
rect -7003 -3274 -6987 -3240
rect -6953 -3274 -6937 -3240
rect -7003 -3290 -6937 -3274
rect -6885 -3240 -6819 -3224
rect -6885 -3274 -6869 -3240
rect -6835 -3274 -6819 -3240
rect -6885 -3290 -6819 -3274
rect -6767 -3240 -6701 -3224
rect -6767 -3274 -6751 -3240
rect -6717 -3274 -6701 -3240
rect -6767 -3290 -6701 -3274
rect -7354 -3312 -7294 -3290
rect -7236 -3312 -7176 -3290
rect -7118 -3312 -7058 -3290
rect -7000 -3312 -6940 -3290
rect -6882 -3312 -6822 -3290
rect -6764 -3312 -6704 -3290
rect -7354 -3734 -7294 -3712
rect -7236 -3734 -7176 -3712
rect -7118 -3734 -7058 -3712
rect -7000 -3734 -6940 -3712
rect -6882 -3734 -6822 -3712
rect -6764 -3734 -6704 -3712
rect -7357 -3750 -7291 -3734
rect -7357 -3784 -7341 -3750
rect -7307 -3784 -7291 -3750
rect -7357 -3800 -7291 -3784
rect -7239 -3750 -7173 -3734
rect -7239 -3784 -7223 -3750
rect -7189 -3784 -7173 -3750
rect -7239 -3800 -7173 -3784
rect -7121 -3750 -7055 -3734
rect -7121 -3784 -7105 -3750
rect -7071 -3784 -7055 -3750
rect -7121 -3800 -7055 -3784
rect -7003 -3750 -6937 -3734
rect -7003 -3784 -6987 -3750
rect -6953 -3784 -6937 -3750
rect -7003 -3800 -6937 -3784
rect -6885 -3750 -6819 -3734
rect -6885 -3784 -6869 -3750
rect -6835 -3784 -6819 -3750
rect -6885 -3800 -6819 -3784
rect -6767 -3750 -6701 -3734
rect -6767 -3784 -6751 -3750
rect -6717 -3784 -6701 -3750
rect -6767 -3800 -6701 -3784
rect 4277 -3038 4343 -3022
rect 4277 -3072 4293 -3038
rect 4327 -3072 4343 -3038
rect 4277 -3088 4343 -3072
rect 4395 -3038 4461 -3022
rect 4395 -3072 4411 -3038
rect 4445 -3072 4461 -3038
rect 4395 -3088 4461 -3072
rect 4513 -3038 4579 -3022
rect 4513 -3072 4529 -3038
rect 4563 -3072 4579 -3038
rect 4513 -3088 4579 -3072
rect 4631 -3038 4697 -3022
rect 4631 -3072 4647 -3038
rect 4681 -3072 4697 -3038
rect 4631 -3088 4697 -3072
rect 4749 -3038 4815 -3022
rect 4749 -3072 4765 -3038
rect 4799 -3072 4815 -3038
rect 4749 -3088 4815 -3072
rect 4867 -3038 4933 -3022
rect 4867 -3072 4883 -3038
rect 4917 -3072 4933 -3038
rect 4867 -3088 4933 -3072
rect 4280 -3110 4340 -3088
rect 4398 -3110 4458 -3088
rect 4516 -3110 4576 -3088
rect 4634 -3110 4694 -3088
rect 4752 -3110 4812 -3088
rect 4870 -3110 4930 -3088
rect 4280 -3532 4340 -3510
rect 4398 -3532 4458 -3510
rect 4516 -3532 4576 -3510
rect 4634 -3532 4694 -3510
rect 4752 -3532 4812 -3510
rect 4870 -3532 4930 -3510
rect 4277 -3548 4343 -3532
rect 4277 -3582 4293 -3548
rect 4327 -3582 4343 -3548
rect 4277 -3598 4343 -3582
rect 4395 -3548 4461 -3532
rect 4395 -3582 4411 -3548
rect 4445 -3582 4461 -3548
rect 4395 -3598 4461 -3582
rect 4513 -3548 4579 -3532
rect 4513 -3582 4529 -3548
rect 4563 -3582 4579 -3548
rect 4513 -3598 4579 -3582
rect 4631 -3548 4697 -3532
rect 4631 -3582 4647 -3548
rect 4681 -3582 4697 -3548
rect 4631 -3598 4697 -3582
rect 4749 -3548 4815 -3532
rect 4749 -3582 4765 -3548
rect 4799 -3582 4815 -3548
rect 4749 -3598 4815 -3582
rect 4867 -3548 4933 -3532
rect 4867 -3582 4883 -3548
rect 4917 -3582 4933 -3548
rect 4867 -3598 4933 -3582
rect 5317 -3038 5383 -3022
rect 5317 -3072 5333 -3038
rect 5367 -3072 5383 -3038
rect 5317 -3088 5383 -3072
rect 5435 -3038 5501 -3022
rect 5435 -3072 5451 -3038
rect 5485 -3072 5501 -3038
rect 5435 -3088 5501 -3072
rect 5553 -3038 5619 -3022
rect 5553 -3072 5569 -3038
rect 5603 -3072 5619 -3038
rect 5553 -3088 5619 -3072
rect 5671 -3038 5737 -3022
rect 5671 -3072 5687 -3038
rect 5721 -3072 5737 -3038
rect 5671 -3088 5737 -3072
rect 5789 -3038 5855 -3022
rect 5789 -3072 5805 -3038
rect 5839 -3072 5855 -3038
rect 5789 -3088 5855 -3072
rect 5907 -3038 5973 -3022
rect 5907 -3072 5923 -3038
rect 5957 -3072 5973 -3038
rect 5907 -3088 5973 -3072
rect 5320 -3110 5380 -3088
rect 5438 -3110 5498 -3088
rect 5556 -3110 5616 -3088
rect 5674 -3110 5734 -3088
rect 5792 -3110 5852 -3088
rect 5910 -3110 5970 -3088
rect 5320 -3532 5380 -3510
rect 5438 -3532 5498 -3510
rect 5556 -3532 5616 -3510
rect 5674 -3532 5734 -3510
rect 5792 -3532 5852 -3510
rect 5910 -3532 5970 -3510
rect 5317 -3548 5383 -3532
rect 5317 -3582 5333 -3548
rect 5367 -3582 5383 -3548
rect 5317 -3598 5383 -3582
rect 5435 -3548 5501 -3532
rect 5435 -3582 5451 -3548
rect 5485 -3582 5501 -3548
rect 5435 -3598 5501 -3582
rect 5553 -3548 5619 -3532
rect 5553 -3582 5569 -3548
rect 5603 -3582 5619 -3548
rect 5553 -3598 5619 -3582
rect 5671 -3548 5737 -3532
rect 5671 -3582 5687 -3548
rect 5721 -3582 5737 -3548
rect 5671 -3598 5737 -3582
rect 5789 -3548 5855 -3532
rect 5789 -3582 5805 -3548
rect 5839 -3582 5855 -3548
rect 5789 -3598 5855 -3582
rect 5907 -3548 5973 -3532
rect 5907 -3582 5923 -3548
rect 5957 -3582 5973 -3548
rect 5907 -3598 5973 -3582
rect 6357 -3038 6423 -3022
rect 6357 -3072 6373 -3038
rect 6407 -3072 6423 -3038
rect 6357 -3088 6423 -3072
rect 6475 -3038 6541 -3022
rect 6475 -3072 6491 -3038
rect 6525 -3072 6541 -3038
rect 6475 -3088 6541 -3072
rect 6593 -3038 6659 -3022
rect 6593 -3072 6609 -3038
rect 6643 -3072 6659 -3038
rect 6593 -3088 6659 -3072
rect 6711 -3038 6777 -3022
rect 6711 -3072 6727 -3038
rect 6761 -3072 6777 -3038
rect 6711 -3088 6777 -3072
rect 6829 -3038 6895 -3022
rect 6829 -3072 6845 -3038
rect 6879 -3072 6895 -3038
rect 6829 -3088 6895 -3072
rect 6947 -3038 7013 -3022
rect 6947 -3072 6963 -3038
rect 6997 -3072 7013 -3038
rect 6947 -3088 7013 -3072
rect 6360 -3110 6420 -3088
rect 6478 -3110 6538 -3088
rect 6596 -3110 6656 -3088
rect 6714 -3110 6774 -3088
rect 6832 -3110 6892 -3088
rect 6950 -3110 7010 -3088
rect 6360 -3532 6420 -3510
rect 6478 -3532 6538 -3510
rect 6596 -3532 6656 -3510
rect 6714 -3532 6774 -3510
rect 6832 -3532 6892 -3510
rect 6950 -3532 7010 -3510
rect 6357 -3548 6423 -3532
rect 6357 -3582 6373 -3548
rect 6407 -3582 6423 -3548
rect 6357 -3598 6423 -3582
rect 6475 -3548 6541 -3532
rect 6475 -3582 6491 -3548
rect 6525 -3582 6541 -3548
rect 6475 -3598 6541 -3582
rect 6593 -3548 6659 -3532
rect 6593 -3582 6609 -3548
rect 6643 -3582 6659 -3548
rect 6593 -3598 6659 -3582
rect 6711 -3548 6777 -3532
rect 6711 -3582 6727 -3548
rect 6761 -3582 6777 -3548
rect 6711 -3598 6777 -3582
rect 6829 -3548 6895 -3532
rect 6829 -3582 6845 -3548
rect 6879 -3582 6895 -3548
rect 6829 -3598 6895 -3582
rect 6947 -3548 7013 -3532
rect 6947 -3582 6963 -3548
rect 6997 -3582 7013 -3548
rect 6947 -3598 7013 -3582
rect 7397 -3038 7463 -3022
rect 7397 -3072 7413 -3038
rect 7447 -3072 7463 -3038
rect 7397 -3088 7463 -3072
rect 7515 -3038 7581 -3022
rect 7515 -3072 7531 -3038
rect 7565 -3072 7581 -3038
rect 7515 -3088 7581 -3072
rect 7633 -3038 7699 -3022
rect 7633 -3072 7649 -3038
rect 7683 -3072 7699 -3038
rect 7633 -3088 7699 -3072
rect 7751 -3038 7817 -3022
rect 7751 -3072 7767 -3038
rect 7801 -3072 7817 -3038
rect 7751 -3088 7817 -3072
rect 7869 -3038 7935 -3022
rect 7869 -3072 7885 -3038
rect 7919 -3072 7935 -3038
rect 7869 -3088 7935 -3072
rect 7987 -3038 8053 -3022
rect 7987 -3072 8003 -3038
rect 8037 -3072 8053 -3038
rect 7987 -3088 8053 -3072
rect 7400 -3110 7460 -3088
rect 7518 -3110 7578 -3088
rect 7636 -3110 7696 -3088
rect 7754 -3110 7814 -3088
rect 7872 -3110 7932 -3088
rect 7990 -3110 8050 -3088
rect 7400 -3532 7460 -3510
rect 7518 -3532 7578 -3510
rect 7636 -3532 7696 -3510
rect 7754 -3532 7814 -3510
rect 7872 -3532 7932 -3510
rect 7990 -3532 8050 -3510
rect 7397 -3548 7463 -3532
rect 7397 -3582 7413 -3548
rect 7447 -3582 7463 -3548
rect 7397 -3598 7463 -3582
rect 7515 -3548 7581 -3532
rect 7515 -3582 7531 -3548
rect 7565 -3582 7581 -3548
rect 7515 -3598 7581 -3582
rect 7633 -3548 7699 -3532
rect 7633 -3582 7649 -3548
rect 7683 -3582 7699 -3548
rect 7633 -3598 7699 -3582
rect 7751 -3548 7817 -3532
rect 7751 -3582 7767 -3548
rect 7801 -3582 7817 -3548
rect 7751 -3598 7817 -3582
rect 7869 -3548 7935 -3532
rect 7869 -3582 7885 -3548
rect 7919 -3582 7935 -3548
rect 7869 -3598 7935 -3582
rect 7987 -3548 8053 -3532
rect 7987 -3582 8003 -3548
rect 8037 -3582 8053 -3548
rect 7987 -3598 8053 -3582
rect 8437 -3038 8503 -3022
rect 8437 -3072 8453 -3038
rect 8487 -3072 8503 -3038
rect 8437 -3088 8503 -3072
rect 8555 -3038 8621 -3022
rect 8555 -3072 8571 -3038
rect 8605 -3072 8621 -3038
rect 8555 -3088 8621 -3072
rect 8673 -3038 8739 -3022
rect 8673 -3072 8689 -3038
rect 8723 -3072 8739 -3038
rect 8673 -3088 8739 -3072
rect 8791 -3038 8857 -3022
rect 8791 -3072 8807 -3038
rect 8841 -3072 8857 -3038
rect 8791 -3088 8857 -3072
rect 8909 -3038 8975 -3022
rect 8909 -3072 8925 -3038
rect 8959 -3072 8975 -3038
rect 8909 -3088 8975 -3072
rect 9027 -3038 9093 -3022
rect 9027 -3072 9043 -3038
rect 9077 -3072 9093 -3038
rect 9027 -3088 9093 -3072
rect 8440 -3110 8500 -3088
rect 8558 -3110 8618 -3088
rect 8676 -3110 8736 -3088
rect 8794 -3110 8854 -3088
rect 8912 -3110 8972 -3088
rect 9030 -3110 9090 -3088
rect 8440 -3532 8500 -3510
rect 8558 -3532 8618 -3510
rect 8676 -3532 8736 -3510
rect 8794 -3532 8854 -3510
rect 8912 -3532 8972 -3510
rect 9030 -3532 9090 -3510
rect 8437 -3548 8503 -3532
rect 8437 -3582 8453 -3548
rect 8487 -3582 8503 -3548
rect 8437 -3598 8503 -3582
rect 8555 -3548 8621 -3532
rect 8555 -3582 8571 -3548
rect 8605 -3582 8621 -3548
rect 8555 -3598 8621 -3582
rect 8673 -3548 8739 -3532
rect 8673 -3582 8689 -3548
rect 8723 -3582 8739 -3548
rect 8673 -3598 8739 -3582
rect 8791 -3548 8857 -3532
rect 8791 -3582 8807 -3548
rect 8841 -3582 8857 -3548
rect 8791 -3598 8857 -3582
rect 8909 -3548 8975 -3532
rect 8909 -3582 8925 -3548
rect 8959 -3582 8975 -3548
rect 8909 -3598 8975 -3582
rect 9027 -3548 9093 -3532
rect 9027 -3582 9043 -3548
rect 9077 -3582 9093 -3548
rect 9027 -3598 9093 -3582
rect 11897 -3038 11963 -3022
rect 11897 -3072 11913 -3038
rect 11947 -3072 11963 -3038
rect 11897 -3088 11963 -3072
rect 12015 -3038 12081 -3022
rect 12015 -3072 12031 -3038
rect 12065 -3072 12081 -3038
rect 12015 -3088 12081 -3072
rect 12133 -3038 12199 -3022
rect 12133 -3072 12149 -3038
rect 12183 -3072 12199 -3038
rect 12133 -3088 12199 -3072
rect 12251 -3038 12317 -3022
rect 12251 -3072 12267 -3038
rect 12301 -3072 12317 -3038
rect 12251 -3088 12317 -3072
rect 12369 -3038 12435 -3022
rect 12369 -3072 12385 -3038
rect 12419 -3072 12435 -3038
rect 12369 -3088 12435 -3072
rect 12487 -3038 12553 -3022
rect 12487 -3072 12503 -3038
rect 12537 -3072 12553 -3038
rect 12487 -3088 12553 -3072
rect 11900 -3110 11960 -3088
rect 12018 -3110 12078 -3088
rect 12136 -3110 12196 -3088
rect 12254 -3110 12314 -3088
rect 12372 -3110 12432 -3088
rect 12490 -3110 12550 -3088
rect 11900 -3532 11960 -3510
rect 12018 -3532 12078 -3510
rect 12136 -3532 12196 -3510
rect 12254 -3532 12314 -3510
rect 12372 -3532 12432 -3510
rect 12490 -3532 12550 -3510
rect 11897 -3548 11963 -3532
rect 11897 -3582 11913 -3548
rect 11947 -3582 11963 -3548
rect 11897 -3598 11963 -3582
rect 12015 -3548 12081 -3532
rect 12015 -3582 12031 -3548
rect 12065 -3582 12081 -3548
rect 12015 -3598 12081 -3582
rect 12133 -3548 12199 -3532
rect 12133 -3582 12149 -3548
rect 12183 -3582 12199 -3548
rect 12133 -3598 12199 -3582
rect 12251 -3548 12317 -3532
rect 12251 -3582 12267 -3548
rect 12301 -3582 12317 -3548
rect 12251 -3598 12317 -3582
rect 12369 -3548 12435 -3532
rect 12369 -3582 12385 -3548
rect 12419 -3582 12435 -3548
rect 12369 -3598 12435 -3582
rect 12487 -3548 12553 -3532
rect 12487 -3582 12503 -3548
rect 12537 -3582 12553 -3548
rect 12487 -3598 12553 -3582
rect 12937 -3038 13003 -3022
rect 12937 -3072 12953 -3038
rect 12987 -3072 13003 -3038
rect 12937 -3088 13003 -3072
rect 13055 -3038 13121 -3022
rect 13055 -3072 13071 -3038
rect 13105 -3072 13121 -3038
rect 13055 -3088 13121 -3072
rect 13173 -3038 13239 -3022
rect 13173 -3072 13189 -3038
rect 13223 -3072 13239 -3038
rect 13173 -3088 13239 -3072
rect 13291 -3038 13357 -3022
rect 13291 -3072 13307 -3038
rect 13341 -3072 13357 -3038
rect 13291 -3088 13357 -3072
rect 13409 -3038 13475 -3022
rect 13409 -3072 13425 -3038
rect 13459 -3072 13475 -3038
rect 13409 -3088 13475 -3072
rect 13527 -3038 13593 -3022
rect 13527 -3072 13543 -3038
rect 13577 -3072 13593 -3038
rect 13527 -3088 13593 -3072
rect 12940 -3110 13000 -3088
rect 13058 -3110 13118 -3088
rect 13176 -3110 13236 -3088
rect 13294 -3110 13354 -3088
rect 13412 -3110 13472 -3088
rect 13530 -3110 13590 -3088
rect 12940 -3532 13000 -3510
rect 13058 -3532 13118 -3510
rect 13176 -3532 13236 -3510
rect 13294 -3532 13354 -3510
rect 13412 -3532 13472 -3510
rect 13530 -3532 13590 -3510
rect 12937 -3548 13003 -3532
rect 12937 -3582 12953 -3548
rect 12987 -3582 13003 -3548
rect 12937 -3598 13003 -3582
rect 13055 -3548 13121 -3532
rect 13055 -3582 13071 -3548
rect 13105 -3582 13121 -3548
rect 13055 -3598 13121 -3582
rect 13173 -3548 13239 -3532
rect 13173 -3582 13189 -3548
rect 13223 -3582 13239 -3548
rect 13173 -3598 13239 -3582
rect 13291 -3548 13357 -3532
rect 13291 -3582 13307 -3548
rect 13341 -3582 13357 -3548
rect 13291 -3598 13357 -3582
rect 13409 -3548 13475 -3532
rect 13409 -3582 13425 -3548
rect 13459 -3582 13475 -3548
rect 13409 -3598 13475 -3582
rect 13527 -3548 13593 -3532
rect 13527 -3582 13543 -3548
rect 13577 -3582 13593 -3548
rect 13527 -3598 13593 -3582
rect 13977 -3038 14043 -3022
rect 13977 -3072 13993 -3038
rect 14027 -3072 14043 -3038
rect 13977 -3088 14043 -3072
rect 14095 -3038 14161 -3022
rect 14095 -3072 14111 -3038
rect 14145 -3072 14161 -3038
rect 14095 -3088 14161 -3072
rect 14213 -3038 14279 -3022
rect 14213 -3072 14229 -3038
rect 14263 -3072 14279 -3038
rect 14213 -3088 14279 -3072
rect 14331 -3038 14397 -3022
rect 14331 -3072 14347 -3038
rect 14381 -3072 14397 -3038
rect 14331 -3088 14397 -3072
rect 14449 -3038 14515 -3022
rect 14449 -3072 14465 -3038
rect 14499 -3072 14515 -3038
rect 14449 -3088 14515 -3072
rect 14567 -3038 14633 -3022
rect 14567 -3072 14583 -3038
rect 14617 -3072 14633 -3038
rect 14567 -3088 14633 -3072
rect 13980 -3110 14040 -3088
rect 14098 -3110 14158 -3088
rect 14216 -3110 14276 -3088
rect 14334 -3110 14394 -3088
rect 14452 -3110 14512 -3088
rect 14570 -3110 14630 -3088
rect 13980 -3532 14040 -3510
rect 14098 -3532 14158 -3510
rect 14216 -3532 14276 -3510
rect 14334 -3532 14394 -3510
rect 14452 -3532 14512 -3510
rect 14570 -3532 14630 -3510
rect 13977 -3548 14043 -3532
rect 13977 -3582 13993 -3548
rect 14027 -3582 14043 -3548
rect 13977 -3598 14043 -3582
rect 14095 -3548 14161 -3532
rect 14095 -3582 14111 -3548
rect 14145 -3582 14161 -3548
rect 14095 -3598 14161 -3582
rect 14213 -3548 14279 -3532
rect 14213 -3582 14229 -3548
rect 14263 -3582 14279 -3548
rect 14213 -3598 14279 -3582
rect 14331 -3548 14397 -3532
rect 14331 -3582 14347 -3548
rect 14381 -3582 14397 -3548
rect 14331 -3598 14397 -3582
rect 14449 -3548 14515 -3532
rect 14449 -3582 14465 -3548
rect 14499 -3582 14515 -3548
rect 14449 -3598 14515 -3582
rect 14567 -3548 14633 -3532
rect 14567 -3582 14583 -3548
rect 14617 -3582 14633 -3548
rect 14567 -3598 14633 -3582
rect 15017 -3038 15083 -3022
rect 15017 -3072 15033 -3038
rect 15067 -3072 15083 -3038
rect 15017 -3088 15083 -3072
rect 15135 -3038 15201 -3022
rect 15135 -3072 15151 -3038
rect 15185 -3072 15201 -3038
rect 15135 -3088 15201 -3072
rect 15253 -3038 15319 -3022
rect 15253 -3072 15269 -3038
rect 15303 -3072 15319 -3038
rect 15253 -3088 15319 -3072
rect 15371 -3038 15437 -3022
rect 15371 -3072 15387 -3038
rect 15421 -3072 15437 -3038
rect 15371 -3088 15437 -3072
rect 15489 -3038 15555 -3022
rect 15489 -3072 15505 -3038
rect 15539 -3072 15555 -3038
rect 15489 -3088 15555 -3072
rect 15607 -3038 15673 -3022
rect 15607 -3072 15623 -3038
rect 15657 -3072 15673 -3038
rect 15607 -3088 15673 -3072
rect 15020 -3110 15080 -3088
rect 15138 -3110 15198 -3088
rect 15256 -3110 15316 -3088
rect 15374 -3110 15434 -3088
rect 15492 -3110 15552 -3088
rect 15610 -3110 15670 -3088
rect 15020 -3532 15080 -3510
rect 15138 -3532 15198 -3510
rect 15256 -3532 15316 -3510
rect 15374 -3532 15434 -3510
rect 15492 -3532 15552 -3510
rect 15610 -3532 15670 -3510
rect 15017 -3548 15083 -3532
rect 15017 -3582 15033 -3548
rect 15067 -3582 15083 -3548
rect 15017 -3598 15083 -3582
rect 15135 -3548 15201 -3532
rect 15135 -3582 15151 -3548
rect 15185 -3582 15201 -3548
rect 15135 -3598 15201 -3582
rect 15253 -3548 15319 -3532
rect 15253 -3582 15269 -3548
rect 15303 -3582 15319 -3548
rect 15253 -3598 15319 -3582
rect 15371 -3548 15437 -3532
rect 15371 -3582 15387 -3548
rect 15421 -3582 15437 -3548
rect 15371 -3598 15437 -3582
rect 15489 -3548 15555 -3532
rect 15489 -3582 15505 -3548
rect 15539 -3582 15555 -3548
rect 15489 -3598 15555 -3582
rect 15607 -3548 15673 -3532
rect 15607 -3582 15623 -3548
rect 15657 -3582 15673 -3548
rect 15607 -3598 15673 -3582
rect 16057 -3038 16123 -3022
rect 16057 -3072 16073 -3038
rect 16107 -3072 16123 -3038
rect 16057 -3088 16123 -3072
rect 16175 -3038 16241 -3022
rect 16175 -3072 16191 -3038
rect 16225 -3072 16241 -3038
rect 16175 -3088 16241 -3072
rect 16293 -3038 16359 -3022
rect 16293 -3072 16309 -3038
rect 16343 -3072 16359 -3038
rect 16293 -3088 16359 -3072
rect 16411 -3038 16477 -3022
rect 16411 -3072 16427 -3038
rect 16461 -3072 16477 -3038
rect 16411 -3088 16477 -3072
rect 16529 -3038 16595 -3022
rect 16529 -3072 16545 -3038
rect 16579 -3072 16595 -3038
rect 16529 -3088 16595 -3072
rect 16647 -3038 16713 -3022
rect 16647 -3072 16663 -3038
rect 16697 -3072 16713 -3038
rect 16647 -3088 16713 -3072
rect 16060 -3110 16120 -3088
rect 16178 -3110 16238 -3088
rect 16296 -3110 16356 -3088
rect 16414 -3110 16474 -3088
rect 16532 -3110 16592 -3088
rect 16650 -3110 16710 -3088
rect 16060 -3532 16120 -3510
rect 16178 -3532 16238 -3510
rect 16296 -3532 16356 -3510
rect 16414 -3532 16474 -3510
rect 16532 -3532 16592 -3510
rect 16650 -3532 16710 -3510
rect 16057 -3548 16123 -3532
rect 16057 -3582 16073 -3548
rect 16107 -3582 16123 -3548
rect 16057 -3598 16123 -3582
rect 16175 -3548 16241 -3532
rect 16175 -3582 16191 -3548
rect 16225 -3582 16241 -3548
rect 16175 -3598 16241 -3582
rect 16293 -3548 16359 -3532
rect 16293 -3582 16309 -3548
rect 16343 -3582 16359 -3548
rect 16293 -3598 16359 -3582
rect 16411 -3548 16477 -3532
rect 16411 -3582 16427 -3548
rect 16461 -3582 16477 -3548
rect 16411 -3598 16477 -3582
rect 16529 -3548 16595 -3532
rect 16529 -3582 16545 -3548
rect 16579 -3582 16595 -3548
rect 16529 -3598 16595 -3582
rect 16647 -3548 16713 -3532
rect 16647 -3582 16663 -3548
rect 16697 -3582 16713 -3548
rect 16647 -3598 16713 -3582
<< polycont >>
rect -886 3648 -852 3682
rect -694 3648 -660 3682
rect -502 3648 -468 3682
rect -310 3648 -276 3682
rect -118 3648 -84 3682
rect -982 3138 -948 3172
rect -790 3138 -756 3172
rect -598 3138 -564 3172
rect -406 3138 -372 3172
rect -214 3138 -180 3172
rect 1914 3648 1948 3682
rect 2106 3648 2140 3682
rect 2298 3648 2332 3682
rect 2490 3648 2524 3682
rect 2682 3648 2716 3682
rect 1818 3138 1852 3172
rect 2010 3138 2044 3172
rect 2202 3138 2236 3172
rect 2394 3138 2428 3172
rect 2586 3138 2620 3172
rect 4482 5502 4516 5536
rect 4674 5502 4708 5536
rect 4866 5502 4900 5536
rect 5058 5502 5092 5536
rect 5250 5502 5284 5536
rect 5442 5502 5476 5536
rect 5634 5502 5668 5536
rect 5826 5502 5860 5536
rect 6018 5502 6052 5536
rect 6210 5502 6244 5536
rect 6402 5502 6436 5536
rect 6594 5502 6628 5536
rect 6786 5502 6820 5536
rect 6978 5502 7012 5536
rect 7170 5502 7204 5536
rect 4578 4992 4612 5026
rect 4770 4992 4804 5026
rect 4962 4992 4996 5026
rect 5154 4992 5188 5026
rect 5346 4992 5380 5026
rect 5538 4992 5572 5026
rect 5730 4992 5764 5026
rect 5922 4992 5956 5026
rect 6114 4992 6148 5026
rect 6306 4992 6340 5026
rect 6498 4992 6532 5026
rect 6690 4992 6724 5026
rect 6882 4992 6916 5026
rect 7074 4992 7108 5026
rect 7266 4992 7300 5026
rect 4578 4884 4612 4918
rect 4770 4884 4804 4918
rect 4962 4884 4996 4918
rect 5154 4884 5188 4918
rect 5346 4884 5380 4918
rect 5538 4884 5572 4918
rect 5730 4884 5764 4918
rect 5922 4884 5956 4918
rect 6114 4884 6148 4918
rect 6306 4884 6340 4918
rect 6498 4884 6532 4918
rect 6690 4884 6724 4918
rect 6882 4884 6916 4918
rect 7074 4884 7108 4918
rect 7266 4884 7300 4918
rect 4482 4374 4516 4408
rect 4674 4374 4708 4408
rect 4866 4374 4900 4408
rect 5058 4374 5092 4408
rect 5250 4374 5284 4408
rect 5442 4374 5476 4408
rect 5634 4374 5668 4408
rect 5826 4374 5860 4408
rect 6018 4374 6052 4408
rect 6210 4374 6244 4408
rect 6402 4374 6436 4408
rect 6594 4374 6628 4408
rect 6786 4374 6820 4408
rect 6978 4374 7012 4408
rect 7170 4374 7204 4408
rect 4482 4266 4516 4300
rect 4674 4266 4708 4300
rect 4866 4266 4900 4300
rect 5058 4266 5092 4300
rect 5250 4266 5284 4300
rect 5442 4266 5476 4300
rect 5634 4266 5668 4300
rect 5826 4266 5860 4300
rect 6018 4266 6052 4300
rect 6210 4266 6244 4300
rect 6402 4266 6436 4300
rect 6594 4266 6628 4300
rect 6786 4266 6820 4300
rect 6978 4266 7012 4300
rect 7170 4266 7204 4300
rect 4578 3756 4612 3790
rect 4770 3756 4804 3790
rect 4962 3756 4996 3790
rect 5154 3756 5188 3790
rect 5346 3756 5380 3790
rect 5538 3756 5572 3790
rect 5730 3756 5764 3790
rect 5922 3756 5956 3790
rect 6114 3756 6148 3790
rect 6306 3756 6340 3790
rect 6498 3756 6532 3790
rect 6690 3756 6724 3790
rect 6882 3756 6916 3790
rect 7074 3756 7108 3790
rect 7266 3756 7300 3790
rect 4578 3648 4612 3682
rect 4770 3648 4804 3682
rect 4962 3648 4996 3682
rect 5154 3648 5188 3682
rect 5346 3648 5380 3682
rect 5538 3648 5572 3682
rect 5730 3648 5764 3682
rect 5922 3648 5956 3682
rect 6114 3648 6148 3682
rect 6306 3648 6340 3682
rect 6498 3648 6532 3682
rect 6690 3648 6724 3682
rect 6882 3648 6916 3682
rect 7074 3648 7108 3682
rect 7266 3648 7300 3682
rect 4482 3138 4516 3172
rect 4674 3138 4708 3172
rect 4866 3138 4900 3172
rect 5058 3138 5092 3172
rect 5250 3138 5284 3172
rect 5442 3138 5476 3172
rect 5634 3138 5668 3172
rect 5826 3138 5860 3172
rect 6018 3138 6052 3172
rect 6210 3138 6244 3172
rect 6402 3138 6436 3172
rect 6594 3138 6628 3172
rect 6786 3138 6820 3172
rect 6978 3138 7012 3172
rect 7170 3138 7204 3172
rect 8122 5502 8156 5536
rect 8314 5502 8348 5536
rect 8506 5502 8540 5536
rect 8698 5502 8732 5536
rect 8890 5502 8924 5536
rect 9082 5502 9116 5536
rect 9274 5502 9308 5536
rect 9466 5502 9500 5536
rect 9658 5502 9692 5536
rect 9850 5502 9884 5536
rect 10042 5502 10076 5536
rect 10234 5502 10268 5536
rect 10426 5502 10460 5536
rect 10618 5502 10652 5536
rect 10810 5502 10844 5536
rect 8218 4992 8252 5026
rect 8410 4992 8444 5026
rect 8602 4992 8636 5026
rect 8794 4992 8828 5026
rect 8986 4992 9020 5026
rect 9178 4992 9212 5026
rect 9370 4992 9404 5026
rect 9562 4992 9596 5026
rect 9754 4992 9788 5026
rect 9946 4992 9980 5026
rect 10138 4992 10172 5026
rect 10330 4992 10364 5026
rect 10522 4992 10556 5026
rect 10714 4992 10748 5026
rect 10906 4992 10940 5026
rect 8218 4884 8252 4918
rect 8410 4884 8444 4918
rect 8602 4884 8636 4918
rect 8794 4884 8828 4918
rect 8986 4884 9020 4918
rect 9178 4884 9212 4918
rect 9370 4884 9404 4918
rect 9562 4884 9596 4918
rect 9754 4884 9788 4918
rect 9946 4884 9980 4918
rect 10138 4884 10172 4918
rect 10330 4884 10364 4918
rect 10522 4884 10556 4918
rect 10714 4884 10748 4918
rect 10906 4884 10940 4918
rect 8122 4374 8156 4408
rect 8314 4374 8348 4408
rect 8506 4374 8540 4408
rect 8698 4374 8732 4408
rect 8890 4374 8924 4408
rect 9082 4374 9116 4408
rect 9274 4374 9308 4408
rect 9466 4374 9500 4408
rect 9658 4374 9692 4408
rect 9850 4374 9884 4408
rect 10042 4374 10076 4408
rect 10234 4374 10268 4408
rect 10426 4374 10460 4408
rect 10618 4374 10652 4408
rect 10810 4374 10844 4408
rect 8122 4266 8156 4300
rect 8314 4266 8348 4300
rect 8506 4266 8540 4300
rect 8698 4266 8732 4300
rect 8890 4266 8924 4300
rect 9082 4266 9116 4300
rect 9274 4266 9308 4300
rect 9466 4266 9500 4300
rect 9658 4266 9692 4300
rect 9850 4266 9884 4300
rect 10042 4266 10076 4300
rect 10234 4266 10268 4300
rect 10426 4266 10460 4300
rect 10618 4266 10652 4300
rect 10810 4266 10844 4300
rect 8218 3756 8252 3790
rect 8410 3756 8444 3790
rect 8602 3756 8636 3790
rect 8794 3756 8828 3790
rect 8986 3756 9020 3790
rect 9178 3756 9212 3790
rect 9370 3756 9404 3790
rect 9562 3756 9596 3790
rect 9754 3756 9788 3790
rect 9946 3756 9980 3790
rect 10138 3756 10172 3790
rect 10330 3756 10364 3790
rect 10522 3756 10556 3790
rect 10714 3756 10748 3790
rect 10906 3756 10940 3790
rect 8218 3648 8252 3682
rect 8410 3648 8444 3682
rect 8602 3648 8636 3682
rect 8794 3648 8828 3682
rect 8986 3648 9020 3682
rect 9178 3648 9212 3682
rect 9370 3648 9404 3682
rect 9562 3648 9596 3682
rect 9754 3648 9788 3682
rect 9946 3648 9980 3682
rect 10138 3648 10172 3682
rect 10330 3648 10364 3682
rect 10522 3648 10556 3682
rect 10714 3648 10748 3682
rect 10906 3648 10940 3682
rect 8122 3138 8156 3172
rect 8314 3138 8348 3172
rect 8506 3138 8540 3172
rect 8698 3138 8732 3172
rect 8890 3138 8924 3172
rect 9082 3138 9116 3172
rect 9274 3138 9308 3172
rect 9466 3138 9500 3172
rect 9658 3138 9692 3172
rect 9850 3138 9884 3172
rect 10042 3138 10076 3172
rect 10234 3138 10268 3172
rect 10426 3138 10460 3172
rect 10618 3138 10652 3172
rect 10810 3138 10844 3172
rect 12102 5502 12136 5536
rect 12294 5502 12328 5536
rect 12486 5502 12520 5536
rect 12678 5502 12712 5536
rect 12870 5502 12904 5536
rect 13062 5502 13096 5536
rect 13254 5502 13288 5536
rect 13446 5502 13480 5536
rect 13638 5502 13672 5536
rect 13830 5502 13864 5536
rect 14022 5502 14056 5536
rect 14214 5502 14248 5536
rect 14406 5502 14440 5536
rect 14598 5502 14632 5536
rect 14790 5502 14824 5536
rect 12198 4992 12232 5026
rect 12390 4992 12424 5026
rect 12582 4992 12616 5026
rect 12774 4992 12808 5026
rect 12966 4992 13000 5026
rect 13158 4992 13192 5026
rect 13350 4992 13384 5026
rect 13542 4992 13576 5026
rect 13734 4992 13768 5026
rect 13926 4992 13960 5026
rect 14118 4992 14152 5026
rect 14310 4992 14344 5026
rect 14502 4992 14536 5026
rect 14694 4992 14728 5026
rect 14886 4992 14920 5026
rect 12198 4884 12232 4918
rect 12390 4884 12424 4918
rect 12582 4884 12616 4918
rect 12774 4884 12808 4918
rect 12966 4884 13000 4918
rect 13158 4884 13192 4918
rect 13350 4884 13384 4918
rect 13542 4884 13576 4918
rect 13734 4884 13768 4918
rect 13926 4884 13960 4918
rect 14118 4884 14152 4918
rect 14310 4884 14344 4918
rect 14502 4884 14536 4918
rect 14694 4884 14728 4918
rect 14886 4884 14920 4918
rect 12102 4374 12136 4408
rect 12294 4374 12328 4408
rect 12486 4374 12520 4408
rect 12678 4374 12712 4408
rect 12870 4374 12904 4408
rect 13062 4374 13096 4408
rect 13254 4374 13288 4408
rect 13446 4374 13480 4408
rect 13638 4374 13672 4408
rect 13830 4374 13864 4408
rect 14022 4374 14056 4408
rect 14214 4374 14248 4408
rect 14406 4374 14440 4408
rect 14598 4374 14632 4408
rect 14790 4374 14824 4408
rect 12102 4266 12136 4300
rect 12294 4266 12328 4300
rect 12486 4266 12520 4300
rect 12678 4266 12712 4300
rect 12870 4266 12904 4300
rect 13062 4266 13096 4300
rect 13254 4266 13288 4300
rect 13446 4266 13480 4300
rect 13638 4266 13672 4300
rect 13830 4266 13864 4300
rect 14022 4266 14056 4300
rect 14214 4266 14248 4300
rect 14406 4266 14440 4300
rect 14598 4266 14632 4300
rect 14790 4266 14824 4300
rect 12198 3756 12232 3790
rect 12390 3756 12424 3790
rect 12582 3756 12616 3790
rect 12774 3756 12808 3790
rect 12966 3756 13000 3790
rect 13158 3756 13192 3790
rect 13350 3756 13384 3790
rect 13542 3756 13576 3790
rect 13734 3756 13768 3790
rect 13926 3756 13960 3790
rect 14118 3756 14152 3790
rect 14310 3756 14344 3790
rect 14502 3756 14536 3790
rect 14694 3756 14728 3790
rect 14886 3756 14920 3790
rect 12198 3648 12232 3682
rect 12390 3648 12424 3682
rect 12582 3648 12616 3682
rect 12774 3648 12808 3682
rect 12966 3648 13000 3682
rect 13158 3648 13192 3682
rect 13350 3648 13384 3682
rect 13542 3648 13576 3682
rect 13734 3648 13768 3682
rect 13926 3648 13960 3682
rect 14118 3648 14152 3682
rect 14310 3648 14344 3682
rect 14502 3648 14536 3682
rect 14694 3648 14728 3682
rect 14886 3648 14920 3682
rect 12102 3138 12136 3172
rect 12294 3138 12328 3172
rect 12486 3138 12520 3172
rect 12678 3138 12712 3172
rect 12870 3138 12904 3172
rect 13062 3138 13096 3172
rect 13254 3138 13288 3172
rect 13446 3138 13480 3172
rect 13638 3138 13672 3172
rect 13830 3138 13864 3172
rect 14022 3138 14056 3172
rect 14214 3138 14248 3172
rect 14406 3138 14440 3172
rect 14598 3138 14632 3172
rect 14790 3138 14824 3172
rect 15742 5502 15776 5536
rect 15934 5502 15968 5536
rect 16126 5502 16160 5536
rect 16318 5502 16352 5536
rect 16510 5502 16544 5536
rect 16702 5502 16736 5536
rect 16894 5502 16928 5536
rect 17086 5502 17120 5536
rect 17278 5502 17312 5536
rect 17470 5502 17504 5536
rect 17662 5502 17696 5536
rect 17854 5502 17888 5536
rect 18046 5502 18080 5536
rect 18238 5502 18272 5536
rect 18430 5502 18464 5536
rect 15838 4992 15872 5026
rect 16030 4992 16064 5026
rect 16222 4992 16256 5026
rect 16414 4992 16448 5026
rect 16606 4992 16640 5026
rect 16798 4992 16832 5026
rect 16990 4992 17024 5026
rect 17182 4992 17216 5026
rect 17374 4992 17408 5026
rect 17566 4992 17600 5026
rect 17758 4992 17792 5026
rect 17950 4992 17984 5026
rect 18142 4992 18176 5026
rect 18334 4992 18368 5026
rect 18526 4992 18560 5026
rect 15838 4884 15872 4918
rect 16030 4884 16064 4918
rect 16222 4884 16256 4918
rect 16414 4884 16448 4918
rect 16606 4884 16640 4918
rect 16798 4884 16832 4918
rect 16990 4884 17024 4918
rect 17182 4884 17216 4918
rect 17374 4884 17408 4918
rect 17566 4884 17600 4918
rect 17758 4884 17792 4918
rect 17950 4884 17984 4918
rect 18142 4884 18176 4918
rect 18334 4884 18368 4918
rect 18526 4884 18560 4918
rect 15742 4374 15776 4408
rect 15934 4374 15968 4408
rect 16126 4374 16160 4408
rect 16318 4374 16352 4408
rect 16510 4374 16544 4408
rect 16702 4374 16736 4408
rect 16894 4374 16928 4408
rect 17086 4374 17120 4408
rect 17278 4374 17312 4408
rect 17470 4374 17504 4408
rect 17662 4374 17696 4408
rect 17854 4374 17888 4408
rect 18046 4374 18080 4408
rect 18238 4374 18272 4408
rect 18430 4374 18464 4408
rect 15742 4266 15776 4300
rect 15934 4266 15968 4300
rect 16126 4266 16160 4300
rect 16318 4266 16352 4300
rect 16510 4266 16544 4300
rect 16702 4266 16736 4300
rect 16894 4266 16928 4300
rect 17086 4266 17120 4300
rect 17278 4266 17312 4300
rect 17470 4266 17504 4300
rect 17662 4266 17696 4300
rect 17854 4266 17888 4300
rect 18046 4266 18080 4300
rect 18238 4266 18272 4300
rect 18430 4266 18464 4300
rect 15838 3756 15872 3790
rect 16030 3756 16064 3790
rect 16222 3756 16256 3790
rect 16414 3756 16448 3790
rect 16606 3756 16640 3790
rect 16798 3756 16832 3790
rect 16990 3756 17024 3790
rect 17182 3756 17216 3790
rect 17374 3756 17408 3790
rect 17566 3756 17600 3790
rect 17758 3756 17792 3790
rect 17950 3756 17984 3790
rect 18142 3756 18176 3790
rect 18334 3756 18368 3790
rect 18526 3756 18560 3790
rect 15838 3648 15872 3682
rect 16030 3648 16064 3682
rect 16222 3648 16256 3682
rect 16414 3648 16448 3682
rect 16606 3648 16640 3682
rect 16798 3648 16832 3682
rect 16990 3648 17024 3682
rect 17182 3648 17216 3682
rect 17374 3648 17408 3682
rect 17566 3648 17600 3682
rect 17758 3648 17792 3682
rect 17950 3648 17984 3682
rect 18142 3648 18176 3682
rect 18334 3648 18368 3682
rect 18526 3648 18560 3682
rect 15742 3138 15776 3172
rect 15934 3138 15968 3172
rect 16126 3138 16160 3172
rect 16318 3138 16352 3172
rect 16510 3138 16544 3172
rect 16702 3138 16736 3172
rect 16894 3138 16928 3172
rect 17086 3138 17120 3172
rect 17278 3138 17312 3172
rect 17470 3138 17504 3172
rect 17662 3138 17696 3172
rect 17854 3138 17888 3172
rect 18046 3138 18080 3172
rect 18238 3138 18272 3172
rect 18430 3138 18464 3172
rect -1522 2670 -1488 2704
rect -1330 2670 -1296 2704
rect -1138 2670 -1104 2704
rect -1426 2160 -1392 2194
rect -1234 2160 -1200 2194
rect -1042 2160 -1008 2194
rect -1426 2052 -1392 2086
rect -1234 2052 -1200 2086
rect -1042 2052 -1008 2086
rect -1522 1542 -1488 1576
rect -1330 1542 -1296 1576
rect -1138 1542 -1104 1576
rect -482 2670 -448 2704
rect -290 2670 -256 2704
rect -98 2670 -64 2704
rect -386 2160 -352 2194
rect -194 2160 -160 2194
rect -2 2160 32 2194
rect -386 2052 -352 2086
rect -194 2052 -160 2086
rect -2 2052 32 2086
rect -482 1542 -448 1576
rect -290 1542 -256 1576
rect -98 1542 -64 1576
rect 558 2670 592 2704
rect 750 2670 784 2704
rect 942 2670 976 2704
rect 654 2160 688 2194
rect 846 2160 880 2194
rect 1038 2160 1072 2194
rect 654 2052 688 2086
rect 846 2052 880 2086
rect 1038 2052 1072 2086
rect 558 1542 592 1576
rect 750 1542 784 1576
rect 942 1542 976 1576
rect 1598 2670 1632 2704
rect 1790 2670 1824 2704
rect 1982 2670 2016 2704
rect 1694 2160 1728 2194
rect 1886 2160 1920 2194
rect 2078 2160 2112 2194
rect 1694 2052 1728 2086
rect 1886 2052 1920 2086
rect 2078 2052 2112 2086
rect 1598 1542 1632 1576
rect 1790 1542 1824 1576
rect 1982 1542 2016 1576
rect 2638 2670 2672 2704
rect 2830 2670 2864 2704
rect 3022 2670 3056 2704
rect 2734 2160 2768 2194
rect 2926 2160 2960 2194
rect 3118 2160 3152 2194
rect 2734 2052 2768 2086
rect 2926 2052 2960 2086
rect 3118 2052 3152 2086
rect 2638 1542 2672 1576
rect 2830 1542 2864 1576
rect 3022 1542 3056 1576
rect 4282 2830 4316 2864
rect 4474 2830 4508 2864
rect 4666 2830 4700 2864
rect 4378 2320 4412 2354
rect 4570 2320 4604 2354
rect 4762 2320 4796 2354
rect 4378 2212 4412 2246
rect 4570 2212 4604 2246
rect 4762 2212 4796 2246
rect 4282 1702 4316 1736
rect 4474 1702 4508 1736
rect 4666 1702 4700 1736
rect 5322 2830 5356 2864
rect 5514 2830 5548 2864
rect 5706 2830 5740 2864
rect 5418 2320 5452 2354
rect 5610 2320 5644 2354
rect 5802 2320 5836 2354
rect 5418 2212 5452 2246
rect 5610 2212 5644 2246
rect 5802 2212 5836 2246
rect 5322 1702 5356 1736
rect 5514 1702 5548 1736
rect 5706 1702 5740 1736
rect 6362 2830 6396 2864
rect 6554 2830 6588 2864
rect 6746 2830 6780 2864
rect 6458 2320 6492 2354
rect 6650 2320 6684 2354
rect 6842 2320 6876 2354
rect 6458 2212 6492 2246
rect 6650 2212 6684 2246
rect 6842 2212 6876 2246
rect 6362 1702 6396 1736
rect 6554 1702 6588 1736
rect 6746 1702 6780 1736
rect 7402 2830 7436 2864
rect 7594 2830 7628 2864
rect 7786 2830 7820 2864
rect 7498 2320 7532 2354
rect 7690 2320 7724 2354
rect 7882 2320 7916 2354
rect 7498 2212 7532 2246
rect 7690 2212 7724 2246
rect 7882 2212 7916 2246
rect 7402 1702 7436 1736
rect 7594 1702 7628 1736
rect 7786 1702 7820 1736
rect 8442 2830 8476 2864
rect 8634 2830 8668 2864
rect 8826 2830 8860 2864
rect 8538 2320 8572 2354
rect 8730 2320 8764 2354
rect 8922 2320 8956 2354
rect 8538 2212 8572 2246
rect 8730 2212 8764 2246
rect 8922 2212 8956 2246
rect 8442 1702 8476 1736
rect 8634 1702 8668 1736
rect 8826 1702 8860 1736
rect 9482 2830 9516 2864
rect 9674 2830 9708 2864
rect 9866 2830 9900 2864
rect 9578 2320 9612 2354
rect 9770 2320 9804 2354
rect 9962 2320 9996 2354
rect 9578 2212 9612 2246
rect 9770 2212 9804 2246
rect 9962 2212 9996 2246
rect 9482 1702 9516 1736
rect 9674 1702 9708 1736
rect 9866 1702 9900 1736
rect 10522 2830 10556 2864
rect 10714 2830 10748 2864
rect 10906 2830 10940 2864
rect 10618 2320 10652 2354
rect 10810 2320 10844 2354
rect 11002 2320 11036 2354
rect 10618 2212 10652 2246
rect 10810 2212 10844 2246
rect 11002 2212 11036 2246
rect 10522 1702 10556 1736
rect 10714 1702 10748 1736
rect 10906 1702 10940 1736
rect 11902 2830 11936 2864
rect 12094 2830 12128 2864
rect 12286 2830 12320 2864
rect 11998 2320 12032 2354
rect 12190 2320 12224 2354
rect 12382 2320 12416 2354
rect 11998 2212 12032 2246
rect 12190 2212 12224 2246
rect 12382 2212 12416 2246
rect 11902 1702 11936 1736
rect 12094 1702 12128 1736
rect 12286 1702 12320 1736
rect 12942 2830 12976 2864
rect 13134 2830 13168 2864
rect 13326 2830 13360 2864
rect 13038 2320 13072 2354
rect 13230 2320 13264 2354
rect 13422 2320 13456 2354
rect 13038 2212 13072 2246
rect 13230 2212 13264 2246
rect 13422 2212 13456 2246
rect 12942 1702 12976 1736
rect 13134 1702 13168 1736
rect 13326 1702 13360 1736
rect 13982 2830 14016 2864
rect 14174 2830 14208 2864
rect 14366 2830 14400 2864
rect 14078 2320 14112 2354
rect 14270 2320 14304 2354
rect 14462 2320 14496 2354
rect 14078 2212 14112 2246
rect 14270 2212 14304 2246
rect 14462 2212 14496 2246
rect 13982 1702 14016 1736
rect 14174 1702 14208 1736
rect 14366 1702 14400 1736
rect 15022 2830 15056 2864
rect 15214 2830 15248 2864
rect 15406 2830 15440 2864
rect 15118 2320 15152 2354
rect 15310 2320 15344 2354
rect 15502 2320 15536 2354
rect 15118 2212 15152 2246
rect 15310 2212 15344 2246
rect 15502 2212 15536 2246
rect 15022 1702 15056 1736
rect 15214 1702 15248 1736
rect 15406 1702 15440 1736
rect 16062 2830 16096 2864
rect 16254 2830 16288 2864
rect 16446 2830 16480 2864
rect 16158 2320 16192 2354
rect 16350 2320 16384 2354
rect 16542 2320 16576 2354
rect 16158 2212 16192 2246
rect 16350 2212 16384 2246
rect 16542 2212 16576 2246
rect 16062 1702 16096 1736
rect 16254 1702 16288 1736
rect 16446 1702 16480 1736
rect 17102 2830 17136 2864
rect 17294 2830 17328 2864
rect 17486 2830 17520 2864
rect 17198 2320 17232 2354
rect 17390 2320 17424 2354
rect 17582 2320 17616 2354
rect 17198 2212 17232 2246
rect 17390 2212 17424 2246
rect 17582 2212 17616 2246
rect 17102 1702 17136 1736
rect 17294 1702 17328 1736
rect 17486 1702 17520 1736
rect 18142 2830 18176 2864
rect 18334 2830 18368 2864
rect 18526 2830 18560 2864
rect 18238 2320 18272 2354
rect 18430 2320 18464 2354
rect 18622 2320 18656 2354
rect 18238 2212 18272 2246
rect 18430 2212 18464 2246
rect 18622 2212 18656 2246
rect 18142 1702 18176 1736
rect 18334 1702 18368 1736
rect 18526 1702 18560 1736
rect -1511 1248 -1477 1282
rect -1393 1248 -1359 1282
rect -1275 1248 -1241 1282
rect -1157 1248 -1123 1282
rect -1039 1248 -1005 1282
rect -921 1248 -887 1282
rect -1511 738 -1477 772
rect -1393 738 -1359 772
rect -1275 738 -1241 772
rect -1157 738 -1123 772
rect -1039 738 -1005 772
rect -921 738 -887 772
rect -471 1248 -437 1282
rect -353 1248 -319 1282
rect -235 1248 -201 1282
rect -117 1248 -83 1282
rect 1 1248 35 1282
rect 119 1248 153 1282
rect -471 738 -437 772
rect -353 738 -319 772
rect -235 738 -201 772
rect -117 738 -83 772
rect 1 738 35 772
rect 119 738 153 772
rect 569 1248 603 1282
rect 687 1248 721 1282
rect 805 1248 839 1282
rect 923 1248 957 1282
rect 1041 1248 1075 1282
rect 1159 1248 1193 1282
rect 569 738 603 772
rect 687 738 721 772
rect 805 738 839 772
rect 923 738 957 772
rect 1041 738 1075 772
rect 1159 738 1193 772
rect 1609 1248 1643 1282
rect 1727 1248 1761 1282
rect 1845 1248 1879 1282
rect 1963 1248 1997 1282
rect 2081 1248 2115 1282
rect 2199 1248 2233 1282
rect 1609 738 1643 772
rect 1727 738 1761 772
rect 1845 738 1879 772
rect 1963 738 1997 772
rect 2081 738 2115 772
rect 2199 738 2233 772
rect 2649 1248 2683 1282
rect 2767 1248 2801 1282
rect 2885 1248 2919 1282
rect 3003 1248 3037 1282
rect 3121 1248 3155 1282
rect 3239 1248 3273 1282
rect 2649 738 2683 772
rect 2767 738 2801 772
rect 2885 738 2919 772
rect 3003 738 3037 772
rect 3121 738 3155 772
rect 3239 738 3273 772
rect 4293 1408 4327 1442
rect 4411 1408 4445 1442
rect 4529 1408 4563 1442
rect 4647 1408 4681 1442
rect 4765 1408 4799 1442
rect 4883 1408 4917 1442
rect 4293 898 4327 932
rect 4411 898 4445 932
rect 4529 898 4563 932
rect 4647 898 4681 932
rect 4765 898 4799 932
rect 4883 898 4917 932
rect 5333 1408 5367 1442
rect 5451 1408 5485 1442
rect 5569 1408 5603 1442
rect 5687 1408 5721 1442
rect 5805 1408 5839 1442
rect 5923 1408 5957 1442
rect 5333 898 5367 932
rect 5451 898 5485 932
rect 5569 898 5603 932
rect 5687 898 5721 932
rect 5805 898 5839 932
rect 5923 898 5957 932
rect 6373 1408 6407 1442
rect 6491 1408 6525 1442
rect 6609 1408 6643 1442
rect 6727 1408 6761 1442
rect 6845 1408 6879 1442
rect 6963 1408 6997 1442
rect 6373 898 6407 932
rect 6491 898 6525 932
rect 6609 898 6643 932
rect 6727 898 6761 932
rect 6845 898 6879 932
rect 6963 898 6997 932
rect 7413 1408 7447 1442
rect 7531 1408 7565 1442
rect 7649 1408 7683 1442
rect 7767 1408 7801 1442
rect 7885 1408 7919 1442
rect 8003 1408 8037 1442
rect 7413 898 7447 932
rect 7531 898 7565 932
rect 7649 898 7683 932
rect 7767 898 7801 932
rect 7885 898 7919 932
rect 8003 898 8037 932
rect 8453 1408 8487 1442
rect 8571 1408 8605 1442
rect 8689 1408 8723 1442
rect 8807 1408 8841 1442
rect 8925 1408 8959 1442
rect 9043 1408 9077 1442
rect 8453 898 8487 932
rect 8571 898 8605 932
rect 8689 898 8723 932
rect 8807 898 8841 932
rect 8925 898 8959 932
rect 9043 898 9077 932
rect 9493 1408 9527 1442
rect 9611 1408 9645 1442
rect 9729 1408 9763 1442
rect 9847 1408 9881 1442
rect 9965 1408 9999 1442
rect 10083 1408 10117 1442
rect 9493 898 9527 932
rect 9611 898 9645 932
rect 9729 898 9763 932
rect 9847 898 9881 932
rect 9965 898 9999 932
rect 10083 898 10117 932
rect 10533 1408 10567 1442
rect 10651 1408 10685 1442
rect 10769 1408 10803 1442
rect 10887 1408 10921 1442
rect 11005 1408 11039 1442
rect 11123 1408 11157 1442
rect 10533 898 10567 932
rect 10651 898 10685 932
rect 10769 898 10803 932
rect 10887 898 10921 932
rect 11005 898 11039 932
rect 11123 898 11157 932
rect 11913 1408 11947 1442
rect 12031 1408 12065 1442
rect 12149 1408 12183 1442
rect 12267 1408 12301 1442
rect 12385 1408 12419 1442
rect 12503 1408 12537 1442
rect 11913 898 11947 932
rect 12031 898 12065 932
rect 12149 898 12183 932
rect 12267 898 12301 932
rect 12385 898 12419 932
rect 12503 898 12537 932
rect 12953 1408 12987 1442
rect 13071 1408 13105 1442
rect 13189 1408 13223 1442
rect 13307 1408 13341 1442
rect 13425 1408 13459 1442
rect 13543 1408 13577 1442
rect 12953 898 12987 932
rect 13071 898 13105 932
rect 13189 898 13223 932
rect 13307 898 13341 932
rect 13425 898 13459 932
rect 13543 898 13577 932
rect 13993 1408 14027 1442
rect 14111 1408 14145 1442
rect 14229 1408 14263 1442
rect 14347 1408 14381 1442
rect 14465 1408 14499 1442
rect 14583 1408 14617 1442
rect 13993 898 14027 932
rect 14111 898 14145 932
rect 14229 898 14263 932
rect 14347 898 14381 932
rect 14465 898 14499 932
rect 14583 898 14617 932
rect 15033 1408 15067 1442
rect 15151 1408 15185 1442
rect 15269 1408 15303 1442
rect 15387 1408 15421 1442
rect 15505 1408 15539 1442
rect 15623 1408 15657 1442
rect 15033 898 15067 932
rect 15151 898 15185 932
rect 15269 898 15303 932
rect 15387 898 15421 932
rect 15505 898 15539 932
rect 15623 898 15657 932
rect 16073 1408 16107 1442
rect 16191 1408 16225 1442
rect 16309 1408 16343 1442
rect 16427 1408 16461 1442
rect 16545 1408 16579 1442
rect 16663 1408 16697 1442
rect 16073 898 16107 932
rect 16191 898 16225 932
rect 16309 898 16343 932
rect 16427 898 16461 932
rect 16545 898 16579 932
rect 16663 898 16697 932
rect 17113 1408 17147 1442
rect 17231 1408 17265 1442
rect 17349 1408 17383 1442
rect 17467 1408 17501 1442
rect 17585 1408 17619 1442
rect 17703 1408 17737 1442
rect 17113 898 17147 932
rect 17231 898 17265 932
rect 17349 898 17383 932
rect 17467 898 17501 932
rect 17585 898 17619 932
rect 17703 898 17737 932
rect 18153 1408 18187 1442
rect 18271 1408 18305 1442
rect 18389 1408 18423 1442
rect 18507 1408 18541 1442
rect 18625 1408 18659 1442
rect 18743 1408 18777 1442
rect 18153 898 18187 932
rect 18271 898 18305 932
rect 18389 898 18423 932
rect 18507 898 18541 932
rect 18625 898 18659 932
rect 18743 898 18777 932
rect -7352 -16 -7318 18
rect -7160 -16 -7126 18
rect -6968 -16 -6934 18
rect -6776 -16 -6742 18
rect -6584 -16 -6550 18
rect -7256 -526 -7222 -492
rect -7064 -526 -7030 -492
rect -6872 -526 -6838 -492
rect -6680 -526 -6646 -492
rect -6488 -526 -6454 -492
rect -7256 -634 -7222 -600
rect -7064 -634 -7030 -600
rect -6872 -634 -6838 -600
rect -6680 -634 -6646 -600
rect -6488 -634 -6454 -600
rect -7352 -1144 -7318 -1110
rect -7160 -1144 -7126 -1110
rect -6968 -1144 -6934 -1110
rect -6776 -1144 -6742 -1110
rect -6584 -1144 -6550 -1110
rect -7352 -1852 -7318 -1818
rect -7160 -1852 -7126 -1818
rect -6968 -1852 -6934 -1818
rect -7256 -2362 -7222 -2328
rect -7064 -2362 -7030 -2328
rect -6872 -2362 -6838 -2328
rect -7256 -2470 -7222 -2436
rect -7064 -2470 -7030 -2436
rect -6872 -2470 -6838 -2436
rect -7352 -2980 -7318 -2946
rect -7160 -2980 -7126 -2946
rect -6968 -2980 -6934 -2946
rect -6072 -1638 -6038 -70
rect -5762 -1638 -5728 -70
rect 4282 590 4316 624
rect 4474 590 4508 624
rect 4666 590 4700 624
rect 4378 80 4412 114
rect 4570 80 4604 114
rect 4762 80 4796 114
rect 4378 -28 4412 6
rect 4570 -28 4604 6
rect 4762 -28 4796 6
rect 4282 -538 4316 -504
rect 4474 -538 4508 -504
rect 4666 -538 4700 -504
rect 5322 590 5356 624
rect 5514 590 5548 624
rect 5706 590 5740 624
rect 5418 80 5452 114
rect 5610 80 5644 114
rect 5802 80 5836 114
rect 5418 -28 5452 6
rect 5610 -28 5644 6
rect 5802 -28 5836 6
rect 5322 -538 5356 -504
rect 5514 -538 5548 -504
rect 5706 -538 5740 -504
rect 6362 590 6396 624
rect 6554 590 6588 624
rect 6746 590 6780 624
rect 6458 80 6492 114
rect 6650 80 6684 114
rect 6842 80 6876 114
rect 6458 -28 6492 6
rect 6650 -28 6684 6
rect 6842 -28 6876 6
rect 6362 -538 6396 -504
rect 6554 -538 6588 -504
rect 6746 -538 6780 -504
rect 7402 590 7436 624
rect 7594 590 7628 624
rect 7786 590 7820 624
rect 7498 80 7532 114
rect 7690 80 7724 114
rect 7882 80 7916 114
rect 7498 -28 7532 6
rect 7690 -28 7724 6
rect 7882 -28 7916 6
rect 7402 -538 7436 -504
rect 7594 -538 7628 -504
rect 7786 -538 7820 -504
rect 8442 590 8476 624
rect 8634 590 8668 624
rect 8826 590 8860 624
rect 8538 80 8572 114
rect 8730 80 8764 114
rect 8922 80 8956 114
rect 8538 -28 8572 6
rect 8730 -28 8764 6
rect 8922 -28 8956 6
rect 8442 -538 8476 -504
rect 8634 -538 8668 -504
rect 8826 -538 8860 -504
rect 9482 590 9516 624
rect 9674 590 9708 624
rect 9866 590 9900 624
rect 9578 80 9612 114
rect 9770 80 9804 114
rect 9962 80 9996 114
rect 9578 -28 9612 6
rect 9770 -28 9804 6
rect 9962 -28 9996 6
rect 9482 -538 9516 -504
rect 9674 -538 9708 -504
rect 9866 -538 9900 -504
rect 10522 590 10556 624
rect 10714 590 10748 624
rect 10906 590 10940 624
rect 10618 80 10652 114
rect 10810 80 10844 114
rect 11002 80 11036 114
rect 10618 -28 10652 6
rect 10810 -28 10844 6
rect 11002 -28 11036 6
rect 10522 -538 10556 -504
rect 10714 -538 10748 -504
rect 10906 -538 10940 -504
rect 11902 590 11936 624
rect 12094 590 12128 624
rect 12286 590 12320 624
rect 11998 80 12032 114
rect 12190 80 12224 114
rect 12382 80 12416 114
rect 11998 -28 12032 6
rect 12190 -28 12224 6
rect 12382 -28 12416 6
rect 11902 -538 11936 -504
rect 12094 -538 12128 -504
rect 12286 -538 12320 -504
rect 12942 590 12976 624
rect 13134 590 13168 624
rect 13326 590 13360 624
rect 13038 80 13072 114
rect 13230 80 13264 114
rect 13422 80 13456 114
rect 13038 -28 13072 6
rect 13230 -28 13264 6
rect 13422 -28 13456 6
rect 12942 -538 12976 -504
rect 13134 -538 13168 -504
rect 13326 -538 13360 -504
rect 13982 590 14016 624
rect 14174 590 14208 624
rect 14366 590 14400 624
rect 14078 80 14112 114
rect 14270 80 14304 114
rect 14462 80 14496 114
rect 14078 -28 14112 6
rect 14270 -28 14304 6
rect 14462 -28 14496 6
rect 13982 -538 14016 -504
rect 14174 -538 14208 -504
rect 14366 -538 14400 -504
rect 15022 590 15056 624
rect 15214 590 15248 624
rect 15406 590 15440 624
rect 15118 80 15152 114
rect 15310 80 15344 114
rect 15502 80 15536 114
rect 15118 -28 15152 6
rect 15310 -28 15344 6
rect 15502 -28 15536 6
rect 15022 -538 15056 -504
rect 15214 -538 15248 -504
rect 15406 -538 15440 -504
rect 16062 590 16096 624
rect 16254 590 16288 624
rect 16446 590 16480 624
rect 16158 80 16192 114
rect 16350 80 16384 114
rect 16542 80 16576 114
rect 16158 -28 16192 6
rect 16350 -28 16384 6
rect 16542 -28 16576 6
rect 16062 -538 16096 -504
rect 16254 -538 16288 -504
rect 16446 -538 16480 -504
rect 17102 590 17136 624
rect 17294 590 17328 624
rect 17486 590 17520 624
rect 17198 80 17232 114
rect 17390 80 17424 114
rect 17582 80 17616 114
rect 17198 -28 17232 6
rect 17390 -28 17424 6
rect 17582 -28 17616 6
rect 17102 -538 17136 -504
rect 17294 -538 17328 -504
rect 17486 -538 17520 -504
rect 18142 590 18176 624
rect 18334 590 18368 624
rect 18526 590 18560 624
rect 18238 80 18272 114
rect 18430 80 18464 114
rect 18622 80 18656 114
rect 18238 -28 18272 6
rect 18430 -28 18464 6
rect 18622 -28 18656 6
rect 18142 -538 18176 -504
rect 18334 -538 18368 -504
rect 18526 -538 18560 -504
rect 4293 -832 4327 -798
rect 4411 -832 4445 -798
rect 4529 -832 4563 -798
rect 4647 -832 4681 -798
rect 4765 -832 4799 -798
rect 4883 -832 4917 -798
rect 4293 -1342 4327 -1308
rect 4411 -1342 4445 -1308
rect 4529 -1342 4563 -1308
rect 4647 -1342 4681 -1308
rect 4765 -1342 4799 -1308
rect 4883 -1342 4917 -1308
rect 5333 -832 5367 -798
rect 5451 -832 5485 -798
rect 5569 -832 5603 -798
rect 5687 -832 5721 -798
rect 5805 -832 5839 -798
rect 5923 -832 5957 -798
rect 5333 -1342 5367 -1308
rect 5451 -1342 5485 -1308
rect 5569 -1342 5603 -1308
rect 5687 -1342 5721 -1308
rect 5805 -1342 5839 -1308
rect 5923 -1342 5957 -1308
rect 6373 -832 6407 -798
rect 6491 -832 6525 -798
rect 6609 -832 6643 -798
rect 6727 -832 6761 -798
rect 6845 -832 6879 -798
rect 6963 -832 6997 -798
rect 6373 -1342 6407 -1308
rect 6491 -1342 6525 -1308
rect 6609 -1342 6643 -1308
rect 6727 -1342 6761 -1308
rect 6845 -1342 6879 -1308
rect 6963 -1342 6997 -1308
rect 7413 -832 7447 -798
rect 7531 -832 7565 -798
rect 7649 -832 7683 -798
rect 7767 -832 7801 -798
rect 7885 -832 7919 -798
rect 8003 -832 8037 -798
rect 7413 -1342 7447 -1308
rect 7531 -1342 7565 -1308
rect 7649 -1342 7683 -1308
rect 7767 -1342 7801 -1308
rect 7885 -1342 7919 -1308
rect 8003 -1342 8037 -1308
rect 8453 -832 8487 -798
rect 8571 -832 8605 -798
rect 8689 -832 8723 -798
rect 8807 -832 8841 -798
rect 8925 -832 8959 -798
rect 9043 -832 9077 -798
rect 8453 -1342 8487 -1308
rect 8571 -1342 8605 -1308
rect 8689 -1342 8723 -1308
rect 8807 -1342 8841 -1308
rect 8925 -1342 8959 -1308
rect 9043 -1342 9077 -1308
rect 9493 -832 9527 -798
rect 9611 -832 9645 -798
rect 9729 -832 9763 -798
rect 9847 -832 9881 -798
rect 9965 -832 9999 -798
rect 10083 -832 10117 -798
rect 9493 -1342 9527 -1308
rect 9611 -1342 9645 -1308
rect 9729 -1342 9763 -1308
rect 9847 -1342 9881 -1308
rect 9965 -1342 9999 -1308
rect 10083 -1342 10117 -1308
rect 10533 -832 10567 -798
rect 10651 -832 10685 -798
rect 10769 -832 10803 -798
rect 10887 -832 10921 -798
rect 11005 -832 11039 -798
rect 11123 -832 11157 -798
rect 10533 -1342 10567 -1308
rect 10651 -1342 10685 -1308
rect 10769 -1342 10803 -1308
rect 10887 -1342 10921 -1308
rect 11005 -1342 11039 -1308
rect 11123 -1342 11157 -1308
rect 11913 -832 11947 -798
rect 12031 -832 12065 -798
rect 12149 -832 12183 -798
rect 12267 -832 12301 -798
rect 12385 -832 12419 -798
rect 12503 -832 12537 -798
rect 11913 -1342 11947 -1308
rect 12031 -1342 12065 -1308
rect 12149 -1342 12183 -1308
rect 12267 -1342 12301 -1308
rect 12385 -1342 12419 -1308
rect 12503 -1342 12537 -1308
rect 12953 -832 12987 -798
rect 13071 -832 13105 -798
rect 13189 -832 13223 -798
rect 13307 -832 13341 -798
rect 13425 -832 13459 -798
rect 13543 -832 13577 -798
rect 12953 -1342 12987 -1308
rect 13071 -1342 13105 -1308
rect 13189 -1342 13223 -1308
rect 13307 -1342 13341 -1308
rect 13425 -1342 13459 -1308
rect 13543 -1342 13577 -1308
rect 13993 -832 14027 -798
rect 14111 -832 14145 -798
rect 14229 -832 14263 -798
rect 14347 -832 14381 -798
rect 14465 -832 14499 -798
rect 14583 -832 14617 -798
rect 13993 -1342 14027 -1308
rect 14111 -1342 14145 -1308
rect 14229 -1342 14263 -1308
rect 14347 -1342 14381 -1308
rect 14465 -1342 14499 -1308
rect 14583 -1342 14617 -1308
rect 15033 -832 15067 -798
rect 15151 -832 15185 -798
rect 15269 -832 15303 -798
rect 15387 -832 15421 -798
rect 15505 -832 15539 -798
rect 15623 -832 15657 -798
rect 15033 -1342 15067 -1308
rect 15151 -1342 15185 -1308
rect 15269 -1342 15303 -1308
rect 15387 -1342 15421 -1308
rect 15505 -1342 15539 -1308
rect 15623 -1342 15657 -1308
rect 16073 -832 16107 -798
rect 16191 -832 16225 -798
rect 16309 -832 16343 -798
rect 16427 -832 16461 -798
rect 16545 -832 16579 -798
rect 16663 -832 16697 -798
rect 16073 -1342 16107 -1308
rect 16191 -1342 16225 -1308
rect 16309 -1342 16343 -1308
rect 16427 -1342 16461 -1308
rect 16545 -1342 16579 -1308
rect 16663 -1342 16697 -1308
rect 17113 -832 17147 -798
rect 17231 -832 17265 -798
rect 17349 -832 17383 -798
rect 17467 -832 17501 -798
rect 17585 -832 17619 -798
rect 17703 -832 17737 -798
rect 17113 -1342 17147 -1308
rect 17231 -1342 17265 -1308
rect 17349 -1342 17383 -1308
rect 17467 -1342 17501 -1308
rect 17585 -1342 17619 -1308
rect 17703 -1342 17737 -1308
rect 18153 -832 18187 -798
rect 18271 -832 18305 -798
rect 18389 -832 18423 -798
rect 18507 -832 18541 -798
rect 18625 -832 18659 -798
rect 18743 -832 18777 -798
rect 18153 -1342 18187 -1308
rect 18271 -1342 18305 -1308
rect 18389 -1342 18423 -1308
rect 18507 -1342 18541 -1308
rect 18625 -1342 18659 -1308
rect 18743 -1342 18777 -1308
rect 4282 -1650 4316 -1616
rect 4474 -1650 4508 -1616
rect 4666 -1650 4700 -1616
rect 4378 -2160 4412 -2126
rect 4570 -2160 4604 -2126
rect 4762 -2160 4796 -2126
rect 4378 -2268 4412 -2234
rect 4570 -2268 4604 -2234
rect 4762 -2268 4796 -2234
rect 4282 -2778 4316 -2744
rect 4474 -2778 4508 -2744
rect 4666 -2778 4700 -2744
rect 5322 -1650 5356 -1616
rect 5514 -1650 5548 -1616
rect 5706 -1650 5740 -1616
rect 5418 -2160 5452 -2126
rect 5610 -2160 5644 -2126
rect 5802 -2160 5836 -2126
rect 5418 -2268 5452 -2234
rect 5610 -2268 5644 -2234
rect 5802 -2268 5836 -2234
rect 5322 -2778 5356 -2744
rect 5514 -2778 5548 -2744
rect 5706 -2778 5740 -2744
rect 6362 -1650 6396 -1616
rect 6554 -1650 6588 -1616
rect 6746 -1650 6780 -1616
rect 6458 -2160 6492 -2126
rect 6650 -2160 6684 -2126
rect 6842 -2160 6876 -2126
rect 6458 -2268 6492 -2234
rect 6650 -2268 6684 -2234
rect 6842 -2268 6876 -2234
rect 6362 -2778 6396 -2744
rect 6554 -2778 6588 -2744
rect 6746 -2778 6780 -2744
rect 7402 -1650 7436 -1616
rect 7594 -1650 7628 -1616
rect 7786 -1650 7820 -1616
rect 7498 -2160 7532 -2126
rect 7690 -2160 7724 -2126
rect 7882 -2160 7916 -2126
rect 7498 -2268 7532 -2234
rect 7690 -2268 7724 -2234
rect 7882 -2268 7916 -2234
rect 7402 -2778 7436 -2744
rect 7594 -2778 7628 -2744
rect 7786 -2778 7820 -2744
rect 8442 -1650 8476 -1616
rect 8634 -1650 8668 -1616
rect 8826 -1650 8860 -1616
rect 8538 -2160 8572 -2126
rect 8730 -2160 8764 -2126
rect 8922 -2160 8956 -2126
rect 8538 -2268 8572 -2234
rect 8730 -2268 8764 -2234
rect 8922 -2268 8956 -2234
rect 8442 -2778 8476 -2744
rect 8634 -2778 8668 -2744
rect 8826 -2778 8860 -2744
rect 11902 -1650 11936 -1616
rect 12094 -1650 12128 -1616
rect 12286 -1650 12320 -1616
rect 11998 -2160 12032 -2126
rect 12190 -2160 12224 -2126
rect 12382 -2160 12416 -2126
rect 11998 -2268 12032 -2234
rect 12190 -2268 12224 -2234
rect 12382 -2268 12416 -2234
rect 11902 -2778 11936 -2744
rect 12094 -2778 12128 -2744
rect 12286 -2778 12320 -2744
rect 12942 -1650 12976 -1616
rect 13134 -1650 13168 -1616
rect 13326 -1650 13360 -1616
rect 13038 -2160 13072 -2126
rect 13230 -2160 13264 -2126
rect 13422 -2160 13456 -2126
rect 13038 -2268 13072 -2234
rect 13230 -2268 13264 -2234
rect 13422 -2268 13456 -2234
rect 12942 -2778 12976 -2744
rect 13134 -2778 13168 -2744
rect 13326 -2778 13360 -2744
rect 13982 -1650 14016 -1616
rect 14174 -1650 14208 -1616
rect 14366 -1650 14400 -1616
rect 14078 -2160 14112 -2126
rect 14270 -2160 14304 -2126
rect 14462 -2160 14496 -2126
rect 14078 -2268 14112 -2234
rect 14270 -2268 14304 -2234
rect 14462 -2268 14496 -2234
rect 13982 -2778 14016 -2744
rect 14174 -2778 14208 -2744
rect 14366 -2778 14400 -2744
rect 15022 -1650 15056 -1616
rect 15214 -1650 15248 -1616
rect 15406 -1650 15440 -1616
rect 15118 -2160 15152 -2126
rect 15310 -2160 15344 -2126
rect 15502 -2160 15536 -2126
rect 15118 -2268 15152 -2234
rect 15310 -2268 15344 -2234
rect 15502 -2268 15536 -2234
rect 15022 -2778 15056 -2744
rect 15214 -2778 15248 -2744
rect 15406 -2778 15440 -2744
rect 16062 -1650 16096 -1616
rect 16254 -1650 16288 -1616
rect 16446 -1650 16480 -1616
rect 16158 -2160 16192 -2126
rect 16350 -2160 16384 -2126
rect 16542 -2160 16576 -2126
rect 16158 -2268 16192 -2234
rect 16350 -2268 16384 -2234
rect 16542 -2268 16576 -2234
rect 16062 -2778 16096 -2744
rect 16254 -2778 16288 -2744
rect 16446 -2778 16480 -2744
rect -7341 -3274 -7307 -3240
rect -7223 -3274 -7189 -3240
rect -7105 -3274 -7071 -3240
rect -6987 -3274 -6953 -3240
rect -6869 -3274 -6835 -3240
rect -6751 -3274 -6717 -3240
rect -7341 -3784 -7307 -3750
rect -7223 -3784 -7189 -3750
rect -7105 -3784 -7071 -3750
rect -6987 -3784 -6953 -3750
rect -6869 -3784 -6835 -3750
rect -6751 -3784 -6717 -3750
rect 4293 -3072 4327 -3038
rect 4411 -3072 4445 -3038
rect 4529 -3072 4563 -3038
rect 4647 -3072 4681 -3038
rect 4765 -3072 4799 -3038
rect 4883 -3072 4917 -3038
rect 4293 -3582 4327 -3548
rect 4411 -3582 4445 -3548
rect 4529 -3582 4563 -3548
rect 4647 -3582 4681 -3548
rect 4765 -3582 4799 -3548
rect 4883 -3582 4917 -3548
rect 5333 -3072 5367 -3038
rect 5451 -3072 5485 -3038
rect 5569 -3072 5603 -3038
rect 5687 -3072 5721 -3038
rect 5805 -3072 5839 -3038
rect 5923 -3072 5957 -3038
rect 5333 -3582 5367 -3548
rect 5451 -3582 5485 -3548
rect 5569 -3582 5603 -3548
rect 5687 -3582 5721 -3548
rect 5805 -3582 5839 -3548
rect 5923 -3582 5957 -3548
rect 6373 -3072 6407 -3038
rect 6491 -3072 6525 -3038
rect 6609 -3072 6643 -3038
rect 6727 -3072 6761 -3038
rect 6845 -3072 6879 -3038
rect 6963 -3072 6997 -3038
rect 6373 -3582 6407 -3548
rect 6491 -3582 6525 -3548
rect 6609 -3582 6643 -3548
rect 6727 -3582 6761 -3548
rect 6845 -3582 6879 -3548
rect 6963 -3582 6997 -3548
rect 7413 -3072 7447 -3038
rect 7531 -3072 7565 -3038
rect 7649 -3072 7683 -3038
rect 7767 -3072 7801 -3038
rect 7885 -3072 7919 -3038
rect 8003 -3072 8037 -3038
rect 7413 -3582 7447 -3548
rect 7531 -3582 7565 -3548
rect 7649 -3582 7683 -3548
rect 7767 -3582 7801 -3548
rect 7885 -3582 7919 -3548
rect 8003 -3582 8037 -3548
rect 8453 -3072 8487 -3038
rect 8571 -3072 8605 -3038
rect 8689 -3072 8723 -3038
rect 8807 -3072 8841 -3038
rect 8925 -3072 8959 -3038
rect 9043 -3072 9077 -3038
rect 8453 -3582 8487 -3548
rect 8571 -3582 8605 -3548
rect 8689 -3582 8723 -3548
rect 8807 -3582 8841 -3548
rect 8925 -3582 8959 -3548
rect 9043 -3582 9077 -3548
rect 11913 -3072 11947 -3038
rect 12031 -3072 12065 -3038
rect 12149 -3072 12183 -3038
rect 12267 -3072 12301 -3038
rect 12385 -3072 12419 -3038
rect 12503 -3072 12537 -3038
rect 11913 -3582 11947 -3548
rect 12031 -3582 12065 -3548
rect 12149 -3582 12183 -3548
rect 12267 -3582 12301 -3548
rect 12385 -3582 12419 -3548
rect 12503 -3582 12537 -3548
rect 12953 -3072 12987 -3038
rect 13071 -3072 13105 -3038
rect 13189 -3072 13223 -3038
rect 13307 -3072 13341 -3038
rect 13425 -3072 13459 -3038
rect 13543 -3072 13577 -3038
rect 12953 -3582 12987 -3548
rect 13071 -3582 13105 -3548
rect 13189 -3582 13223 -3548
rect 13307 -3582 13341 -3548
rect 13425 -3582 13459 -3548
rect 13543 -3582 13577 -3548
rect 13993 -3072 14027 -3038
rect 14111 -3072 14145 -3038
rect 14229 -3072 14263 -3038
rect 14347 -3072 14381 -3038
rect 14465 -3072 14499 -3038
rect 14583 -3072 14617 -3038
rect 13993 -3582 14027 -3548
rect 14111 -3582 14145 -3548
rect 14229 -3582 14263 -3548
rect 14347 -3582 14381 -3548
rect 14465 -3582 14499 -3548
rect 14583 -3582 14617 -3548
rect 15033 -3072 15067 -3038
rect 15151 -3072 15185 -3038
rect 15269 -3072 15303 -3038
rect 15387 -3072 15421 -3038
rect 15505 -3072 15539 -3038
rect 15623 -3072 15657 -3038
rect 15033 -3582 15067 -3548
rect 15151 -3582 15185 -3548
rect 15269 -3582 15303 -3548
rect 15387 -3582 15421 -3548
rect 15505 -3582 15539 -3548
rect 15623 -3582 15657 -3548
rect 16073 -3072 16107 -3038
rect 16191 -3072 16225 -3038
rect 16309 -3072 16343 -3038
rect 16427 -3072 16461 -3038
rect 16545 -3072 16579 -3038
rect 16663 -3072 16697 -3038
rect 16073 -3582 16107 -3548
rect 16191 -3582 16225 -3548
rect 16309 -3582 16343 -3548
rect 16427 -3582 16461 -3548
rect 16545 -3582 16579 -3548
rect 16663 -3582 16697 -3548
<< xpolycontact >>
rect -1434 6170 -1152 6602
rect -1434 5338 -1152 5770
rect -1056 6170 -774 6602
rect -1056 5338 -774 5770
rect -678 6170 -396 6602
rect -678 5338 -396 5770
rect -300 6170 -18 6602
rect -300 5338 -18 5770
rect 78 6170 360 6602
rect 78 5338 360 5770
rect -1434 4802 -1152 5234
rect -1434 3970 -1152 4402
rect -1056 4802 -774 5234
rect -1056 3970 -774 4402
rect -678 4802 -396 5234
rect -678 3970 -396 4402
rect -300 4802 -18 5234
rect -300 3970 -18 4402
rect 78 4802 360 5234
rect 78 3970 360 4402
rect 1366 6170 1648 6602
rect 1366 5338 1648 5770
rect 1744 6170 2026 6602
rect 1744 5338 2026 5770
rect 2122 6170 2404 6602
rect 2122 5338 2404 5770
rect 2500 6170 2782 6602
rect 2500 5338 2782 5770
rect 2878 6170 3160 6602
rect 2878 5338 3160 5770
rect 1366 4802 1648 5234
rect 1366 3970 1648 4402
rect 1744 4802 2026 5234
rect 1744 3970 2026 4402
rect 2122 4802 2404 5234
rect 2122 3970 2404 4402
rect 2500 4802 2782 5234
rect 2500 3970 2782 4402
rect 2878 4802 3160 5234
rect 2878 3970 3160 4402
<< xpolyres >>
rect -1434 5770 -1152 6170
rect -1056 5770 -774 6170
rect -678 5770 -396 6170
rect -300 5770 -18 6170
rect 78 5770 360 6170
rect -1434 4402 -1152 4802
rect -1056 4402 -774 4802
rect -678 4402 -396 4802
rect -300 4402 -18 4802
rect 78 4402 360 4802
rect 1366 5770 1648 6170
rect 1744 5770 2026 6170
rect 2122 5770 2404 6170
rect 2500 5770 2782 6170
rect 2878 5770 3160 6170
rect 1366 4402 1648 4802
rect 1744 4402 2026 4802
rect 2122 4402 2404 4802
rect 2500 4402 2782 4802
rect 2878 4402 3160 4802
<< locali >>
rect -1564 6698 -1468 6732
rect 394 6698 490 6732
rect -1564 6636 -1530 6698
rect 456 6636 490 6698
rect -1564 3874 -1530 3936
rect 456 3874 490 3936
rect -1564 3840 -1468 3874
rect 394 3840 490 3874
rect 1236 6698 1332 6732
rect 3194 6698 3290 6732
rect 1236 6636 1270 6698
rect 3256 6636 3290 6698
rect 1236 3874 1270 3936
rect 3256 3874 3290 3936
rect 1236 3840 1332 3874
rect 3194 3840 3290 3874
rect 4320 5604 4416 5638
rect 7366 5604 7462 5638
rect 4320 5542 4354 5604
rect -1136 3784 68 3840
rect 1664 3784 2868 3840
rect -1144 3750 -1048 3784
rect -18 3750 78 3784
rect -1144 3688 -1110 3750
rect 44 3688 78 3750
rect -902 3648 -886 3682
rect -852 3648 -836 3682
rect -710 3648 -694 3682
rect -660 3648 -644 3682
rect -518 3648 -502 3682
rect -468 3648 -452 3682
rect -326 3648 -310 3682
rect -276 3648 -260 3682
rect -134 3648 -118 3682
rect -84 3648 -68 3682
rect -1030 3598 -996 3614
rect -1030 3206 -996 3222
rect -934 3598 -900 3614
rect -934 3206 -900 3222
rect -838 3598 -804 3614
rect -838 3206 -804 3222
rect -742 3598 -708 3614
rect -742 3206 -708 3222
rect -646 3598 -612 3614
rect -646 3206 -612 3222
rect -550 3598 -516 3614
rect -550 3206 -516 3222
rect -454 3598 -420 3614
rect -454 3206 -420 3222
rect -358 3598 -324 3614
rect -358 3206 -324 3222
rect -262 3598 -228 3614
rect -262 3206 -228 3222
rect -166 3598 -132 3614
rect -166 3206 -132 3222
rect -70 3598 -36 3614
rect -70 3206 -36 3222
rect -998 3138 -982 3172
rect -948 3138 -932 3172
rect -806 3138 -790 3172
rect -756 3138 -740 3172
rect -614 3138 -598 3172
rect -564 3138 -548 3172
rect -422 3138 -406 3172
rect -372 3138 -356 3172
rect -230 3138 -214 3172
rect -180 3138 -164 3172
rect -1144 3070 -1110 3132
rect 44 3070 78 3132
rect -1144 3060 -1048 3070
rect -1160 3036 -1048 3060
rect -18 3036 78 3070
rect 1656 3750 1752 3784
rect 2782 3750 2878 3784
rect 1656 3688 1690 3750
rect 2844 3688 2878 3750
rect 1898 3648 1914 3682
rect 1948 3648 1964 3682
rect 2090 3648 2106 3682
rect 2140 3648 2156 3682
rect 2282 3648 2298 3682
rect 2332 3648 2348 3682
rect 2474 3648 2490 3682
rect 2524 3648 2540 3682
rect 2666 3648 2682 3682
rect 2716 3648 2732 3682
rect 1770 3598 1804 3614
rect 1770 3206 1804 3222
rect 1866 3598 1900 3614
rect 1866 3206 1900 3222
rect 1962 3598 1996 3614
rect 1962 3206 1996 3222
rect 2058 3598 2092 3614
rect 2058 3206 2092 3222
rect 2154 3598 2188 3614
rect 2154 3206 2188 3222
rect 2250 3598 2284 3614
rect 2250 3206 2284 3222
rect 2346 3598 2380 3614
rect 2346 3206 2380 3222
rect 2442 3598 2476 3614
rect 2442 3206 2476 3222
rect 2538 3598 2572 3614
rect 2538 3206 2572 3222
rect 2634 3598 2668 3614
rect 2634 3206 2668 3222
rect 2730 3598 2764 3614
rect 2730 3206 2764 3222
rect 1802 3138 1818 3172
rect 1852 3138 1868 3172
rect 1994 3138 2010 3172
rect 2044 3138 2060 3172
rect 2186 3138 2202 3172
rect 2236 3138 2252 3172
rect 2378 3138 2394 3172
rect 2428 3138 2444 3172
rect 2570 3138 2586 3172
rect 2620 3138 2636 3172
rect 1656 3070 1690 3132
rect 2844 3070 2878 3132
rect 1656 3036 1752 3070
rect 2782 3036 2878 3070
rect 7428 5542 7462 5604
rect 4466 5502 4482 5536
rect 4516 5502 4532 5536
rect 4658 5502 4674 5536
rect 4708 5502 4724 5536
rect 4850 5502 4866 5536
rect 4900 5502 4916 5536
rect 5042 5502 5058 5536
rect 5092 5502 5108 5536
rect 5234 5502 5250 5536
rect 5284 5502 5300 5536
rect 5426 5502 5442 5536
rect 5476 5502 5492 5536
rect 5618 5502 5634 5536
rect 5668 5502 5684 5536
rect 5810 5502 5826 5536
rect 5860 5502 5876 5536
rect 6002 5502 6018 5536
rect 6052 5502 6068 5536
rect 6194 5502 6210 5536
rect 6244 5502 6260 5536
rect 6386 5502 6402 5536
rect 6436 5502 6452 5536
rect 6578 5502 6594 5536
rect 6628 5502 6644 5536
rect 6770 5502 6786 5536
rect 6820 5502 6836 5536
rect 6962 5502 6978 5536
rect 7012 5502 7028 5536
rect 7154 5502 7170 5536
rect 7204 5502 7220 5536
rect 4434 5452 4468 5468
rect 4434 5060 4468 5076
rect 4530 5452 4564 5468
rect 4530 5060 4564 5076
rect 4626 5452 4660 5468
rect 4626 5060 4660 5076
rect 4722 5452 4756 5468
rect 4722 5060 4756 5076
rect 4818 5452 4852 5468
rect 4818 5060 4852 5076
rect 4914 5452 4948 5468
rect 4914 5060 4948 5076
rect 5010 5452 5044 5468
rect 5010 5060 5044 5076
rect 5106 5452 5140 5468
rect 5106 5060 5140 5076
rect 5202 5452 5236 5468
rect 5202 5060 5236 5076
rect 5298 5452 5332 5468
rect 5298 5060 5332 5076
rect 5394 5452 5428 5468
rect 5394 5060 5428 5076
rect 5490 5452 5524 5468
rect 5490 5060 5524 5076
rect 5586 5452 5620 5468
rect 5586 5060 5620 5076
rect 5682 5452 5716 5468
rect 5682 5060 5716 5076
rect 5778 5452 5812 5468
rect 5778 5060 5812 5076
rect 5874 5452 5908 5468
rect 5874 5060 5908 5076
rect 5970 5452 6004 5468
rect 5970 5060 6004 5076
rect 6066 5452 6100 5468
rect 6066 5060 6100 5076
rect 6162 5452 6196 5468
rect 6162 5060 6196 5076
rect 6258 5452 6292 5468
rect 6258 5060 6292 5076
rect 6354 5452 6388 5468
rect 6354 5060 6388 5076
rect 6450 5452 6484 5468
rect 6450 5060 6484 5076
rect 6546 5452 6580 5468
rect 6546 5060 6580 5076
rect 6642 5452 6676 5468
rect 6642 5060 6676 5076
rect 6738 5452 6772 5468
rect 6738 5060 6772 5076
rect 6834 5452 6868 5468
rect 6834 5060 6868 5076
rect 6930 5452 6964 5468
rect 6930 5060 6964 5076
rect 7026 5452 7060 5468
rect 7026 5060 7060 5076
rect 7122 5452 7156 5468
rect 7122 5060 7156 5076
rect 7218 5452 7252 5468
rect 7218 5060 7252 5076
rect 7314 5452 7348 5468
rect 7314 5060 7348 5076
rect 4562 4992 4578 5026
rect 4612 4992 4628 5026
rect 4754 4992 4770 5026
rect 4804 4992 4820 5026
rect 4946 4992 4962 5026
rect 4996 4992 5012 5026
rect 5138 4992 5154 5026
rect 5188 4992 5204 5026
rect 5330 4992 5346 5026
rect 5380 4992 5396 5026
rect 5522 4992 5538 5026
rect 5572 4992 5588 5026
rect 5714 4992 5730 5026
rect 5764 4992 5780 5026
rect 5906 4992 5922 5026
rect 5956 4992 5972 5026
rect 6098 4992 6114 5026
rect 6148 4992 6164 5026
rect 6290 4992 6306 5026
rect 6340 4992 6356 5026
rect 6482 4992 6498 5026
rect 6532 4992 6548 5026
rect 6674 4992 6690 5026
rect 6724 4992 6740 5026
rect 6866 4992 6882 5026
rect 6916 4992 6932 5026
rect 7058 4992 7074 5026
rect 7108 4992 7124 5026
rect 7250 4992 7266 5026
rect 7300 4992 7316 5026
rect 4562 4884 4578 4918
rect 4612 4884 4628 4918
rect 4754 4884 4770 4918
rect 4804 4884 4820 4918
rect 4946 4884 4962 4918
rect 4996 4884 5012 4918
rect 5138 4884 5154 4918
rect 5188 4884 5204 4918
rect 5330 4884 5346 4918
rect 5380 4884 5396 4918
rect 5522 4884 5538 4918
rect 5572 4884 5588 4918
rect 5714 4884 5730 4918
rect 5764 4884 5780 4918
rect 5906 4884 5922 4918
rect 5956 4884 5972 4918
rect 6098 4884 6114 4918
rect 6148 4884 6164 4918
rect 6290 4884 6306 4918
rect 6340 4884 6356 4918
rect 6482 4884 6498 4918
rect 6532 4884 6548 4918
rect 6674 4884 6690 4918
rect 6724 4884 6740 4918
rect 6866 4884 6882 4918
rect 6916 4884 6932 4918
rect 7058 4884 7074 4918
rect 7108 4884 7124 4918
rect 7250 4884 7266 4918
rect 7300 4884 7316 4918
rect 4434 4834 4468 4850
rect 4434 4442 4468 4458
rect 4530 4834 4564 4850
rect 4530 4442 4564 4458
rect 4626 4834 4660 4850
rect 4626 4442 4660 4458
rect 4722 4834 4756 4850
rect 4722 4442 4756 4458
rect 4818 4834 4852 4850
rect 4818 4442 4852 4458
rect 4914 4834 4948 4850
rect 4914 4442 4948 4458
rect 5010 4834 5044 4850
rect 5010 4442 5044 4458
rect 5106 4834 5140 4850
rect 5106 4442 5140 4458
rect 5202 4834 5236 4850
rect 5202 4442 5236 4458
rect 5298 4834 5332 4850
rect 5298 4442 5332 4458
rect 5394 4834 5428 4850
rect 5394 4442 5428 4458
rect 5490 4834 5524 4850
rect 5490 4442 5524 4458
rect 5586 4834 5620 4850
rect 5586 4442 5620 4458
rect 5682 4834 5716 4850
rect 5682 4442 5716 4458
rect 5778 4834 5812 4850
rect 5778 4442 5812 4458
rect 5874 4834 5908 4850
rect 5874 4442 5908 4458
rect 5970 4834 6004 4850
rect 5970 4442 6004 4458
rect 6066 4834 6100 4850
rect 6066 4442 6100 4458
rect 6162 4834 6196 4850
rect 6162 4442 6196 4458
rect 6258 4834 6292 4850
rect 6258 4442 6292 4458
rect 6354 4834 6388 4850
rect 6354 4442 6388 4458
rect 6450 4834 6484 4850
rect 6450 4442 6484 4458
rect 6546 4834 6580 4850
rect 6546 4442 6580 4458
rect 6642 4834 6676 4850
rect 6642 4442 6676 4458
rect 6738 4834 6772 4850
rect 6738 4442 6772 4458
rect 6834 4834 6868 4850
rect 6834 4442 6868 4458
rect 6930 4834 6964 4850
rect 6930 4442 6964 4458
rect 7026 4834 7060 4850
rect 7026 4442 7060 4458
rect 7122 4834 7156 4850
rect 7122 4442 7156 4458
rect 7218 4834 7252 4850
rect 7218 4442 7252 4458
rect 7314 4834 7348 4850
rect 7314 4442 7348 4458
rect 4466 4374 4482 4408
rect 4516 4374 4532 4408
rect 4658 4374 4674 4408
rect 4708 4374 4724 4408
rect 4850 4374 4866 4408
rect 4900 4374 4916 4408
rect 5042 4374 5058 4408
rect 5092 4374 5108 4408
rect 5234 4374 5250 4408
rect 5284 4374 5300 4408
rect 5426 4374 5442 4408
rect 5476 4374 5492 4408
rect 5618 4374 5634 4408
rect 5668 4374 5684 4408
rect 5810 4374 5826 4408
rect 5860 4374 5876 4408
rect 6002 4374 6018 4408
rect 6052 4374 6068 4408
rect 6194 4374 6210 4408
rect 6244 4374 6260 4408
rect 6386 4374 6402 4408
rect 6436 4374 6452 4408
rect 6578 4374 6594 4408
rect 6628 4374 6644 4408
rect 6770 4374 6786 4408
rect 6820 4374 6836 4408
rect 6962 4374 6978 4408
rect 7012 4374 7028 4408
rect 7154 4374 7170 4408
rect 7204 4374 7220 4408
rect 4466 4266 4482 4300
rect 4516 4266 4532 4300
rect 4658 4266 4674 4300
rect 4708 4266 4724 4300
rect 4850 4266 4866 4300
rect 4900 4266 4916 4300
rect 5042 4266 5058 4300
rect 5092 4266 5108 4300
rect 5234 4266 5250 4300
rect 5284 4266 5300 4300
rect 5426 4266 5442 4300
rect 5476 4266 5492 4300
rect 5618 4266 5634 4300
rect 5668 4266 5684 4300
rect 5810 4266 5826 4300
rect 5860 4266 5876 4300
rect 6002 4266 6018 4300
rect 6052 4266 6068 4300
rect 6194 4266 6210 4300
rect 6244 4266 6260 4300
rect 6386 4266 6402 4300
rect 6436 4266 6452 4300
rect 6578 4266 6594 4300
rect 6628 4266 6644 4300
rect 6770 4266 6786 4300
rect 6820 4266 6836 4300
rect 6962 4266 6978 4300
rect 7012 4266 7028 4300
rect 7154 4266 7170 4300
rect 7204 4266 7220 4300
rect 4434 4216 4468 4232
rect 4434 3824 4468 3840
rect 4530 4216 4564 4232
rect 4530 3824 4564 3840
rect 4626 4216 4660 4232
rect 4626 3824 4660 3840
rect 4722 4216 4756 4232
rect 4722 3824 4756 3840
rect 4818 4216 4852 4232
rect 4818 3824 4852 3840
rect 4914 4216 4948 4232
rect 4914 3824 4948 3840
rect 5010 4216 5044 4232
rect 5010 3824 5044 3840
rect 5106 4216 5140 4232
rect 5106 3824 5140 3840
rect 5202 4216 5236 4232
rect 5202 3824 5236 3840
rect 5298 4216 5332 4232
rect 5298 3824 5332 3840
rect 5394 4216 5428 4232
rect 5394 3824 5428 3840
rect 5490 4216 5524 4232
rect 5490 3824 5524 3840
rect 5586 4216 5620 4232
rect 5586 3824 5620 3840
rect 5682 4216 5716 4232
rect 5682 3824 5716 3840
rect 5778 4216 5812 4232
rect 5778 3824 5812 3840
rect 5874 4216 5908 4232
rect 5874 3824 5908 3840
rect 5970 4216 6004 4232
rect 5970 3824 6004 3840
rect 6066 4216 6100 4232
rect 6066 3824 6100 3840
rect 6162 4216 6196 4232
rect 6162 3824 6196 3840
rect 6258 4216 6292 4232
rect 6258 3824 6292 3840
rect 6354 4216 6388 4232
rect 6354 3824 6388 3840
rect 6450 4216 6484 4232
rect 6450 3824 6484 3840
rect 6546 4216 6580 4232
rect 6546 3824 6580 3840
rect 6642 4216 6676 4232
rect 6642 3824 6676 3840
rect 6738 4216 6772 4232
rect 6738 3824 6772 3840
rect 6834 4216 6868 4232
rect 6834 3824 6868 3840
rect 6930 4216 6964 4232
rect 6930 3824 6964 3840
rect 7026 4216 7060 4232
rect 7026 3824 7060 3840
rect 7122 4216 7156 4232
rect 7122 3824 7156 3840
rect 7218 4216 7252 4232
rect 7218 3824 7252 3840
rect 7314 4216 7348 4232
rect 7314 3824 7348 3840
rect 4562 3756 4578 3790
rect 4612 3756 4628 3790
rect 4754 3756 4770 3790
rect 4804 3756 4820 3790
rect 4946 3756 4962 3790
rect 4996 3756 5012 3790
rect 5138 3756 5154 3790
rect 5188 3756 5204 3790
rect 5330 3756 5346 3790
rect 5380 3756 5396 3790
rect 5522 3756 5538 3790
rect 5572 3756 5588 3790
rect 5714 3756 5730 3790
rect 5764 3756 5780 3790
rect 5906 3756 5922 3790
rect 5956 3756 5972 3790
rect 6098 3756 6114 3790
rect 6148 3756 6164 3790
rect 6290 3756 6306 3790
rect 6340 3756 6356 3790
rect 6482 3756 6498 3790
rect 6532 3756 6548 3790
rect 6674 3756 6690 3790
rect 6724 3756 6740 3790
rect 6866 3756 6882 3790
rect 6916 3756 6932 3790
rect 7058 3756 7074 3790
rect 7108 3756 7124 3790
rect 7250 3756 7266 3790
rect 7300 3756 7316 3790
rect 4562 3648 4578 3682
rect 4612 3648 4628 3682
rect 4754 3648 4770 3682
rect 4804 3648 4820 3682
rect 4946 3648 4962 3682
rect 4996 3648 5012 3682
rect 5138 3648 5154 3682
rect 5188 3648 5204 3682
rect 5330 3648 5346 3682
rect 5380 3648 5396 3682
rect 5522 3648 5538 3682
rect 5572 3648 5588 3682
rect 5714 3648 5730 3682
rect 5764 3648 5780 3682
rect 5906 3648 5922 3682
rect 5956 3648 5972 3682
rect 6098 3648 6114 3682
rect 6148 3648 6164 3682
rect 6290 3648 6306 3682
rect 6340 3648 6356 3682
rect 6482 3648 6498 3682
rect 6532 3648 6548 3682
rect 6674 3648 6690 3682
rect 6724 3648 6740 3682
rect 6866 3648 6882 3682
rect 6916 3648 6932 3682
rect 7058 3648 7074 3682
rect 7108 3648 7124 3682
rect 7250 3648 7266 3682
rect 7300 3648 7316 3682
rect 4434 3598 4468 3614
rect 4434 3206 4468 3222
rect 4530 3598 4564 3614
rect 4530 3206 4564 3222
rect 4626 3598 4660 3614
rect 4626 3206 4660 3222
rect 4722 3598 4756 3614
rect 4722 3206 4756 3222
rect 4818 3598 4852 3614
rect 4818 3206 4852 3222
rect 4914 3598 4948 3614
rect 4914 3206 4948 3222
rect 5010 3598 5044 3614
rect 5010 3206 5044 3222
rect 5106 3598 5140 3614
rect 5106 3206 5140 3222
rect 5202 3598 5236 3614
rect 5202 3206 5236 3222
rect 5298 3598 5332 3614
rect 5298 3206 5332 3222
rect 5394 3598 5428 3614
rect 5394 3206 5428 3222
rect 5490 3598 5524 3614
rect 5490 3206 5524 3222
rect 5586 3598 5620 3614
rect 5586 3206 5620 3222
rect 5682 3598 5716 3614
rect 5682 3206 5716 3222
rect 5778 3598 5812 3614
rect 5778 3206 5812 3222
rect 5874 3598 5908 3614
rect 5874 3206 5908 3222
rect 5970 3598 6004 3614
rect 5970 3206 6004 3222
rect 6066 3598 6100 3614
rect 6066 3206 6100 3222
rect 6162 3598 6196 3614
rect 6162 3206 6196 3222
rect 6258 3598 6292 3614
rect 6258 3206 6292 3222
rect 6354 3598 6388 3614
rect 6354 3206 6388 3222
rect 6450 3598 6484 3614
rect 6450 3206 6484 3222
rect 6546 3598 6580 3614
rect 6546 3206 6580 3222
rect 6642 3598 6676 3614
rect 6642 3206 6676 3222
rect 6738 3598 6772 3614
rect 6738 3206 6772 3222
rect 6834 3598 6868 3614
rect 6834 3206 6868 3222
rect 6930 3598 6964 3614
rect 6930 3206 6964 3222
rect 7026 3598 7060 3614
rect 7026 3206 7060 3222
rect 7122 3598 7156 3614
rect 7122 3206 7156 3222
rect 7218 3598 7252 3614
rect 7218 3206 7252 3222
rect 7314 3598 7348 3614
rect 7314 3206 7348 3222
rect 4466 3138 4482 3172
rect 4516 3138 4532 3172
rect 4658 3138 4674 3172
rect 4708 3138 4724 3172
rect 4850 3138 4866 3172
rect 4900 3138 4916 3172
rect 5042 3138 5058 3172
rect 5092 3138 5108 3172
rect 5234 3138 5250 3172
rect 5284 3138 5300 3172
rect 5426 3138 5442 3172
rect 5476 3138 5492 3172
rect 5618 3138 5634 3172
rect 5668 3138 5684 3172
rect 5810 3138 5826 3172
rect 5860 3138 5876 3172
rect 6002 3138 6018 3172
rect 6052 3138 6068 3172
rect 6194 3138 6210 3172
rect 6244 3138 6260 3172
rect 6386 3138 6402 3172
rect 6436 3138 6452 3172
rect 6578 3138 6594 3172
rect 6628 3138 6644 3172
rect 6770 3138 6786 3172
rect 6820 3138 6836 3172
rect 6962 3138 6978 3172
rect 7012 3138 7028 3172
rect 7154 3138 7170 3172
rect 7204 3138 7220 3172
rect 4320 3070 4354 3132
rect 7428 3070 7462 3132
rect 4320 3036 4416 3070
rect 7366 3060 7462 3070
rect 7960 5604 8056 5638
rect 11006 5604 11102 5638
rect 7960 5542 7994 5604
rect 11068 5542 11102 5604
rect 8106 5502 8122 5536
rect 8156 5502 8172 5536
rect 8298 5502 8314 5536
rect 8348 5502 8364 5536
rect 8490 5502 8506 5536
rect 8540 5502 8556 5536
rect 8682 5502 8698 5536
rect 8732 5502 8748 5536
rect 8874 5502 8890 5536
rect 8924 5502 8940 5536
rect 9066 5502 9082 5536
rect 9116 5502 9132 5536
rect 9258 5502 9274 5536
rect 9308 5502 9324 5536
rect 9450 5502 9466 5536
rect 9500 5502 9516 5536
rect 9642 5502 9658 5536
rect 9692 5502 9708 5536
rect 9834 5502 9850 5536
rect 9884 5502 9900 5536
rect 10026 5502 10042 5536
rect 10076 5502 10092 5536
rect 10218 5502 10234 5536
rect 10268 5502 10284 5536
rect 10410 5502 10426 5536
rect 10460 5502 10476 5536
rect 10602 5502 10618 5536
rect 10652 5502 10668 5536
rect 10794 5502 10810 5536
rect 10844 5502 10860 5536
rect 8074 5452 8108 5468
rect 8074 5060 8108 5076
rect 8170 5452 8204 5468
rect 8170 5060 8204 5076
rect 8266 5452 8300 5468
rect 8266 5060 8300 5076
rect 8362 5452 8396 5468
rect 8362 5060 8396 5076
rect 8458 5452 8492 5468
rect 8458 5060 8492 5076
rect 8554 5452 8588 5468
rect 8554 5060 8588 5076
rect 8650 5452 8684 5468
rect 8650 5060 8684 5076
rect 8746 5452 8780 5468
rect 8746 5060 8780 5076
rect 8842 5452 8876 5468
rect 8842 5060 8876 5076
rect 8938 5452 8972 5468
rect 8938 5060 8972 5076
rect 9034 5452 9068 5468
rect 9034 5060 9068 5076
rect 9130 5452 9164 5468
rect 9130 5060 9164 5076
rect 9226 5452 9260 5468
rect 9226 5060 9260 5076
rect 9322 5452 9356 5468
rect 9322 5060 9356 5076
rect 9418 5452 9452 5468
rect 9418 5060 9452 5076
rect 9514 5452 9548 5468
rect 9514 5060 9548 5076
rect 9610 5452 9644 5468
rect 9610 5060 9644 5076
rect 9706 5452 9740 5468
rect 9706 5060 9740 5076
rect 9802 5452 9836 5468
rect 9802 5060 9836 5076
rect 9898 5452 9932 5468
rect 9898 5060 9932 5076
rect 9994 5452 10028 5468
rect 9994 5060 10028 5076
rect 10090 5452 10124 5468
rect 10090 5060 10124 5076
rect 10186 5452 10220 5468
rect 10186 5060 10220 5076
rect 10282 5452 10316 5468
rect 10282 5060 10316 5076
rect 10378 5452 10412 5468
rect 10378 5060 10412 5076
rect 10474 5452 10508 5468
rect 10474 5060 10508 5076
rect 10570 5452 10604 5468
rect 10570 5060 10604 5076
rect 10666 5452 10700 5468
rect 10666 5060 10700 5076
rect 10762 5452 10796 5468
rect 10762 5060 10796 5076
rect 10858 5452 10892 5468
rect 10858 5060 10892 5076
rect 10954 5452 10988 5468
rect 10954 5060 10988 5076
rect 8202 4992 8218 5026
rect 8252 4992 8268 5026
rect 8394 4992 8410 5026
rect 8444 4992 8460 5026
rect 8586 4992 8602 5026
rect 8636 4992 8652 5026
rect 8778 4992 8794 5026
rect 8828 4992 8844 5026
rect 8970 4992 8986 5026
rect 9020 4992 9036 5026
rect 9162 4992 9178 5026
rect 9212 4992 9228 5026
rect 9354 4992 9370 5026
rect 9404 4992 9420 5026
rect 9546 4992 9562 5026
rect 9596 4992 9612 5026
rect 9738 4992 9754 5026
rect 9788 4992 9804 5026
rect 9930 4992 9946 5026
rect 9980 4992 9996 5026
rect 10122 4992 10138 5026
rect 10172 4992 10188 5026
rect 10314 4992 10330 5026
rect 10364 4992 10380 5026
rect 10506 4992 10522 5026
rect 10556 4992 10572 5026
rect 10698 4992 10714 5026
rect 10748 4992 10764 5026
rect 10890 4992 10906 5026
rect 10940 4992 10956 5026
rect 8202 4884 8218 4918
rect 8252 4884 8268 4918
rect 8394 4884 8410 4918
rect 8444 4884 8460 4918
rect 8586 4884 8602 4918
rect 8636 4884 8652 4918
rect 8778 4884 8794 4918
rect 8828 4884 8844 4918
rect 8970 4884 8986 4918
rect 9020 4884 9036 4918
rect 9162 4884 9178 4918
rect 9212 4884 9228 4918
rect 9354 4884 9370 4918
rect 9404 4884 9420 4918
rect 9546 4884 9562 4918
rect 9596 4884 9612 4918
rect 9738 4884 9754 4918
rect 9788 4884 9804 4918
rect 9930 4884 9946 4918
rect 9980 4884 9996 4918
rect 10122 4884 10138 4918
rect 10172 4884 10188 4918
rect 10314 4884 10330 4918
rect 10364 4884 10380 4918
rect 10506 4884 10522 4918
rect 10556 4884 10572 4918
rect 10698 4884 10714 4918
rect 10748 4884 10764 4918
rect 10890 4884 10906 4918
rect 10940 4884 10956 4918
rect 8074 4834 8108 4850
rect 8074 4442 8108 4458
rect 8170 4834 8204 4850
rect 8170 4442 8204 4458
rect 8266 4834 8300 4850
rect 8266 4442 8300 4458
rect 8362 4834 8396 4850
rect 8362 4442 8396 4458
rect 8458 4834 8492 4850
rect 8458 4442 8492 4458
rect 8554 4834 8588 4850
rect 8554 4442 8588 4458
rect 8650 4834 8684 4850
rect 8650 4442 8684 4458
rect 8746 4834 8780 4850
rect 8746 4442 8780 4458
rect 8842 4834 8876 4850
rect 8842 4442 8876 4458
rect 8938 4834 8972 4850
rect 8938 4442 8972 4458
rect 9034 4834 9068 4850
rect 9034 4442 9068 4458
rect 9130 4834 9164 4850
rect 9130 4442 9164 4458
rect 9226 4834 9260 4850
rect 9226 4442 9260 4458
rect 9322 4834 9356 4850
rect 9322 4442 9356 4458
rect 9418 4834 9452 4850
rect 9418 4442 9452 4458
rect 9514 4834 9548 4850
rect 9514 4442 9548 4458
rect 9610 4834 9644 4850
rect 9610 4442 9644 4458
rect 9706 4834 9740 4850
rect 9706 4442 9740 4458
rect 9802 4834 9836 4850
rect 9802 4442 9836 4458
rect 9898 4834 9932 4850
rect 9898 4442 9932 4458
rect 9994 4834 10028 4850
rect 9994 4442 10028 4458
rect 10090 4834 10124 4850
rect 10090 4442 10124 4458
rect 10186 4834 10220 4850
rect 10186 4442 10220 4458
rect 10282 4834 10316 4850
rect 10282 4442 10316 4458
rect 10378 4834 10412 4850
rect 10378 4442 10412 4458
rect 10474 4834 10508 4850
rect 10474 4442 10508 4458
rect 10570 4834 10604 4850
rect 10570 4442 10604 4458
rect 10666 4834 10700 4850
rect 10666 4442 10700 4458
rect 10762 4834 10796 4850
rect 10762 4442 10796 4458
rect 10858 4834 10892 4850
rect 10858 4442 10892 4458
rect 10954 4834 10988 4850
rect 10954 4442 10988 4458
rect 8106 4374 8122 4408
rect 8156 4374 8172 4408
rect 8298 4374 8314 4408
rect 8348 4374 8364 4408
rect 8490 4374 8506 4408
rect 8540 4374 8556 4408
rect 8682 4374 8698 4408
rect 8732 4374 8748 4408
rect 8874 4374 8890 4408
rect 8924 4374 8940 4408
rect 9066 4374 9082 4408
rect 9116 4374 9132 4408
rect 9258 4374 9274 4408
rect 9308 4374 9324 4408
rect 9450 4374 9466 4408
rect 9500 4374 9516 4408
rect 9642 4374 9658 4408
rect 9692 4374 9708 4408
rect 9834 4374 9850 4408
rect 9884 4374 9900 4408
rect 10026 4374 10042 4408
rect 10076 4374 10092 4408
rect 10218 4374 10234 4408
rect 10268 4374 10284 4408
rect 10410 4374 10426 4408
rect 10460 4374 10476 4408
rect 10602 4374 10618 4408
rect 10652 4374 10668 4408
rect 10794 4374 10810 4408
rect 10844 4374 10860 4408
rect 8106 4266 8122 4300
rect 8156 4266 8172 4300
rect 8298 4266 8314 4300
rect 8348 4266 8364 4300
rect 8490 4266 8506 4300
rect 8540 4266 8556 4300
rect 8682 4266 8698 4300
rect 8732 4266 8748 4300
rect 8874 4266 8890 4300
rect 8924 4266 8940 4300
rect 9066 4266 9082 4300
rect 9116 4266 9132 4300
rect 9258 4266 9274 4300
rect 9308 4266 9324 4300
rect 9450 4266 9466 4300
rect 9500 4266 9516 4300
rect 9642 4266 9658 4300
rect 9692 4266 9708 4300
rect 9834 4266 9850 4300
rect 9884 4266 9900 4300
rect 10026 4266 10042 4300
rect 10076 4266 10092 4300
rect 10218 4266 10234 4300
rect 10268 4266 10284 4300
rect 10410 4266 10426 4300
rect 10460 4266 10476 4300
rect 10602 4266 10618 4300
rect 10652 4266 10668 4300
rect 10794 4266 10810 4300
rect 10844 4266 10860 4300
rect 8074 4216 8108 4232
rect 8074 3824 8108 3840
rect 8170 4216 8204 4232
rect 8170 3824 8204 3840
rect 8266 4216 8300 4232
rect 8266 3824 8300 3840
rect 8362 4216 8396 4232
rect 8362 3824 8396 3840
rect 8458 4216 8492 4232
rect 8458 3824 8492 3840
rect 8554 4216 8588 4232
rect 8554 3824 8588 3840
rect 8650 4216 8684 4232
rect 8650 3824 8684 3840
rect 8746 4216 8780 4232
rect 8746 3824 8780 3840
rect 8842 4216 8876 4232
rect 8842 3824 8876 3840
rect 8938 4216 8972 4232
rect 8938 3824 8972 3840
rect 9034 4216 9068 4232
rect 9034 3824 9068 3840
rect 9130 4216 9164 4232
rect 9130 3824 9164 3840
rect 9226 4216 9260 4232
rect 9226 3824 9260 3840
rect 9322 4216 9356 4232
rect 9322 3824 9356 3840
rect 9418 4216 9452 4232
rect 9418 3824 9452 3840
rect 9514 4216 9548 4232
rect 9514 3824 9548 3840
rect 9610 4216 9644 4232
rect 9610 3824 9644 3840
rect 9706 4216 9740 4232
rect 9706 3824 9740 3840
rect 9802 4216 9836 4232
rect 9802 3824 9836 3840
rect 9898 4216 9932 4232
rect 9898 3824 9932 3840
rect 9994 4216 10028 4232
rect 9994 3824 10028 3840
rect 10090 4216 10124 4232
rect 10090 3824 10124 3840
rect 10186 4216 10220 4232
rect 10186 3824 10220 3840
rect 10282 4216 10316 4232
rect 10282 3824 10316 3840
rect 10378 4216 10412 4232
rect 10378 3824 10412 3840
rect 10474 4216 10508 4232
rect 10474 3824 10508 3840
rect 10570 4216 10604 4232
rect 10570 3824 10604 3840
rect 10666 4216 10700 4232
rect 10666 3824 10700 3840
rect 10762 4216 10796 4232
rect 10762 3824 10796 3840
rect 10858 4216 10892 4232
rect 10858 3824 10892 3840
rect 10954 4216 10988 4232
rect 10954 3824 10988 3840
rect 8202 3756 8218 3790
rect 8252 3756 8268 3790
rect 8394 3756 8410 3790
rect 8444 3756 8460 3790
rect 8586 3756 8602 3790
rect 8636 3756 8652 3790
rect 8778 3756 8794 3790
rect 8828 3756 8844 3790
rect 8970 3756 8986 3790
rect 9020 3756 9036 3790
rect 9162 3756 9178 3790
rect 9212 3756 9228 3790
rect 9354 3756 9370 3790
rect 9404 3756 9420 3790
rect 9546 3756 9562 3790
rect 9596 3756 9612 3790
rect 9738 3756 9754 3790
rect 9788 3756 9804 3790
rect 9930 3756 9946 3790
rect 9980 3756 9996 3790
rect 10122 3756 10138 3790
rect 10172 3756 10188 3790
rect 10314 3756 10330 3790
rect 10364 3756 10380 3790
rect 10506 3756 10522 3790
rect 10556 3756 10572 3790
rect 10698 3756 10714 3790
rect 10748 3756 10764 3790
rect 10890 3756 10906 3790
rect 10940 3756 10956 3790
rect 8202 3648 8218 3682
rect 8252 3648 8268 3682
rect 8394 3648 8410 3682
rect 8444 3648 8460 3682
rect 8586 3648 8602 3682
rect 8636 3648 8652 3682
rect 8778 3648 8794 3682
rect 8828 3648 8844 3682
rect 8970 3648 8986 3682
rect 9020 3648 9036 3682
rect 9162 3648 9178 3682
rect 9212 3648 9228 3682
rect 9354 3648 9370 3682
rect 9404 3648 9420 3682
rect 9546 3648 9562 3682
rect 9596 3648 9612 3682
rect 9738 3648 9754 3682
rect 9788 3648 9804 3682
rect 9930 3648 9946 3682
rect 9980 3648 9996 3682
rect 10122 3648 10138 3682
rect 10172 3648 10188 3682
rect 10314 3648 10330 3682
rect 10364 3648 10380 3682
rect 10506 3648 10522 3682
rect 10556 3648 10572 3682
rect 10698 3648 10714 3682
rect 10748 3648 10764 3682
rect 10890 3648 10906 3682
rect 10940 3648 10956 3682
rect 8074 3598 8108 3614
rect 8074 3206 8108 3222
rect 8170 3598 8204 3614
rect 8170 3206 8204 3222
rect 8266 3598 8300 3614
rect 8266 3206 8300 3222
rect 8362 3598 8396 3614
rect 8362 3206 8396 3222
rect 8458 3598 8492 3614
rect 8458 3206 8492 3222
rect 8554 3598 8588 3614
rect 8554 3206 8588 3222
rect 8650 3598 8684 3614
rect 8650 3206 8684 3222
rect 8746 3598 8780 3614
rect 8746 3206 8780 3222
rect 8842 3598 8876 3614
rect 8842 3206 8876 3222
rect 8938 3598 8972 3614
rect 8938 3206 8972 3222
rect 9034 3598 9068 3614
rect 9034 3206 9068 3222
rect 9130 3598 9164 3614
rect 9130 3206 9164 3222
rect 9226 3598 9260 3614
rect 9226 3206 9260 3222
rect 9322 3598 9356 3614
rect 9322 3206 9356 3222
rect 9418 3598 9452 3614
rect 9418 3206 9452 3222
rect 9514 3598 9548 3614
rect 9514 3206 9548 3222
rect 9610 3598 9644 3614
rect 9610 3206 9644 3222
rect 9706 3598 9740 3614
rect 9706 3206 9740 3222
rect 9802 3598 9836 3614
rect 9802 3206 9836 3222
rect 9898 3598 9932 3614
rect 9898 3206 9932 3222
rect 9994 3598 10028 3614
rect 9994 3206 10028 3222
rect 10090 3598 10124 3614
rect 10090 3206 10124 3222
rect 10186 3598 10220 3614
rect 10186 3206 10220 3222
rect 10282 3598 10316 3614
rect 10282 3206 10316 3222
rect 10378 3598 10412 3614
rect 10378 3206 10412 3222
rect 10474 3598 10508 3614
rect 10474 3206 10508 3222
rect 10570 3598 10604 3614
rect 10570 3206 10604 3222
rect 10666 3598 10700 3614
rect 10666 3206 10700 3222
rect 10762 3598 10796 3614
rect 10762 3206 10796 3222
rect 10858 3598 10892 3614
rect 10858 3206 10892 3222
rect 10954 3598 10988 3614
rect 10954 3206 10988 3222
rect 8106 3138 8122 3172
rect 8156 3138 8172 3172
rect 8298 3138 8314 3172
rect 8348 3138 8364 3172
rect 8490 3138 8506 3172
rect 8540 3138 8556 3172
rect 8682 3138 8698 3172
rect 8732 3138 8748 3172
rect 8874 3138 8890 3172
rect 8924 3138 8940 3172
rect 9066 3138 9082 3172
rect 9116 3138 9132 3172
rect 9258 3138 9274 3172
rect 9308 3138 9324 3172
rect 9450 3138 9466 3172
rect 9500 3138 9516 3172
rect 9642 3138 9658 3172
rect 9692 3138 9708 3172
rect 9834 3138 9850 3172
rect 9884 3138 9900 3172
rect 10026 3138 10042 3172
rect 10076 3138 10092 3172
rect 10218 3138 10234 3172
rect 10268 3138 10284 3172
rect 10410 3138 10426 3172
rect 10460 3138 10476 3172
rect 10602 3138 10618 3172
rect 10652 3138 10668 3172
rect 10794 3138 10810 3172
rect 10844 3138 10860 3172
rect 7960 3070 7994 3132
rect 11068 3070 11102 3132
rect 7960 3060 8056 3070
rect 7366 3036 8056 3060
rect 11006 3060 11102 3070
rect 11940 5604 12036 5638
rect 14986 5604 15082 5638
rect 11940 5542 11974 5604
rect 15048 5542 15082 5604
rect 12086 5502 12102 5536
rect 12136 5502 12152 5536
rect 12278 5502 12294 5536
rect 12328 5502 12344 5536
rect 12470 5502 12486 5536
rect 12520 5502 12536 5536
rect 12662 5502 12678 5536
rect 12712 5502 12728 5536
rect 12854 5502 12870 5536
rect 12904 5502 12920 5536
rect 13046 5502 13062 5536
rect 13096 5502 13112 5536
rect 13238 5502 13254 5536
rect 13288 5502 13304 5536
rect 13430 5502 13446 5536
rect 13480 5502 13496 5536
rect 13622 5502 13638 5536
rect 13672 5502 13688 5536
rect 13814 5502 13830 5536
rect 13864 5502 13880 5536
rect 14006 5502 14022 5536
rect 14056 5502 14072 5536
rect 14198 5502 14214 5536
rect 14248 5502 14264 5536
rect 14390 5502 14406 5536
rect 14440 5502 14456 5536
rect 14582 5502 14598 5536
rect 14632 5502 14648 5536
rect 14774 5502 14790 5536
rect 14824 5502 14840 5536
rect 12054 5452 12088 5468
rect 12054 5060 12088 5076
rect 12150 5452 12184 5468
rect 12150 5060 12184 5076
rect 12246 5452 12280 5468
rect 12246 5060 12280 5076
rect 12342 5452 12376 5468
rect 12342 5060 12376 5076
rect 12438 5452 12472 5468
rect 12438 5060 12472 5076
rect 12534 5452 12568 5468
rect 12534 5060 12568 5076
rect 12630 5452 12664 5468
rect 12630 5060 12664 5076
rect 12726 5452 12760 5468
rect 12726 5060 12760 5076
rect 12822 5452 12856 5468
rect 12822 5060 12856 5076
rect 12918 5452 12952 5468
rect 12918 5060 12952 5076
rect 13014 5452 13048 5468
rect 13014 5060 13048 5076
rect 13110 5452 13144 5468
rect 13110 5060 13144 5076
rect 13206 5452 13240 5468
rect 13206 5060 13240 5076
rect 13302 5452 13336 5468
rect 13302 5060 13336 5076
rect 13398 5452 13432 5468
rect 13398 5060 13432 5076
rect 13494 5452 13528 5468
rect 13494 5060 13528 5076
rect 13590 5452 13624 5468
rect 13590 5060 13624 5076
rect 13686 5452 13720 5468
rect 13686 5060 13720 5076
rect 13782 5452 13816 5468
rect 13782 5060 13816 5076
rect 13878 5452 13912 5468
rect 13878 5060 13912 5076
rect 13974 5452 14008 5468
rect 13974 5060 14008 5076
rect 14070 5452 14104 5468
rect 14070 5060 14104 5076
rect 14166 5452 14200 5468
rect 14166 5060 14200 5076
rect 14262 5452 14296 5468
rect 14262 5060 14296 5076
rect 14358 5452 14392 5468
rect 14358 5060 14392 5076
rect 14454 5452 14488 5468
rect 14454 5060 14488 5076
rect 14550 5452 14584 5468
rect 14550 5060 14584 5076
rect 14646 5452 14680 5468
rect 14646 5060 14680 5076
rect 14742 5452 14776 5468
rect 14742 5060 14776 5076
rect 14838 5452 14872 5468
rect 14838 5060 14872 5076
rect 14934 5452 14968 5468
rect 14934 5060 14968 5076
rect 12182 4992 12198 5026
rect 12232 4992 12248 5026
rect 12374 4992 12390 5026
rect 12424 4992 12440 5026
rect 12566 4992 12582 5026
rect 12616 4992 12632 5026
rect 12758 4992 12774 5026
rect 12808 4992 12824 5026
rect 12950 4992 12966 5026
rect 13000 4992 13016 5026
rect 13142 4992 13158 5026
rect 13192 4992 13208 5026
rect 13334 4992 13350 5026
rect 13384 4992 13400 5026
rect 13526 4992 13542 5026
rect 13576 4992 13592 5026
rect 13718 4992 13734 5026
rect 13768 4992 13784 5026
rect 13910 4992 13926 5026
rect 13960 4992 13976 5026
rect 14102 4992 14118 5026
rect 14152 4992 14168 5026
rect 14294 4992 14310 5026
rect 14344 4992 14360 5026
rect 14486 4992 14502 5026
rect 14536 4992 14552 5026
rect 14678 4992 14694 5026
rect 14728 4992 14744 5026
rect 14870 4992 14886 5026
rect 14920 4992 14936 5026
rect 12182 4884 12198 4918
rect 12232 4884 12248 4918
rect 12374 4884 12390 4918
rect 12424 4884 12440 4918
rect 12566 4884 12582 4918
rect 12616 4884 12632 4918
rect 12758 4884 12774 4918
rect 12808 4884 12824 4918
rect 12950 4884 12966 4918
rect 13000 4884 13016 4918
rect 13142 4884 13158 4918
rect 13192 4884 13208 4918
rect 13334 4884 13350 4918
rect 13384 4884 13400 4918
rect 13526 4884 13542 4918
rect 13576 4884 13592 4918
rect 13718 4884 13734 4918
rect 13768 4884 13784 4918
rect 13910 4884 13926 4918
rect 13960 4884 13976 4918
rect 14102 4884 14118 4918
rect 14152 4884 14168 4918
rect 14294 4884 14310 4918
rect 14344 4884 14360 4918
rect 14486 4884 14502 4918
rect 14536 4884 14552 4918
rect 14678 4884 14694 4918
rect 14728 4884 14744 4918
rect 14870 4884 14886 4918
rect 14920 4884 14936 4918
rect 12054 4834 12088 4850
rect 12054 4442 12088 4458
rect 12150 4834 12184 4850
rect 12150 4442 12184 4458
rect 12246 4834 12280 4850
rect 12246 4442 12280 4458
rect 12342 4834 12376 4850
rect 12342 4442 12376 4458
rect 12438 4834 12472 4850
rect 12438 4442 12472 4458
rect 12534 4834 12568 4850
rect 12534 4442 12568 4458
rect 12630 4834 12664 4850
rect 12630 4442 12664 4458
rect 12726 4834 12760 4850
rect 12726 4442 12760 4458
rect 12822 4834 12856 4850
rect 12822 4442 12856 4458
rect 12918 4834 12952 4850
rect 12918 4442 12952 4458
rect 13014 4834 13048 4850
rect 13014 4442 13048 4458
rect 13110 4834 13144 4850
rect 13110 4442 13144 4458
rect 13206 4834 13240 4850
rect 13206 4442 13240 4458
rect 13302 4834 13336 4850
rect 13302 4442 13336 4458
rect 13398 4834 13432 4850
rect 13398 4442 13432 4458
rect 13494 4834 13528 4850
rect 13494 4442 13528 4458
rect 13590 4834 13624 4850
rect 13590 4442 13624 4458
rect 13686 4834 13720 4850
rect 13686 4442 13720 4458
rect 13782 4834 13816 4850
rect 13782 4442 13816 4458
rect 13878 4834 13912 4850
rect 13878 4442 13912 4458
rect 13974 4834 14008 4850
rect 13974 4442 14008 4458
rect 14070 4834 14104 4850
rect 14070 4442 14104 4458
rect 14166 4834 14200 4850
rect 14166 4442 14200 4458
rect 14262 4834 14296 4850
rect 14262 4442 14296 4458
rect 14358 4834 14392 4850
rect 14358 4442 14392 4458
rect 14454 4834 14488 4850
rect 14454 4442 14488 4458
rect 14550 4834 14584 4850
rect 14550 4442 14584 4458
rect 14646 4834 14680 4850
rect 14646 4442 14680 4458
rect 14742 4834 14776 4850
rect 14742 4442 14776 4458
rect 14838 4834 14872 4850
rect 14838 4442 14872 4458
rect 14934 4834 14968 4850
rect 14934 4442 14968 4458
rect 12086 4374 12102 4408
rect 12136 4374 12152 4408
rect 12278 4374 12294 4408
rect 12328 4374 12344 4408
rect 12470 4374 12486 4408
rect 12520 4374 12536 4408
rect 12662 4374 12678 4408
rect 12712 4374 12728 4408
rect 12854 4374 12870 4408
rect 12904 4374 12920 4408
rect 13046 4374 13062 4408
rect 13096 4374 13112 4408
rect 13238 4374 13254 4408
rect 13288 4374 13304 4408
rect 13430 4374 13446 4408
rect 13480 4374 13496 4408
rect 13622 4374 13638 4408
rect 13672 4374 13688 4408
rect 13814 4374 13830 4408
rect 13864 4374 13880 4408
rect 14006 4374 14022 4408
rect 14056 4374 14072 4408
rect 14198 4374 14214 4408
rect 14248 4374 14264 4408
rect 14390 4374 14406 4408
rect 14440 4374 14456 4408
rect 14582 4374 14598 4408
rect 14632 4374 14648 4408
rect 14774 4374 14790 4408
rect 14824 4374 14840 4408
rect 12086 4266 12102 4300
rect 12136 4266 12152 4300
rect 12278 4266 12294 4300
rect 12328 4266 12344 4300
rect 12470 4266 12486 4300
rect 12520 4266 12536 4300
rect 12662 4266 12678 4300
rect 12712 4266 12728 4300
rect 12854 4266 12870 4300
rect 12904 4266 12920 4300
rect 13046 4266 13062 4300
rect 13096 4266 13112 4300
rect 13238 4266 13254 4300
rect 13288 4266 13304 4300
rect 13430 4266 13446 4300
rect 13480 4266 13496 4300
rect 13622 4266 13638 4300
rect 13672 4266 13688 4300
rect 13814 4266 13830 4300
rect 13864 4266 13880 4300
rect 14006 4266 14022 4300
rect 14056 4266 14072 4300
rect 14198 4266 14214 4300
rect 14248 4266 14264 4300
rect 14390 4266 14406 4300
rect 14440 4266 14456 4300
rect 14582 4266 14598 4300
rect 14632 4266 14648 4300
rect 14774 4266 14790 4300
rect 14824 4266 14840 4300
rect 12054 4216 12088 4232
rect 12054 3824 12088 3840
rect 12150 4216 12184 4232
rect 12150 3824 12184 3840
rect 12246 4216 12280 4232
rect 12246 3824 12280 3840
rect 12342 4216 12376 4232
rect 12342 3824 12376 3840
rect 12438 4216 12472 4232
rect 12438 3824 12472 3840
rect 12534 4216 12568 4232
rect 12534 3824 12568 3840
rect 12630 4216 12664 4232
rect 12630 3824 12664 3840
rect 12726 4216 12760 4232
rect 12726 3824 12760 3840
rect 12822 4216 12856 4232
rect 12822 3824 12856 3840
rect 12918 4216 12952 4232
rect 12918 3824 12952 3840
rect 13014 4216 13048 4232
rect 13014 3824 13048 3840
rect 13110 4216 13144 4232
rect 13110 3824 13144 3840
rect 13206 4216 13240 4232
rect 13206 3824 13240 3840
rect 13302 4216 13336 4232
rect 13302 3824 13336 3840
rect 13398 4216 13432 4232
rect 13398 3824 13432 3840
rect 13494 4216 13528 4232
rect 13494 3824 13528 3840
rect 13590 4216 13624 4232
rect 13590 3824 13624 3840
rect 13686 4216 13720 4232
rect 13686 3824 13720 3840
rect 13782 4216 13816 4232
rect 13782 3824 13816 3840
rect 13878 4216 13912 4232
rect 13878 3824 13912 3840
rect 13974 4216 14008 4232
rect 13974 3824 14008 3840
rect 14070 4216 14104 4232
rect 14070 3824 14104 3840
rect 14166 4216 14200 4232
rect 14166 3824 14200 3840
rect 14262 4216 14296 4232
rect 14262 3824 14296 3840
rect 14358 4216 14392 4232
rect 14358 3824 14392 3840
rect 14454 4216 14488 4232
rect 14454 3824 14488 3840
rect 14550 4216 14584 4232
rect 14550 3824 14584 3840
rect 14646 4216 14680 4232
rect 14646 3824 14680 3840
rect 14742 4216 14776 4232
rect 14742 3824 14776 3840
rect 14838 4216 14872 4232
rect 14838 3824 14872 3840
rect 14934 4216 14968 4232
rect 14934 3824 14968 3840
rect 12182 3756 12198 3790
rect 12232 3756 12248 3790
rect 12374 3756 12390 3790
rect 12424 3756 12440 3790
rect 12566 3756 12582 3790
rect 12616 3756 12632 3790
rect 12758 3756 12774 3790
rect 12808 3756 12824 3790
rect 12950 3756 12966 3790
rect 13000 3756 13016 3790
rect 13142 3756 13158 3790
rect 13192 3756 13208 3790
rect 13334 3756 13350 3790
rect 13384 3756 13400 3790
rect 13526 3756 13542 3790
rect 13576 3756 13592 3790
rect 13718 3756 13734 3790
rect 13768 3756 13784 3790
rect 13910 3756 13926 3790
rect 13960 3756 13976 3790
rect 14102 3756 14118 3790
rect 14152 3756 14168 3790
rect 14294 3756 14310 3790
rect 14344 3756 14360 3790
rect 14486 3756 14502 3790
rect 14536 3756 14552 3790
rect 14678 3756 14694 3790
rect 14728 3756 14744 3790
rect 14870 3756 14886 3790
rect 14920 3756 14936 3790
rect 12182 3648 12198 3682
rect 12232 3648 12248 3682
rect 12374 3648 12390 3682
rect 12424 3648 12440 3682
rect 12566 3648 12582 3682
rect 12616 3648 12632 3682
rect 12758 3648 12774 3682
rect 12808 3648 12824 3682
rect 12950 3648 12966 3682
rect 13000 3648 13016 3682
rect 13142 3648 13158 3682
rect 13192 3648 13208 3682
rect 13334 3648 13350 3682
rect 13384 3648 13400 3682
rect 13526 3648 13542 3682
rect 13576 3648 13592 3682
rect 13718 3648 13734 3682
rect 13768 3648 13784 3682
rect 13910 3648 13926 3682
rect 13960 3648 13976 3682
rect 14102 3648 14118 3682
rect 14152 3648 14168 3682
rect 14294 3648 14310 3682
rect 14344 3648 14360 3682
rect 14486 3648 14502 3682
rect 14536 3648 14552 3682
rect 14678 3648 14694 3682
rect 14728 3648 14744 3682
rect 14870 3648 14886 3682
rect 14920 3648 14936 3682
rect 12054 3598 12088 3614
rect 12054 3206 12088 3222
rect 12150 3598 12184 3614
rect 12150 3206 12184 3222
rect 12246 3598 12280 3614
rect 12246 3206 12280 3222
rect 12342 3598 12376 3614
rect 12342 3206 12376 3222
rect 12438 3598 12472 3614
rect 12438 3206 12472 3222
rect 12534 3598 12568 3614
rect 12534 3206 12568 3222
rect 12630 3598 12664 3614
rect 12630 3206 12664 3222
rect 12726 3598 12760 3614
rect 12726 3206 12760 3222
rect 12822 3598 12856 3614
rect 12822 3206 12856 3222
rect 12918 3598 12952 3614
rect 12918 3206 12952 3222
rect 13014 3598 13048 3614
rect 13014 3206 13048 3222
rect 13110 3598 13144 3614
rect 13110 3206 13144 3222
rect 13206 3598 13240 3614
rect 13206 3206 13240 3222
rect 13302 3598 13336 3614
rect 13302 3206 13336 3222
rect 13398 3598 13432 3614
rect 13398 3206 13432 3222
rect 13494 3598 13528 3614
rect 13494 3206 13528 3222
rect 13590 3598 13624 3614
rect 13590 3206 13624 3222
rect 13686 3598 13720 3614
rect 13686 3206 13720 3222
rect 13782 3598 13816 3614
rect 13782 3206 13816 3222
rect 13878 3598 13912 3614
rect 13878 3206 13912 3222
rect 13974 3598 14008 3614
rect 13974 3206 14008 3222
rect 14070 3598 14104 3614
rect 14070 3206 14104 3222
rect 14166 3598 14200 3614
rect 14166 3206 14200 3222
rect 14262 3598 14296 3614
rect 14262 3206 14296 3222
rect 14358 3598 14392 3614
rect 14358 3206 14392 3222
rect 14454 3598 14488 3614
rect 14454 3206 14488 3222
rect 14550 3598 14584 3614
rect 14550 3206 14584 3222
rect 14646 3598 14680 3614
rect 14646 3206 14680 3222
rect 14742 3598 14776 3614
rect 14742 3206 14776 3222
rect 14838 3598 14872 3614
rect 14838 3206 14872 3222
rect 14934 3598 14968 3614
rect 14934 3206 14968 3222
rect 12086 3138 12102 3172
rect 12136 3138 12152 3172
rect 12278 3138 12294 3172
rect 12328 3138 12344 3172
rect 12470 3138 12486 3172
rect 12520 3138 12536 3172
rect 12662 3138 12678 3172
rect 12712 3138 12728 3172
rect 12854 3138 12870 3172
rect 12904 3138 12920 3172
rect 13046 3138 13062 3172
rect 13096 3138 13112 3172
rect 13238 3138 13254 3172
rect 13288 3138 13304 3172
rect 13430 3138 13446 3172
rect 13480 3138 13496 3172
rect 13622 3138 13638 3172
rect 13672 3138 13688 3172
rect 13814 3138 13830 3172
rect 13864 3138 13880 3172
rect 14006 3138 14022 3172
rect 14056 3138 14072 3172
rect 14198 3138 14214 3172
rect 14248 3138 14264 3172
rect 14390 3138 14406 3172
rect 14440 3138 14456 3172
rect 14582 3138 14598 3172
rect 14632 3138 14648 3172
rect 14774 3138 14790 3172
rect 14824 3138 14840 3172
rect 11940 3070 11974 3132
rect 15048 3070 15082 3132
rect 11006 3036 11104 3060
rect 11940 3036 12036 3070
rect 14986 3060 15082 3070
rect 15580 5604 15676 5638
rect 18626 5604 18722 5638
rect 15580 5542 15614 5604
rect 18688 5542 18722 5604
rect 15726 5502 15742 5536
rect 15776 5502 15792 5536
rect 15918 5502 15934 5536
rect 15968 5502 15984 5536
rect 16110 5502 16126 5536
rect 16160 5502 16176 5536
rect 16302 5502 16318 5536
rect 16352 5502 16368 5536
rect 16494 5502 16510 5536
rect 16544 5502 16560 5536
rect 16686 5502 16702 5536
rect 16736 5502 16752 5536
rect 16878 5502 16894 5536
rect 16928 5502 16944 5536
rect 17070 5502 17086 5536
rect 17120 5502 17136 5536
rect 17262 5502 17278 5536
rect 17312 5502 17328 5536
rect 17454 5502 17470 5536
rect 17504 5502 17520 5536
rect 17646 5502 17662 5536
rect 17696 5502 17712 5536
rect 17838 5502 17854 5536
rect 17888 5502 17904 5536
rect 18030 5502 18046 5536
rect 18080 5502 18096 5536
rect 18222 5502 18238 5536
rect 18272 5502 18288 5536
rect 18414 5502 18430 5536
rect 18464 5502 18480 5536
rect 15694 5452 15728 5468
rect 15694 5060 15728 5076
rect 15790 5452 15824 5468
rect 15790 5060 15824 5076
rect 15886 5452 15920 5468
rect 15886 5060 15920 5076
rect 15982 5452 16016 5468
rect 15982 5060 16016 5076
rect 16078 5452 16112 5468
rect 16078 5060 16112 5076
rect 16174 5452 16208 5468
rect 16174 5060 16208 5076
rect 16270 5452 16304 5468
rect 16270 5060 16304 5076
rect 16366 5452 16400 5468
rect 16366 5060 16400 5076
rect 16462 5452 16496 5468
rect 16462 5060 16496 5076
rect 16558 5452 16592 5468
rect 16558 5060 16592 5076
rect 16654 5452 16688 5468
rect 16654 5060 16688 5076
rect 16750 5452 16784 5468
rect 16750 5060 16784 5076
rect 16846 5452 16880 5468
rect 16846 5060 16880 5076
rect 16942 5452 16976 5468
rect 16942 5060 16976 5076
rect 17038 5452 17072 5468
rect 17038 5060 17072 5076
rect 17134 5452 17168 5468
rect 17134 5060 17168 5076
rect 17230 5452 17264 5468
rect 17230 5060 17264 5076
rect 17326 5452 17360 5468
rect 17326 5060 17360 5076
rect 17422 5452 17456 5468
rect 17422 5060 17456 5076
rect 17518 5452 17552 5468
rect 17518 5060 17552 5076
rect 17614 5452 17648 5468
rect 17614 5060 17648 5076
rect 17710 5452 17744 5468
rect 17710 5060 17744 5076
rect 17806 5452 17840 5468
rect 17806 5060 17840 5076
rect 17902 5452 17936 5468
rect 17902 5060 17936 5076
rect 17998 5452 18032 5468
rect 17998 5060 18032 5076
rect 18094 5452 18128 5468
rect 18094 5060 18128 5076
rect 18190 5452 18224 5468
rect 18190 5060 18224 5076
rect 18286 5452 18320 5468
rect 18286 5060 18320 5076
rect 18382 5452 18416 5468
rect 18382 5060 18416 5076
rect 18478 5452 18512 5468
rect 18478 5060 18512 5076
rect 18574 5452 18608 5468
rect 18574 5060 18608 5076
rect 15822 4992 15838 5026
rect 15872 4992 15888 5026
rect 16014 4992 16030 5026
rect 16064 4992 16080 5026
rect 16206 4992 16222 5026
rect 16256 4992 16272 5026
rect 16398 4992 16414 5026
rect 16448 4992 16464 5026
rect 16590 4992 16606 5026
rect 16640 4992 16656 5026
rect 16782 4992 16798 5026
rect 16832 4992 16848 5026
rect 16974 4992 16990 5026
rect 17024 4992 17040 5026
rect 17166 4992 17182 5026
rect 17216 4992 17232 5026
rect 17358 4992 17374 5026
rect 17408 4992 17424 5026
rect 17550 4992 17566 5026
rect 17600 4992 17616 5026
rect 17742 4992 17758 5026
rect 17792 4992 17808 5026
rect 17934 4992 17950 5026
rect 17984 4992 18000 5026
rect 18126 4992 18142 5026
rect 18176 4992 18192 5026
rect 18318 4992 18334 5026
rect 18368 4992 18384 5026
rect 18510 4992 18526 5026
rect 18560 4992 18576 5026
rect 15822 4884 15838 4918
rect 15872 4884 15888 4918
rect 16014 4884 16030 4918
rect 16064 4884 16080 4918
rect 16206 4884 16222 4918
rect 16256 4884 16272 4918
rect 16398 4884 16414 4918
rect 16448 4884 16464 4918
rect 16590 4884 16606 4918
rect 16640 4884 16656 4918
rect 16782 4884 16798 4918
rect 16832 4884 16848 4918
rect 16974 4884 16990 4918
rect 17024 4884 17040 4918
rect 17166 4884 17182 4918
rect 17216 4884 17232 4918
rect 17358 4884 17374 4918
rect 17408 4884 17424 4918
rect 17550 4884 17566 4918
rect 17600 4884 17616 4918
rect 17742 4884 17758 4918
rect 17792 4884 17808 4918
rect 17934 4884 17950 4918
rect 17984 4884 18000 4918
rect 18126 4884 18142 4918
rect 18176 4884 18192 4918
rect 18318 4884 18334 4918
rect 18368 4884 18384 4918
rect 18510 4884 18526 4918
rect 18560 4884 18576 4918
rect 15694 4834 15728 4850
rect 15694 4442 15728 4458
rect 15790 4834 15824 4850
rect 15790 4442 15824 4458
rect 15886 4834 15920 4850
rect 15886 4442 15920 4458
rect 15982 4834 16016 4850
rect 15982 4442 16016 4458
rect 16078 4834 16112 4850
rect 16078 4442 16112 4458
rect 16174 4834 16208 4850
rect 16174 4442 16208 4458
rect 16270 4834 16304 4850
rect 16270 4442 16304 4458
rect 16366 4834 16400 4850
rect 16366 4442 16400 4458
rect 16462 4834 16496 4850
rect 16462 4442 16496 4458
rect 16558 4834 16592 4850
rect 16558 4442 16592 4458
rect 16654 4834 16688 4850
rect 16654 4442 16688 4458
rect 16750 4834 16784 4850
rect 16750 4442 16784 4458
rect 16846 4834 16880 4850
rect 16846 4442 16880 4458
rect 16942 4834 16976 4850
rect 16942 4442 16976 4458
rect 17038 4834 17072 4850
rect 17038 4442 17072 4458
rect 17134 4834 17168 4850
rect 17134 4442 17168 4458
rect 17230 4834 17264 4850
rect 17230 4442 17264 4458
rect 17326 4834 17360 4850
rect 17326 4442 17360 4458
rect 17422 4834 17456 4850
rect 17422 4442 17456 4458
rect 17518 4834 17552 4850
rect 17518 4442 17552 4458
rect 17614 4834 17648 4850
rect 17614 4442 17648 4458
rect 17710 4834 17744 4850
rect 17710 4442 17744 4458
rect 17806 4834 17840 4850
rect 17806 4442 17840 4458
rect 17902 4834 17936 4850
rect 17902 4442 17936 4458
rect 17998 4834 18032 4850
rect 17998 4442 18032 4458
rect 18094 4834 18128 4850
rect 18094 4442 18128 4458
rect 18190 4834 18224 4850
rect 18190 4442 18224 4458
rect 18286 4834 18320 4850
rect 18286 4442 18320 4458
rect 18382 4834 18416 4850
rect 18382 4442 18416 4458
rect 18478 4834 18512 4850
rect 18478 4442 18512 4458
rect 18574 4834 18608 4850
rect 18574 4442 18608 4458
rect 15726 4374 15742 4408
rect 15776 4374 15792 4408
rect 15918 4374 15934 4408
rect 15968 4374 15984 4408
rect 16110 4374 16126 4408
rect 16160 4374 16176 4408
rect 16302 4374 16318 4408
rect 16352 4374 16368 4408
rect 16494 4374 16510 4408
rect 16544 4374 16560 4408
rect 16686 4374 16702 4408
rect 16736 4374 16752 4408
rect 16878 4374 16894 4408
rect 16928 4374 16944 4408
rect 17070 4374 17086 4408
rect 17120 4374 17136 4408
rect 17262 4374 17278 4408
rect 17312 4374 17328 4408
rect 17454 4374 17470 4408
rect 17504 4374 17520 4408
rect 17646 4374 17662 4408
rect 17696 4374 17712 4408
rect 17838 4374 17854 4408
rect 17888 4374 17904 4408
rect 18030 4374 18046 4408
rect 18080 4374 18096 4408
rect 18222 4374 18238 4408
rect 18272 4374 18288 4408
rect 18414 4374 18430 4408
rect 18464 4374 18480 4408
rect 15726 4266 15742 4300
rect 15776 4266 15792 4300
rect 15918 4266 15934 4300
rect 15968 4266 15984 4300
rect 16110 4266 16126 4300
rect 16160 4266 16176 4300
rect 16302 4266 16318 4300
rect 16352 4266 16368 4300
rect 16494 4266 16510 4300
rect 16544 4266 16560 4300
rect 16686 4266 16702 4300
rect 16736 4266 16752 4300
rect 16878 4266 16894 4300
rect 16928 4266 16944 4300
rect 17070 4266 17086 4300
rect 17120 4266 17136 4300
rect 17262 4266 17278 4300
rect 17312 4266 17328 4300
rect 17454 4266 17470 4300
rect 17504 4266 17520 4300
rect 17646 4266 17662 4300
rect 17696 4266 17712 4300
rect 17838 4266 17854 4300
rect 17888 4266 17904 4300
rect 18030 4266 18046 4300
rect 18080 4266 18096 4300
rect 18222 4266 18238 4300
rect 18272 4266 18288 4300
rect 18414 4266 18430 4300
rect 18464 4266 18480 4300
rect 15694 4216 15728 4232
rect 15694 3824 15728 3840
rect 15790 4216 15824 4232
rect 15790 3824 15824 3840
rect 15886 4216 15920 4232
rect 15886 3824 15920 3840
rect 15982 4216 16016 4232
rect 15982 3824 16016 3840
rect 16078 4216 16112 4232
rect 16078 3824 16112 3840
rect 16174 4216 16208 4232
rect 16174 3824 16208 3840
rect 16270 4216 16304 4232
rect 16270 3824 16304 3840
rect 16366 4216 16400 4232
rect 16366 3824 16400 3840
rect 16462 4216 16496 4232
rect 16462 3824 16496 3840
rect 16558 4216 16592 4232
rect 16558 3824 16592 3840
rect 16654 4216 16688 4232
rect 16654 3824 16688 3840
rect 16750 4216 16784 4232
rect 16750 3824 16784 3840
rect 16846 4216 16880 4232
rect 16846 3824 16880 3840
rect 16942 4216 16976 4232
rect 16942 3824 16976 3840
rect 17038 4216 17072 4232
rect 17038 3824 17072 3840
rect 17134 4216 17168 4232
rect 17134 3824 17168 3840
rect 17230 4216 17264 4232
rect 17230 3824 17264 3840
rect 17326 4216 17360 4232
rect 17326 3824 17360 3840
rect 17422 4216 17456 4232
rect 17422 3824 17456 3840
rect 17518 4216 17552 4232
rect 17518 3824 17552 3840
rect 17614 4216 17648 4232
rect 17614 3824 17648 3840
rect 17710 4216 17744 4232
rect 17710 3824 17744 3840
rect 17806 4216 17840 4232
rect 17806 3824 17840 3840
rect 17902 4216 17936 4232
rect 17902 3824 17936 3840
rect 17998 4216 18032 4232
rect 17998 3824 18032 3840
rect 18094 4216 18128 4232
rect 18094 3824 18128 3840
rect 18190 4216 18224 4232
rect 18190 3824 18224 3840
rect 18286 4216 18320 4232
rect 18286 3824 18320 3840
rect 18382 4216 18416 4232
rect 18382 3824 18416 3840
rect 18478 4216 18512 4232
rect 18478 3824 18512 3840
rect 18574 4216 18608 4232
rect 18574 3824 18608 3840
rect 15822 3756 15838 3790
rect 15872 3756 15888 3790
rect 16014 3756 16030 3790
rect 16064 3756 16080 3790
rect 16206 3756 16222 3790
rect 16256 3756 16272 3790
rect 16398 3756 16414 3790
rect 16448 3756 16464 3790
rect 16590 3756 16606 3790
rect 16640 3756 16656 3790
rect 16782 3756 16798 3790
rect 16832 3756 16848 3790
rect 16974 3756 16990 3790
rect 17024 3756 17040 3790
rect 17166 3756 17182 3790
rect 17216 3756 17232 3790
rect 17358 3756 17374 3790
rect 17408 3756 17424 3790
rect 17550 3756 17566 3790
rect 17600 3756 17616 3790
rect 17742 3756 17758 3790
rect 17792 3756 17808 3790
rect 17934 3756 17950 3790
rect 17984 3756 18000 3790
rect 18126 3756 18142 3790
rect 18176 3756 18192 3790
rect 18318 3756 18334 3790
rect 18368 3756 18384 3790
rect 18510 3756 18526 3790
rect 18560 3756 18576 3790
rect 15822 3648 15838 3682
rect 15872 3648 15888 3682
rect 16014 3648 16030 3682
rect 16064 3648 16080 3682
rect 16206 3648 16222 3682
rect 16256 3648 16272 3682
rect 16398 3648 16414 3682
rect 16448 3648 16464 3682
rect 16590 3648 16606 3682
rect 16640 3648 16656 3682
rect 16782 3648 16798 3682
rect 16832 3648 16848 3682
rect 16974 3648 16990 3682
rect 17024 3648 17040 3682
rect 17166 3648 17182 3682
rect 17216 3648 17232 3682
rect 17358 3648 17374 3682
rect 17408 3648 17424 3682
rect 17550 3648 17566 3682
rect 17600 3648 17616 3682
rect 17742 3648 17758 3682
rect 17792 3648 17808 3682
rect 17934 3648 17950 3682
rect 17984 3648 18000 3682
rect 18126 3648 18142 3682
rect 18176 3648 18192 3682
rect 18318 3648 18334 3682
rect 18368 3648 18384 3682
rect 18510 3648 18526 3682
rect 18560 3648 18576 3682
rect 15694 3598 15728 3614
rect 15694 3206 15728 3222
rect 15790 3598 15824 3614
rect 15790 3206 15824 3222
rect 15886 3598 15920 3614
rect 15886 3206 15920 3222
rect 15982 3598 16016 3614
rect 15982 3206 16016 3222
rect 16078 3598 16112 3614
rect 16078 3206 16112 3222
rect 16174 3598 16208 3614
rect 16174 3206 16208 3222
rect 16270 3598 16304 3614
rect 16270 3206 16304 3222
rect 16366 3598 16400 3614
rect 16366 3206 16400 3222
rect 16462 3598 16496 3614
rect 16462 3206 16496 3222
rect 16558 3598 16592 3614
rect 16558 3206 16592 3222
rect 16654 3598 16688 3614
rect 16654 3206 16688 3222
rect 16750 3598 16784 3614
rect 16750 3206 16784 3222
rect 16846 3598 16880 3614
rect 16846 3206 16880 3222
rect 16942 3598 16976 3614
rect 16942 3206 16976 3222
rect 17038 3598 17072 3614
rect 17038 3206 17072 3222
rect 17134 3598 17168 3614
rect 17134 3206 17168 3222
rect 17230 3598 17264 3614
rect 17230 3206 17264 3222
rect 17326 3598 17360 3614
rect 17326 3206 17360 3222
rect 17422 3598 17456 3614
rect 17422 3206 17456 3222
rect 17518 3598 17552 3614
rect 17518 3206 17552 3222
rect 17614 3598 17648 3614
rect 17614 3206 17648 3222
rect 17710 3598 17744 3614
rect 17710 3206 17744 3222
rect 17806 3598 17840 3614
rect 17806 3206 17840 3222
rect 17902 3598 17936 3614
rect 17902 3206 17936 3222
rect 17998 3598 18032 3614
rect 17998 3206 18032 3222
rect 18094 3598 18128 3614
rect 18094 3206 18128 3222
rect 18190 3598 18224 3614
rect 18190 3206 18224 3222
rect 18286 3598 18320 3614
rect 18286 3206 18320 3222
rect 18382 3598 18416 3614
rect 18382 3206 18416 3222
rect 18478 3598 18512 3614
rect 18478 3206 18512 3222
rect 18574 3598 18608 3614
rect 18574 3206 18608 3222
rect 15726 3138 15742 3172
rect 15776 3138 15792 3172
rect 15918 3138 15934 3172
rect 15968 3138 15984 3172
rect 16110 3138 16126 3172
rect 16160 3138 16176 3172
rect 16302 3138 16318 3172
rect 16352 3138 16368 3172
rect 16494 3138 16510 3172
rect 16544 3138 16560 3172
rect 16686 3138 16702 3172
rect 16736 3138 16752 3172
rect 16878 3138 16894 3172
rect 16928 3138 16944 3172
rect 17070 3138 17086 3172
rect 17120 3138 17136 3172
rect 17262 3138 17278 3172
rect 17312 3138 17328 3172
rect 17454 3138 17470 3172
rect 17504 3138 17520 3172
rect 17646 3138 17662 3172
rect 17696 3138 17712 3172
rect 17838 3138 17854 3172
rect 17888 3138 17904 3172
rect 18030 3138 18046 3172
rect 18080 3138 18096 3172
rect 18222 3138 18238 3172
rect 18272 3138 18288 3172
rect 18414 3138 18430 3172
rect 18464 3138 18480 3172
rect 15580 3070 15614 3132
rect 18688 3070 18722 3132
rect 15580 3060 15676 3070
rect 14986 3036 15676 3060
rect 18626 3060 18722 3070
rect 18626 3036 18724 3060
rect -1160 2806 12 3036
rect 1660 2806 2868 3036
rect 4344 2966 11104 3036
rect 11964 2966 18724 3036
rect 4120 2932 4216 2966
rect 4862 2960 5256 2966
rect 4862 2932 4958 2960
rect 4120 2870 4154 2932
rect -1684 2772 -1588 2806
rect -942 2792 -548 2806
rect -942 2772 -846 2792
rect -1684 2710 -1650 2772
rect -880 2710 -846 2772
rect -736 2772 -548 2792
rect 98 2772 194 2806
rect -736 2760 -610 2772
rect -1538 2670 -1522 2704
rect -1488 2670 -1472 2704
rect -1346 2670 -1330 2704
rect -1296 2670 -1280 2704
rect -1154 2670 -1138 2704
rect -1104 2670 -1088 2704
rect -1570 2620 -1536 2636
rect -1570 2228 -1536 2244
rect -1474 2620 -1440 2636
rect -1474 2228 -1440 2244
rect -1378 2620 -1344 2636
rect -1378 2228 -1344 2244
rect -1282 2620 -1248 2636
rect -1282 2228 -1248 2244
rect -1186 2620 -1152 2636
rect -1186 2228 -1152 2244
rect -1090 2620 -1056 2636
rect -1090 2228 -1056 2244
rect -994 2620 -960 2636
rect -994 2228 -960 2244
rect -1442 2160 -1426 2194
rect -1392 2160 -1376 2194
rect -1250 2160 -1234 2194
rect -1200 2160 -1184 2194
rect -1058 2160 -1042 2194
rect -1008 2160 -992 2194
rect -1442 2052 -1426 2086
rect -1392 2052 -1376 2086
rect -1250 2052 -1234 2086
rect -1200 2052 -1184 2086
rect -1058 2052 -1042 2086
rect -1008 2052 -992 2086
rect -1570 2002 -1536 2018
rect -1570 1610 -1536 1626
rect -1474 2002 -1440 2018
rect -1474 1610 -1440 1626
rect -1378 2002 -1344 2018
rect -1378 1610 -1344 1626
rect -1282 2002 -1248 2018
rect -1282 1610 -1248 1626
rect -1186 2002 -1152 2018
rect -1186 1610 -1152 1626
rect -1090 2002 -1056 2018
rect -1090 1610 -1056 1626
rect -994 2002 -960 2018
rect -994 1610 -960 1626
rect -1538 1542 -1522 1576
rect -1488 1542 -1472 1576
rect -1346 1542 -1330 1576
rect -1296 1542 -1280 1576
rect -1154 1542 -1138 1576
rect -1104 1542 -1088 1576
rect -1684 1474 -1650 1536
rect -644 2710 -610 2760
rect -880 1474 -846 1536
rect -1684 1440 -1588 1474
rect -942 1452 -846 1474
rect -736 1536 -644 2008
rect 160 2710 194 2772
rect -498 2670 -482 2704
rect -448 2670 -432 2704
rect -306 2670 -290 2704
rect -256 2670 -240 2704
rect -114 2670 -98 2704
rect -64 2670 -48 2704
rect -530 2620 -496 2636
rect -530 2228 -496 2244
rect -434 2620 -400 2636
rect -434 2228 -400 2244
rect -338 2620 -304 2636
rect -338 2228 -304 2244
rect -242 2620 -208 2636
rect -242 2228 -208 2244
rect -146 2620 -112 2636
rect -146 2228 -112 2244
rect -50 2620 -16 2636
rect -50 2228 -16 2244
rect 46 2620 80 2636
rect 46 2228 80 2244
rect -402 2160 -386 2194
rect -352 2160 -336 2194
rect -210 2160 -194 2194
rect -160 2160 -144 2194
rect -18 2160 -2 2194
rect 32 2160 48 2194
rect -402 2052 -386 2086
rect -352 2052 -336 2086
rect -210 2052 -194 2086
rect -160 2052 -144 2086
rect -18 2052 -2 2086
rect 32 2052 48 2086
rect -530 2002 -496 2018
rect -530 1610 -496 1626
rect -434 2002 -400 2018
rect -434 1610 -400 1626
rect -338 2002 -304 2018
rect -338 1610 -304 1626
rect -242 2002 -208 2018
rect -242 1610 -208 1626
rect -146 2002 -112 2018
rect -146 1610 -112 1626
rect -50 2002 -16 2018
rect -50 1610 -16 1626
rect 46 2002 80 2018
rect 46 1610 80 1626
rect -498 1542 -482 1576
rect -448 1542 -432 1576
rect -306 1542 -290 1576
rect -256 1542 -240 1576
rect -114 1542 -98 1576
rect -64 1542 -48 1576
rect -736 1474 -610 1536
rect 160 1474 194 1536
rect -942 1440 -844 1452
rect -1684 1384 -844 1440
rect -736 1440 -548 1474
rect 98 1452 194 1474
rect 396 2772 492 2806
rect 1138 2772 1234 2806
rect 396 2710 430 2772
rect 1200 2710 1234 2772
rect 542 2670 558 2704
rect 592 2670 608 2704
rect 734 2670 750 2704
rect 784 2670 800 2704
rect 926 2670 942 2704
rect 976 2670 992 2704
rect 510 2620 544 2636
rect 510 2228 544 2244
rect 606 2620 640 2636
rect 606 2228 640 2244
rect 702 2620 736 2636
rect 702 2228 736 2244
rect 798 2620 832 2636
rect 798 2228 832 2244
rect 894 2620 928 2636
rect 894 2228 928 2244
rect 990 2620 1024 2636
rect 990 2228 1024 2244
rect 1086 2620 1120 2636
rect 1086 2228 1120 2244
rect 638 2160 654 2194
rect 688 2160 704 2194
rect 830 2160 846 2194
rect 880 2160 896 2194
rect 1022 2160 1038 2194
rect 1072 2160 1088 2194
rect 638 2052 654 2086
rect 688 2052 704 2086
rect 830 2052 846 2086
rect 880 2052 896 2086
rect 1022 2052 1038 2086
rect 1072 2052 1088 2086
rect 510 2002 544 2018
rect 510 1610 544 1626
rect 606 2002 640 2018
rect 606 1610 640 1626
rect 702 2002 736 2018
rect 702 1610 736 1626
rect 798 2002 832 2018
rect 798 1610 832 1626
rect 894 2002 928 2018
rect 894 1610 928 1626
rect 990 2002 1024 2018
rect 990 1610 1024 1626
rect 1086 2002 1120 2018
rect 1086 1610 1120 1626
rect 542 1542 558 1576
rect 592 1542 608 1576
rect 734 1542 750 1576
rect 784 1542 800 1576
rect 926 1542 942 1576
rect 976 1542 992 1576
rect 396 1474 430 1536
rect 1200 1474 1234 1536
rect 98 1440 196 1452
rect -736 1384 196 1440
rect 396 1440 492 1474
rect 1138 1452 1234 1474
rect 1436 2772 1532 2806
rect 2178 2796 2572 2806
rect 2178 2772 2274 2796
rect 1436 2710 1470 2772
rect 2240 2710 2274 2772
rect 2376 2772 2572 2796
rect 3218 2772 3314 2806
rect 2376 2760 2510 2772
rect 1582 2670 1598 2704
rect 1632 2670 1648 2704
rect 1774 2670 1790 2704
rect 1824 2670 1840 2704
rect 1966 2670 1982 2704
rect 2016 2670 2032 2704
rect 1550 2620 1584 2636
rect 1550 2228 1584 2244
rect 1646 2620 1680 2636
rect 1646 2228 1680 2244
rect 1742 2620 1776 2636
rect 1742 2228 1776 2244
rect 1838 2620 1872 2636
rect 1838 2228 1872 2244
rect 1934 2620 1968 2636
rect 1934 2228 1968 2244
rect 2030 2620 2064 2636
rect 2030 2228 2064 2244
rect 2126 2620 2160 2636
rect 2126 2228 2160 2244
rect 1678 2160 1694 2194
rect 1728 2160 1744 2194
rect 1870 2160 1886 2194
rect 1920 2160 1936 2194
rect 2062 2160 2078 2194
rect 2112 2160 2128 2194
rect 1678 2052 1694 2086
rect 1728 2052 1744 2086
rect 1870 2052 1886 2086
rect 1920 2052 1936 2086
rect 2062 2052 2078 2086
rect 2112 2052 2128 2086
rect 1550 2002 1584 2018
rect 1550 1610 1584 1626
rect 1646 2002 1680 2018
rect 1646 1610 1680 1626
rect 1742 2002 1776 2018
rect 1742 1610 1776 1626
rect 1838 2002 1872 2018
rect 1838 1610 1872 1626
rect 1934 2002 1968 2018
rect 1934 1610 1968 1626
rect 2030 2002 2064 2018
rect 2030 1610 2064 1626
rect 2126 2002 2160 2018
rect 2126 1610 2160 1626
rect 1582 1542 1598 1576
rect 1632 1542 1648 1576
rect 1774 1542 1790 1576
rect 1824 1542 1840 1576
rect 1966 1542 1982 1576
rect 2016 1542 2032 1576
rect 1436 1474 1470 1536
rect 2476 2710 2510 2760
rect 2240 1474 2274 1536
rect 1138 1440 1236 1452
rect 396 1384 1236 1440
rect 1436 1440 1532 1474
rect 2178 1452 2274 1474
rect 2376 1536 2476 2008
rect 3280 2710 3314 2772
rect 2622 2670 2638 2704
rect 2672 2670 2688 2704
rect 2814 2670 2830 2704
rect 2864 2670 2880 2704
rect 3006 2670 3022 2704
rect 3056 2670 3072 2704
rect 2590 2620 2624 2636
rect 2590 2228 2624 2244
rect 2686 2620 2720 2636
rect 2686 2228 2720 2244
rect 2782 2620 2816 2636
rect 2782 2228 2816 2244
rect 2878 2620 2912 2636
rect 2878 2228 2912 2244
rect 2974 2620 3008 2636
rect 2974 2228 3008 2244
rect 3070 2620 3104 2636
rect 3070 2228 3104 2244
rect 3166 2620 3200 2636
rect 3166 2228 3200 2244
rect 2718 2160 2734 2194
rect 2768 2160 2784 2194
rect 2910 2160 2926 2194
rect 2960 2160 2976 2194
rect 3102 2160 3118 2194
rect 3152 2160 3168 2194
rect 2718 2052 2734 2086
rect 2768 2052 2784 2086
rect 2910 2052 2926 2086
rect 2960 2052 2976 2086
rect 3102 2052 3118 2086
rect 3152 2052 3168 2086
rect 2590 2002 2624 2018
rect 2590 1610 2624 1626
rect 2686 2002 2720 2018
rect 2686 1610 2720 1626
rect 2782 2002 2816 2018
rect 2782 1610 2816 1626
rect 2878 2002 2912 2018
rect 2878 1610 2912 1626
rect 2974 2002 3008 2018
rect 2974 1610 3008 1626
rect 3070 2002 3104 2018
rect 3070 1610 3104 1626
rect 3166 2002 3200 2018
rect 3166 1610 3200 1626
rect 2622 1542 2638 1576
rect 2672 1542 2688 1576
rect 2814 1542 2830 1576
rect 2864 1542 2880 1576
rect 3006 1542 3022 1576
rect 3056 1542 3072 1576
rect 2376 1474 2510 1536
rect 3280 1474 3314 1536
rect 2178 1440 2276 1452
rect 1436 1384 2276 1440
rect 2376 1440 2572 1474
rect 3218 1452 3314 1474
rect 4924 2870 4958 2932
rect 4266 2830 4282 2864
rect 4316 2830 4332 2864
rect 4458 2830 4474 2864
rect 4508 2830 4524 2864
rect 4650 2830 4666 2864
rect 4700 2830 4716 2864
rect 4234 2780 4268 2796
rect 4234 2388 4268 2404
rect 4330 2780 4364 2796
rect 4330 2388 4364 2404
rect 4426 2780 4460 2796
rect 4426 2388 4460 2404
rect 4522 2780 4556 2796
rect 4522 2388 4556 2404
rect 4618 2780 4652 2796
rect 4618 2388 4652 2404
rect 4714 2780 4748 2796
rect 4714 2388 4748 2404
rect 4810 2780 4844 2796
rect 4810 2388 4844 2404
rect 4362 2320 4378 2354
rect 4412 2320 4428 2354
rect 4554 2320 4570 2354
rect 4604 2320 4620 2354
rect 4746 2320 4762 2354
rect 4796 2320 4812 2354
rect 4362 2212 4378 2246
rect 4412 2212 4428 2246
rect 4554 2212 4570 2246
rect 4604 2212 4620 2246
rect 4746 2212 4762 2246
rect 4796 2212 4812 2246
rect 4234 2162 4268 2178
rect 4234 1770 4268 1786
rect 4330 2162 4364 2178
rect 4330 1770 4364 1786
rect 4426 2162 4460 2178
rect 4426 1770 4460 1786
rect 4522 2162 4556 2178
rect 4522 1770 4556 1786
rect 4618 2162 4652 2178
rect 4618 1770 4652 1786
rect 4714 2162 4748 2178
rect 4714 1770 4748 1786
rect 4810 2162 4844 2178
rect 4810 1770 4844 1786
rect 4266 1702 4282 1736
rect 4316 1702 4332 1736
rect 4458 1702 4474 1736
rect 4508 1702 4524 1736
rect 4650 1702 4666 1736
rect 4700 1702 4716 1736
rect 4120 1634 4154 1696
rect 4924 1634 4958 1696
rect 4120 1600 4216 1634
rect 4862 1612 4958 1634
rect 5160 2932 5256 2960
rect 5902 2960 6296 2966
rect 5902 2932 5998 2960
rect 5160 2870 5194 2932
rect 5964 2870 5998 2932
rect 5306 2830 5322 2864
rect 5356 2830 5372 2864
rect 5498 2830 5514 2864
rect 5548 2830 5564 2864
rect 5690 2830 5706 2864
rect 5740 2830 5756 2864
rect 5274 2780 5308 2796
rect 5274 2388 5308 2404
rect 5370 2780 5404 2796
rect 5370 2388 5404 2404
rect 5466 2780 5500 2796
rect 5466 2388 5500 2404
rect 5562 2780 5596 2796
rect 5562 2388 5596 2404
rect 5658 2780 5692 2796
rect 5658 2388 5692 2404
rect 5754 2780 5788 2796
rect 5754 2388 5788 2404
rect 5850 2780 5884 2796
rect 5850 2388 5884 2404
rect 5402 2320 5418 2354
rect 5452 2320 5468 2354
rect 5594 2320 5610 2354
rect 5644 2320 5660 2354
rect 5786 2320 5802 2354
rect 5836 2320 5852 2354
rect 5402 2212 5418 2246
rect 5452 2212 5468 2246
rect 5594 2212 5610 2246
rect 5644 2212 5660 2246
rect 5786 2212 5802 2246
rect 5836 2212 5852 2246
rect 5274 2162 5308 2178
rect 5274 1770 5308 1786
rect 5370 2162 5404 2178
rect 5370 1770 5404 1786
rect 5466 2162 5500 2178
rect 5466 1770 5500 1786
rect 5562 2162 5596 2178
rect 5562 1770 5596 1786
rect 5658 2162 5692 2178
rect 5658 1770 5692 1786
rect 5754 2162 5788 2178
rect 5754 1770 5788 1786
rect 5850 2162 5884 2178
rect 5850 1770 5884 1786
rect 5306 1702 5322 1736
rect 5356 1702 5372 1736
rect 5498 1702 5514 1736
rect 5548 1702 5564 1736
rect 5690 1702 5706 1736
rect 5740 1702 5756 1736
rect 5160 1634 5194 1696
rect 5964 1634 5998 1696
rect 4862 1600 4960 1612
rect 4120 1544 4960 1600
rect 5160 1600 5256 1634
rect 5902 1612 5998 1634
rect 6200 2932 6296 2960
rect 6942 2960 7336 2966
rect 6942 2932 7038 2960
rect 6200 2870 6234 2932
rect 7004 2870 7038 2932
rect 6346 2830 6362 2864
rect 6396 2830 6412 2864
rect 6538 2830 6554 2864
rect 6588 2830 6604 2864
rect 6730 2830 6746 2864
rect 6780 2830 6796 2864
rect 6314 2780 6348 2796
rect 6314 2388 6348 2404
rect 6410 2780 6444 2796
rect 6410 2388 6444 2404
rect 6506 2780 6540 2796
rect 6506 2388 6540 2404
rect 6602 2780 6636 2796
rect 6602 2388 6636 2404
rect 6698 2780 6732 2796
rect 6698 2388 6732 2404
rect 6794 2780 6828 2796
rect 6794 2388 6828 2404
rect 6890 2780 6924 2796
rect 6890 2388 6924 2404
rect 6442 2320 6458 2354
rect 6492 2320 6508 2354
rect 6634 2320 6650 2354
rect 6684 2320 6700 2354
rect 6826 2320 6842 2354
rect 6876 2320 6892 2354
rect 6442 2212 6458 2246
rect 6492 2212 6508 2246
rect 6634 2212 6650 2246
rect 6684 2212 6700 2246
rect 6826 2212 6842 2246
rect 6876 2212 6892 2246
rect 6314 2162 6348 2178
rect 6314 1770 6348 1786
rect 6410 2162 6444 2178
rect 6410 1770 6444 1786
rect 6506 2162 6540 2178
rect 6506 1770 6540 1786
rect 6602 2162 6636 2178
rect 6602 1770 6636 1786
rect 6698 2162 6732 2178
rect 6698 1770 6732 1786
rect 6794 2162 6828 2178
rect 6794 1770 6828 1786
rect 6890 2162 6924 2178
rect 6890 1770 6924 1786
rect 6346 1702 6362 1736
rect 6396 1702 6412 1736
rect 6538 1702 6554 1736
rect 6588 1702 6604 1736
rect 6730 1702 6746 1736
rect 6780 1702 6796 1736
rect 6200 1634 6234 1696
rect 7004 1634 7038 1696
rect 5902 1600 6000 1612
rect 5160 1544 6000 1600
rect 6200 1600 6296 1634
rect 6942 1612 7038 1634
rect 7240 2932 7336 2960
rect 7982 2960 8376 2966
rect 7982 2932 8078 2960
rect 7240 2870 7274 2932
rect 8044 2870 8078 2932
rect 7386 2830 7402 2864
rect 7436 2830 7452 2864
rect 7578 2830 7594 2864
rect 7628 2830 7644 2864
rect 7770 2830 7786 2864
rect 7820 2830 7836 2864
rect 7354 2780 7388 2796
rect 7354 2388 7388 2404
rect 7450 2780 7484 2796
rect 7450 2388 7484 2404
rect 7546 2780 7580 2796
rect 7546 2388 7580 2404
rect 7642 2780 7676 2796
rect 7642 2388 7676 2404
rect 7738 2780 7772 2796
rect 7738 2388 7772 2404
rect 7834 2780 7868 2796
rect 7834 2388 7868 2404
rect 7930 2780 7964 2796
rect 7930 2388 7964 2404
rect 7482 2320 7498 2354
rect 7532 2320 7548 2354
rect 7674 2320 7690 2354
rect 7724 2320 7740 2354
rect 7866 2320 7882 2354
rect 7916 2320 7932 2354
rect 7482 2212 7498 2246
rect 7532 2212 7548 2246
rect 7674 2212 7690 2246
rect 7724 2212 7740 2246
rect 7866 2212 7882 2246
rect 7916 2212 7932 2246
rect 7354 2162 7388 2178
rect 7354 1770 7388 1786
rect 7450 2162 7484 2178
rect 7450 1770 7484 1786
rect 7546 2162 7580 2178
rect 7546 1770 7580 1786
rect 7642 2162 7676 2178
rect 7642 1770 7676 1786
rect 7738 2162 7772 2178
rect 7738 1770 7772 1786
rect 7834 2162 7868 2178
rect 7834 1770 7868 1786
rect 7930 2162 7964 2178
rect 7930 1770 7964 1786
rect 7386 1702 7402 1736
rect 7436 1702 7452 1736
rect 7578 1702 7594 1736
rect 7628 1702 7644 1736
rect 7770 1702 7786 1736
rect 7820 1702 7836 1736
rect 7240 1634 7274 1696
rect 8044 1634 8078 1696
rect 6942 1600 7040 1612
rect 6200 1544 7040 1600
rect 7240 1600 7336 1634
rect 7982 1612 8078 1634
rect 8280 2932 8376 2960
rect 9022 2960 9416 2966
rect 9022 2932 9118 2960
rect 8280 2870 8314 2932
rect 9084 2870 9118 2932
rect 8426 2830 8442 2864
rect 8476 2830 8492 2864
rect 8618 2830 8634 2864
rect 8668 2830 8684 2864
rect 8810 2830 8826 2864
rect 8860 2830 8876 2864
rect 8394 2780 8428 2796
rect 8394 2388 8428 2404
rect 8490 2780 8524 2796
rect 8490 2388 8524 2404
rect 8586 2780 8620 2796
rect 8586 2388 8620 2404
rect 8682 2780 8716 2796
rect 8682 2388 8716 2404
rect 8778 2780 8812 2796
rect 8778 2388 8812 2404
rect 8874 2780 8908 2796
rect 8874 2388 8908 2404
rect 8970 2780 9004 2796
rect 8970 2388 9004 2404
rect 8522 2320 8538 2354
rect 8572 2320 8588 2354
rect 8714 2320 8730 2354
rect 8764 2320 8780 2354
rect 8906 2320 8922 2354
rect 8956 2320 8972 2354
rect 8522 2212 8538 2246
rect 8572 2212 8588 2246
rect 8714 2212 8730 2246
rect 8764 2212 8780 2246
rect 8906 2212 8922 2246
rect 8956 2212 8972 2246
rect 8394 2162 8428 2178
rect 8394 1770 8428 1786
rect 8490 2162 8524 2178
rect 8490 1770 8524 1786
rect 8586 2162 8620 2178
rect 8586 1770 8620 1786
rect 8682 2162 8716 2178
rect 8682 1770 8716 1786
rect 8778 2162 8812 2178
rect 8778 1770 8812 1786
rect 8874 2162 8908 2178
rect 8874 1770 8908 1786
rect 8970 2162 9004 2178
rect 8970 1770 9004 1786
rect 8426 1702 8442 1736
rect 8476 1702 8492 1736
rect 8618 1702 8634 1736
rect 8668 1702 8684 1736
rect 8810 1702 8826 1736
rect 8860 1702 8876 1736
rect 8280 1634 8314 1696
rect 9084 1634 9118 1696
rect 7982 1600 8080 1612
rect 7240 1544 8080 1600
rect 8280 1600 8376 1634
rect 9022 1612 9118 1634
rect 9320 2932 9416 2960
rect 10062 2960 10456 2966
rect 10062 2932 10158 2960
rect 9320 2870 9354 2932
rect 10124 2870 10158 2932
rect 9466 2830 9482 2864
rect 9516 2830 9532 2864
rect 9658 2830 9674 2864
rect 9708 2830 9724 2864
rect 9850 2830 9866 2864
rect 9900 2830 9916 2864
rect 9434 2780 9468 2796
rect 9434 2388 9468 2404
rect 9530 2780 9564 2796
rect 9530 2388 9564 2404
rect 9626 2780 9660 2796
rect 9626 2388 9660 2404
rect 9722 2780 9756 2796
rect 9722 2388 9756 2404
rect 9818 2780 9852 2796
rect 9818 2388 9852 2404
rect 9914 2780 9948 2796
rect 9914 2388 9948 2404
rect 10010 2780 10044 2796
rect 10010 2388 10044 2404
rect 9562 2320 9578 2354
rect 9612 2320 9628 2354
rect 9754 2320 9770 2354
rect 9804 2320 9820 2354
rect 9946 2320 9962 2354
rect 9996 2320 10012 2354
rect 9562 2212 9578 2246
rect 9612 2212 9628 2246
rect 9754 2212 9770 2246
rect 9804 2212 9820 2246
rect 9946 2212 9962 2246
rect 9996 2212 10012 2246
rect 9434 2162 9468 2178
rect 9434 1770 9468 1786
rect 9530 2162 9564 2178
rect 9530 1770 9564 1786
rect 9626 2162 9660 2178
rect 9626 1770 9660 1786
rect 9722 2162 9756 2178
rect 9722 1770 9756 1786
rect 9818 2162 9852 2178
rect 9818 1770 9852 1786
rect 9914 2162 9948 2178
rect 9914 1770 9948 1786
rect 10010 2162 10044 2178
rect 10010 1770 10044 1786
rect 9466 1702 9482 1736
rect 9516 1702 9532 1736
rect 9658 1702 9674 1736
rect 9708 1702 9724 1736
rect 9850 1702 9866 1736
rect 9900 1702 9916 1736
rect 9320 1634 9354 1696
rect 10124 1634 10158 1696
rect 9022 1600 9120 1612
rect 8280 1544 9120 1600
rect 9320 1600 9416 1634
rect 10062 1612 10158 1634
rect 10360 2932 10456 2960
rect 11102 2932 11198 2966
rect 10360 2870 10394 2932
rect 11164 2870 11198 2932
rect 10506 2830 10522 2864
rect 10556 2830 10572 2864
rect 10698 2830 10714 2864
rect 10748 2830 10764 2864
rect 10890 2830 10906 2864
rect 10940 2830 10956 2864
rect 10474 2780 10508 2796
rect 10474 2388 10508 2404
rect 10570 2780 10604 2796
rect 10570 2388 10604 2404
rect 10666 2780 10700 2796
rect 10666 2388 10700 2404
rect 10762 2780 10796 2796
rect 10762 2388 10796 2404
rect 10858 2780 10892 2796
rect 10858 2388 10892 2404
rect 10954 2780 10988 2796
rect 10954 2388 10988 2404
rect 11050 2780 11084 2796
rect 11050 2388 11084 2404
rect 10602 2320 10618 2354
rect 10652 2320 10668 2354
rect 10794 2320 10810 2354
rect 10844 2320 10860 2354
rect 10986 2320 11002 2354
rect 11036 2320 11052 2354
rect 10602 2212 10618 2246
rect 10652 2212 10668 2246
rect 10794 2212 10810 2246
rect 10844 2212 10860 2246
rect 10986 2212 11002 2246
rect 11036 2212 11052 2246
rect 10474 2162 10508 2178
rect 10474 1770 10508 1786
rect 10570 2162 10604 2178
rect 10570 1770 10604 1786
rect 10666 2162 10700 2178
rect 10666 1770 10700 1786
rect 10762 2162 10796 2178
rect 10762 1770 10796 1786
rect 10858 2162 10892 2178
rect 10858 1770 10892 1786
rect 10954 2162 10988 2178
rect 10954 1770 10988 1786
rect 11050 2162 11084 2178
rect 11050 1770 11084 1786
rect 10506 1702 10522 1736
rect 10556 1702 10572 1736
rect 10698 1702 10714 1736
rect 10748 1702 10764 1736
rect 10890 1702 10906 1736
rect 10940 1702 10956 1736
rect 10360 1634 10394 1696
rect 11164 1634 11198 1696
rect 10062 1600 10160 1612
rect 9320 1544 10160 1600
rect 10360 1600 10456 1634
rect 11102 1612 11198 1634
rect 11740 2932 11836 2966
rect 12482 2960 12876 2966
rect 12482 2932 12578 2960
rect 11740 2870 11774 2932
rect 12544 2870 12578 2932
rect 11886 2830 11902 2864
rect 11936 2830 11952 2864
rect 12078 2830 12094 2864
rect 12128 2830 12144 2864
rect 12270 2830 12286 2864
rect 12320 2830 12336 2864
rect 11854 2780 11888 2796
rect 11854 2388 11888 2404
rect 11950 2780 11984 2796
rect 11950 2388 11984 2404
rect 12046 2780 12080 2796
rect 12046 2388 12080 2404
rect 12142 2780 12176 2796
rect 12142 2388 12176 2404
rect 12238 2780 12272 2796
rect 12238 2388 12272 2404
rect 12334 2780 12368 2796
rect 12334 2388 12368 2404
rect 12430 2780 12464 2796
rect 12430 2388 12464 2404
rect 11982 2320 11998 2354
rect 12032 2320 12048 2354
rect 12174 2320 12190 2354
rect 12224 2320 12240 2354
rect 12366 2320 12382 2354
rect 12416 2320 12432 2354
rect 11982 2212 11998 2246
rect 12032 2212 12048 2246
rect 12174 2212 12190 2246
rect 12224 2212 12240 2246
rect 12366 2212 12382 2246
rect 12416 2212 12432 2246
rect 11854 2162 11888 2178
rect 11854 1770 11888 1786
rect 11950 2162 11984 2178
rect 11950 1770 11984 1786
rect 12046 2162 12080 2178
rect 12046 1770 12080 1786
rect 12142 2162 12176 2178
rect 12142 1770 12176 1786
rect 12238 2162 12272 2178
rect 12238 1770 12272 1786
rect 12334 2162 12368 2178
rect 12334 1770 12368 1786
rect 12430 2162 12464 2178
rect 12430 1770 12464 1786
rect 11886 1702 11902 1736
rect 11936 1702 11952 1736
rect 12078 1702 12094 1736
rect 12128 1702 12144 1736
rect 12270 1702 12286 1736
rect 12320 1702 12336 1736
rect 11740 1634 11774 1696
rect 12544 1634 12578 1696
rect 11102 1600 11200 1612
rect 10360 1544 11200 1600
rect 11740 1600 11836 1634
rect 12482 1612 12578 1634
rect 12780 2932 12876 2960
rect 13522 2960 13916 2966
rect 13522 2932 13618 2960
rect 12780 2870 12814 2932
rect 13584 2870 13618 2932
rect 12926 2830 12942 2864
rect 12976 2830 12992 2864
rect 13118 2830 13134 2864
rect 13168 2830 13184 2864
rect 13310 2830 13326 2864
rect 13360 2830 13376 2864
rect 12894 2780 12928 2796
rect 12894 2388 12928 2404
rect 12990 2780 13024 2796
rect 12990 2388 13024 2404
rect 13086 2780 13120 2796
rect 13086 2388 13120 2404
rect 13182 2780 13216 2796
rect 13182 2388 13216 2404
rect 13278 2780 13312 2796
rect 13278 2388 13312 2404
rect 13374 2780 13408 2796
rect 13374 2388 13408 2404
rect 13470 2780 13504 2796
rect 13470 2388 13504 2404
rect 13022 2320 13038 2354
rect 13072 2320 13088 2354
rect 13214 2320 13230 2354
rect 13264 2320 13280 2354
rect 13406 2320 13422 2354
rect 13456 2320 13472 2354
rect 13022 2212 13038 2246
rect 13072 2212 13088 2246
rect 13214 2212 13230 2246
rect 13264 2212 13280 2246
rect 13406 2212 13422 2246
rect 13456 2212 13472 2246
rect 12894 2162 12928 2178
rect 12894 1770 12928 1786
rect 12990 2162 13024 2178
rect 12990 1770 13024 1786
rect 13086 2162 13120 2178
rect 13086 1770 13120 1786
rect 13182 2162 13216 2178
rect 13182 1770 13216 1786
rect 13278 2162 13312 2178
rect 13278 1770 13312 1786
rect 13374 2162 13408 2178
rect 13374 1770 13408 1786
rect 13470 2162 13504 2178
rect 13470 1770 13504 1786
rect 12926 1702 12942 1736
rect 12976 1702 12992 1736
rect 13118 1702 13134 1736
rect 13168 1702 13184 1736
rect 13310 1702 13326 1736
rect 13360 1702 13376 1736
rect 12780 1634 12814 1696
rect 13584 1634 13618 1696
rect 12482 1600 12580 1612
rect 11740 1544 12580 1600
rect 12780 1600 12876 1634
rect 13522 1612 13618 1634
rect 13820 2932 13916 2960
rect 14562 2960 14956 2966
rect 14562 2932 14658 2960
rect 13820 2870 13854 2932
rect 14624 2870 14658 2932
rect 13966 2830 13982 2864
rect 14016 2830 14032 2864
rect 14158 2830 14174 2864
rect 14208 2830 14224 2864
rect 14350 2830 14366 2864
rect 14400 2830 14416 2864
rect 13934 2780 13968 2796
rect 13934 2388 13968 2404
rect 14030 2780 14064 2796
rect 14030 2388 14064 2404
rect 14126 2780 14160 2796
rect 14126 2388 14160 2404
rect 14222 2780 14256 2796
rect 14222 2388 14256 2404
rect 14318 2780 14352 2796
rect 14318 2388 14352 2404
rect 14414 2780 14448 2796
rect 14414 2388 14448 2404
rect 14510 2780 14544 2796
rect 14510 2388 14544 2404
rect 14062 2320 14078 2354
rect 14112 2320 14128 2354
rect 14254 2320 14270 2354
rect 14304 2320 14320 2354
rect 14446 2320 14462 2354
rect 14496 2320 14512 2354
rect 14062 2212 14078 2246
rect 14112 2212 14128 2246
rect 14254 2212 14270 2246
rect 14304 2212 14320 2246
rect 14446 2212 14462 2246
rect 14496 2212 14512 2246
rect 13934 2162 13968 2178
rect 13934 1770 13968 1786
rect 14030 2162 14064 2178
rect 14030 1770 14064 1786
rect 14126 2162 14160 2178
rect 14126 1770 14160 1786
rect 14222 2162 14256 2178
rect 14222 1770 14256 1786
rect 14318 2162 14352 2178
rect 14318 1770 14352 1786
rect 14414 2162 14448 2178
rect 14414 1770 14448 1786
rect 14510 2162 14544 2178
rect 14510 1770 14544 1786
rect 13966 1702 13982 1736
rect 14016 1702 14032 1736
rect 14158 1702 14174 1736
rect 14208 1702 14224 1736
rect 14350 1702 14366 1736
rect 14400 1702 14416 1736
rect 13820 1634 13854 1696
rect 14624 1634 14658 1696
rect 13522 1600 13620 1612
rect 12780 1544 13620 1600
rect 13820 1600 13916 1634
rect 14562 1612 14658 1634
rect 14860 2932 14956 2960
rect 15602 2960 15996 2966
rect 15602 2932 15698 2960
rect 14860 2870 14894 2932
rect 15664 2870 15698 2932
rect 15006 2830 15022 2864
rect 15056 2830 15072 2864
rect 15198 2830 15214 2864
rect 15248 2830 15264 2864
rect 15390 2830 15406 2864
rect 15440 2830 15456 2864
rect 14974 2780 15008 2796
rect 14974 2388 15008 2404
rect 15070 2780 15104 2796
rect 15070 2388 15104 2404
rect 15166 2780 15200 2796
rect 15166 2388 15200 2404
rect 15262 2780 15296 2796
rect 15262 2388 15296 2404
rect 15358 2780 15392 2796
rect 15358 2388 15392 2404
rect 15454 2780 15488 2796
rect 15454 2388 15488 2404
rect 15550 2780 15584 2796
rect 15550 2388 15584 2404
rect 15102 2320 15118 2354
rect 15152 2320 15168 2354
rect 15294 2320 15310 2354
rect 15344 2320 15360 2354
rect 15486 2320 15502 2354
rect 15536 2320 15552 2354
rect 15102 2212 15118 2246
rect 15152 2212 15168 2246
rect 15294 2212 15310 2246
rect 15344 2212 15360 2246
rect 15486 2212 15502 2246
rect 15536 2212 15552 2246
rect 14974 2162 15008 2178
rect 14974 1770 15008 1786
rect 15070 2162 15104 2178
rect 15070 1770 15104 1786
rect 15166 2162 15200 2178
rect 15166 1770 15200 1786
rect 15262 2162 15296 2178
rect 15262 1770 15296 1786
rect 15358 2162 15392 2178
rect 15358 1770 15392 1786
rect 15454 2162 15488 2178
rect 15454 1770 15488 1786
rect 15550 2162 15584 2178
rect 15550 1770 15584 1786
rect 15006 1702 15022 1736
rect 15056 1702 15072 1736
rect 15198 1702 15214 1736
rect 15248 1702 15264 1736
rect 15390 1702 15406 1736
rect 15440 1702 15456 1736
rect 14860 1634 14894 1696
rect 15664 1634 15698 1696
rect 14562 1600 14660 1612
rect 13820 1544 14660 1600
rect 14860 1600 14956 1634
rect 15602 1612 15698 1634
rect 15900 2932 15996 2960
rect 16642 2960 17036 2966
rect 16642 2932 16738 2960
rect 15900 2870 15934 2932
rect 16704 2870 16738 2932
rect 16046 2830 16062 2864
rect 16096 2830 16112 2864
rect 16238 2830 16254 2864
rect 16288 2830 16304 2864
rect 16430 2830 16446 2864
rect 16480 2830 16496 2864
rect 16014 2780 16048 2796
rect 16014 2388 16048 2404
rect 16110 2780 16144 2796
rect 16110 2388 16144 2404
rect 16206 2780 16240 2796
rect 16206 2388 16240 2404
rect 16302 2780 16336 2796
rect 16302 2388 16336 2404
rect 16398 2780 16432 2796
rect 16398 2388 16432 2404
rect 16494 2780 16528 2796
rect 16494 2388 16528 2404
rect 16590 2780 16624 2796
rect 16590 2388 16624 2404
rect 16142 2320 16158 2354
rect 16192 2320 16208 2354
rect 16334 2320 16350 2354
rect 16384 2320 16400 2354
rect 16526 2320 16542 2354
rect 16576 2320 16592 2354
rect 16142 2212 16158 2246
rect 16192 2212 16208 2246
rect 16334 2212 16350 2246
rect 16384 2212 16400 2246
rect 16526 2212 16542 2246
rect 16576 2212 16592 2246
rect 16014 2162 16048 2178
rect 16014 1770 16048 1786
rect 16110 2162 16144 2178
rect 16110 1770 16144 1786
rect 16206 2162 16240 2178
rect 16206 1770 16240 1786
rect 16302 2162 16336 2178
rect 16302 1770 16336 1786
rect 16398 2162 16432 2178
rect 16398 1770 16432 1786
rect 16494 2162 16528 2178
rect 16494 1770 16528 1786
rect 16590 2162 16624 2178
rect 16590 1770 16624 1786
rect 16046 1702 16062 1736
rect 16096 1702 16112 1736
rect 16238 1702 16254 1736
rect 16288 1702 16304 1736
rect 16430 1702 16446 1736
rect 16480 1702 16496 1736
rect 15900 1634 15934 1696
rect 16704 1634 16738 1696
rect 15602 1600 15700 1612
rect 14860 1544 15700 1600
rect 15900 1600 15996 1634
rect 16642 1612 16738 1634
rect 16940 2932 17036 2960
rect 17682 2960 18076 2966
rect 17682 2932 17778 2960
rect 16940 2870 16974 2932
rect 17744 2870 17778 2932
rect 17086 2830 17102 2864
rect 17136 2830 17152 2864
rect 17278 2830 17294 2864
rect 17328 2830 17344 2864
rect 17470 2830 17486 2864
rect 17520 2830 17536 2864
rect 17054 2780 17088 2796
rect 17054 2388 17088 2404
rect 17150 2780 17184 2796
rect 17150 2388 17184 2404
rect 17246 2780 17280 2796
rect 17246 2388 17280 2404
rect 17342 2780 17376 2796
rect 17342 2388 17376 2404
rect 17438 2780 17472 2796
rect 17438 2388 17472 2404
rect 17534 2780 17568 2796
rect 17534 2388 17568 2404
rect 17630 2780 17664 2796
rect 17630 2388 17664 2404
rect 17182 2320 17198 2354
rect 17232 2320 17248 2354
rect 17374 2320 17390 2354
rect 17424 2320 17440 2354
rect 17566 2320 17582 2354
rect 17616 2320 17632 2354
rect 17182 2212 17198 2246
rect 17232 2212 17248 2246
rect 17374 2212 17390 2246
rect 17424 2212 17440 2246
rect 17566 2212 17582 2246
rect 17616 2212 17632 2246
rect 17054 2162 17088 2178
rect 17054 1770 17088 1786
rect 17150 2162 17184 2178
rect 17150 1770 17184 1786
rect 17246 2162 17280 2178
rect 17246 1770 17280 1786
rect 17342 2162 17376 2178
rect 17342 1770 17376 1786
rect 17438 2162 17472 2178
rect 17438 1770 17472 1786
rect 17534 2162 17568 2178
rect 17534 1770 17568 1786
rect 17630 2162 17664 2178
rect 17630 1770 17664 1786
rect 17086 1702 17102 1736
rect 17136 1702 17152 1736
rect 17278 1702 17294 1736
rect 17328 1702 17344 1736
rect 17470 1702 17486 1736
rect 17520 1702 17536 1736
rect 16940 1634 16974 1696
rect 17744 1634 17778 1696
rect 16642 1600 16740 1612
rect 15900 1544 16740 1600
rect 16940 1600 17036 1634
rect 17682 1612 17778 1634
rect 17980 2932 18076 2960
rect 18722 2932 18818 2966
rect 17980 2870 18014 2932
rect 18784 2870 18818 2932
rect 18126 2830 18142 2864
rect 18176 2830 18192 2864
rect 18318 2830 18334 2864
rect 18368 2830 18384 2864
rect 18510 2830 18526 2864
rect 18560 2830 18576 2864
rect 18094 2780 18128 2796
rect 18094 2388 18128 2404
rect 18190 2780 18224 2796
rect 18190 2388 18224 2404
rect 18286 2780 18320 2796
rect 18286 2388 18320 2404
rect 18382 2780 18416 2796
rect 18382 2388 18416 2404
rect 18478 2780 18512 2796
rect 18478 2388 18512 2404
rect 18574 2780 18608 2796
rect 18574 2388 18608 2404
rect 18670 2780 18704 2796
rect 18670 2388 18704 2404
rect 18222 2320 18238 2354
rect 18272 2320 18288 2354
rect 18414 2320 18430 2354
rect 18464 2320 18480 2354
rect 18606 2320 18622 2354
rect 18656 2320 18672 2354
rect 18222 2212 18238 2246
rect 18272 2212 18288 2246
rect 18414 2212 18430 2246
rect 18464 2212 18480 2246
rect 18606 2212 18622 2246
rect 18656 2212 18672 2246
rect 18094 2162 18128 2178
rect 18094 1770 18128 1786
rect 18190 2162 18224 2178
rect 18190 1770 18224 1786
rect 18286 2162 18320 2178
rect 18286 1770 18320 1786
rect 18382 2162 18416 2178
rect 18382 1770 18416 1786
rect 18478 2162 18512 2178
rect 18478 1770 18512 1786
rect 18574 2162 18608 2178
rect 18574 1770 18608 1786
rect 18670 2162 18704 2178
rect 18670 1770 18704 1786
rect 18126 1702 18142 1736
rect 18176 1702 18192 1736
rect 18318 1702 18334 1736
rect 18368 1702 18384 1736
rect 18510 1702 18526 1736
rect 18560 1702 18576 1736
rect 17980 1634 18014 1696
rect 18784 1634 18818 1696
rect 17682 1600 17780 1612
rect 16940 1544 17780 1600
rect 17980 1600 18076 1634
rect 18722 1612 18818 1634
rect 18722 1600 18820 1612
rect 17980 1544 18820 1600
rect 4120 1510 4216 1544
rect 4994 1510 5090 1544
rect 3218 1440 3316 1452
rect 2376 1384 3316 1440
rect 4120 1448 4154 1510
rect -1684 1350 -1588 1384
rect -810 1350 -548 1384
rect 230 1350 326 1384
rect -1684 1288 -1650 1350
rect -748 1288 -610 1350
rect -1527 1248 -1511 1282
rect -1477 1248 -1461 1282
rect -1409 1248 -1393 1282
rect -1359 1248 -1343 1282
rect -1291 1248 -1275 1282
rect -1241 1248 -1225 1282
rect -1173 1248 -1157 1282
rect -1123 1248 -1107 1282
rect -1055 1248 -1039 1282
rect -1005 1248 -989 1282
rect -937 1248 -921 1282
rect -887 1248 -871 1282
rect -1570 1198 -1536 1214
rect -1570 806 -1536 822
rect -1452 1198 -1418 1214
rect -1452 806 -1418 822
rect -1334 1198 -1300 1214
rect -1334 806 -1300 822
rect -1216 1198 -1182 1214
rect -1216 806 -1182 822
rect -1098 1198 -1064 1214
rect -1098 806 -1064 822
rect -980 1198 -946 1214
rect -980 806 -946 822
rect -862 1198 -828 1214
rect -862 806 -828 822
rect -1527 738 -1511 772
rect -1477 738 -1461 772
rect -1409 738 -1393 772
rect -1359 738 -1343 772
rect -1291 738 -1275 772
rect -1241 738 -1225 772
rect -1173 738 -1157 772
rect -1123 738 -1107 772
rect -1055 738 -1039 772
rect -1005 738 -989 772
rect -937 738 -921 772
rect -887 738 -871 772
rect -1684 670 -1650 732
rect -714 732 -644 1288
rect 292 1288 326 1350
rect -487 1248 -471 1282
rect -437 1248 -421 1282
rect -369 1248 -353 1282
rect -319 1248 -303 1282
rect -251 1248 -235 1282
rect -201 1248 -185 1282
rect -133 1248 -117 1282
rect -83 1248 -67 1282
rect -15 1248 1 1282
rect 35 1248 51 1282
rect 103 1248 119 1282
rect 153 1248 169 1282
rect -530 1198 -496 1214
rect -530 806 -496 822
rect -412 1198 -378 1214
rect -412 806 -378 822
rect -294 1198 -260 1214
rect -294 806 -260 822
rect -176 1198 -142 1214
rect -176 806 -142 822
rect -58 1198 -24 1214
rect -58 806 -24 822
rect 60 1198 94 1214
rect 60 806 94 822
rect 178 1198 212 1214
rect 178 806 212 822
rect -487 738 -471 772
rect -437 738 -421 772
rect -369 738 -353 772
rect -319 738 -303 772
rect -251 738 -235 772
rect -201 738 -185 772
rect -133 738 -117 772
rect -83 738 -67 772
rect -15 738 1 772
rect 35 738 51 772
rect 103 738 119 772
rect 153 738 169 772
rect -748 670 -610 732
rect 396 1350 492 1384
rect 1270 1350 1366 1384
rect 396 1288 430 1350
rect 326 788 396 1252
rect 292 670 326 732
rect -1684 652 -1588 670
rect -1688 636 -1588 652
rect -810 636 -548 670
rect 230 652 326 670
rect 1332 1288 1366 1350
rect 553 1248 569 1282
rect 603 1248 619 1282
rect 671 1248 687 1282
rect 721 1248 737 1282
rect 789 1248 805 1282
rect 839 1248 855 1282
rect 907 1248 923 1282
rect 957 1248 973 1282
rect 1025 1248 1041 1282
rect 1075 1248 1091 1282
rect 1143 1248 1159 1282
rect 1193 1248 1209 1282
rect 510 1198 544 1214
rect 510 806 544 822
rect 628 1198 662 1214
rect 628 806 662 822
rect 746 1198 780 1214
rect 746 806 780 822
rect 864 1198 898 1214
rect 864 806 898 822
rect 982 1198 1016 1214
rect 982 806 1016 822
rect 1100 1198 1134 1214
rect 1100 806 1134 822
rect 1218 1198 1252 1214
rect 1218 806 1252 822
rect 553 738 569 772
rect 603 738 619 772
rect 671 738 687 772
rect 721 738 737 772
rect 789 738 805 772
rect 839 738 855 772
rect 907 738 923 772
rect 957 738 973 772
rect 1025 738 1041 772
rect 1075 738 1091 772
rect 1143 738 1159 772
rect 1193 738 1209 772
rect 396 670 430 732
rect 1436 1350 1532 1384
rect 2310 1350 2572 1384
rect 3350 1350 3446 1384
rect 1436 1288 1470 1350
rect 1366 796 1436 1260
rect 1332 670 1366 732
rect 396 652 492 670
rect 230 636 492 652
rect 1270 636 1366 670
rect 2372 1288 2510 1350
rect 1593 1248 1609 1282
rect 1643 1248 1659 1282
rect 1711 1248 1727 1282
rect 1761 1248 1777 1282
rect 1829 1248 1845 1282
rect 1879 1248 1895 1282
rect 1947 1248 1963 1282
rect 1997 1248 2013 1282
rect 2065 1248 2081 1282
rect 2115 1248 2131 1282
rect 2183 1248 2199 1282
rect 2233 1248 2249 1282
rect 1550 1198 1584 1214
rect 1550 806 1584 822
rect 1668 1198 1702 1214
rect 1668 806 1702 822
rect 1786 1198 1820 1214
rect 1786 806 1820 822
rect 1904 1198 1938 1214
rect 1904 806 1938 822
rect 2022 1198 2056 1214
rect 2022 806 2056 822
rect 2140 1198 2174 1214
rect 2140 806 2174 822
rect 2258 1198 2292 1214
rect 2258 806 2292 822
rect 1593 738 1609 772
rect 1643 738 1659 772
rect 1711 738 1727 772
rect 1761 738 1777 772
rect 1829 738 1845 772
rect 1879 738 1895 772
rect 1947 738 1963 772
rect 1997 738 2013 772
rect 2065 738 2081 772
rect 2115 738 2131 772
rect 2183 738 2199 772
rect 2233 738 2249 772
rect 1436 670 1470 732
rect 2406 732 2476 1288
rect 3412 1288 3446 1350
rect 2633 1248 2649 1282
rect 2683 1248 2699 1282
rect 2751 1248 2767 1282
rect 2801 1248 2817 1282
rect 2869 1248 2885 1282
rect 2919 1248 2935 1282
rect 2987 1248 3003 1282
rect 3037 1248 3053 1282
rect 3105 1248 3121 1282
rect 3155 1248 3171 1282
rect 3223 1248 3239 1282
rect 3273 1248 3289 1282
rect 2590 1198 2624 1214
rect 2590 806 2624 822
rect 2708 1198 2742 1214
rect 2708 806 2742 822
rect 2826 1198 2860 1214
rect 2826 806 2860 822
rect 2944 1198 2978 1214
rect 2944 806 2978 822
rect 3062 1198 3096 1214
rect 3062 806 3096 822
rect 3180 1198 3214 1214
rect 3180 806 3214 822
rect 3298 1198 3332 1214
rect 3298 806 3332 822
rect 2633 738 2649 772
rect 2683 738 2699 772
rect 2751 738 2767 772
rect 2801 738 2817 772
rect 2869 738 2885 772
rect 2919 738 2935 772
rect 2987 738 3003 772
rect 3037 738 3053 772
rect 3105 738 3121 772
rect 3155 738 3171 772
rect 3223 738 3239 772
rect 3273 738 3289 772
rect 2372 670 2510 732
rect 5056 1448 5090 1510
rect 4277 1408 4293 1442
rect 4327 1408 4343 1442
rect 4395 1408 4411 1442
rect 4445 1408 4461 1442
rect 4513 1408 4529 1442
rect 4563 1408 4579 1442
rect 4631 1408 4647 1442
rect 4681 1408 4697 1442
rect 4749 1408 4765 1442
rect 4799 1408 4815 1442
rect 4867 1408 4883 1442
rect 4917 1408 4933 1442
rect 4234 1358 4268 1374
rect 4234 966 4268 982
rect 4352 1358 4386 1374
rect 4352 966 4386 982
rect 4470 1358 4504 1374
rect 4470 966 4504 982
rect 4588 1358 4622 1374
rect 4588 966 4622 982
rect 4706 1358 4740 1374
rect 4706 966 4740 982
rect 4824 1358 4858 1374
rect 4824 966 4858 982
rect 4942 1358 4976 1374
rect 4942 966 4976 982
rect 4277 898 4293 932
rect 4327 898 4343 932
rect 4395 898 4411 932
rect 4445 898 4461 932
rect 4513 898 4529 932
rect 4563 898 4579 932
rect 4631 898 4647 932
rect 4681 898 4697 932
rect 4749 898 4765 932
rect 4799 898 4815 932
rect 4867 898 4883 932
rect 4917 898 4933 932
rect 4120 830 4154 892
rect 5056 830 5090 892
rect 4120 796 4216 830
rect 4994 796 5090 830
rect 5160 1510 5256 1544
rect 6034 1510 6130 1544
rect 5160 1448 5194 1510
rect 6096 1448 6130 1510
rect 5317 1408 5333 1442
rect 5367 1408 5383 1442
rect 5435 1408 5451 1442
rect 5485 1408 5501 1442
rect 5553 1408 5569 1442
rect 5603 1408 5619 1442
rect 5671 1408 5687 1442
rect 5721 1408 5737 1442
rect 5789 1408 5805 1442
rect 5839 1408 5855 1442
rect 5907 1408 5923 1442
rect 5957 1408 5973 1442
rect 5274 1358 5308 1374
rect 5274 966 5308 982
rect 5392 1358 5426 1374
rect 5392 966 5426 982
rect 5510 1358 5544 1374
rect 5510 966 5544 982
rect 5628 1358 5662 1374
rect 5628 966 5662 982
rect 5746 1358 5780 1374
rect 5746 966 5780 982
rect 5864 1358 5898 1374
rect 5864 966 5898 982
rect 5982 1358 6016 1374
rect 5982 966 6016 982
rect 5317 898 5333 932
rect 5367 898 5383 932
rect 5435 898 5451 932
rect 5485 898 5501 932
rect 5553 898 5569 932
rect 5603 898 5619 932
rect 5671 898 5687 932
rect 5721 898 5737 932
rect 5789 898 5805 932
rect 5839 898 5855 932
rect 5907 898 5923 932
rect 5957 898 5973 932
rect 5160 830 5194 892
rect 6096 830 6130 892
rect 5160 796 5256 830
rect 6034 796 6130 830
rect 6200 1510 6296 1544
rect 7074 1510 7170 1544
rect 6200 1448 6234 1510
rect 7136 1448 7170 1510
rect 6357 1408 6373 1442
rect 6407 1408 6423 1442
rect 6475 1408 6491 1442
rect 6525 1408 6541 1442
rect 6593 1408 6609 1442
rect 6643 1408 6659 1442
rect 6711 1408 6727 1442
rect 6761 1408 6777 1442
rect 6829 1408 6845 1442
rect 6879 1408 6895 1442
rect 6947 1408 6963 1442
rect 6997 1408 7013 1442
rect 6314 1358 6348 1374
rect 6314 966 6348 982
rect 6432 1358 6466 1374
rect 6432 966 6466 982
rect 6550 1358 6584 1374
rect 6550 966 6584 982
rect 6668 1358 6702 1374
rect 6668 966 6702 982
rect 6786 1358 6820 1374
rect 6786 966 6820 982
rect 6904 1358 6938 1374
rect 6904 966 6938 982
rect 7022 1358 7056 1374
rect 7022 966 7056 982
rect 6357 898 6373 932
rect 6407 898 6423 932
rect 6475 898 6491 932
rect 6525 898 6541 932
rect 6593 898 6609 932
rect 6643 898 6659 932
rect 6711 898 6727 932
rect 6761 898 6777 932
rect 6829 898 6845 932
rect 6879 898 6895 932
rect 6947 898 6963 932
rect 6997 898 7013 932
rect 6200 830 6234 892
rect 7136 830 7170 892
rect 6200 796 6296 830
rect 7074 796 7170 830
rect 7240 1510 7336 1544
rect 8114 1510 8210 1544
rect 7240 1448 7274 1510
rect 8176 1448 8210 1510
rect 7397 1408 7413 1442
rect 7447 1408 7463 1442
rect 7515 1408 7531 1442
rect 7565 1408 7581 1442
rect 7633 1408 7649 1442
rect 7683 1408 7699 1442
rect 7751 1408 7767 1442
rect 7801 1408 7817 1442
rect 7869 1408 7885 1442
rect 7919 1408 7935 1442
rect 7987 1408 8003 1442
rect 8037 1408 8053 1442
rect 7354 1358 7388 1374
rect 7354 966 7388 982
rect 7472 1358 7506 1374
rect 7472 966 7506 982
rect 7590 1358 7624 1374
rect 7590 966 7624 982
rect 7708 1358 7742 1374
rect 7708 966 7742 982
rect 7826 1358 7860 1374
rect 7826 966 7860 982
rect 7944 1358 7978 1374
rect 7944 966 7978 982
rect 8062 1358 8096 1374
rect 8062 966 8096 982
rect 7397 898 7413 932
rect 7447 898 7463 932
rect 7515 898 7531 932
rect 7565 898 7581 932
rect 7633 898 7649 932
rect 7683 898 7699 932
rect 7751 898 7767 932
rect 7801 898 7817 932
rect 7869 898 7885 932
rect 7919 898 7935 932
rect 7987 898 8003 932
rect 8037 898 8053 932
rect 7240 830 7274 892
rect 8176 830 8210 892
rect 7240 796 7336 830
rect 8114 796 8210 830
rect 8280 1510 8376 1544
rect 9154 1510 9250 1544
rect 8280 1448 8314 1510
rect 9216 1448 9250 1510
rect 8437 1408 8453 1442
rect 8487 1408 8503 1442
rect 8555 1408 8571 1442
rect 8605 1408 8621 1442
rect 8673 1408 8689 1442
rect 8723 1408 8739 1442
rect 8791 1408 8807 1442
rect 8841 1408 8857 1442
rect 8909 1408 8925 1442
rect 8959 1408 8975 1442
rect 9027 1408 9043 1442
rect 9077 1408 9093 1442
rect 8394 1358 8428 1374
rect 8394 966 8428 982
rect 8512 1358 8546 1374
rect 8512 966 8546 982
rect 8630 1358 8664 1374
rect 8630 966 8664 982
rect 8748 1358 8782 1374
rect 8748 966 8782 982
rect 8866 1358 8900 1374
rect 8866 966 8900 982
rect 8984 1358 9018 1374
rect 8984 966 9018 982
rect 9102 1358 9136 1374
rect 9102 966 9136 982
rect 8437 898 8453 932
rect 8487 898 8503 932
rect 8555 898 8571 932
rect 8605 898 8621 932
rect 8673 898 8689 932
rect 8723 898 8739 932
rect 8791 898 8807 932
rect 8841 898 8857 932
rect 8909 898 8925 932
rect 8959 898 8975 932
rect 9027 898 9043 932
rect 9077 898 9093 932
rect 8280 830 8314 892
rect 9216 830 9250 892
rect 8280 796 8376 830
rect 9154 796 9250 830
rect 9320 1510 9416 1544
rect 10194 1510 10290 1544
rect 9320 1448 9354 1510
rect 10256 1448 10290 1510
rect 9477 1408 9493 1442
rect 9527 1408 9543 1442
rect 9595 1408 9611 1442
rect 9645 1408 9661 1442
rect 9713 1408 9729 1442
rect 9763 1408 9779 1442
rect 9831 1408 9847 1442
rect 9881 1408 9897 1442
rect 9949 1408 9965 1442
rect 9999 1408 10015 1442
rect 10067 1408 10083 1442
rect 10117 1408 10133 1442
rect 9434 1358 9468 1374
rect 9434 966 9468 982
rect 9552 1358 9586 1374
rect 9552 966 9586 982
rect 9670 1358 9704 1374
rect 9670 966 9704 982
rect 9788 1358 9822 1374
rect 9788 966 9822 982
rect 9906 1358 9940 1374
rect 9906 966 9940 982
rect 10024 1358 10058 1374
rect 10024 966 10058 982
rect 10142 1358 10176 1374
rect 10142 966 10176 982
rect 9477 898 9493 932
rect 9527 898 9543 932
rect 9595 898 9611 932
rect 9645 898 9661 932
rect 9713 898 9729 932
rect 9763 898 9779 932
rect 9831 898 9847 932
rect 9881 898 9897 932
rect 9949 898 9965 932
rect 9999 898 10015 932
rect 10067 898 10083 932
rect 10117 898 10133 932
rect 9320 830 9354 892
rect 10256 830 10290 892
rect 9320 796 9416 830
rect 10194 796 10290 830
rect 10360 1510 10456 1544
rect 11234 1510 11330 1544
rect 10360 1448 10394 1510
rect 11296 1448 11330 1510
rect 10517 1408 10533 1442
rect 10567 1408 10583 1442
rect 10635 1408 10651 1442
rect 10685 1408 10701 1442
rect 10753 1408 10769 1442
rect 10803 1408 10819 1442
rect 10871 1408 10887 1442
rect 10921 1408 10937 1442
rect 10989 1408 11005 1442
rect 11039 1408 11055 1442
rect 11107 1408 11123 1442
rect 11157 1408 11173 1442
rect 10474 1358 10508 1374
rect 10474 966 10508 982
rect 10592 1358 10626 1374
rect 10592 966 10626 982
rect 10710 1358 10744 1374
rect 10710 966 10744 982
rect 10828 1358 10862 1374
rect 10828 966 10862 982
rect 10946 1358 10980 1374
rect 10946 966 10980 982
rect 11064 1358 11098 1374
rect 11064 966 11098 982
rect 11182 1358 11216 1374
rect 11182 966 11216 982
rect 10517 898 10533 932
rect 10567 898 10583 932
rect 10635 898 10651 932
rect 10685 898 10701 932
rect 10753 898 10769 932
rect 10803 898 10819 932
rect 10871 898 10887 932
rect 10921 898 10937 932
rect 10989 898 11005 932
rect 11039 898 11055 932
rect 11107 898 11123 932
rect 11157 898 11173 932
rect 10360 830 10394 892
rect 11296 830 11330 892
rect 10360 796 10456 830
rect 11234 796 11330 830
rect 11740 1510 11836 1544
rect 12614 1510 12710 1544
rect 11740 1448 11774 1510
rect 12676 1448 12710 1510
rect 11897 1408 11913 1442
rect 11947 1408 11963 1442
rect 12015 1408 12031 1442
rect 12065 1408 12081 1442
rect 12133 1408 12149 1442
rect 12183 1408 12199 1442
rect 12251 1408 12267 1442
rect 12301 1408 12317 1442
rect 12369 1408 12385 1442
rect 12419 1408 12435 1442
rect 12487 1408 12503 1442
rect 12537 1408 12553 1442
rect 11854 1358 11888 1374
rect 11854 966 11888 982
rect 11972 1358 12006 1374
rect 11972 966 12006 982
rect 12090 1358 12124 1374
rect 12090 966 12124 982
rect 12208 1358 12242 1374
rect 12208 966 12242 982
rect 12326 1358 12360 1374
rect 12326 966 12360 982
rect 12444 1358 12478 1374
rect 12444 966 12478 982
rect 12562 1358 12596 1374
rect 12562 966 12596 982
rect 11897 898 11913 932
rect 11947 898 11963 932
rect 12015 898 12031 932
rect 12065 898 12081 932
rect 12133 898 12149 932
rect 12183 898 12199 932
rect 12251 898 12267 932
rect 12301 898 12317 932
rect 12369 898 12385 932
rect 12419 898 12435 932
rect 12487 898 12503 932
rect 12537 898 12553 932
rect 11740 830 11774 892
rect 12676 830 12710 892
rect 11740 796 11836 830
rect 12614 796 12710 830
rect 12780 1510 12876 1544
rect 13654 1510 13750 1544
rect 12780 1448 12814 1510
rect 13716 1448 13750 1510
rect 12937 1408 12953 1442
rect 12987 1408 13003 1442
rect 13055 1408 13071 1442
rect 13105 1408 13121 1442
rect 13173 1408 13189 1442
rect 13223 1408 13239 1442
rect 13291 1408 13307 1442
rect 13341 1408 13357 1442
rect 13409 1408 13425 1442
rect 13459 1408 13475 1442
rect 13527 1408 13543 1442
rect 13577 1408 13593 1442
rect 12894 1358 12928 1374
rect 12894 966 12928 982
rect 13012 1358 13046 1374
rect 13012 966 13046 982
rect 13130 1358 13164 1374
rect 13130 966 13164 982
rect 13248 1358 13282 1374
rect 13248 966 13282 982
rect 13366 1358 13400 1374
rect 13366 966 13400 982
rect 13484 1358 13518 1374
rect 13484 966 13518 982
rect 13602 1358 13636 1374
rect 13602 966 13636 982
rect 12937 898 12953 932
rect 12987 898 13003 932
rect 13055 898 13071 932
rect 13105 898 13121 932
rect 13173 898 13189 932
rect 13223 898 13239 932
rect 13291 898 13307 932
rect 13341 898 13357 932
rect 13409 898 13425 932
rect 13459 898 13475 932
rect 13527 898 13543 932
rect 13577 898 13593 932
rect 12780 830 12814 892
rect 13716 830 13750 892
rect 12780 796 12876 830
rect 13654 796 13750 830
rect 13820 1510 13916 1544
rect 14694 1510 14790 1544
rect 13820 1448 13854 1510
rect 14756 1448 14790 1510
rect 13977 1408 13993 1442
rect 14027 1408 14043 1442
rect 14095 1408 14111 1442
rect 14145 1408 14161 1442
rect 14213 1408 14229 1442
rect 14263 1408 14279 1442
rect 14331 1408 14347 1442
rect 14381 1408 14397 1442
rect 14449 1408 14465 1442
rect 14499 1408 14515 1442
rect 14567 1408 14583 1442
rect 14617 1408 14633 1442
rect 13934 1358 13968 1374
rect 13934 966 13968 982
rect 14052 1358 14086 1374
rect 14052 966 14086 982
rect 14170 1358 14204 1374
rect 14170 966 14204 982
rect 14288 1358 14322 1374
rect 14288 966 14322 982
rect 14406 1358 14440 1374
rect 14406 966 14440 982
rect 14524 1358 14558 1374
rect 14524 966 14558 982
rect 14642 1358 14676 1374
rect 14642 966 14676 982
rect 13977 898 13993 932
rect 14027 898 14043 932
rect 14095 898 14111 932
rect 14145 898 14161 932
rect 14213 898 14229 932
rect 14263 898 14279 932
rect 14331 898 14347 932
rect 14381 898 14397 932
rect 14449 898 14465 932
rect 14499 898 14515 932
rect 14567 898 14583 932
rect 14617 898 14633 932
rect 13820 830 13854 892
rect 14756 830 14790 892
rect 13820 796 13916 830
rect 14694 796 14790 830
rect 14860 1510 14956 1544
rect 15734 1510 15830 1544
rect 14860 1448 14894 1510
rect 15796 1448 15830 1510
rect 15017 1408 15033 1442
rect 15067 1408 15083 1442
rect 15135 1408 15151 1442
rect 15185 1408 15201 1442
rect 15253 1408 15269 1442
rect 15303 1408 15319 1442
rect 15371 1408 15387 1442
rect 15421 1408 15437 1442
rect 15489 1408 15505 1442
rect 15539 1408 15555 1442
rect 15607 1408 15623 1442
rect 15657 1408 15673 1442
rect 14974 1358 15008 1374
rect 14974 966 15008 982
rect 15092 1358 15126 1374
rect 15092 966 15126 982
rect 15210 1358 15244 1374
rect 15210 966 15244 982
rect 15328 1358 15362 1374
rect 15328 966 15362 982
rect 15446 1358 15480 1374
rect 15446 966 15480 982
rect 15564 1358 15598 1374
rect 15564 966 15598 982
rect 15682 1358 15716 1374
rect 15682 966 15716 982
rect 15017 898 15033 932
rect 15067 898 15083 932
rect 15135 898 15151 932
rect 15185 898 15201 932
rect 15253 898 15269 932
rect 15303 898 15319 932
rect 15371 898 15387 932
rect 15421 898 15437 932
rect 15489 898 15505 932
rect 15539 898 15555 932
rect 15607 898 15623 932
rect 15657 898 15673 932
rect 14860 830 14894 892
rect 15796 830 15830 892
rect 14860 796 14956 830
rect 15734 796 15830 830
rect 15900 1510 15996 1544
rect 16774 1510 16870 1544
rect 15900 1448 15934 1510
rect 16836 1448 16870 1510
rect 16057 1408 16073 1442
rect 16107 1408 16123 1442
rect 16175 1408 16191 1442
rect 16225 1408 16241 1442
rect 16293 1408 16309 1442
rect 16343 1408 16359 1442
rect 16411 1408 16427 1442
rect 16461 1408 16477 1442
rect 16529 1408 16545 1442
rect 16579 1408 16595 1442
rect 16647 1408 16663 1442
rect 16697 1408 16713 1442
rect 16014 1358 16048 1374
rect 16014 966 16048 982
rect 16132 1358 16166 1374
rect 16132 966 16166 982
rect 16250 1358 16284 1374
rect 16250 966 16284 982
rect 16368 1358 16402 1374
rect 16368 966 16402 982
rect 16486 1358 16520 1374
rect 16486 966 16520 982
rect 16604 1358 16638 1374
rect 16604 966 16638 982
rect 16722 1358 16756 1374
rect 16722 966 16756 982
rect 16057 898 16073 932
rect 16107 898 16123 932
rect 16175 898 16191 932
rect 16225 898 16241 932
rect 16293 898 16309 932
rect 16343 898 16359 932
rect 16411 898 16427 932
rect 16461 898 16477 932
rect 16529 898 16545 932
rect 16579 898 16595 932
rect 16647 898 16663 932
rect 16697 898 16713 932
rect 15900 830 15934 892
rect 16836 830 16870 892
rect 15900 796 15996 830
rect 16774 796 16870 830
rect 16940 1510 17036 1544
rect 17814 1510 17910 1544
rect 16940 1448 16974 1510
rect 17876 1448 17910 1510
rect 17097 1408 17113 1442
rect 17147 1408 17163 1442
rect 17215 1408 17231 1442
rect 17265 1408 17281 1442
rect 17333 1408 17349 1442
rect 17383 1408 17399 1442
rect 17451 1408 17467 1442
rect 17501 1408 17517 1442
rect 17569 1408 17585 1442
rect 17619 1408 17635 1442
rect 17687 1408 17703 1442
rect 17737 1408 17753 1442
rect 17054 1358 17088 1374
rect 17054 966 17088 982
rect 17172 1358 17206 1374
rect 17172 966 17206 982
rect 17290 1358 17324 1374
rect 17290 966 17324 982
rect 17408 1358 17442 1374
rect 17408 966 17442 982
rect 17526 1358 17560 1374
rect 17526 966 17560 982
rect 17644 1358 17678 1374
rect 17644 966 17678 982
rect 17762 1358 17796 1374
rect 17762 966 17796 982
rect 17097 898 17113 932
rect 17147 898 17163 932
rect 17215 898 17231 932
rect 17265 898 17281 932
rect 17333 898 17349 932
rect 17383 898 17399 932
rect 17451 898 17467 932
rect 17501 898 17517 932
rect 17569 898 17585 932
rect 17619 898 17635 932
rect 17687 898 17703 932
rect 17737 898 17753 932
rect 16940 830 16974 892
rect 17876 830 17910 892
rect 16940 796 17036 830
rect 17814 796 17910 830
rect 17980 1510 18076 1544
rect 18854 1510 18950 1544
rect 17980 1448 18014 1510
rect 18916 1448 18950 1510
rect 18137 1408 18153 1442
rect 18187 1408 18203 1442
rect 18255 1408 18271 1442
rect 18305 1408 18321 1442
rect 18373 1408 18389 1442
rect 18423 1408 18439 1442
rect 18491 1408 18507 1442
rect 18541 1408 18557 1442
rect 18609 1408 18625 1442
rect 18659 1408 18675 1442
rect 18727 1408 18743 1442
rect 18777 1408 18793 1442
rect 18094 1358 18128 1374
rect 18094 966 18128 982
rect 18212 1358 18246 1374
rect 18212 966 18246 982
rect 18330 1358 18364 1374
rect 18330 966 18364 982
rect 18448 1358 18482 1374
rect 18448 966 18482 982
rect 18566 1358 18600 1374
rect 18566 966 18600 982
rect 18684 1358 18718 1374
rect 18684 966 18718 982
rect 18802 1358 18836 1374
rect 18802 966 18836 982
rect 18137 898 18153 932
rect 18187 898 18203 932
rect 18255 898 18271 932
rect 18305 898 18321 932
rect 18373 898 18389 932
rect 18423 898 18439 932
rect 18491 898 18507 932
rect 18541 898 18557 932
rect 18609 898 18625 932
rect 18659 898 18675 932
rect 18727 898 18743 932
rect 18777 898 18793 932
rect 17980 830 18014 892
rect 18916 830 18950 892
rect 17980 796 18076 830
rect 18854 796 18950 830
rect 3412 670 3446 732
rect 4124 726 4944 796
rect 5184 726 5984 796
rect 6224 726 6964 796
rect 7264 726 8004 796
rect 8304 726 9024 796
rect 9344 726 10064 796
rect 11744 726 12564 796
rect 12804 726 13604 796
rect 13844 726 14584 796
rect 14884 726 15624 796
rect 15924 726 16644 796
rect 16964 726 17684 796
rect 1436 636 1532 670
rect 2310 636 2572 670
rect 3350 636 3446 670
rect 4120 692 4216 726
rect 4862 692 4958 726
rect -1688 540 1356 636
rect -1376 476 -1072 540
rect -1376 412 -1308 476
rect -1128 412 -1072 476
rect -1376 400 -1072 412
rect 2764 492 3132 636
rect 2764 408 2800 492
rect 3068 408 3132 492
rect 4120 630 4154 692
rect -6302 120 -6150 122
rect -7514 86 -7418 120
rect -6388 106 -6150 120
rect -6388 86 -6078 106
rect -7514 24 -7480 86
rect -6326 72 -6078 86
rect -5722 72 -5626 106
rect -6326 24 -6140 72
rect -7368 -16 -7352 18
rect -7318 -16 -7302 18
rect -7176 -16 -7160 18
rect -7126 -16 -7110 18
rect -6984 -16 -6968 18
rect -6934 -16 -6918 18
rect -6792 -16 -6776 18
rect -6742 -16 -6726 18
rect -6600 -16 -6584 18
rect -6550 -16 -6534 18
rect -7400 -66 -7366 -50
rect -7400 -458 -7366 -442
rect -7304 -66 -7270 -50
rect -7304 -458 -7270 -442
rect -7208 -66 -7174 -50
rect -7208 -458 -7174 -442
rect -7112 -66 -7078 -50
rect -7112 -458 -7078 -442
rect -7016 -66 -6982 -50
rect -7016 -458 -6982 -442
rect -6920 -66 -6886 -50
rect -6920 -458 -6886 -442
rect -6824 -66 -6790 -50
rect -6824 -458 -6790 -442
rect -6728 -66 -6694 -50
rect -6728 -458 -6694 -442
rect -6632 -66 -6598 -50
rect -6632 -458 -6598 -442
rect -6536 -66 -6502 -50
rect -6536 -458 -6502 -442
rect -6440 -66 -6406 -50
rect -6440 -458 -6406 -442
rect -7272 -526 -7256 -492
rect -7222 -526 -7206 -492
rect -7080 -526 -7064 -492
rect -7030 -526 -7014 -492
rect -6888 -526 -6872 -492
rect -6838 -526 -6822 -492
rect -6696 -526 -6680 -492
rect -6646 -526 -6630 -492
rect -6504 -526 -6488 -492
rect -6454 -526 -6438 -492
rect -7272 -634 -7256 -600
rect -7222 -634 -7206 -600
rect -7080 -634 -7064 -600
rect -7030 -634 -7014 -600
rect -6888 -634 -6872 -600
rect -6838 -634 -6822 -600
rect -6696 -634 -6680 -600
rect -6646 -634 -6630 -600
rect -6504 -634 -6488 -600
rect -6454 -634 -6438 -600
rect -7400 -684 -7366 -668
rect -7400 -1076 -7366 -1060
rect -7304 -684 -7270 -668
rect -7304 -1076 -7270 -1060
rect -7208 -684 -7174 -668
rect -7208 -1076 -7174 -1060
rect -7112 -684 -7078 -668
rect -7112 -1076 -7078 -1060
rect -7016 -684 -6982 -668
rect -7016 -1076 -6982 -1060
rect -6920 -684 -6886 -668
rect -6920 -1076 -6886 -1060
rect -6824 -684 -6790 -668
rect -6824 -1076 -6790 -1060
rect -6728 -684 -6694 -668
rect -6728 -1076 -6694 -1060
rect -6632 -684 -6598 -668
rect -6632 -1076 -6598 -1060
rect -6536 -684 -6502 -668
rect -6536 -1076 -6502 -1060
rect -6440 -684 -6406 -668
rect -6440 -1076 -6406 -1060
rect -7368 -1144 -7352 -1110
rect -7318 -1144 -7302 -1110
rect -7176 -1144 -7160 -1110
rect -7126 -1144 -7110 -1110
rect -6984 -1144 -6968 -1110
rect -6934 -1144 -6918 -1110
rect -6792 -1144 -6776 -1110
rect -6742 -1144 -6726 -1110
rect -6600 -1144 -6584 -1110
rect -6550 -1144 -6534 -1110
rect -7514 -1212 -7480 -1150
rect -6292 10 -6140 24
rect -6292 -1150 -6174 10
rect -6326 -1212 -6174 -1150
rect -7514 -1246 -7418 -1212
rect -6388 -1246 -6174 -1212
rect -7514 -1750 -7418 -1716
rect -6772 -1750 -6676 -1716
rect -7514 -1812 -7480 -1750
rect -6710 -1812 -6676 -1750
rect -7368 -1852 -7352 -1818
rect -7318 -1852 -7302 -1818
rect -7176 -1852 -7160 -1818
rect -7126 -1852 -7110 -1818
rect -6984 -1852 -6968 -1818
rect -6934 -1852 -6918 -1818
rect -7400 -1902 -7366 -1886
rect -7400 -2294 -7366 -2278
rect -7304 -1902 -7270 -1886
rect -7304 -2294 -7270 -2278
rect -7208 -1902 -7174 -1886
rect -7208 -2294 -7174 -2278
rect -7112 -1902 -7078 -1886
rect -7112 -2294 -7078 -2278
rect -7016 -1902 -6982 -1886
rect -7016 -2294 -6982 -2278
rect -6920 -1902 -6886 -1886
rect -6920 -2294 -6886 -2278
rect -6824 -1902 -6790 -1886
rect -6824 -2294 -6790 -2278
rect -7272 -2362 -7256 -2328
rect -7222 -2362 -7206 -2328
rect -7080 -2362 -7064 -2328
rect -7030 -2362 -7014 -2328
rect -6888 -2362 -6872 -2328
rect -6838 -2362 -6822 -2328
rect -7272 -2470 -7256 -2436
rect -7222 -2470 -7206 -2436
rect -7080 -2470 -7064 -2436
rect -7030 -2470 -7014 -2436
rect -6888 -2470 -6872 -2436
rect -6838 -2470 -6822 -2436
rect -7400 -2520 -7366 -2504
rect -7400 -2912 -7366 -2896
rect -7304 -2520 -7270 -2504
rect -7304 -2912 -7270 -2896
rect -7208 -2520 -7174 -2504
rect -7208 -2912 -7174 -2896
rect -7112 -2520 -7078 -2504
rect -7112 -2912 -7078 -2896
rect -7016 -2520 -6982 -2504
rect -7016 -2912 -6982 -2896
rect -6920 -2520 -6886 -2504
rect -6920 -2912 -6886 -2896
rect -6824 -2520 -6790 -2504
rect -6824 -2912 -6790 -2896
rect -7368 -2980 -7352 -2946
rect -7318 -2980 -7302 -2946
rect -7176 -2980 -7160 -2946
rect -7126 -2980 -7110 -2946
rect -6984 -2980 -6968 -2946
rect -6934 -2980 -6918 -2946
rect -7514 -3048 -7480 -2986
rect -6310 -1718 -6174 -1246
rect -5660 10 -5626 72
rect -6004 -42 -5988 -8
rect -5812 -42 -5796 -8
rect -6072 -70 -6038 -54
rect -6140 -1718 -6134 -1226
rect -6072 -1654 -6038 -1638
rect -5762 -70 -5728 -54
rect -5762 -1654 -5728 -1638
rect -6004 -1700 -5988 -1666
rect -5812 -1700 -5796 -1666
rect -6310 -1754 -6134 -1718
rect 4924 630 4958 692
rect 4266 590 4282 624
rect 4316 590 4332 624
rect 4458 590 4474 624
rect 4508 590 4524 624
rect 4650 590 4666 624
rect 4700 590 4716 624
rect 4234 540 4268 556
rect 4234 148 4268 164
rect 4330 540 4364 556
rect 4330 148 4364 164
rect 4426 540 4460 556
rect 4426 148 4460 164
rect 4522 540 4556 556
rect 4522 148 4556 164
rect 4618 540 4652 556
rect 4618 148 4652 164
rect 4714 540 4748 556
rect 4714 148 4748 164
rect 4810 540 4844 556
rect 4810 148 4844 164
rect 4362 80 4378 114
rect 4412 80 4428 114
rect 4554 80 4570 114
rect 4604 80 4620 114
rect 4746 80 4762 114
rect 4796 80 4812 114
rect 4362 -28 4378 6
rect 4412 -28 4428 6
rect 4554 -28 4570 6
rect 4604 -28 4620 6
rect 4746 -28 4762 6
rect 4796 -28 4812 6
rect 4234 -78 4268 -62
rect 4234 -470 4268 -454
rect 4330 -78 4364 -62
rect 4330 -470 4364 -454
rect 4426 -78 4460 -62
rect 4426 -470 4460 -454
rect 4522 -78 4556 -62
rect 4522 -470 4556 -454
rect 4618 -78 4652 -62
rect 4618 -470 4652 -454
rect 4714 -78 4748 -62
rect 4714 -470 4748 -454
rect 4810 -78 4844 -62
rect 4810 -470 4844 -454
rect 4266 -538 4282 -504
rect 4316 -538 4332 -504
rect 4458 -538 4474 -504
rect 4508 -538 4524 -504
rect 4650 -538 4666 -504
rect 4700 -538 4716 -504
rect 4120 -606 4154 -544
rect 4924 -606 4958 -544
rect 4120 -640 4216 -606
rect 4862 -628 4958 -606
rect 5160 692 5256 726
rect 5902 692 5998 726
rect 5160 630 5194 692
rect 5964 630 5998 692
rect 5306 590 5322 624
rect 5356 590 5372 624
rect 5498 590 5514 624
rect 5548 590 5564 624
rect 5690 590 5706 624
rect 5740 590 5756 624
rect 5274 540 5308 556
rect 5274 148 5308 164
rect 5370 540 5404 556
rect 5370 148 5404 164
rect 5466 540 5500 556
rect 5466 148 5500 164
rect 5562 540 5596 556
rect 5562 148 5596 164
rect 5658 540 5692 556
rect 5658 148 5692 164
rect 5754 540 5788 556
rect 5754 148 5788 164
rect 5850 540 5884 556
rect 5850 148 5884 164
rect 5402 80 5418 114
rect 5452 80 5468 114
rect 5594 80 5610 114
rect 5644 80 5660 114
rect 5786 80 5802 114
rect 5836 80 5852 114
rect 5402 -28 5418 6
rect 5452 -28 5468 6
rect 5594 -28 5610 6
rect 5644 -28 5660 6
rect 5786 -28 5802 6
rect 5836 -28 5852 6
rect 5274 -78 5308 -62
rect 5274 -470 5308 -454
rect 5370 -78 5404 -62
rect 5370 -470 5404 -454
rect 5466 -78 5500 -62
rect 5466 -470 5500 -454
rect 5562 -78 5596 -62
rect 5562 -470 5596 -454
rect 5658 -78 5692 -62
rect 5658 -470 5692 -454
rect 5754 -78 5788 -62
rect 5754 -470 5788 -454
rect 5850 -78 5884 -62
rect 5850 -470 5884 -454
rect 5306 -538 5322 -504
rect 5356 -538 5372 -504
rect 5498 -538 5514 -504
rect 5548 -538 5564 -504
rect 5690 -538 5706 -504
rect 5740 -538 5756 -504
rect 5160 -606 5194 -544
rect 5964 -606 5998 -544
rect 4862 -640 4960 -628
rect 4120 -696 4960 -640
rect 5160 -640 5256 -606
rect 5902 -628 5998 -606
rect 6200 692 6296 726
rect 6942 692 7038 726
rect 6200 630 6234 692
rect 7004 630 7038 692
rect 6346 590 6362 624
rect 6396 590 6412 624
rect 6538 590 6554 624
rect 6588 590 6604 624
rect 6730 590 6746 624
rect 6780 590 6796 624
rect 6314 540 6348 556
rect 6314 148 6348 164
rect 6410 540 6444 556
rect 6410 148 6444 164
rect 6506 540 6540 556
rect 6506 148 6540 164
rect 6602 540 6636 556
rect 6602 148 6636 164
rect 6698 540 6732 556
rect 6698 148 6732 164
rect 6794 540 6828 556
rect 6794 148 6828 164
rect 6890 540 6924 556
rect 6890 148 6924 164
rect 6442 80 6458 114
rect 6492 80 6508 114
rect 6634 80 6650 114
rect 6684 80 6700 114
rect 6826 80 6842 114
rect 6876 80 6892 114
rect 6442 -28 6458 6
rect 6492 -28 6508 6
rect 6634 -28 6650 6
rect 6684 -28 6700 6
rect 6826 -28 6842 6
rect 6876 -28 6892 6
rect 6314 -78 6348 -62
rect 6314 -470 6348 -454
rect 6410 -78 6444 -62
rect 6410 -470 6444 -454
rect 6506 -78 6540 -62
rect 6506 -470 6540 -454
rect 6602 -78 6636 -62
rect 6602 -470 6636 -454
rect 6698 -78 6732 -62
rect 6698 -470 6732 -454
rect 6794 -78 6828 -62
rect 6794 -470 6828 -454
rect 6890 -78 6924 -62
rect 6890 -470 6924 -454
rect 6346 -538 6362 -504
rect 6396 -538 6412 -504
rect 6538 -538 6554 -504
rect 6588 -538 6604 -504
rect 6730 -538 6746 -504
rect 6780 -538 6796 -504
rect 6200 -606 6234 -544
rect 7004 -606 7038 -544
rect 5902 -640 6000 -628
rect 5160 -696 6000 -640
rect 6200 -640 6296 -606
rect 6942 -628 7038 -606
rect 7240 692 7336 726
rect 7982 692 8078 726
rect 7240 630 7274 692
rect 8044 630 8078 692
rect 7386 590 7402 624
rect 7436 590 7452 624
rect 7578 590 7594 624
rect 7628 590 7644 624
rect 7770 590 7786 624
rect 7820 590 7836 624
rect 7354 540 7388 556
rect 7354 148 7388 164
rect 7450 540 7484 556
rect 7450 148 7484 164
rect 7546 540 7580 556
rect 7546 148 7580 164
rect 7642 540 7676 556
rect 7642 148 7676 164
rect 7738 540 7772 556
rect 7738 148 7772 164
rect 7834 540 7868 556
rect 7834 148 7868 164
rect 7930 540 7964 556
rect 7930 148 7964 164
rect 7482 80 7498 114
rect 7532 80 7548 114
rect 7674 80 7690 114
rect 7724 80 7740 114
rect 7866 80 7882 114
rect 7916 80 7932 114
rect 7482 -28 7498 6
rect 7532 -28 7548 6
rect 7674 -28 7690 6
rect 7724 -28 7740 6
rect 7866 -28 7882 6
rect 7916 -28 7932 6
rect 7354 -78 7388 -62
rect 7354 -470 7388 -454
rect 7450 -78 7484 -62
rect 7450 -470 7484 -454
rect 7546 -78 7580 -62
rect 7546 -470 7580 -454
rect 7642 -78 7676 -62
rect 7642 -470 7676 -454
rect 7738 -78 7772 -62
rect 7738 -470 7772 -454
rect 7834 -78 7868 -62
rect 7834 -470 7868 -454
rect 7930 -78 7964 -62
rect 7930 -470 7964 -454
rect 7386 -538 7402 -504
rect 7436 -538 7452 -504
rect 7578 -538 7594 -504
rect 7628 -538 7644 -504
rect 7770 -538 7786 -504
rect 7820 -538 7836 -504
rect 7240 -606 7274 -544
rect 8044 -606 8078 -544
rect 6942 -640 7040 -628
rect 6200 -696 7040 -640
rect 7240 -640 7336 -606
rect 7982 -628 8078 -606
rect 8280 692 8376 726
rect 9022 692 9118 726
rect 8280 630 8314 692
rect 9084 630 9118 692
rect 8426 590 8442 624
rect 8476 590 8492 624
rect 8618 590 8634 624
rect 8668 590 8684 624
rect 8810 590 8826 624
rect 8860 590 8876 624
rect 8394 540 8428 556
rect 8394 148 8428 164
rect 8490 540 8524 556
rect 8490 148 8524 164
rect 8586 540 8620 556
rect 8586 148 8620 164
rect 8682 540 8716 556
rect 8682 148 8716 164
rect 8778 540 8812 556
rect 8778 148 8812 164
rect 8874 540 8908 556
rect 8874 148 8908 164
rect 8970 540 9004 556
rect 8970 148 9004 164
rect 8522 80 8538 114
rect 8572 80 8588 114
rect 8714 80 8730 114
rect 8764 80 8780 114
rect 8906 80 8922 114
rect 8956 80 8972 114
rect 8522 -28 8538 6
rect 8572 -28 8588 6
rect 8714 -28 8730 6
rect 8764 -28 8780 6
rect 8906 -28 8922 6
rect 8956 -28 8972 6
rect 8394 -78 8428 -62
rect 8394 -470 8428 -454
rect 8490 -78 8524 -62
rect 8490 -470 8524 -454
rect 8586 -78 8620 -62
rect 8586 -470 8620 -454
rect 8682 -78 8716 -62
rect 8682 -470 8716 -454
rect 8778 -78 8812 -62
rect 8778 -470 8812 -454
rect 8874 -78 8908 -62
rect 8874 -470 8908 -454
rect 8970 -78 9004 -62
rect 8970 -470 9004 -454
rect 8426 -538 8442 -504
rect 8476 -538 8492 -504
rect 8618 -538 8634 -504
rect 8668 -538 8684 -504
rect 8810 -538 8826 -504
rect 8860 -538 8876 -504
rect 8280 -606 8314 -544
rect 9084 -606 9118 -544
rect 7982 -640 8080 -628
rect 7240 -696 8080 -640
rect 8280 -640 8376 -606
rect 9022 -628 9118 -606
rect 9320 692 9416 726
rect 10062 692 10158 726
rect 9320 630 9354 692
rect 10124 630 10158 692
rect 9466 590 9482 624
rect 9516 590 9532 624
rect 9658 590 9674 624
rect 9708 590 9724 624
rect 9850 590 9866 624
rect 9900 590 9916 624
rect 9434 540 9468 556
rect 9434 148 9468 164
rect 9530 540 9564 556
rect 9530 148 9564 164
rect 9626 540 9660 556
rect 9626 148 9660 164
rect 9722 540 9756 556
rect 9722 148 9756 164
rect 9818 540 9852 556
rect 9818 148 9852 164
rect 9914 540 9948 556
rect 9914 148 9948 164
rect 10010 540 10044 556
rect 10010 148 10044 164
rect 9562 80 9578 114
rect 9612 80 9628 114
rect 9754 80 9770 114
rect 9804 80 9820 114
rect 9946 80 9962 114
rect 9996 80 10012 114
rect 9562 -28 9578 6
rect 9612 -28 9628 6
rect 9754 -28 9770 6
rect 9804 -28 9820 6
rect 9946 -28 9962 6
rect 9996 -28 10012 6
rect 9434 -78 9468 -62
rect 9434 -470 9468 -454
rect 9530 -78 9564 -62
rect 9530 -470 9564 -454
rect 9626 -78 9660 -62
rect 9626 -470 9660 -454
rect 9722 -78 9756 -62
rect 9722 -470 9756 -454
rect 9818 -78 9852 -62
rect 9818 -470 9852 -454
rect 9914 -78 9948 -62
rect 9914 -470 9948 -454
rect 10010 -78 10044 -62
rect 10010 -470 10044 -454
rect 9466 -538 9482 -504
rect 9516 -538 9532 -504
rect 9658 -538 9674 -504
rect 9708 -538 9724 -504
rect 9850 -538 9866 -504
rect 9900 -538 9916 -504
rect 9320 -606 9354 -544
rect 10124 -606 10158 -544
rect 9022 -640 9120 -628
rect 8280 -696 9120 -640
rect 9320 -640 9416 -606
rect 10062 -628 10158 -606
rect 10360 692 10456 726
rect 11102 692 11198 726
rect 10360 630 10394 692
rect 11164 630 11198 692
rect 10506 590 10522 624
rect 10556 590 10572 624
rect 10698 590 10714 624
rect 10748 590 10764 624
rect 10890 590 10906 624
rect 10940 590 10956 624
rect 10474 540 10508 556
rect 10474 148 10508 164
rect 10570 540 10604 556
rect 10570 148 10604 164
rect 10666 540 10700 556
rect 10666 148 10700 164
rect 10762 540 10796 556
rect 10762 148 10796 164
rect 10858 540 10892 556
rect 10858 148 10892 164
rect 10954 540 10988 556
rect 10954 148 10988 164
rect 11050 540 11084 556
rect 11050 148 11084 164
rect 10602 80 10618 114
rect 10652 80 10668 114
rect 10794 80 10810 114
rect 10844 80 10860 114
rect 10986 80 11002 114
rect 11036 80 11052 114
rect 10602 -28 10618 6
rect 10652 -28 10668 6
rect 10794 -28 10810 6
rect 10844 -28 10860 6
rect 10986 -28 11002 6
rect 11036 -28 11052 6
rect 10474 -78 10508 -62
rect 10474 -470 10508 -454
rect 10570 -78 10604 -62
rect 10570 -470 10604 -454
rect 10666 -78 10700 -62
rect 10666 -470 10700 -454
rect 10762 -78 10796 -62
rect 10762 -470 10796 -454
rect 10858 -78 10892 -62
rect 10858 -470 10892 -454
rect 10954 -78 10988 -62
rect 10954 -470 10988 -454
rect 11050 -78 11084 -62
rect 11050 -470 11084 -454
rect 10506 -538 10522 -504
rect 10556 -538 10572 -504
rect 10698 -538 10714 -504
rect 10748 -538 10764 -504
rect 10890 -538 10906 -504
rect 10940 -538 10956 -504
rect 10360 -606 10394 -544
rect 11164 -606 11198 -544
rect 10062 -640 10160 -628
rect 9320 -696 10160 -640
rect 10360 -640 10456 -606
rect 11102 -628 11198 -606
rect 11740 692 11836 726
rect 12482 692 12578 726
rect 11740 630 11774 692
rect 12544 630 12578 692
rect 11886 590 11902 624
rect 11936 590 11952 624
rect 12078 590 12094 624
rect 12128 590 12144 624
rect 12270 590 12286 624
rect 12320 590 12336 624
rect 11854 540 11888 556
rect 11854 148 11888 164
rect 11950 540 11984 556
rect 11950 148 11984 164
rect 12046 540 12080 556
rect 12046 148 12080 164
rect 12142 540 12176 556
rect 12142 148 12176 164
rect 12238 540 12272 556
rect 12238 148 12272 164
rect 12334 540 12368 556
rect 12334 148 12368 164
rect 12430 540 12464 556
rect 12430 148 12464 164
rect 11982 80 11998 114
rect 12032 80 12048 114
rect 12174 80 12190 114
rect 12224 80 12240 114
rect 12366 80 12382 114
rect 12416 80 12432 114
rect 11982 -28 11998 6
rect 12032 -28 12048 6
rect 12174 -28 12190 6
rect 12224 -28 12240 6
rect 12366 -28 12382 6
rect 12416 -28 12432 6
rect 11854 -78 11888 -62
rect 11854 -470 11888 -454
rect 11950 -78 11984 -62
rect 11950 -470 11984 -454
rect 12046 -78 12080 -62
rect 12046 -470 12080 -454
rect 12142 -78 12176 -62
rect 12142 -470 12176 -454
rect 12238 -78 12272 -62
rect 12238 -470 12272 -454
rect 12334 -78 12368 -62
rect 12334 -470 12368 -454
rect 12430 -78 12464 -62
rect 12430 -470 12464 -454
rect 11886 -538 11902 -504
rect 11936 -538 11952 -504
rect 12078 -538 12094 -504
rect 12128 -538 12144 -504
rect 12270 -538 12286 -504
rect 12320 -538 12336 -504
rect 11740 -606 11774 -544
rect 12544 -606 12578 -544
rect 11102 -640 11200 -628
rect 10360 -696 11200 -640
rect 11740 -640 11836 -606
rect 12482 -628 12578 -606
rect 12780 692 12876 726
rect 13522 692 13618 726
rect 12780 630 12814 692
rect 13584 630 13618 692
rect 12926 590 12942 624
rect 12976 590 12992 624
rect 13118 590 13134 624
rect 13168 590 13184 624
rect 13310 590 13326 624
rect 13360 590 13376 624
rect 12894 540 12928 556
rect 12894 148 12928 164
rect 12990 540 13024 556
rect 12990 148 13024 164
rect 13086 540 13120 556
rect 13086 148 13120 164
rect 13182 540 13216 556
rect 13182 148 13216 164
rect 13278 540 13312 556
rect 13278 148 13312 164
rect 13374 540 13408 556
rect 13374 148 13408 164
rect 13470 540 13504 556
rect 13470 148 13504 164
rect 13022 80 13038 114
rect 13072 80 13088 114
rect 13214 80 13230 114
rect 13264 80 13280 114
rect 13406 80 13422 114
rect 13456 80 13472 114
rect 13022 -28 13038 6
rect 13072 -28 13088 6
rect 13214 -28 13230 6
rect 13264 -28 13280 6
rect 13406 -28 13422 6
rect 13456 -28 13472 6
rect 12894 -78 12928 -62
rect 12894 -470 12928 -454
rect 12990 -78 13024 -62
rect 12990 -470 13024 -454
rect 13086 -78 13120 -62
rect 13086 -470 13120 -454
rect 13182 -78 13216 -62
rect 13182 -470 13216 -454
rect 13278 -78 13312 -62
rect 13278 -470 13312 -454
rect 13374 -78 13408 -62
rect 13374 -470 13408 -454
rect 13470 -78 13504 -62
rect 13470 -470 13504 -454
rect 12926 -538 12942 -504
rect 12976 -538 12992 -504
rect 13118 -538 13134 -504
rect 13168 -538 13184 -504
rect 13310 -538 13326 -504
rect 13360 -538 13376 -504
rect 12780 -606 12814 -544
rect 13584 -606 13618 -544
rect 12482 -640 12580 -628
rect 11740 -696 12580 -640
rect 12780 -640 12876 -606
rect 13522 -628 13618 -606
rect 13820 692 13916 726
rect 14562 692 14658 726
rect 13820 630 13854 692
rect 14624 630 14658 692
rect 13966 590 13982 624
rect 14016 590 14032 624
rect 14158 590 14174 624
rect 14208 590 14224 624
rect 14350 590 14366 624
rect 14400 590 14416 624
rect 13934 540 13968 556
rect 13934 148 13968 164
rect 14030 540 14064 556
rect 14030 148 14064 164
rect 14126 540 14160 556
rect 14126 148 14160 164
rect 14222 540 14256 556
rect 14222 148 14256 164
rect 14318 540 14352 556
rect 14318 148 14352 164
rect 14414 540 14448 556
rect 14414 148 14448 164
rect 14510 540 14544 556
rect 14510 148 14544 164
rect 14062 80 14078 114
rect 14112 80 14128 114
rect 14254 80 14270 114
rect 14304 80 14320 114
rect 14446 80 14462 114
rect 14496 80 14512 114
rect 14062 -28 14078 6
rect 14112 -28 14128 6
rect 14254 -28 14270 6
rect 14304 -28 14320 6
rect 14446 -28 14462 6
rect 14496 -28 14512 6
rect 13934 -78 13968 -62
rect 13934 -470 13968 -454
rect 14030 -78 14064 -62
rect 14030 -470 14064 -454
rect 14126 -78 14160 -62
rect 14126 -470 14160 -454
rect 14222 -78 14256 -62
rect 14222 -470 14256 -454
rect 14318 -78 14352 -62
rect 14318 -470 14352 -454
rect 14414 -78 14448 -62
rect 14414 -470 14448 -454
rect 14510 -78 14544 -62
rect 14510 -470 14544 -454
rect 13966 -538 13982 -504
rect 14016 -538 14032 -504
rect 14158 -538 14174 -504
rect 14208 -538 14224 -504
rect 14350 -538 14366 -504
rect 14400 -538 14416 -504
rect 13820 -606 13854 -544
rect 14624 -606 14658 -544
rect 13522 -640 13620 -628
rect 12780 -696 13620 -640
rect 13820 -640 13916 -606
rect 14562 -628 14658 -606
rect 14860 692 14956 726
rect 15602 692 15698 726
rect 14860 630 14894 692
rect 15664 630 15698 692
rect 15006 590 15022 624
rect 15056 590 15072 624
rect 15198 590 15214 624
rect 15248 590 15264 624
rect 15390 590 15406 624
rect 15440 590 15456 624
rect 14974 540 15008 556
rect 14974 148 15008 164
rect 15070 540 15104 556
rect 15070 148 15104 164
rect 15166 540 15200 556
rect 15166 148 15200 164
rect 15262 540 15296 556
rect 15262 148 15296 164
rect 15358 540 15392 556
rect 15358 148 15392 164
rect 15454 540 15488 556
rect 15454 148 15488 164
rect 15550 540 15584 556
rect 15550 148 15584 164
rect 15102 80 15118 114
rect 15152 80 15168 114
rect 15294 80 15310 114
rect 15344 80 15360 114
rect 15486 80 15502 114
rect 15536 80 15552 114
rect 15102 -28 15118 6
rect 15152 -28 15168 6
rect 15294 -28 15310 6
rect 15344 -28 15360 6
rect 15486 -28 15502 6
rect 15536 -28 15552 6
rect 14974 -78 15008 -62
rect 14974 -470 15008 -454
rect 15070 -78 15104 -62
rect 15070 -470 15104 -454
rect 15166 -78 15200 -62
rect 15166 -470 15200 -454
rect 15262 -78 15296 -62
rect 15262 -470 15296 -454
rect 15358 -78 15392 -62
rect 15358 -470 15392 -454
rect 15454 -78 15488 -62
rect 15454 -470 15488 -454
rect 15550 -78 15584 -62
rect 15550 -470 15584 -454
rect 15006 -538 15022 -504
rect 15056 -538 15072 -504
rect 15198 -538 15214 -504
rect 15248 -538 15264 -504
rect 15390 -538 15406 -504
rect 15440 -538 15456 -504
rect 14860 -606 14894 -544
rect 15664 -606 15698 -544
rect 14562 -640 14660 -628
rect 13820 -696 14660 -640
rect 14860 -640 14956 -606
rect 15602 -628 15698 -606
rect 15900 692 15996 726
rect 16642 692 16738 726
rect 15900 630 15934 692
rect 16704 630 16738 692
rect 16046 590 16062 624
rect 16096 590 16112 624
rect 16238 590 16254 624
rect 16288 590 16304 624
rect 16430 590 16446 624
rect 16480 590 16496 624
rect 16014 540 16048 556
rect 16014 148 16048 164
rect 16110 540 16144 556
rect 16110 148 16144 164
rect 16206 540 16240 556
rect 16206 148 16240 164
rect 16302 540 16336 556
rect 16302 148 16336 164
rect 16398 540 16432 556
rect 16398 148 16432 164
rect 16494 540 16528 556
rect 16494 148 16528 164
rect 16590 540 16624 556
rect 16590 148 16624 164
rect 16142 80 16158 114
rect 16192 80 16208 114
rect 16334 80 16350 114
rect 16384 80 16400 114
rect 16526 80 16542 114
rect 16576 80 16592 114
rect 16142 -28 16158 6
rect 16192 -28 16208 6
rect 16334 -28 16350 6
rect 16384 -28 16400 6
rect 16526 -28 16542 6
rect 16576 -28 16592 6
rect 16014 -78 16048 -62
rect 16014 -470 16048 -454
rect 16110 -78 16144 -62
rect 16110 -470 16144 -454
rect 16206 -78 16240 -62
rect 16206 -470 16240 -454
rect 16302 -78 16336 -62
rect 16302 -470 16336 -454
rect 16398 -78 16432 -62
rect 16398 -470 16432 -454
rect 16494 -78 16528 -62
rect 16494 -470 16528 -454
rect 16590 -78 16624 -62
rect 16590 -470 16624 -454
rect 16046 -538 16062 -504
rect 16096 -538 16112 -504
rect 16238 -538 16254 -504
rect 16288 -538 16304 -504
rect 16430 -538 16446 -504
rect 16480 -538 16496 -504
rect 15900 -606 15934 -544
rect 16704 -606 16738 -544
rect 15602 -640 15700 -628
rect 14860 -696 15700 -640
rect 15900 -640 15996 -606
rect 16642 -628 16738 -606
rect 16940 692 17036 726
rect 17682 692 17778 726
rect 16940 630 16974 692
rect 17744 630 17778 692
rect 17086 590 17102 624
rect 17136 590 17152 624
rect 17278 590 17294 624
rect 17328 590 17344 624
rect 17470 590 17486 624
rect 17520 590 17536 624
rect 17054 540 17088 556
rect 17054 148 17088 164
rect 17150 540 17184 556
rect 17150 148 17184 164
rect 17246 540 17280 556
rect 17246 148 17280 164
rect 17342 540 17376 556
rect 17342 148 17376 164
rect 17438 540 17472 556
rect 17438 148 17472 164
rect 17534 540 17568 556
rect 17534 148 17568 164
rect 17630 540 17664 556
rect 17630 148 17664 164
rect 17182 80 17198 114
rect 17232 80 17248 114
rect 17374 80 17390 114
rect 17424 80 17440 114
rect 17566 80 17582 114
rect 17616 80 17632 114
rect 17182 -28 17198 6
rect 17232 -28 17248 6
rect 17374 -28 17390 6
rect 17424 -28 17440 6
rect 17566 -28 17582 6
rect 17616 -28 17632 6
rect 17054 -78 17088 -62
rect 17054 -470 17088 -454
rect 17150 -78 17184 -62
rect 17150 -470 17184 -454
rect 17246 -78 17280 -62
rect 17246 -470 17280 -454
rect 17342 -78 17376 -62
rect 17342 -470 17376 -454
rect 17438 -78 17472 -62
rect 17438 -470 17472 -454
rect 17534 -78 17568 -62
rect 17534 -470 17568 -454
rect 17630 -78 17664 -62
rect 17630 -470 17664 -454
rect 17086 -538 17102 -504
rect 17136 -538 17152 -504
rect 17278 -538 17294 -504
rect 17328 -538 17344 -504
rect 17470 -538 17486 -504
rect 17520 -538 17536 -504
rect 16940 -606 16974 -544
rect 17744 -606 17778 -544
rect 16642 -640 16740 -628
rect 15900 -696 16740 -640
rect 16940 -640 17036 -606
rect 17682 -628 17778 -606
rect 17980 692 18076 726
rect 18722 692 18818 726
rect 17980 630 18014 692
rect 18784 630 18818 692
rect 18126 590 18142 624
rect 18176 590 18192 624
rect 18318 590 18334 624
rect 18368 590 18384 624
rect 18510 590 18526 624
rect 18560 590 18576 624
rect 18094 540 18128 556
rect 18094 148 18128 164
rect 18190 540 18224 556
rect 18190 148 18224 164
rect 18286 540 18320 556
rect 18286 148 18320 164
rect 18382 540 18416 556
rect 18382 148 18416 164
rect 18478 540 18512 556
rect 18478 148 18512 164
rect 18574 540 18608 556
rect 18574 148 18608 164
rect 18670 540 18704 556
rect 18670 148 18704 164
rect 18222 80 18238 114
rect 18272 80 18288 114
rect 18414 80 18430 114
rect 18464 80 18480 114
rect 18606 80 18622 114
rect 18656 80 18672 114
rect 18222 -28 18238 6
rect 18272 -28 18288 6
rect 18414 -28 18430 6
rect 18464 -28 18480 6
rect 18606 -28 18622 6
rect 18656 -28 18672 6
rect 18094 -78 18128 -62
rect 18094 -470 18128 -454
rect 18190 -78 18224 -62
rect 18190 -470 18224 -454
rect 18286 -78 18320 -62
rect 18286 -470 18320 -454
rect 18382 -78 18416 -62
rect 18382 -470 18416 -454
rect 18478 -78 18512 -62
rect 18478 -470 18512 -454
rect 18574 -78 18608 -62
rect 18574 -470 18608 -454
rect 18670 -78 18704 -62
rect 18670 -470 18704 -454
rect 18126 -538 18142 -504
rect 18176 -538 18192 -504
rect 18318 -538 18334 -504
rect 18368 -538 18384 -504
rect 18510 -538 18526 -504
rect 18560 -538 18576 -504
rect 17980 -606 18014 -544
rect 18784 -606 18818 -544
rect 17682 -640 17780 -628
rect 16940 -696 17780 -640
rect 17980 -640 18076 -606
rect 18722 -628 18818 -606
rect 18722 -640 18820 -628
rect 17980 -696 18820 -640
rect 4120 -730 4216 -696
rect 4994 -700 5090 -696
rect 5160 -700 5256 -696
rect 4994 -730 5256 -700
rect 6034 -700 6130 -696
rect 6200 -700 6296 -696
rect 6034 -730 6296 -700
rect 7074 -700 7170 -696
rect 7240 -700 7336 -696
rect 7074 -730 7336 -700
rect 8114 -700 8210 -696
rect 8280 -700 8376 -696
rect 8114 -730 8376 -700
rect 9154 -700 9250 -696
rect 9320 -700 9416 -696
rect 9154 -730 9416 -700
rect 10194 -730 10290 -696
rect 4120 -792 4154 -730
rect 5056 -792 5194 -730
rect 4277 -832 4293 -798
rect 4327 -832 4343 -798
rect 4395 -832 4411 -798
rect 4445 -832 4461 -798
rect 4513 -832 4529 -798
rect 4563 -832 4579 -798
rect 4631 -832 4647 -798
rect 4681 -832 4697 -798
rect 4749 -832 4765 -798
rect 4799 -832 4815 -798
rect 4867 -832 4883 -798
rect 4917 -832 4933 -798
rect 4234 -882 4268 -866
rect 4234 -1274 4268 -1258
rect 4352 -882 4386 -866
rect 4352 -1274 4386 -1258
rect 4470 -882 4504 -866
rect 4470 -1274 4504 -1258
rect 4588 -882 4622 -866
rect 4588 -1274 4622 -1258
rect 4706 -882 4740 -866
rect 4706 -1274 4740 -1258
rect 4824 -882 4858 -866
rect 4824 -1274 4858 -1258
rect 4942 -882 4976 -866
rect 4942 -1274 4976 -1258
rect 4277 -1342 4293 -1308
rect 4327 -1342 4343 -1308
rect 4395 -1342 4411 -1308
rect 4445 -1342 4461 -1308
rect 4513 -1342 4529 -1308
rect 4563 -1342 4579 -1308
rect 4631 -1342 4647 -1308
rect 4681 -1342 4697 -1308
rect 4749 -1342 4765 -1308
rect 4799 -1342 4815 -1308
rect 4867 -1342 4883 -1308
rect 4917 -1342 4933 -1308
rect 4120 -1410 4154 -1348
rect 5090 -1348 5160 -792
rect 6096 -792 6234 -730
rect 5317 -832 5333 -798
rect 5367 -832 5383 -798
rect 5435 -832 5451 -798
rect 5485 -832 5501 -798
rect 5553 -832 5569 -798
rect 5603 -832 5619 -798
rect 5671 -832 5687 -798
rect 5721 -832 5737 -798
rect 5789 -832 5805 -798
rect 5839 -832 5855 -798
rect 5907 -832 5923 -798
rect 5957 -832 5973 -798
rect 5274 -882 5308 -866
rect 5274 -1274 5308 -1258
rect 5392 -882 5426 -866
rect 5392 -1274 5426 -1258
rect 5510 -882 5544 -866
rect 5510 -1274 5544 -1258
rect 5628 -882 5662 -866
rect 5628 -1274 5662 -1258
rect 5746 -882 5780 -866
rect 5746 -1274 5780 -1258
rect 5864 -882 5898 -866
rect 5864 -1274 5898 -1258
rect 5982 -882 6016 -866
rect 5982 -1274 6016 -1258
rect 5317 -1342 5333 -1308
rect 5367 -1342 5383 -1308
rect 5435 -1342 5451 -1308
rect 5485 -1342 5501 -1308
rect 5553 -1342 5569 -1308
rect 5603 -1342 5619 -1308
rect 5671 -1342 5687 -1308
rect 5721 -1342 5737 -1308
rect 5789 -1342 5805 -1308
rect 5839 -1342 5855 -1308
rect 5907 -1342 5923 -1308
rect 5957 -1342 5973 -1308
rect 5056 -1410 5194 -1348
rect 6130 -1348 6200 -792
rect 7136 -792 7274 -730
rect 6357 -832 6373 -798
rect 6407 -832 6423 -798
rect 6475 -832 6491 -798
rect 6525 -832 6541 -798
rect 6593 -832 6609 -798
rect 6643 -832 6659 -798
rect 6711 -832 6727 -798
rect 6761 -832 6777 -798
rect 6829 -832 6845 -798
rect 6879 -832 6895 -798
rect 6947 -832 6963 -798
rect 6997 -832 7013 -798
rect 6314 -882 6348 -866
rect 6314 -1274 6348 -1258
rect 6432 -882 6466 -866
rect 6432 -1274 6466 -1258
rect 6550 -882 6584 -866
rect 6550 -1274 6584 -1258
rect 6668 -882 6702 -866
rect 6668 -1274 6702 -1258
rect 6786 -882 6820 -866
rect 6786 -1274 6820 -1258
rect 6904 -882 6938 -866
rect 6904 -1274 6938 -1258
rect 7022 -882 7056 -866
rect 7022 -1274 7056 -1258
rect 6357 -1342 6373 -1308
rect 6407 -1342 6423 -1308
rect 6475 -1342 6491 -1308
rect 6525 -1342 6541 -1308
rect 6593 -1342 6609 -1308
rect 6643 -1342 6659 -1308
rect 6711 -1342 6727 -1308
rect 6761 -1342 6777 -1308
rect 6829 -1342 6845 -1308
rect 6879 -1342 6895 -1308
rect 6947 -1342 6963 -1308
rect 6997 -1342 7013 -1308
rect 6096 -1410 6234 -1348
rect 7170 -1348 7240 -792
rect 8176 -792 8314 -730
rect 7397 -832 7413 -798
rect 7447 -832 7463 -798
rect 7515 -832 7531 -798
rect 7565 -832 7581 -798
rect 7633 -832 7649 -798
rect 7683 -832 7699 -798
rect 7751 -832 7767 -798
rect 7801 -832 7817 -798
rect 7869 -832 7885 -798
rect 7919 -832 7935 -798
rect 7987 -832 8003 -798
rect 8037 -832 8053 -798
rect 7354 -882 7388 -866
rect 7354 -1274 7388 -1258
rect 7472 -882 7506 -866
rect 7472 -1274 7506 -1258
rect 7590 -882 7624 -866
rect 7590 -1274 7624 -1258
rect 7708 -882 7742 -866
rect 7708 -1274 7742 -1258
rect 7826 -882 7860 -866
rect 7826 -1274 7860 -1258
rect 7944 -882 7978 -866
rect 7944 -1274 7978 -1258
rect 8062 -882 8096 -866
rect 8062 -1274 8096 -1258
rect 7397 -1342 7413 -1308
rect 7447 -1342 7463 -1308
rect 7515 -1342 7531 -1308
rect 7565 -1342 7581 -1308
rect 7633 -1342 7649 -1308
rect 7683 -1342 7699 -1308
rect 7751 -1342 7767 -1308
rect 7801 -1342 7817 -1308
rect 7869 -1342 7885 -1308
rect 7919 -1342 7935 -1308
rect 7987 -1342 8003 -1308
rect 8037 -1342 8053 -1308
rect 7136 -1410 7274 -1348
rect 8210 -1348 8280 -792
rect 9216 -792 9354 -730
rect 8437 -832 8453 -798
rect 8487 -832 8503 -798
rect 8555 -832 8571 -798
rect 8605 -832 8621 -798
rect 8673 -832 8689 -798
rect 8723 -832 8739 -798
rect 8791 -832 8807 -798
rect 8841 -832 8857 -798
rect 8909 -832 8925 -798
rect 8959 -832 8975 -798
rect 9027 -832 9043 -798
rect 9077 -832 9093 -798
rect 8394 -882 8428 -866
rect 8394 -1274 8428 -1258
rect 8512 -882 8546 -866
rect 8512 -1274 8546 -1258
rect 8630 -882 8664 -866
rect 8630 -1274 8664 -1258
rect 8748 -882 8782 -866
rect 8748 -1274 8782 -1258
rect 8866 -882 8900 -866
rect 8866 -1274 8900 -1258
rect 8984 -882 9018 -866
rect 8984 -1274 9018 -1258
rect 9102 -882 9136 -866
rect 9102 -1274 9136 -1258
rect 8437 -1342 8453 -1308
rect 8487 -1342 8503 -1308
rect 8555 -1342 8571 -1308
rect 8605 -1342 8621 -1308
rect 8673 -1342 8689 -1308
rect 8723 -1342 8739 -1308
rect 8791 -1342 8807 -1308
rect 8841 -1342 8857 -1308
rect 8909 -1342 8925 -1308
rect 8959 -1342 8975 -1308
rect 9027 -1342 9043 -1308
rect 9077 -1342 9093 -1308
rect 8176 -1410 8314 -1348
rect 9250 -1348 9320 -792
rect 10256 -792 10290 -730
rect 9477 -832 9493 -798
rect 9527 -832 9543 -798
rect 9595 -832 9611 -798
rect 9645 -832 9661 -798
rect 9713 -832 9729 -798
rect 9763 -832 9779 -798
rect 9831 -832 9847 -798
rect 9881 -832 9897 -798
rect 9949 -832 9965 -798
rect 9999 -832 10015 -798
rect 10067 -832 10083 -798
rect 10117 -832 10133 -798
rect 9434 -882 9468 -866
rect 9434 -1274 9468 -1258
rect 9552 -882 9586 -866
rect 9552 -1274 9586 -1258
rect 9670 -882 9704 -866
rect 9670 -1274 9704 -1258
rect 9788 -882 9822 -866
rect 9788 -1274 9822 -1258
rect 9906 -882 9940 -866
rect 9906 -1274 9940 -1258
rect 10024 -882 10058 -866
rect 10024 -1274 10058 -1258
rect 10142 -882 10176 -866
rect 10142 -1274 10176 -1258
rect 9477 -1342 9493 -1308
rect 9527 -1342 9543 -1308
rect 9595 -1342 9611 -1308
rect 9645 -1342 9661 -1308
rect 9713 -1342 9729 -1308
rect 9763 -1342 9779 -1308
rect 9831 -1342 9847 -1308
rect 9881 -1342 9897 -1308
rect 9949 -1342 9965 -1308
rect 9999 -1342 10015 -1308
rect 10067 -1342 10083 -1308
rect 10117 -1342 10133 -1308
rect 9216 -1410 9354 -1348
rect 10256 -1410 10290 -1348
rect 4120 -1444 4216 -1410
rect 4994 -1440 5256 -1410
rect 4994 -1444 5090 -1440
rect 5160 -1444 5256 -1440
rect 6034 -1440 6296 -1410
rect 6034 -1444 6130 -1440
rect 6200 -1444 6296 -1440
rect 7074 -1440 7336 -1410
rect 7074 -1444 7170 -1440
rect 7240 -1444 7336 -1440
rect 8114 -1440 8376 -1410
rect 8114 -1444 8210 -1440
rect 8280 -1444 8376 -1440
rect 9154 -1440 9416 -1410
rect 9154 -1444 9250 -1440
rect 9320 -1444 9416 -1440
rect 10194 -1444 10290 -1410
rect 10360 -730 10456 -696
rect 11234 -730 11330 -696
rect 10360 -792 10394 -730
rect 11296 -792 11330 -730
rect 10517 -832 10533 -798
rect 10567 -832 10583 -798
rect 10635 -832 10651 -798
rect 10685 -832 10701 -798
rect 10753 -832 10769 -798
rect 10803 -832 10819 -798
rect 10871 -832 10887 -798
rect 10921 -832 10937 -798
rect 10989 -832 11005 -798
rect 11039 -832 11055 -798
rect 11107 -832 11123 -798
rect 11157 -832 11173 -798
rect 10474 -882 10508 -866
rect 10474 -1274 10508 -1258
rect 10592 -882 10626 -866
rect 10592 -1274 10626 -1258
rect 10710 -882 10744 -866
rect 10710 -1274 10744 -1258
rect 10828 -882 10862 -866
rect 10828 -1274 10862 -1258
rect 10946 -882 10980 -866
rect 10946 -1274 10980 -1258
rect 11064 -882 11098 -866
rect 11064 -1274 11098 -1258
rect 11182 -882 11216 -866
rect 11182 -1274 11216 -1258
rect 10517 -1342 10533 -1308
rect 10567 -1342 10583 -1308
rect 10635 -1342 10651 -1308
rect 10685 -1342 10701 -1308
rect 10753 -1342 10769 -1308
rect 10803 -1342 10819 -1308
rect 10871 -1342 10887 -1308
rect 10921 -1342 10937 -1308
rect 10989 -1342 11005 -1308
rect 11039 -1342 11055 -1308
rect 11107 -1342 11123 -1308
rect 11157 -1342 11173 -1308
rect 10360 -1410 10394 -1348
rect 11296 -1410 11330 -1348
rect 10360 -1444 10456 -1410
rect 11234 -1444 11330 -1410
rect 11740 -730 11836 -696
rect 12614 -700 12710 -696
rect 12780 -700 12876 -696
rect 12614 -730 12876 -700
rect 13654 -700 13750 -696
rect 13820 -700 13916 -696
rect 13654 -730 13916 -700
rect 14694 -700 14790 -696
rect 14860 -700 14956 -696
rect 14694 -730 14956 -700
rect 15734 -700 15830 -696
rect 15900 -700 15996 -696
rect 15734 -730 15996 -700
rect 16774 -700 16870 -696
rect 16940 -700 17036 -696
rect 16774 -730 17036 -700
rect 17814 -730 17910 -696
rect 11740 -792 11774 -730
rect 12676 -792 12814 -730
rect 11897 -832 11913 -798
rect 11947 -832 11963 -798
rect 12015 -832 12031 -798
rect 12065 -832 12081 -798
rect 12133 -832 12149 -798
rect 12183 -832 12199 -798
rect 12251 -832 12267 -798
rect 12301 -832 12317 -798
rect 12369 -832 12385 -798
rect 12419 -832 12435 -798
rect 12487 -832 12503 -798
rect 12537 -832 12553 -798
rect 11854 -882 11888 -866
rect 11854 -1274 11888 -1258
rect 11972 -882 12006 -866
rect 11972 -1274 12006 -1258
rect 12090 -882 12124 -866
rect 12090 -1274 12124 -1258
rect 12208 -882 12242 -866
rect 12208 -1274 12242 -1258
rect 12326 -882 12360 -866
rect 12326 -1274 12360 -1258
rect 12444 -882 12478 -866
rect 12444 -1274 12478 -1258
rect 12562 -882 12596 -866
rect 12562 -1274 12596 -1258
rect 11897 -1342 11913 -1308
rect 11947 -1342 11963 -1308
rect 12015 -1342 12031 -1308
rect 12065 -1342 12081 -1308
rect 12133 -1342 12149 -1308
rect 12183 -1342 12199 -1308
rect 12251 -1342 12267 -1308
rect 12301 -1342 12317 -1308
rect 12369 -1342 12385 -1308
rect 12419 -1342 12435 -1308
rect 12487 -1342 12503 -1308
rect 12537 -1342 12553 -1308
rect 11740 -1410 11774 -1348
rect 12710 -1348 12780 -792
rect 13716 -792 13854 -730
rect 12937 -832 12953 -798
rect 12987 -832 13003 -798
rect 13055 -832 13071 -798
rect 13105 -832 13121 -798
rect 13173 -832 13189 -798
rect 13223 -832 13239 -798
rect 13291 -832 13307 -798
rect 13341 -832 13357 -798
rect 13409 -832 13425 -798
rect 13459 -832 13475 -798
rect 13527 -832 13543 -798
rect 13577 -832 13593 -798
rect 12894 -882 12928 -866
rect 12894 -1274 12928 -1258
rect 13012 -882 13046 -866
rect 13012 -1274 13046 -1258
rect 13130 -882 13164 -866
rect 13130 -1274 13164 -1258
rect 13248 -882 13282 -866
rect 13248 -1274 13282 -1258
rect 13366 -882 13400 -866
rect 13366 -1274 13400 -1258
rect 13484 -882 13518 -866
rect 13484 -1274 13518 -1258
rect 13602 -882 13636 -866
rect 13602 -1274 13636 -1258
rect 12937 -1342 12953 -1308
rect 12987 -1342 13003 -1308
rect 13055 -1342 13071 -1308
rect 13105 -1342 13121 -1308
rect 13173 -1342 13189 -1308
rect 13223 -1342 13239 -1308
rect 13291 -1342 13307 -1308
rect 13341 -1342 13357 -1308
rect 13409 -1342 13425 -1308
rect 13459 -1342 13475 -1308
rect 13527 -1342 13543 -1308
rect 13577 -1342 13593 -1308
rect 12676 -1410 12814 -1348
rect 13750 -1348 13820 -792
rect 14756 -792 14894 -730
rect 13977 -832 13993 -798
rect 14027 -832 14043 -798
rect 14095 -832 14111 -798
rect 14145 -832 14161 -798
rect 14213 -832 14229 -798
rect 14263 -832 14279 -798
rect 14331 -832 14347 -798
rect 14381 -832 14397 -798
rect 14449 -832 14465 -798
rect 14499 -832 14515 -798
rect 14567 -832 14583 -798
rect 14617 -832 14633 -798
rect 13934 -882 13968 -866
rect 13934 -1274 13968 -1258
rect 14052 -882 14086 -866
rect 14052 -1274 14086 -1258
rect 14170 -882 14204 -866
rect 14170 -1274 14204 -1258
rect 14288 -882 14322 -866
rect 14288 -1274 14322 -1258
rect 14406 -882 14440 -866
rect 14406 -1274 14440 -1258
rect 14524 -882 14558 -866
rect 14524 -1274 14558 -1258
rect 14642 -882 14676 -866
rect 14642 -1274 14676 -1258
rect 13977 -1342 13993 -1308
rect 14027 -1342 14043 -1308
rect 14095 -1342 14111 -1308
rect 14145 -1342 14161 -1308
rect 14213 -1342 14229 -1308
rect 14263 -1342 14279 -1308
rect 14331 -1342 14347 -1308
rect 14381 -1342 14397 -1308
rect 14449 -1342 14465 -1308
rect 14499 -1342 14515 -1308
rect 14567 -1342 14583 -1308
rect 14617 -1342 14633 -1308
rect 13716 -1410 13854 -1348
rect 14790 -1348 14860 -792
rect 15796 -792 15934 -730
rect 15017 -832 15033 -798
rect 15067 -832 15083 -798
rect 15135 -832 15151 -798
rect 15185 -832 15201 -798
rect 15253 -832 15269 -798
rect 15303 -832 15319 -798
rect 15371 -832 15387 -798
rect 15421 -832 15437 -798
rect 15489 -832 15505 -798
rect 15539 -832 15555 -798
rect 15607 -832 15623 -798
rect 15657 -832 15673 -798
rect 14974 -882 15008 -866
rect 14974 -1274 15008 -1258
rect 15092 -882 15126 -866
rect 15092 -1274 15126 -1258
rect 15210 -882 15244 -866
rect 15210 -1274 15244 -1258
rect 15328 -882 15362 -866
rect 15328 -1274 15362 -1258
rect 15446 -882 15480 -866
rect 15446 -1274 15480 -1258
rect 15564 -882 15598 -866
rect 15564 -1274 15598 -1258
rect 15682 -882 15716 -866
rect 15682 -1274 15716 -1258
rect 15017 -1342 15033 -1308
rect 15067 -1342 15083 -1308
rect 15135 -1342 15151 -1308
rect 15185 -1342 15201 -1308
rect 15253 -1342 15269 -1308
rect 15303 -1342 15319 -1308
rect 15371 -1342 15387 -1308
rect 15421 -1342 15437 -1308
rect 15489 -1342 15505 -1308
rect 15539 -1342 15555 -1308
rect 15607 -1342 15623 -1308
rect 15657 -1342 15673 -1308
rect 14756 -1410 14894 -1348
rect 15830 -1348 15900 -792
rect 16836 -792 16974 -730
rect 16057 -832 16073 -798
rect 16107 -832 16123 -798
rect 16175 -832 16191 -798
rect 16225 -832 16241 -798
rect 16293 -832 16309 -798
rect 16343 -832 16359 -798
rect 16411 -832 16427 -798
rect 16461 -832 16477 -798
rect 16529 -832 16545 -798
rect 16579 -832 16595 -798
rect 16647 -832 16663 -798
rect 16697 -832 16713 -798
rect 16014 -882 16048 -866
rect 16014 -1274 16048 -1258
rect 16132 -882 16166 -866
rect 16132 -1274 16166 -1258
rect 16250 -882 16284 -866
rect 16250 -1274 16284 -1258
rect 16368 -882 16402 -866
rect 16368 -1274 16402 -1258
rect 16486 -882 16520 -866
rect 16486 -1274 16520 -1258
rect 16604 -882 16638 -866
rect 16604 -1274 16638 -1258
rect 16722 -882 16756 -866
rect 16722 -1274 16756 -1258
rect 16057 -1342 16073 -1308
rect 16107 -1342 16123 -1308
rect 16175 -1342 16191 -1308
rect 16225 -1342 16241 -1308
rect 16293 -1342 16309 -1308
rect 16343 -1342 16359 -1308
rect 16411 -1342 16427 -1308
rect 16461 -1342 16477 -1308
rect 16529 -1342 16545 -1308
rect 16579 -1342 16595 -1308
rect 16647 -1342 16663 -1308
rect 16697 -1342 16713 -1308
rect 15796 -1410 15934 -1348
rect 16870 -1348 16940 -792
rect 17876 -792 17910 -730
rect 17097 -832 17113 -798
rect 17147 -832 17163 -798
rect 17215 -832 17231 -798
rect 17265 -832 17281 -798
rect 17333 -832 17349 -798
rect 17383 -832 17399 -798
rect 17451 -832 17467 -798
rect 17501 -832 17517 -798
rect 17569 -832 17585 -798
rect 17619 -832 17635 -798
rect 17687 -832 17703 -798
rect 17737 -832 17753 -798
rect 17054 -882 17088 -866
rect 17054 -1274 17088 -1258
rect 17172 -882 17206 -866
rect 17172 -1274 17206 -1258
rect 17290 -882 17324 -866
rect 17290 -1274 17324 -1258
rect 17408 -882 17442 -866
rect 17408 -1274 17442 -1258
rect 17526 -882 17560 -866
rect 17526 -1274 17560 -1258
rect 17644 -882 17678 -866
rect 17644 -1274 17678 -1258
rect 17762 -882 17796 -866
rect 17762 -1274 17796 -1258
rect 17097 -1342 17113 -1308
rect 17147 -1342 17163 -1308
rect 17215 -1342 17231 -1308
rect 17265 -1342 17281 -1308
rect 17333 -1342 17349 -1308
rect 17383 -1342 17399 -1308
rect 17451 -1342 17467 -1308
rect 17501 -1342 17517 -1308
rect 17569 -1342 17585 -1308
rect 17619 -1342 17635 -1308
rect 17687 -1342 17703 -1308
rect 17737 -1342 17753 -1308
rect 16836 -1410 16974 -1348
rect 17876 -1410 17910 -1348
rect 11740 -1444 11836 -1410
rect 12614 -1440 12876 -1410
rect 12614 -1444 12710 -1440
rect 12780 -1444 12876 -1440
rect 13654 -1440 13916 -1410
rect 13654 -1444 13750 -1440
rect 13820 -1444 13916 -1440
rect 14694 -1440 14956 -1410
rect 14694 -1444 14790 -1440
rect 14860 -1444 14956 -1440
rect 15734 -1440 15996 -1410
rect 15734 -1444 15830 -1440
rect 15900 -1444 15996 -1440
rect 16774 -1440 17036 -1410
rect 16774 -1444 16870 -1440
rect 16940 -1444 17036 -1440
rect 17814 -1444 17910 -1410
rect 17980 -730 18076 -696
rect 18854 -730 18950 -696
rect 17980 -792 18014 -730
rect 18916 -792 18950 -730
rect 18137 -832 18153 -798
rect 18187 -832 18203 -798
rect 18255 -832 18271 -798
rect 18305 -832 18321 -798
rect 18373 -832 18389 -798
rect 18423 -832 18439 -798
rect 18491 -832 18507 -798
rect 18541 -832 18557 -798
rect 18609 -832 18625 -798
rect 18659 -832 18675 -798
rect 18727 -832 18743 -798
rect 18777 -832 18793 -798
rect 18094 -882 18128 -866
rect 18094 -1274 18128 -1258
rect 18212 -882 18246 -866
rect 18212 -1274 18246 -1258
rect 18330 -882 18364 -866
rect 18330 -1274 18364 -1258
rect 18448 -882 18482 -866
rect 18448 -1274 18482 -1258
rect 18566 -882 18600 -866
rect 18566 -1274 18600 -1258
rect 18684 -882 18718 -866
rect 18684 -1274 18718 -1258
rect 18802 -882 18836 -866
rect 18802 -1274 18836 -1258
rect 18137 -1342 18153 -1308
rect 18187 -1342 18203 -1308
rect 18255 -1342 18271 -1308
rect 18305 -1342 18321 -1308
rect 18373 -1342 18389 -1308
rect 18423 -1342 18439 -1308
rect 18491 -1342 18507 -1308
rect 18541 -1342 18557 -1308
rect 18609 -1342 18625 -1308
rect 18659 -1342 18675 -1308
rect 18727 -1342 18743 -1308
rect 18777 -1342 18793 -1308
rect 17980 -1410 18014 -1348
rect 18916 -1410 18950 -1348
rect 17980 -1444 18076 -1410
rect 18854 -1444 18950 -1410
rect 4184 -1514 4904 -1444
rect 5224 -1514 5944 -1444
rect 6224 -1514 6944 -1444
rect 7264 -1514 7984 -1444
rect 8324 -1514 9044 -1444
rect 11804 -1514 12524 -1444
rect 12844 -1514 13564 -1444
rect 13844 -1514 14564 -1444
rect 14884 -1514 15604 -1444
rect 15944 -1514 16664 -1444
rect -6310 -1834 -6186 -1754
rect -5660 -1780 -5626 -1718
rect -5722 -1814 -5626 -1780
rect 4120 -1548 4216 -1514
rect 4862 -1548 4958 -1514
rect 4120 -1610 4154 -1548
rect -6710 -3048 -6676 -2986
rect -7514 -3082 -7418 -3048
rect -6772 -3070 -6676 -3048
rect 4924 -1610 4958 -1548
rect 4266 -1650 4282 -1616
rect 4316 -1650 4332 -1616
rect 4458 -1650 4474 -1616
rect 4508 -1650 4524 -1616
rect 4650 -1650 4666 -1616
rect 4700 -1650 4716 -1616
rect 4234 -1700 4268 -1684
rect 4234 -2092 4268 -2076
rect 4330 -1700 4364 -1684
rect 4330 -2092 4364 -2076
rect 4426 -1700 4460 -1684
rect 4426 -2092 4460 -2076
rect 4522 -1700 4556 -1684
rect 4522 -2092 4556 -2076
rect 4618 -1700 4652 -1684
rect 4618 -2092 4652 -2076
rect 4714 -1700 4748 -1684
rect 4714 -2092 4748 -2076
rect 4810 -1700 4844 -1684
rect 4810 -2092 4844 -2076
rect 4362 -2160 4378 -2126
rect 4412 -2160 4428 -2126
rect 4554 -2160 4570 -2126
rect 4604 -2160 4620 -2126
rect 4746 -2160 4762 -2126
rect 4796 -2160 4812 -2126
rect 4362 -2268 4378 -2234
rect 4412 -2268 4428 -2234
rect 4554 -2268 4570 -2234
rect 4604 -2268 4620 -2234
rect 4746 -2268 4762 -2234
rect 4796 -2268 4812 -2234
rect 4234 -2318 4268 -2302
rect 4234 -2710 4268 -2694
rect 4330 -2318 4364 -2302
rect 4330 -2710 4364 -2694
rect 4426 -2318 4460 -2302
rect 4426 -2710 4460 -2694
rect 4522 -2318 4556 -2302
rect 4522 -2710 4556 -2694
rect 4618 -2318 4652 -2302
rect 4618 -2710 4652 -2694
rect 4714 -2318 4748 -2302
rect 4714 -2710 4748 -2694
rect 4810 -2318 4844 -2302
rect 4810 -2710 4844 -2694
rect 4266 -2778 4282 -2744
rect 4316 -2778 4332 -2744
rect 4458 -2778 4474 -2744
rect 4508 -2778 4524 -2744
rect 4650 -2778 4666 -2744
rect 4700 -2778 4716 -2744
rect 4120 -2846 4154 -2784
rect 4924 -2846 4958 -2784
rect 4120 -2880 4216 -2846
rect 4862 -2868 4958 -2846
rect 5160 -1548 5256 -1514
rect 5902 -1548 5998 -1514
rect 5160 -1610 5194 -1548
rect 5964 -1610 5998 -1548
rect 5306 -1650 5322 -1616
rect 5356 -1650 5372 -1616
rect 5498 -1650 5514 -1616
rect 5548 -1650 5564 -1616
rect 5690 -1650 5706 -1616
rect 5740 -1650 5756 -1616
rect 5274 -1700 5308 -1684
rect 5274 -2092 5308 -2076
rect 5370 -1700 5404 -1684
rect 5370 -2092 5404 -2076
rect 5466 -1700 5500 -1684
rect 5466 -2092 5500 -2076
rect 5562 -1700 5596 -1684
rect 5562 -2092 5596 -2076
rect 5658 -1700 5692 -1684
rect 5658 -2092 5692 -2076
rect 5754 -1700 5788 -1684
rect 5754 -2092 5788 -2076
rect 5850 -1700 5884 -1684
rect 5850 -2092 5884 -2076
rect 5402 -2160 5418 -2126
rect 5452 -2160 5468 -2126
rect 5594 -2160 5610 -2126
rect 5644 -2160 5660 -2126
rect 5786 -2160 5802 -2126
rect 5836 -2160 5852 -2126
rect 5402 -2268 5418 -2234
rect 5452 -2268 5468 -2234
rect 5594 -2268 5610 -2234
rect 5644 -2268 5660 -2234
rect 5786 -2268 5802 -2234
rect 5836 -2268 5852 -2234
rect 5274 -2318 5308 -2302
rect 5274 -2710 5308 -2694
rect 5370 -2318 5404 -2302
rect 5370 -2710 5404 -2694
rect 5466 -2318 5500 -2302
rect 5466 -2710 5500 -2694
rect 5562 -2318 5596 -2302
rect 5562 -2710 5596 -2694
rect 5658 -2318 5692 -2302
rect 5658 -2710 5692 -2694
rect 5754 -2318 5788 -2302
rect 5754 -2710 5788 -2694
rect 5850 -2318 5884 -2302
rect 5850 -2710 5884 -2694
rect 5306 -2778 5322 -2744
rect 5356 -2778 5372 -2744
rect 5498 -2778 5514 -2744
rect 5548 -2778 5564 -2744
rect 5690 -2778 5706 -2744
rect 5740 -2778 5756 -2744
rect 5160 -2846 5194 -2784
rect 5964 -2846 5998 -2784
rect 4862 -2880 4960 -2868
rect 4120 -2936 4960 -2880
rect 5160 -2880 5256 -2846
rect 5902 -2868 5998 -2846
rect 6200 -1548 6296 -1514
rect 6942 -1548 7038 -1514
rect 6200 -1610 6234 -1548
rect 7004 -1610 7038 -1548
rect 6346 -1650 6362 -1616
rect 6396 -1650 6412 -1616
rect 6538 -1650 6554 -1616
rect 6588 -1650 6604 -1616
rect 6730 -1650 6746 -1616
rect 6780 -1650 6796 -1616
rect 6314 -1700 6348 -1684
rect 6314 -2092 6348 -2076
rect 6410 -1700 6444 -1684
rect 6410 -2092 6444 -2076
rect 6506 -1700 6540 -1684
rect 6506 -2092 6540 -2076
rect 6602 -1700 6636 -1684
rect 6602 -2092 6636 -2076
rect 6698 -1700 6732 -1684
rect 6698 -2092 6732 -2076
rect 6794 -1700 6828 -1684
rect 6794 -2092 6828 -2076
rect 6890 -1700 6924 -1684
rect 6890 -2092 6924 -2076
rect 6442 -2160 6458 -2126
rect 6492 -2160 6508 -2126
rect 6634 -2160 6650 -2126
rect 6684 -2160 6700 -2126
rect 6826 -2160 6842 -2126
rect 6876 -2160 6892 -2126
rect 6442 -2268 6458 -2234
rect 6492 -2268 6508 -2234
rect 6634 -2268 6650 -2234
rect 6684 -2268 6700 -2234
rect 6826 -2268 6842 -2234
rect 6876 -2268 6892 -2234
rect 6314 -2318 6348 -2302
rect 6314 -2710 6348 -2694
rect 6410 -2318 6444 -2302
rect 6410 -2710 6444 -2694
rect 6506 -2318 6540 -2302
rect 6506 -2710 6540 -2694
rect 6602 -2318 6636 -2302
rect 6602 -2710 6636 -2694
rect 6698 -2318 6732 -2302
rect 6698 -2710 6732 -2694
rect 6794 -2318 6828 -2302
rect 6794 -2710 6828 -2694
rect 6890 -2318 6924 -2302
rect 6890 -2710 6924 -2694
rect 6346 -2778 6362 -2744
rect 6396 -2778 6412 -2744
rect 6538 -2778 6554 -2744
rect 6588 -2778 6604 -2744
rect 6730 -2778 6746 -2744
rect 6780 -2778 6796 -2744
rect 6200 -2846 6234 -2784
rect 7004 -2846 7038 -2784
rect 5902 -2880 6000 -2868
rect 5160 -2936 6000 -2880
rect 6200 -2880 6296 -2846
rect 6942 -2868 7038 -2846
rect 7240 -1548 7336 -1514
rect 7982 -1548 8078 -1514
rect 7240 -1610 7274 -1548
rect 8044 -1610 8078 -1548
rect 7386 -1650 7402 -1616
rect 7436 -1650 7452 -1616
rect 7578 -1650 7594 -1616
rect 7628 -1650 7644 -1616
rect 7770 -1650 7786 -1616
rect 7820 -1650 7836 -1616
rect 7354 -1700 7388 -1684
rect 7354 -2092 7388 -2076
rect 7450 -1700 7484 -1684
rect 7450 -2092 7484 -2076
rect 7546 -1700 7580 -1684
rect 7546 -2092 7580 -2076
rect 7642 -1700 7676 -1684
rect 7642 -2092 7676 -2076
rect 7738 -1700 7772 -1684
rect 7738 -2092 7772 -2076
rect 7834 -1700 7868 -1684
rect 7834 -2092 7868 -2076
rect 7930 -1700 7964 -1684
rect 7930 -2092 7964 -2076
rect 7482 -2160 7498 -2126
rect 7532 -2160 7548 -2126
rect 7674 -2160 7690 -2126
rect 7724 -2160 7740 -2126
rect 7866 -2160 7882 -2126
rect 7916 -2160 7932 -2126
rect 7482 -2268 7498 -2234
rect 7532 -2268 7548 -2234
rect 7674 -2268 7690 -2234
rect 7724 -2268 7740 -2234
rect 7866 -2268 7882 -2234
rect 7916 -2268 7932 -2234
rect 7354 -2318 7388 -2302
rect 7354 -2710 7388 -2694
rect 7450 -2318 7484 -2302
rect 7450 -2710 7484 -2694
rect 7546 -2318 7580 -2302
rect 7546 -2710 7580 -2694
rect 7642 -2318 7676 -2302
rect 7642 -2710 7676 -2694
rect 7738 -2318 7772 -2302
rect 7738 -2710 7772 -2694
rect 7834 -2318 7868 -2302
rect 7834 -2710 7868 -2694
rect 7930 -2318 7964 -2302
rect 7930 -2710 7964 -2694
rect 7386 -2778 7402 -2744
rect 7436 -2778 7452 -2744
rect 7578 -2778 7594 -2744
rect 7628 -2778 7644 -2744
rect 7770 -2778 7786 -2744
rect 7820 -2778 7836 -2744
rect 7240 -2846 7274 -2784
rect 8044 -2846 8078 -2784
rect 6942 -2880 7040 -2868
rect 6200 -2936 7040 -2880
rect 7240 -2880 7336 -2846
rect 7982 -2868 8078 -2846
rect 8280 -1548 8376 -1514
rect 9022 -1548 9118 -1514
rect 8280 -1610 8314 -1548
rect 9084 -1610 9118 -1548
rect 8426 -1650 8442 -1616
rect 8476 -1650 8492 -1616
rect 8618 -1650 8634 -1616
rect 8668 -1650 8684 -1616
rect 8810 -1650 8826 -1616
rect 8860 -1650 8876 -1616
rect 8394 -1700 8428 -1684
rect 8394 -2092 8428 -2076
rect 8490 -1700 8524 -1684
rect 8490 -2092 8524 -2076
rect 8586 -1700 8620 -1684
rect 8586 -2092 8620 -2076
rect 8682 -1700 8716 -1684
rect 8682 -2092 8716 -2076
rect 8778 -1700 8812 -1684
rect 8778 -2092 8812 -2076
rect 8874 -1700 8908 -1684
rect 8874 -2092 8908 -2076
rect 8970 -1700 9004 -1684
rect 8970 -2092 9004 -2076
rect 8522 -2160 8538 -2126
rect 8572 -2160 8588 -2126
rect 8714 -2160 8730 -2126
rect 8764 -2160 8780 -2126
rect 8906 -2160 8922 -2126
rect 8956 -2160 8972 -2126
rect 8522 -2268 8538 -2234
rect 8572 -2268 8588 -2234
rect 8714 -2268 8730 -2234
rect 8764 -2268 8780 -2234
rect 8906 -2268 8922 -2234
rect 8956 -2268 8972 -2234
rect 8394 -2318 8428 -2302
rect 8394 -2710 8428 -2694
rect 8490 -2318 8524 -2302
rect 8490 -2710 8524 -2694
rect 8586 -2318 8620 -2302
rect 8586 -2710 8620 -2694
rect 8682 -2318 8716 -2302
rect 8682 -2710 8716 -2694
rect 8778 -2318 8812 -2302
rect 8778 -2710 8812 -2694
rect 8874 -2318 8908 -2302
rect 8874 -2710 8908 -2694
rect 8970 -2318 9004 -2302
rect 8970 -2710 9004 -2694
rect 8426 -2778 8442 -2744
rect 8476 -2778 8492 -2744
rect 8618 -2778 8634 -2744
rect 8668 -2778 8684 -2744
rect 8810 -2778 8826 -2744
rect 8860 -2778 8876 -2744
rect 8280 -2846 8314 -2784
rect 9084 -2846 9118 -2784
rect 7982 -2880 8080 -2868
rect 7240 -2936 8080 -2880
rect 8280 -2880 8376 -2846
rect 9022 -2868 9118 -2846
rect 11740 -1548 11836 -1514
rect 12482 -1548 12578 -1514
rect 11740 -1610 11774 -1548
rect 12544 -1610 12578 -1548
rect 11886 -1650 11902 -1616
rect 11936 -1650 11952 -1616
rect 12078 -1650 12094 -1616
rect 12128 -1650 12144 -1616
rect 12270 -1650 12286 -1616
rect 12320 -1650 12336 -1616
rect 11854 -1700 11888 -1684
rect 11854 -2092 11888 -2076
rect 11950 -1700 11984 -1684
rect 11950 -2092 11984 -2076
rect 12046 -1700 12080 -1684
rect 12046 -2092 12080 -2076
rect 12142 -1700 12176 -1684
rect 12142 -2092 12176 -2076
rect 12238 -1700 12272 -1684
rect 12238 -2092 12272 -2076
rect 12334 -1700 12368 -1684
rect 12334 -2092 12368 -2076
rect 12430 -1700 12464 -1684
rect 12430 -2092 12464 -2076
rect 11982 -2160 11998 -2126
rect 12032 -2160 12048 -2126
rect 12174 -2160 12190 -2126
rect 12224 -2160 12240 -2126
rect 12366 -2160 12382 -2126
rect 12416 -2160 12432 -2126
rect 11982 -2268 11998 -2234
rect 12032 -2268 12048 -2234
rect 12174 -2268 12190 -2234
rect 12224 -2268 12240 -2234
rect 12366 -2268 12382 -2234
rect 12416 -2268 12432 -2234
rect 11854 -2318 11888 -2302
rect 11854 -2710 11888 -2694
rect 11950 -2318 11984 -2302
rect 11950 -2710 11984 -2694
rect 12046 -2318 12080 -2302
rect 12046 -2710 12080 -2694
rect 12142 -2318 12176 -2302
rect 12142 -2710 12176 -2694
rect 12238 -2318 12272 -2302
rect 12238 -2710 12272 -2694
rect 12334 -2318 12368 -2302
rect 12334 -2710 12368 -2694
rect 12430 -2318 12464 -2302
rect 12430 -2710 12464 -2694
rect 11886 -2778 11902 -2744
rect 11936 -2778 11952 -2744
rect 12078 -2778 12094 -2744
rect 12128 -2778 12144 -2744
rect 12270 -2778 12286 -2744
rect 12320 -2778 12336 -2744
rect 11740 -2846 11774 -2784
rect 12544 -2846 12578 -2784
rect 9022 -2880 9120 -2868
rect 8280 -2936 9120 -2880
rect 11740 -2880 11836 -2846
rect 12482 -2868 12578 -2846
rect 12780 -1548 12876 -1514
rect 13522 -1548 13618 -1514
rect 12780 -1610 12814 -1548
rect 13584 -1610 13618 -1548
rect 12926 -1650 12942 -1616
rect 12976 -1650 12992 -1616
rect 13118 -1650 13134 -1616
rect 13168 -1650 13184 -1616
rect 13310 -1650 13326 -1616
rect 13360 -1650 13376 -1616
rect 12894 -1700 12928 -1684
rect 12894 -2092 12928 -2076
rect 12990 -1700 13024 -1684
rect 12990 -2092 13024 -2076
rect 13086 -1700 13120 -1684
rect 13086 -2092 13120 -2076
rect 13182 -1700 13216 -1684
rect 13182 -2092 13216 -2076
rect 13278 -1700 13312 -1684
rect 13278 -2092 13312 -2076
rect 13374 -1700 13408 -1684
rect 13374 -2092 13408 -2076
rect 13470 -1700 13504 -1684
rect 13470 -2092 13504 -2076
rect 13022 -2160 13038 -2126
rect 13072 -2160 13088 -2126
rect 13214 -2160 13230 -2126
rect 13264 -2160 13280 -2126
rect 13406 -2160 13422 -2126
rect 13456 -2160 13472 -2126
rect 13022 -2268 13038 -2234
rect 13072 -2268 13088 -2234
rect 13214 -2268 13230 -2234
rect 13264 -2268 13280 -2234
rect 13406 -2268 13422 -2234
rect 13456 -2268 13472 -2234
rect 12894 -2318 12928 -2302
rect 12894 -2710 12928 -2694
rect 12990 -2318 13024 -2302
rect 12990 -2710 13024 -2694
rect 13086 -2318 13120 -2302
rect 13086 -2710 13120 -2694
rect 13182 -2318 13216 -2302
rect 13182 -2710 13216 -2694
rect 13278 -2318 13312 -2302
rect 13278 -2710 13312 -2694
rect 13374 -2318 13408 -2302
rect 13374 -2710 13408 -2694
rect 13470 -2318 13504 -2302
rect 13470 -2710 13504 -2694
rect 12926 -2778 12942 -2744
rect 12976 -2778 12992 -2744
rect 13118 -2778 13134 -2744
rect 13168 -2778 13184 -2744
rect 13310 -2778 13326 -2744
rect 13360 -2778 13376 -2744
rect 12780 -2846 12814 -2784
rect 13584 -2846 13618 -2784
rect 12482 -2880 12580 -2868
rect 11740 -2936 12580 -2880
rect 12780 -2880 12876 -2846
rect 13522 -2868 13618 -2846
rect 13820 -1548 13916 -1514
rect 14562 -1548 14658 -1514
rect 13820 -1610 13854 -1548
rect 14624 -1610 14658 -1548
rect 13966 -1650 13982 -1616
rect 14016 -1650 14032 -1616
rect 14158 -1650 14174 -1616
rect 14208 -1650 14224 -1616
rect 14350 -1650 14366 -1616
rect 14400 -1650 14416 -1616
rect 13934 -1700 13968 -1684
rect 13934 -2092 13968 -2076
rect 14030 -1700 14064 -1684
rect 14030 -2092 14064 -2076
rect 14126 -1700 14160 -1684
rect 14126 -2092 14160 -2076
rect 14222 -1700 14256 -1684
rect 14222 -2092 14256 -2076
rect 14318 -1700 14352 -1684
rect 14318 -2092 14352 -2076
rect 14414 -1700 14448 -1684
rect 14414 -2092 14448 -2076
rect 14510 -1700 14544 -1684
rect 14510 -2092 14544 -2076
rect 14062 -2160 14078 -2126
rect 14112 -2160 14128 -2126
rect 14254 -2160 14270 -2126
rect 14304 -2160 14320 -2126
rect 14446 -2160 14462 -2126
rect 14496 -2160 14512 -2126
rect 14062 -2268 14078 -2234
rect 14112 -2268 14128 -2234
rect 14254 -2268 14270 -2234
rect 14304 -2268 14320 -2234
rect 14446 -2268 14462 -2234
rect 14496 -2268 14512 -2234
rect 13934 -2318 13968 -2302
rect 13934 -2710 13968 -2694
rect 14030 -2318 14064 -2302
rect 14030 -2710 14064 -2694
rect 14126 -2318 14160 -2302
rect 14126 -2710 14160 -2694
rect 14222 -2318 14256 -2302
rect 14222 -2710 14256 -2694
rect 14318 -2318 14352 -2302
rect 14318 -2710 14352 -2694
rect 14414 -2318 14448 -2302
rect 14414 -2710 14448 -2694
rect 14510 -2318 14544 -2302
rect 14510 -2710 14544 -2694
rect 13966 -2778 13982 -2744
rect 14016 -2778 14032 -2744
rect 14158 -2778 14174 -2744
rect 14208 -2778 14224 -2744
rect 14350 -2778 14366 -2744
rect 14400 -2778 14416 -2744
rect 13820 -2846 13854 -2784
rect 14624 -2846 14658 -2784
rect 13522 -2880 13620 -2868
rect 12780 -2936 13620 -2880
rect 13820 -2880 13916 -2846
rect 14562 -2868 14658 -2846
rect 14860 -1548 14956 -1514
rect 15602 -1548 15698 -1514
rect 14860 -1610 14894 -1548
rect 15664 -1610 15698 -1548
rect 15006 -1650 15022 -1616
rect 15056 -1650 15072 -1616
rect 15198 -1650 15214 -1616
rect 15248 -1650 15264 -1616
rect 15390 -1650 15406 -1616
rect 15440 -1650 15456 -1616
rect 14974 -1700 15008 -1684
rect 14974 -2092 15008 -2076
rect 15070 -1700 15104 -1684
rect 15070 -2092 15104 -2076
rect 15166 -1700 15200 -1684
rect 15166 -2092 15200 -2076
rect 15262 -1700 15296 -1684
rect 15262 -2092 15296 -2076
rect 15358 -1700 15392 -1684
rect 15358 -2092 15392 -2076
rect 15454 -1700 15488 -1684
rect 15454 -2092 15488 -2076
rect 15550 -1700 15584 -1684
rect 15550 -2092 15584 -2076
rect 15102 -2160 15118 -2126
rect 15152 -2160 15168 -2126
rect 15294 -2160 15310 -2126
rect 15344 -2160 15360 -2126
rect 15486 -2160 15502 -2126
rect 15536 -2160 15552 -2126
rect 15102 -2268 15118 -2234
rect 15152 -2268 15168 -2234
rect 15294 -2268 15310 -2234
rect 15344 -2268 15360 -2234
rect 15486 -2268 15502 -2234
rect 15536 -2268 15552 -2234
rect 14974 -2318 15008 -2302
rect 14974 -2710 15008 -2694
rect 15070 -2318 15104 -2302
rect 15070 -2710 15104 -2694
rect 15166 -2318 15200 -2302
rect 15166 -2710 15200 -2694
rect 15262 -2318 15296 -2302
rect 15262 -2710 15296 -2694
rect 15358 -2318 15392 -2302
rect 15358 -2710 15392 -2694
rect 15454 -2318 15488 -2302
rect 15454 -2710 15488 -2694
rect 15550 -2318 15584 -2302
rect 15550 -2710 15584 -2694
rect 15006 -2778 15022 -2744
rect 15056 -2778 15072 -2744
rect 15198 -2778 15214 -2744
rect 15248 -2778 15264 -2744
rect 15390 -2778 15406 -2744
rect 15440 -2778 15456 -2744
rect 14860 -2846 14894 -2784
rect 15664 -2846 15698 -2784
rect 14562 -2880 14660 -2868
rect 13820 -2936 14660 -2880
rect 14860 -2880 14956 -2846
rect 15602 -2868 15698 -2846
rect 15900 -1548 15996 -1514
rect 16642 -1548 16738 -1514
rect 15900 -1610 15934 -1548
rect 16704 -1610 16738 -1548
rect 16046 -1650 16062 -1616
rect 16096 -1650 16112 -1616
rect 16238 -1650 16254 -1616
rect 16288 -1650 16304 -1616
rect 16430 -1650 16446 -1616
rect 16480 -1650 16496 -1616
rect 16014 -1700 16048 -1684
rect 16014 -2092 16048 -2076
rect 16110 -1700 16144 -1684
rect 16110 -2092 16144 -2076
rect 16206 -1700 16240 -1684
rect 16206 -2092 16240 -2076
rect 16302 -1700 16336 -1684
rect 16302 -2092 16336 -2076
rect 16398 -1700 16432 -1684
rect 16398 -2092 16432 -2076
rect 16494 -1700 16528 -1684
rect 16494 -2092 16528 -2076
rect 16590 -1700 16624 -1684
rect 16590 -2092 16624 -2076
rect 16142 -2160 16158 -2126
rect 16192 -2160 16208 -2126
rect 16334 -2160 16350 -2126
rect 16384 -2160 16400 -2126
rect 16526 -2160 16542 -2126
rect 16576 -2160 16592 -2126
rect 16142 -2268 16158 -2234
rect 16192 -2268 16208 -2234
rect 16334 -2268 16350 -2234
rect 16384 -2268 16400 -2234
rect 16526 -2268 16542 -2234
rect 16576 -2268 16592 -2234
rect 16014 -2318 16048 -2302
rect 16014 -2710 16048 -2694
rect 16110 -2318 16144 -2302
rect 16110 -2710 16144 -2694
rect 16206 -2318 16240 -2302
rect 16206 -2710 16240 -2694
rect 16302 -2318 16336 -2302
rect 16302 -2710 16336 -2694
rect 16398 -2318 16432 -2302
rect 16398 -2710 16432 -2694
rect 16494 -2318 16528 -2302
rect 16494 -2710 16528 -2694
rect 16590 -2318 16624 -2302
rect 16590 -2710 16624 -2694
rect 16046 -2778 16062 -2744
rect 16096 -2778 16112 -2744
rect 16238 -2778 16254 -2744
rect 16288 -2778 16304 -2744
rect 16430 -2778 16446 -2744
rect 16480 -2778 16496 -2744
rect 15900 -2846 15934 -2784
rect 16704 -2846 16738 -2784
rect 15602 -2880 15700 -2868
rect 14860 -2936 15700 -2880
rect 15900 -2880 15996 -2846
rect 16642 -2868 16738 -2846
rect 16642 -2880 16740 -2868
rect 15900 -2936 16740 -2880
rect 4120 -2970 4216 -2936
rect 4994 -2970 5090 -2936
rect 4120 -3032 4154 -2970
rect -6772 -3082 -6674 -3070
rect -7514 -3138 -6674 -3082
rect -7514 -3172 -7418 -3138
rect -6640 -3172 -6544 -3138
rect -7514 -3234 -7480 -3172
rect -6578 -3234 -6544 -3172
rect -7357 -3274 -7341 -3240
rect -7307 -3274 -7291 -3240
rect -7239 -3274 -7223 -3240
rect -7189 -3274 -7173 -3240
rect -7121 -3274 -7105 -3240
rect -7071 -3274 -7055 -3240
rect -7003 -3274 -6987 -3240
rect -6953 -3274 -6937 -3240
rect -6885 -3274 -6869 -3240
rect -6835 -3274 -6819 -3240
rect -6767 -3274 -6751 -3240
rect -6717 -3274 -6701 -3240
rect -7400 -3324 -7366 -3308
rect -7400 -3716 -7366 -3700
rect -7282 -3324 -7248 -3308
rect -7282 -3716 -7248 -3700
rect -7164 -3324 -7130 -3308
rect -7164 -3716 -7130 -3700
rect -7046 -3324 -7012 -3308
rect -7046 -3716 -7012 -3700
rect -6928 -3324 -6894 -3308
rect -6928 -3716 -6894 -3700
rect -6810 -3324 -6776 -3308
rect -6810 -3716 -6776 -3700
rect -6692 -3324 -6658 -3308
rect -6692 -3716 -6658 -3700
rect -7357 -3784 -7341 -3750
rect -7307 -3784 -7291 -3750
rect -7239 -3784 -7223 -3750
rect -7189 -3784 -7173 -3750
rect -7121 -3784 -7105 -3750
rect -7071 -3784 -7055 -3750
rect -7003 -3784 -6987 -3750
rect -6953 -3784 -6937 -3750
rect -6885 -3784 -6869 -3750
rect -6835 -3784 -6819 -3750
rect -6767 -3784 -6751 -3750
rect -6717 -3784 -6701 -3750
rect -7514 -3852 -7480 -3790
rect 5056 -3032 5090 -2970
rect 4277 -3072 4293 -3038
rect 4327 -3072 4343 -3038
rect 4395 -3072 4411 -3038
rect 4445 -3072 4461 -3038
rect 4513 -3072 4529 -3038
rect 4563 -3072 4579 -3038
rect 4631 -3072 4647 -3038
rect 4681 -3072 4697 -3038
rect 4749 -3072 4765 -3038
rect 4799 -3072 4815 -3038
rect 4867 -3072 4883 -3038
rect 4917 -3072 4933 -3038
rect 4234 -3122 4268 -3106
rect 4234 -3514 4268 -3498
rect 4352 -3122 4386 -3106
rect 4352 -3514 4386 -3498
rect 4470 -3122 4504 -3106
rect 4470 -3514 4504 -3498
rect 4588 -3122 4622 -3106
rect 4588 -3514 4622 -3498
rect 4706 -3122 4740 -3106
rect 4706 -3514 4740 -3498
rect 4824 -3122 4858 -3106
rect 4824 -3514 4858 -3498
rect 4942 -3122 4976 -3106
rect 4942 -3514 4976 -3498
rect 4277 -3582 4293 -3548
rect 4327 -3582 4343 -3548
rect 4395 -3582 4411 -3548
rect 4445 -3582 4461 -3548
rect 4513 -3582 4529 -3548
rect 4563 -3582 4579 -3548
rect 4631 -3582 4647 -3548
rect 4681 -3582 4697 -3548
rect 4749 -3582 4765 -3548
rect 4799 -3582 4815 -3548
rect 4867 -3582 4883 -3548
rect 4917 -3582 4933 -3548
rect 4120 -3650 4154 -3588
rect 5056 -3650 5090 -3588
rect 4120 -3684 4216 -3650
rect 4994 -3660 5090 -3650
rect 5160 -2970 5256 -2936
rect 6034 -2970 6130 -2936
rect 5160 -3032 5194 -2970
rect 6096 -3032 6130 -2970
rect 5317 -3072 5333 -3038
rect 5367 -3072 5383 -3038
rect 5435 -3072 5451 -3038
rect 5485 -3072 5501 -3038
rect 5553 -3072 5569 -3038
rect 5603 -3072 5619 -3038
rect 5671 -3072 5687 -3038
rect 5721 -3072 5737 -3038
rect 5789 -3072 5805 -3038
rect 5839 -3072 5855 -3038
rect 5907 -3072 5923 -3038
rect 5957 -3072 5973 -3038
rect 5274 -3122 5308 -3106
rect 5274 -3514 5308 -3498
rect 5392 -3122 5426 -3106
rect 5392 -3514 5426 -3498
rect 5510 -3122 5544 -3106
rect 5510 -3514 5544 -3498
rect 5628 -3122 5662 -3106
rect 5628 -3514 5662 -3498
rect 5746 -3122 5780 -3106
rect 5746 -3514 5780 -3498
rect 5864 -3122 5898 -3106
rect 5864 -3514 5898 -3498
rect 5982 -3122 6016 -3106
rect 5982 -3514 6016 -3498
rect 5317 -3582 5333 -3548
rect 5367 -3582 5383 -3548
rect 5435 -3582 5451 -3548
rect 5485 -3582 5501 -3548
rect 5553 -3582 5569 -3548
rect 5603 -3582 5619 -3548
rect 5671 -3582 5687 -3548
rect 5721 -3582 5737 -3548
rect 5789 -3582 5805 -3548
rect 5839 -3582 5855 -3548
rect 5907 -3582 5923 -3548
rect 5957 -3582 5973 -3548
rect 5160 -3650 5194 -3588
rect 6096 -3650 6130 -3588
rect 5160 -3660 5256 -3650
rect 4994 -3684 5256 -3660
rect 6034 -3660 6130 -3650
rect 6200 -2970 6296 -2936
rect 7074 -2970 7170 -2936
rect 6200 -3032 6234 -2970
rect 7136 -3032 7170 -2970
rect 6357 -3072 6373 -3038
rect 6407 -3072 6423 -3038
rect 6475 -3072 6491 -3038
rect 6525 -3072 6541 -3038
rect 6593 -3072 6609 -3038
rect 6643 -3072 6659 -3038
rect 6711 -3072 6727 -3038
rect 6761 -3072 6777 -3038
rect 6829 -3072 6845 -3038
rect 6879 -3072 6895 -3038
rect 6947 -3072 6963 -3038
rect 6997 -3072 7013 -3038
rect 6314 -3122 6348 -3106
rect 6314 -3514 6348 -3498
rect 6432 -3122 6466 -3106
rect 6432 -3514 6466 -3498
rect 6550 -3122 6584 -3106
rect 6550 -3514 6584 -3498
rect 6668 -3122 6702 -3106
rect 6668 -3514 6702 -3498
rect 6786 -3122 6820 -3106
rect 6786 -3514 6820 -3498
rect 6904 -3122 6938 -3106
rect 6904 -3514 6938 -3498
rect 7022 -3122 7056 -3106
rect 7022 -3514 7056 -3498
rect 6357 -3582 6373 -3548
rect 6407 -3582 6423 -3548
rect 6475 -3582 6491 -3548
rect 6525 -3582 6541 -3548
rect 6593 -3582 6609 -3548
rect 6643 -3582 6659 -3548
rect 6711 -3582 6727 -3548
rect 6761 -3582 6777 -3548
rect 6829 -3582 6845 -3548
rect 6879 -3582 6895 -3548
rect 6947 -3582 6963 -3548
rect 6997 -3582 7013 -3548
rect 6200 -3650 6234 -3588
rect 7136 -3650 7170 -3588
rect 6200 -3660 6296 -3650
rect 6034 -3684 6296 -3660
rect 7074 -3660 7170 -3650
rect 7240 -2970 7336 -2936
rect 8114 -2970 8210 -2936
rect 7240 -3032 7274 -2970
rect 8176 -3032 8210 -2970
rect 7397 -3072 7413 -3038
rect 7447 -3072 7463 -3038
rect 7515 -3072 7531 -3038
rect 7565 -3072 7581 -3038
rect 7633 -3072 7649 -3038
rect 7683 -3072 7699 -3038
rect 7751 -3072 7767 -3038
rect 7801 -3072 7817 -3038
rect 7869 -3072 7885 -3038
rect 7919 -3072 7935 -3038
rect 7987 -3072 8003 -3038
rect 8037 -3072 8053 -3038
rect 7354 -3122 7388 -3106
rect 7354 -3514 7388 -3498
rect 7472 -3122 7506 -3106
rect 7472 -3514 7506 -3498
rect 7590 -3122 7624 -3106
rect 7590 -3514 7624 -3498
rect 7708 -3122 7742 -3106
rect 7708 -3514 7742 -3498
rect 7826 -3122 7860 -3106
rect 7826 -3514 7860 -3498
rect 7944 -3122 7978 -3106
rect 7944 -3514 7978 -3498
rect 8062 -3122 8096 -3106
rect 8062 -3514 8096 -3498
rect 7397 -3582 7413 -3548
rect 7447 -3582 7463 -3548
rect 7515 -3582 7531 -3548
rect 7565 -3582 7581 -3548
rect 7633 -3582 7649 -3548
rect 7683 -3582 7699 -3548
rect 7751 -3582 7767 -3548
rect 7801 -3582 7817 -3548
rect 7869 -3582 7885 -3548
rect 7919 -3582 7935 -3548
rect 7987 -3582 8003 -3548
rect 8037 -3582 8053 -3548
rect 7240 -3650 7274 -3588
rect 8176 -3650 8210 -3588
rect 7240 -3660 7336 -3650
rect 7074 -3684 7336 -3660
rect 8114 -3660 8210 -3650
rect 8280 -2970 8376 -2936
rect 9154 -2970 9250 -2936
rect 8280 -3032 8314 -2970
rect 9216 -3032 9250 -2970
rect 8437 -3072 8453 -3038
rect 8487 -3072 8503 -3038
rect 8555 -3072 8571 -3038
rect 8605 -3072 8621 -3038
rect 8673 -3072 8689 -3038
rect 8723 -3072 8739 -3038
rect 8791 -3072 8807 -3038
rect 8841 -3072 8857 -3038
rect 8909 -3072 8925 -3038
rect 8959 -3072 8975 -3038
rect 9027 -3072 9043 -3038
rect 9077 -3072 9093 -3038
rect 8394 -3122 8428 -3106
rect 8394 -3514 8428 -3498
rect 8512 -3122 8546 -3106
rect 8512 -3514 8546 -3498
rect 8630 -3122 8664 -3106
rect 8630 -3514 8664 -3498
rect 8748 -3122 8782 -3106
rect 8748 -3514 8782 -3498
rect 8866 -3122 8900 -3106
rect 8866 -3514 8900 -3498
rect 8984 -3122 9018 -3106
rect 8984 -3514 9018 -3498
rect 9102 -3122 9136 -3106
rect 9102 -3514 9136 -3498
rect 8437 -3582 8453 -3548
rect 8487 -3582 8503 -3548
rect 8555 -3582 8571 -3548
rect 8605 -3582 8621 -3548
rect 8673 -3582 8689 -3548
rect 8723 -3582 8739 -3548
rect 8791 -3582 8807 -3548
rect 8841 -3582 8857 -3548
rect 8909 -3582 8925 -3548
rect 8959 -3582 8975 -3548
rect 9027 -3582 9043 -3548
rect 9077 -3582 9093 -3548
rect 8280 -3650 8314 -3588
rect 9216 -3650 9250 -3588
rect 8280 -3660 8376 -3650
rect 8114 -3684 8376 -3660
rect 9154 -3684 9250 -3650
rect 11740 -2970 11836 -2936
rect 12614 -2970 12710 -2936
rect 11740 -3032 11774 -2970
rect 12676 -3032 12710 -2970
rect 11897 -3072 11913 -3038
rect 11947 -3072 11963 -3038
rect 12015 -3072 12031 -3038
rect 12065 -3072 12081 -3038
rect 12133 -3072 12149 -3038
rect 12183 -3072 12199 -3038
rect 12251 -3072 12267 -3038
rect 12301 -3072 12317 -3038
rect 12369 -3072 12385 -3038
rect 12419 -3072 12435 -3038
rect 12487 -3072 12503 -3038
rect 12537 -3072 12553 -3038
rect 11854 -3122 11888 -3106
rect 11854 -3514 11888 -3498
rect 11972 -3122 12006 -3106
rect 11972 -3514 12006 -3498
rect 12090 -3122 12124 -3106
rect 12090 -3514 12124 -3498
rect 12208 -3122 12242 -3106
rect 12208 -3514 12242 -3498
rect 12326 -3122 12360 -3106
rect 12326 -3514 12360 -3498
rect 12444 -3122 12478 -3106
rect 12444 -3514 12478 -3498
rect 12562 -3122 12596 -3106
rect 12562 -3514 12596 -3498
rect 11897 -3582 11913 -3548
rect 11947 -3582 11963 -3548
rect 12015 -3582 12031 -3548
rect 12065 -3582 12081 -3548
rect 12133 -3582 12149 -3548
rect 12183 -3582 12199 -3548
rect 12251 -3582 12267 -3548
rect 12301 -3582 12317 -3548
rect 12369 -3582 12385 -3548
rect 12419 -3582 12435 -3548
rect 12487 -3582 12503 -3548
rect 12537 -3582 12553 -3548
rect 11740 -3650 11774 -3588
rect 12676 -3650 12710 -3588
rect 11740 -3684 11836 -3650
rect 12614 -3660 12710 -3650
rect 12780 -2970 12876 -2936
rect 13654 -2970 13750 -2936
rect 12780 -3032 12814 -2970
rect 13716 -3032 13750 -2970
rect 12937 -3072 12953 -3038
rect 12987 -3072 13003 -3038
rect 13055 -3072 13071 -3038
rect 13105 -3072 13121 -3038
rect 13173 -3072 13189 -3038
rect 13223 -3072 13239 -3038
rect 13291 -3072 13307 -3038
rect 13341 -3072 13357 -3038
rect 13409 -3072 13425 -3038
rect 13459 -3072 13475 -3038
rect 13527 -3072 13543 -3038
rect 13577 -3072 13593 -3038
rect 12894 -3122 12928 -3106
rect 12894 -3514 12928 -3498
rect 13012 -3122 13046 -3106
rect 13012 -3514 13046 -3498
rect 13130 -3122 13164 -3106
rect 13130 -3514 13164 -3498
rect 13248 -3122 13282 -3106
rect 13248 -3514 13282 -3498
rect 13366 -3122 13400 -3106
rect 13366 -3514 13400 -3498
rect 13484 -3122 13518 -3106
rect 13484 -3514 13518 -3498
rect 13602 -3122 13636 -3106
rect 13602 -3514 13636 -3498
rect 12937 -3582 12953 -3548
rect 12987 -3582 13003 -3548
rect 13055 -3582 13071 -3548
rect 13105 -3582 13121 -3548
rect 13173 -3582 13189 -3548
rect 13223 -3582 13239 -3548
rect 13291 -3582 13307 -3548
rect 13341 -3582 13357 -3548
rect 13409 -3582 13425 -3548
rect 13459 -3582 13475 -3548
rect 13527 -3582 13543 -3548
rect 13577 -3582 13593 -3548
rect 12780 -3650 12814 -3588
rect 13716 -3650 13750 -3588
rect 12780 -3660 12876 -3650
rect 12614 -3684 12876 -3660
rect 13654 -3660 13750 -3650
rect 13820 -2970 13916 -2936
rect 14694 -2970 14790 -2936
rect 13820 -3032 13854 -2970
rect 14756 -3032 14790 -2970
rect 13977 -3072 13993 -3038
rect 14027 -3072 14043 -3038
rect 14095 -3072 14111 -3038
rect 14145 -3072 14161 -3038
rect 14213 -3072 14229 -3038
rect 14263 -3072 14279 -3038
rect 14331 -3072 14347 -3038
rect 14381 -3072 14397 -3038
rect 14449 -3072 14465 -3038
rect 14499 -3072 14515 -3038
rect 14567 -3072 14583 -3038
rect 14617 -3072 14633 -3038
rect 13934 -3122 13968 -3106
rect 13934 -3514 13968 -3498
rect 14052 -3122 14086 -3106
rect 14052 -3514 14086 -3498
rect 14170 -3122 14204 -3106
rect 14170 -3514 14204 -3498
rect 14288 -3122 14322 -3106
rect 14288 -3514 14322 -3498
rect 14406 -3122 14440 -3106
rect 14406 -3514 14440 -3498
rect 14524 -3122 14558 -3106
rect 14524 -3514 14558 -3498
rect 14642 -3122 14676 -3106
rect 14642 -3514 14676 -3498
rect 13977 -3582 13993 -3548
rect 14027 -3582 14043 -3548
rect 14095 -3582 14111 -3548
rect 14145 -3582 14161 -3548
rect 14213 -3582 14229 -3548
rect 14263 -3582 14279 -3548
rect 14331 -3582 14347 -3548
rect 14381 -3582 14397 -3548
rect 14449 -3582 14465 -3548
rect 14499 -3582 14515 -3548
rect 14567 -3582 14583 -3548
rect 14617 -3582 14633 -3548
rect 13820 -3650 13854 -3588
rect 14756 -3650 14790 -3588
rect 13820 -3660 13916 -3650
rect 13654 -3684 13916 -3660
rect 14694 -3660 14790 -3650
rect 14860 -2970 14956 -2936
rect 15734 -2970 15830 -2936
rect 14860 -3032 14894 -2970
rect 15796 -3032 15830 -2970
rect 15017 -3072 15033 -3038
rect 15067 -3072 15083 -3038
rect 15135 -3072 15151 -3038
rect 15185 -3072 15201 -3038
rect 15253 -3072 15269 -3038
rect 15303 -3072 15319 -3038
rect 15371 -3072 15387 -3038
rect 15421 -3072 15437 -3038
rect 15489 -3072 15505 -3038
rect 15539 -3072 15555 -3038
rect 15607 -3072 15623 -3038
rect 15657 -3072 15673 -3038
rect 14974 -3122 15008 -3106
rect 14974 -3514 15008 -3498
rect 15092 -3122 15126 -3106
rect 15092 -3514 15126 -3498
rect 15210 -3122 15244 -3106
rect 15210 -3514 15244 -3498
rect 15328 -3122 15362 -3106
rect 15328 -3514 15362 -3498
rect 15446 -3122 15480 -3106
rect 15446 -3514 15480 -3498
rect 15564 -3122 15598 -3106
rect 15564 -3514 15598 -3498
rect 15682 -3122 15716 -3106
rect 15682 -3514 15716 -3498
rect 15017 -3582 15033 -3548
rect 15067 -3582 15083 -3548
rect 15135 -3582 15151 -3548
rect 15185 -3582 15201 -3548
rect 15253 -3582 15269 -3548
rect 15303 -3582 15319 -3548
rect 15371 -3582 15387 -3548
rect 15421 -3582 15437 -3548
rect 15489 -3582 15505 -3548
rect 15539 -3582 15555 -3548
rect 15607 -3582 15623 -3548
rect 15657 -3582 15673 -3548
rect 14860 -3650 14894 -3588
rect 15796 -3650 15830 -3588
rect 14860 -3660 14956 -3650
rect 14694 -3684 14956 -3660
rect 15734 -3660 15830 -3650
rect 15900 -2970 15996 -2936
rect 16774 -2970 16870 -2936
rect 15900 -3032 15934 -2970
rect 16836 -3032 16870 -2970
rect 16057 -3072 16073 -3038
rect 16107 -3072 16123 -3038
rect 16175 -3072 16191 -3038
rect 16225 -3072 16241 -3038
rect 16293 -3072 16309 -3038
rect 16343 -3072 16359 -3038
rect 16411 -3072 16427 -3038
rect 16461 -3072 16477 -3038
rect 16529 -3072 16545 -3038
rect 16579 -3072 16595 -3038
rect 16647 -3072 16663 -3038
rect 16697 -3072 16713 -3038
rect 16014 -3122 16048 -3106
rect 16014 -3514 16048 -3498
rect 16132 -3122 16166 -3106
rect 16132 -3514 16166 -3498
rect 16250 -3122 16284 -3106
rect 16250 -3514 16284 -3498
rect 16368 -3122 16402 -3106
rect 16368 -3514 16402 -3498
rect 16486 -3122 16520 -3106
rect 16486 -3514 16520 -3498
rect 16604 -3122 16638 -3106
rect 16604 -3514 16638 -3498
rect 16722 -3122 16756 -3106
rect 16722 -3514 16756 -3498
rect 16057 -3582 16073 -3548
rect 16107 -3582 16123 -3548
rect 16175 -3582 16191 -3548
rect 16225 -3582 16241 -3548
rect 16293 -3582 16309 -3548
rect 16343 -3582 16359 -3548
rect 16411 -3582 16427 -3548
rect 16461 -3582 16477 -3548
rect 16529 -3582 16545 -3548
rect 16579 -3582 16595 -3548
rect 16647 -3582 16663 -3548
rect 16697 -3582 16713 -3548
rect 15900 -3650 15934 -3588
rect 16836 -3650 16870 -3588
rect 15900 -3660 15996 -3650
rect 15734 -3684 15996 -3660
rect 16774 -3684 16870 -3650
rect 4124 -3720 9244 -3684
rect 4124 -3760 4924 -3720
rect -6578 -3852 -6544 -3790
rect 5224 -3760 8564 -3720
rect 8864 -3760 9244 -3720
rect 11744 -3720 16864 -3684
rect 11744 -3760 12544 -3720
rect 12844 -3760 16184 -3720
rect 16484 -3760 16864 -3720
rect -7514 -3886 -7418 -3852
rect -6640 -3886 -6544 -3852
<< viali >>
rect -1418 6187 -1168 6584
rect -1040 6187 -790 6584
rect -662 6187 -412 6584
rect -284 6187 -34 6584
rect 94 6187 344 6584
rect -1418 5356 -1168 5753
rect -1040 5356 -790 5753
rect -662 5356 -412 5753
rect -284 5356 -34 5753
rect 94 5356 344 5753
rect -1418 4819 -1168 5216
rect -1040 4819 -790 5216
rect -662 4819 -412 5216
rect -284 4819 -34 5216
rect 94 4819 344 5216
rect -1418 3988 -1168 4385
rect -1040 3988 -790 4385
rect -662 3988 -412 4385
rect -284 3988 -34 4385
rect 94 3988 344 4385
rect 1382 6187 1632 6584
rect 1760 6187 2010 6584
rect 2138 6187 2388 6584
rect 2516 6187 2766 6584
rect 2894 6187 3144 6584
rect 1382 5356 1632 5753
rect 1760 5356 2010 5753
rect 2138 5356 2388 5753
rect 2516 5356 2766 5753
rect 2894 5356 3144 5753
rect 1382 4819 1632 5216
rect 1760 4819 2010 5216
rect 2138 4819 2388 5216
rect 2516 4819 2766 5216
rect 2894 4819 3144 5216
rect 1382 3988 1632 4385
rect 1760 3988 2010 4385
rect 2138 3988 2388 4385
rect 2516 3988 2766 4385
rect 2894 3988 3144 4385
rect -886 3648 -852 3682
rect -694 3648 -660 3682
rect -502 3648 -468 3682
rect -310 3648 -276 3682
rect -118 3648 -84 3682
rect -1030 3222 -996 3598
rect -934 3222 -900 3598
rect -838 3222 -804 3598
rect -742 3222 -708 3598
rect -646 3222 -612 3598
rect -550 3222 -516 3598
rect -454 3222 -420 3598
rect -358 3222 -324 3598
rect -262 3222 -228 3598
rect -166 3222 -132 3598
rect -70 3222 -36 3598
rect -982 3138 -948 3172
rect -790 3138 -756 3172
rect -598 3138 -564 3172
rect -406 3138 -372 3172
rect -214 3138 -180 3172
rect 1914 3648 1948 3682
rect 2106 3648 2140 3682
rect 2298 3648 2332 3682
rect 2490 3648 2524 3682
rect 2682 3648 2716 3682
rect 1770 3222 1804 3598
rect 1866 3222 1900 3598
rect 1962 3222 1996 3598
rect 2058 3222 2092 3598
rect 2154 3222 2188 3598
rect 2250 3222 2284 3598
rect 2346 3222 2380 3598
rect 2442 3222 2476 3598
rect 2538 3222 2572 3598
rect 2634 3222 2668 3598
rect 2730 3222 2764 3598
rect 1818 3138 1852 3172
rect 2010 3138 2044 3172
rect 2202 3138 2236 3172
rect 2394 3138 2428 3172
rect 2586 3138 2620 3172
rect 4482 5502 4516 5536
rect 4674 5502 4708 5536
rect 4866 5502 4900 5536
rect 5058 5502 5092 5536
rect 5250 5502 5284 5536
rect 5442 5502 5476 5536
rect 5634 5502 5668 5536
rect 5826 5502 5860 5536
rect 6018 5502 6052 5536
rect 6210 5502 6244 5536
rect 6402 5502 6436 5536
rect 6594 5502 6628 5536
rect 6786 5502 6820 5536
rect 6978 5502 7012 5536
rect 7170 5502 7204 5536
rect 4434 5076 4468 5452
rect 4530 5076 4564 5452
rect 4626 5076 4660 5452
rect 4722 5076 4756 5452
rect 4818 5076 4852 5452
rect 4914 5076 4948 5452
rect 5010 5076 5044 5452
rect 5106 5076 5140 5452
rect 5202 5076 5236 5452
rect 5298 5076 5332 5452
rect 5394 5076 5428 5452
rect 5490 5076 5524 5452
rect 5586 5076 5620 5452
rect 5682 5076 5716 5452
rect 5778 5076 5812 5452
rect 5874 5076 5908 5452
rect 5970 5076 6004 5452
rect 6066 5076 6100 5452
rect 6162 5076 6196 5452
rect 6258 5076 6292 5452
rect 6354 5076 6388 5452
rect 6450 5076 6484 5452
rect 6546 5076 6580 5452
rect 6642 5076 6676 5452
rect 6738 5076 6772 5452
rect 6834 5076 6868 5452
rect 6930 5076 6964 5452
rect 7026 5076 7060 5452
rect 7122 5076 7156 5452
rect 7218 5076 7252 5452
rect 7314 5076 7348 5452
rect 4578 4992 4612 5026
rect 4770 4992 4804 5026
rect 4962 4992 4996 5026
rect 5154 4992 5188 5026
rect 5346 4992 5380 5026
rect 5538 4992 5572 5026
rect 5730 4992 5764 5026
rect 5922 4992 5956 5026
rect 6114 4992 6148 5026
rect 6306 4992 6340 5026
rect 6498 4992 6532 5026
rect 6690 4992 6724 5026
rect 6882 4992 6916 5026
rect 7074 4992 7108 5026
rect 7266 4992 7300 5026
rect 4578 4884 4612 4918
rect 4770 4884 4804 4918
rect 4962 4884 4996 4918
rect 5154 4884 5188 4918
rect 5346 4884 5380 4918
rect 5538 4884 5572 4918
rect 5730 4884 5764 4918
rect 5922 4884 5956 4918
rect 6114 4884 6148 4918
rect 6306 4884 6340 4918
rect 6498 4884 6532 4918
rect 6690 4884 6724 4918
rect 6882 4884 6916 4918
rect 7074 4884 7108 4918
rect 7266 4884 7300 4918
rect 4434 4458 4468 4834
rect 4530 4458 4564 4834
rect 4626 4458 4660 4834
rect 4722 4458 4756 4834
rect 4818 4458 4852 4834
rect 4914 4458 4948 4834
rect 5010 4458 5044 4834
rect 5106 4458 5140 4834
rect 5202 4458 5236 4834
rect 5298 4458 5332 4834
rect 5394 4458 5428 4834
rect 5490 4458 5524 4834
rect 5586 4458 5620 4834
rect 5682 4458 5716 4834
rect 5778 4458 5812 4834
rect 5874 4458 5908 4834
rect 5970 4458 6004 4834
rect 6066 4458 6100 4834
rect 6162 4458 6196 4834
rect 6258 4458 6292 4834
rect 6354 4458 6388 4834
rect 6450 4458 6484 4834
rect 6546 4458 6580 4834
rect 6642 4458 6676 4834
rect 6738 4458 6772 4834
rect 6834 4458 6868 4834
rect 6930 4458 6964 4834
rect 7026 4458 7060 4834
rect 7122 4458 7156 4834
rect 7218 4458 7252 4834
rect 7314 4458 7348 4834
rect 4482 4374 4516 4408
rect 4674 4374 4708 4408
rect 4866 4374 4900 4408
rect 5058 4374 5092 4408
rect 5250 4374 5284 4408
rect 5442 4374 5476 4408
rect 5634 4374 5668 4408
rect 5826 4374 5860 4408
rect 6018 4374 6052 4408
rect 6210 4374 6244 4408
rect 6402 4374 6436 4408
rect 6594 4374 6628 4408
rect 6786 4374 6820 4408
rect 6978 4374 7012 4408
rect 7170 4374 7204 4408
rect 4482 4266 4516 4300
rect 4674 4266 4708 4300
rect 4866 4266 4900 4300
rect 5058 4266 5092 4300
rect 5250 4266 5284 4300
rect 5442 4266 5476 4300
rect 5634 4266 5668 4300
rect 5826 4266 5860 4300
rect 6018 4266 6052 4300
rect 6210 4266 6244 4300
rect 6402 4266 6436 4300
rect 6594 4266 6628 4300
rect 6786 4266 6820 4300
rect 6978 4266 7012 4300
rect 7170 4266 7204 4300
rect 4434 3840 4468 4216
rect 4530 3840 4564 4216
rect 4626 3840 4660 4216
rect 4722 3840 4756 4216
rect 4818 3840 4852 4216
rect 4914 3840 4948 4216
rect 5010 3840 5044 4216
rect 5106 3840 5140 4216
rect 5202 3840 5236 4216
rect 5298 3840 5332 4216
rect 5394 3840 5428 4216
rect 5490 3840 5524 4216
rect 5586 3840 5620 4216
rect 5682 3840 5716 4216
rect 5778 3840 5812 4216
rect 5874 3840 5908 4216
rect 5970 3840 6004 4216
rect 6066 3840 6100 4216
rect 6162 3840 6196 4216
rect 6258 3840 6292 4216
rect 6354 3840 6388 4216
rect 6450 3840 6484 4216
rect 6546 3840 6580 4216
rect 6642 3840 6676 4216
rect 6738 3840 6772 4216
rect 6834 3840 6868 4216
rect 6930 3840 6964 4216
rect 7026 3840 7060 4216
rect 7122 3840 7156 4216
rect 7218 3840 7252 4216
rect 7314 3840 7348 4216
rect 4578 3756 4612 3790
rect 4770 3756 4804 3790
rect 4962 3756 4996 3790
rect 5154 3756 5188 3790
rect 5346 3756 5380 3790
rect 5538 3756 5572 3790
rect 5730 3756 5764 3790
rect 5922 3756 5956 3790
rect 6114 3756 6148 3790
rect 6306 3756 6340 3790
rect 6498 3756 6532 3790
rect 6690 3756 6724 3790
rect 6882 3756 6916 3790
rect 7074 3756 7108 3790
rect 7266 3756 7300 3790
rect 4578 3648 4612 3682
rect 4770 3648 4804 3682
rect 4962 3648 4996 3682
rect 5154 3648 5188 3682
rect 5346 3648 5380 3682
rect 5538 3648 5572 3682
rect 5730 3648 5764 3682
rect 5922 3648 5956 3682
rect 6114 3648 6148 3682
rect 6306 3648 6340 3682
rect 6498 3648 6532 3682
rect 6690 3648 6724 3682
rect 6882 3648 6916 3682
rect 7074 3648 7108 3682
rect 7266 3648 7300 3682
rect 4434 3222 4468 3598
rect 4530 3222 4564 3598
rect 4626 3222 4660 3598
rect 4722 3222 4756 3598
rect 4818 3222 4852 3598
rect 4914 3222 4948 3598
rect 5010 3222 5044 3598
rect 5106 3222 5140 3598
rect 5202 3222 5236 3598
rect 5298 3222 5332 3598
rect 5394 3222 5428 3598
rect 5490 3222 5524 3598
rect 5586 3222 5620 3598
rect 5682 3222 5716 3598
rect 5778 3222 5812 3598
rect 5874 3222 5908 3598
rect 5970 3222 6004 3598
rect 6066 3222 6100 3598
rect 6162 3222 6196 3598
rect 6258 3222 6292 3598
rect 6354 3222 6388 3598
rect 6450 3222 6484 3598
rect 6546 3222 6580 3598
rect 6642 3222 6676 3598
rect 6738 3222 6772 3598
rect 6834 3222 6868 3598
rect 6930 3222 6964 3598
rect 7026 3222 7060 3598
rect 7122 3222 7156 3598
rect 7218 3222 7252 3598
rect 7314 3222 7348 3598
rect 4482 3138 4516 3172
rect 4674 3138 4708 3172
rect 4866 3138 4900 3172
rect 5058 3138 5092 3172
rect 5250 3138 5284 3172
rect 5442 3138 5476 3172
rect 5634 3138 5668 3172
rect 5826 3138 5860 3172
rect 6018 3138 6052 3172
rect 6210 3138 6244 3172
rect 6402 3138 6436 3172
rect 6594 3138 6628 3172
rect 6786 3138 6820 3172
rect 6978 3138 7012 3172
rect 7170 3138 7204 3172
rect 8122 5502 8156 5536
rect 8314 5502 8348 5536
rect 8506 5502 8540 5536
rect 8698 5502 8732 5536
rect 8890 5502 8924 5536
rect 9082 5502 9116 5536
rect 9274 5502 9308 5536
rect 9466 5502 9500 5536
rect 9658 5502 9692 5536
rect 9850 5502 9884 5536
rect 10042 5502 10076 5536
rect 10234 5502 10268 5536
rect 10426 5502 10460 5536
rect 10618 5502 10652 5536
rect 10810 5502 10844 5536
rect 8074 5076 8108 5452
rect 8170 5076 8204 5452
rect 8266 5076 8300 5452
rect 8362 5076 8396 5452
rect 8458 5076 8492 5452
rect 8554 5076 8588 5452
rect 8650 5076 8684 5452
rect 8746 5076 8780 5452
rect 8842 5076 8876 5452
rect 8938 5076 8972 5452
rect 9034 5076 9068 5452
rect 9130 5076 9164 5452
rect 9226 5076 9260 5452
rect 9322 5076 9356 5452
rect 9418 5076 9452 5452
rect 9514 5076 9548 5452
rect 9610 5076 9644 5452
rect 9706 5076 9740 5452
rect 9802 5076 9836 5452
rect 9898 5076 9932 5452
rect 9994 5076 10028 5452
rect 10090 5076 10124 5452
rect 10186 5076 10220 5452
rect 10282 5076 10316 5452
rect 10378 5076 10412 5452
rect 10474 5076 10508 5452
rect 10570 5076 10604 5452
rect 10666 5076 10700 5452
rect 10762 5076 10796 5452
rect 10858 5076 10892 5452
rect 10954 5076 10988 5452
rect 8218 4992 8252 5026
rect 8410 4992 8444 5026
rect 8602 4992 8636 5026
rect 8794 4992 8828 5026
rect 8986 4992 9020 5026
rect 9178 4992 9212 5026
rect 9370 4992 9404 5026
rect 9562 4992 9596 5026
rect 9754 4992 9788 5026
rect 9946 4992 9980 5026
rect 10138 4992 10172 5026
rect 10330 4992 10364 5026
rect 10522 4992 10556 5026
rect 10714 4992 10748 5026
rect 10906 4992 10940 5026
rect 8218 4884 8252 4918
rect 8410 4884 8444 4918
rect 8602 4884 8636 4918
rect 8794 4884 8828 4918
rect 8986 4884 9020 4918
rect 9178 4884 9212 4918
rect 9370 4884 9404 4918
rect 9562 4884 9596 4918
rect 9754 4884 9788 4918
rect 9946 4884 9980 4918
rect 10138 4884 10172 4918
rect 10330 4884 10364 4918
rect 10522 4884 10556 4918
rect 10714 4884 10748 4918
rect 10906 4884 10940 4918
rect 8074 4458 8108 4834
rect 8170 4458 8204 4834
rect 8266 4458 8300 4834
rect 8362 4458 8396 4834
rect 8458 4458 8492 4834
rect 8554 4458 8588 4834
rect 8650 4458 8684 4834
rect 8746 4458 8780 4834
rect 8842 4458 8876 4834
rect 8938 4458 8972 4834
rect 9034 4458 9068 4834
rect 9130 4458 9164 4834
rect 9226 4458 9260 4834
rect 9322 4458 9356 4834
rect 9418 4458 9452 4834
rect 9514 4458 9548 4834
rect 9610 4458 9644 4834
rect 9706 4458 9740 4834
rect 9802 4458 9836 4834
rect 9898 4458 9932 4834
rect 9994 4458 10028 4834
rect 10090 4458 10124 4834
rect 10186 4458 10220 4834
rect 10282 4458 10316 4834
rect 10378 4458 10412 4834
rect 10474 4458 10508 4834
rect 10570 4458 10604 4834
rect 10666 4458 10700 4834
rect 10762 4458 10796 4834
rect 10858 4458 10892 4834
rect 10954 4458 10988 4834
rect 8122 4374 8156 4408
rect 8314 4374 8348 4408
rect 8506 4374 8540 4408
rect 8698 4374 8732 4408
rect 8890 4374 8924 4408
rect 9082 4374 9116 4408
rect 9274 4374 9308 4408
rect 9466 4374 9500 4408
rect 9658 4374 9692 4408
rect 9850 4374 9884 4408
rect 10042 4374 10076 4408
rect 10234 4374 10268 4408
rect 10426 4374 10460 4408
rect 10618 4374 10652 4408
rect 10810 4374 10844 4408
rect 8122 4266 8156 4300
rect 8314 4266 8348 4300
rect 8506 4266 8540 4300
rect 8698 4266 8732 4300
rect 8890 4266 8924 4300
rect 9082 4266 9116 4300
rect 9274 4266 9308 4300
rect 9466 4266 9500 4300
rect 9658 4266 9692 4300
rect 9850 4266 9884 4300
rect 10042 4266 10076 4300
rect 10234 4266 10268 4300
rect 10426 4266 10460 4300
rect 10618 4266 10652 4300
rect 10810 4266 10844 4300
rect 8074 3840 8108 4216
rect 8170 3840 8204 4216
rect 8266 3840 8300 4216
rect 8362 3840 8396 4216
rect 8458 3840 8492 4216
rect 8554 3840 8588 4216
rect 8650 3840 8684 4216
rect 8746 3840 8780 4216
rect 8842 3840 8876 4216
rect 8938 3840 8972 4216
rect 9034 3840 9068 4216
rect 9130 3840 9164 4216
rect 9226 3840 9260 4216
rect 9322 3840 9356 4216
rect 9418 3840 9452 4216
rect 9514 3840 9548 4216
rect 9610 3840 9644 4216
rect 9706 3840 9740 4216
rect 9802 3840 9836 4216
rect 9898 3840 9932 4216
rect 9994 3840 10028 4216
rect 10090 3840 10124 4216
rect 10186 3840 10220 4216
rect 10282 3840 10316 4216
rect 10378 3840 10412 4216
rect 10474 3840 10508 4216
rect 10570 3840 10604 4216
rect 10666 3840 10700 4216
rect 10762 3840 10796 4216
rect 10858 3840 10892 4216
rect 10954 3840 10988 4216
rect 8218 3756 8252 3790
rect 8410 3756 8444 3790
rect 8602 3756 8636 3790
rect 8794 3756 8828 3790
rect 8986 3756 9020 3790
rect 9178 3756 9212 3790
rect 9370 3756 9404 3790
rect 9562 3756 9596 3790
rect 9754 3756 9788 3790
rect 9946 3756 9980 3790
rect 10138 3756 10172 3790
rect 10330 3756 10364 3790
rect 10522 3756 10556 3790
rect 10714 3756 10748 3790
rect 10906 3756 10940 3790
rect 8218 3648 8252 3682
rect 8410 3648 8444 3682
rect 8602 3648 8636 3682
rect 8794 3648 8828 3682
rect 8986 3648 9020 3682
rect 9178 3648 9212 3682
rect 9370 3648 9404 3682
rect 9562 3648 9596 3682
rect 9754 3648 9788 3682
rect 9946 3648 9980 3682
rect 10138 3648 10172 3682
rect 10330 3648 10364 3682
rect 10522 3648 10556 3682
rect 10714 3648 10748 3682
rect 10906 3648 10940 3682
rect 8074 3222 8108 3598
rect 8170 3222 8204 3598
rect 8266 3222 8300 3598
rect 8362 3222 8396 3598
rect 8458 3222 8492 3598
rect 8554 3222 8588 3598
rect 8650 3222 8684 3598
rect 8746 3222 8780 3598
rect 8842 3222 8876 3598
rect 8938 3222 8972 3598
rect 9034 3222 9068 3598
rect 9130 3222 9164 3598
rect 9226 3222 9260 3598
rect 9322 3222 9356 3598
rect 9418 3222 9452 3598
rect 9514 3222 9548 3598
rect 9610 3222 9644 3598
rect 9706 3222 9740 3598
rect 9802 3222 9836 3598
rect 9898 3222 9932 3598
rect 9994 3222 10028 3598
rect 10090 3222 10124 3598
rect 10186 3222 10220 3598
rect 10282 3222 10316 3598
rect 10378 3222 10412 3598
rect 10474 3222 10508 3598
rect 10570 3222 10604 3598
rect 10666 3222 10700 3598
rect 10762 3222 10796 3598
rect 10858 3222 10892 3598
rect 10954 3222 10988 3598
rect 8122 3138 8156 3172
rect 8314 3138 8348 3172
rect 8506 3138 8540 3172
rect 8698 3138 8732 3172
rect 8890 3138 8924 3172
rect 9082 3138 9116 3172
rect 9274 3138 9308 3172
rect 9466 3138 9500 3172
rect 9658 3138 9692 3172
rect 9850 3138 9884 3172
rect 10042 3138 10076 3172
rect 10234 3138 10268 3172
rect 10426 3138 10460 3172
rect 10618 3138 10652 3172
rect 10810 3138 10844 3172
rect 12102 5502 12136 5536
rect 12294 5502 12328 5536
rect 12486 5502 12520 5536
rect 12678 5502 12712 5536
rect 12870 5502 12904 5536
rect 13062 5502 13096 5536
rect 13254 5502 13288 5536
rect 13446 5502 13480 5536
rect 13638 5502 13672 5536
rect 13830 5502 13864 5536
rect 14022 5502 14056 5536
rect 14214 5502 14248 5536
rect 14406 5502 14440 5536
rect 14598 5502 14632 5536
rect 14790 5502 14824 5536
rect 12054 5076 12088 5452
rect 12150 5076 12184 5452
rect 12246 5076 12280 5452
rect 12342 5076 12376 5452
rect 12438 5076 12472 5452
rect 12534 5076 12568 5452
rect 12630 5076 12664 5452
rect 12726 5076 12760 5452
rect 12822 5076 12856 5452
rect 12918 5076 12952 5452
rect 13014 5076 13048 5452
rect 13110 5076 13144 5452
rect 13206 5076 13240 5452
rect 13302 5076 13336 5452
rect 13398 5076 13432 5452
rect 13494 5076 13528 5452
rect 13590 5076 13624 5452
rect 13686 5076 13720 5452
rect 13782 5076 13816 5452
rect 13878 5076 13912 5452
rect 13974 5076 14008 5452
rect 14070 5076 14104 5452
rect 14166 5076 14200 5452
rect 14262 5076 14296 5452
rect 14358 5076 14392 5452
rect 14454 5076 14488 5452
rect 14550 5076 14584 5452
rect 14646 5076 14680 5452
rect 14742 5076 14776 5452
rect 14838 5076 14872 5452
rect 14934 5076 14968 5452
rect 12198 4992 12232 5026
rect 12390 4992 12424 5026
rect 12582 4992 12616 5026
rect 12774 4992 12808 5026
rect 12966 4992 13000 5026
rect 13158 4992 13192 5026
rect 13350 4992 13384 5026
rect 13542 4992 13576 5026
rect 13734 4992 13768 5026
rect 13926 4992 13960 5026
rect 14118 4992 14152 5026
rect 14310 4992 14344 5026
rect 14502 4992 14536 5026
rect 14694 4992 14728 5026
rect 14886 4992 14920 5026
rect 12198 4884 12232 4918
rect 12390 4884 12424 4918
rect 12582 4884 12616 4918
rect 12774 4884 12808 4918
rect 12966 4884 13000 4918
rect 13158 4884 13192 4918
rect 13350 4884 13384 4918
rect 13542 4884 13576 4918
rect 13734 4884 13768 4918
rect 13926 4884 13960 4918
rect 14118 4884 14152 4918
rect 14310 4884 14344 4918
rect 14502 4884 14536 4918
rect 14694 4884 14728 4918
rect 14886 4884 14920 4918
rect 12054 4458 12088 4834
rect 12150 4458 12184 4834
rect 12246 4458 12280 4834
rect 12342 4458 12376 4834
rect 12438 4458 12472 4834
rect 12534 4458 12568 4834
rect 12630 4458 12664 4834
rect 12726 4458 12760 4834
rect 12822 4458 12856 4834
rect 12918 4458 12952 4834
rect 13014 4458 13048 4834
rect 13110 4458 13144 4834
rect 13206 4458 13240 4834
rect 13302 4458 13336 4834
rect 13398 4458 13432 4834
rect 13494 4458 13528 4834
rect 13590 4458 13624 4834
rect 13686 4458 13720 4834
rect 13782 4458 13816 4834
rect 13878 4458 13912 4834
rect 13974 4458 14008 4834
rect 14070 4458 14104 4834
rect 14166 4458 14200 4834
rect 14262 4458 14296 4834
rect 14358 4458 14392 4834
rect 14454 4458 14488 4834
rect 14550 4458 14584 4834
rect 14646 4458 14680 4834
rect 14742 4458 14776 4834
rect 14838 4458 14872 4834
rect 14934 4458 14968 4834
rect 12102 4374 12136 4408
rect 12294 4374 12328 4408
rect 12486 4374 12520 4408
rect 12678 4374 12712 4408
rect 12870 4374 12904 4408
rect 13062 4374 13096 4408
rect 13254 4374 13288 4408
rect 13446 4374 13480 4408
rect 13638 4374 13672 4408
rect 13830 4374 13864 4408
rect 14022 4374 14056 4408
rect 14214 4374 14248 4408
rect 14406 4374 14440 4408
rect 14598 4374 14632 4408
rect 14790 4374 14824 4408
rect 12102 4266 12136 4300
rect 12294 4266 12328 4300
rect 12486 4266 12520 4300
rect 12678 4266 12712 4300
rect 12870 4266 12904 4300
rect 13062 4266 13096 4300
rect 13254 4266 13288 4300
rect 13446 4266 13480 4300
rect 13638 4266 13672 4300
rect 13830 4266 13864 4300
rect 14022 4266 14056 4300
rect 14214 4266 14248 4300
rect 14406 4266 14440 4300
rect 14598 4266 14632 4300
rect 14790 4266 14824 4300
rect 12054 3840 12088 4216
rect 12150 3840 12184 4216
rect 12246 3840 12280 4216
rect 12342 3840 12376 4216
rect 12438 3840 12472 4216
rect 12534 3840 12568 4216
rect 12630 3840 12664 4216
rect 12726 3840 12760 4216
rect 12822 3840 12856 4216
rect 12918 3840 12952 4216
rect 13014 3840 13048 4216
rect 13110 3840 13144 4216
rect 13206 3840 13240 4216
rect 13302 3840 13336 4216
rect 13398 3840 13432 4216
rect 13494 3840 13528 4216
rect 13590 3840 13624 4216
rect 13686 3840 13720 4216
rect 13782 3840 13816 4216
rect 13878 3840 13912 4216
rect 13974 3840 14008 4216
rect 14070 3840 14104 4216
rect 14166 3840 14200 4216
rect 14262 3840 14296 4216
rect 14358 3840 14392 4216
rect 14454 3840 14488 4216
rect 14550 3840 14584 4216
rect 14646 3840 14680 4216
rect 14742 3840 14776 4216
rect 14838 3840 14872 4216
rect 14934 3840 14968 4216
rect 12198 3756 12232 3790
rect 12390 3756 12424 3790
rect 12582 3756 12616 3790
rect 12774 3756 12808 3790
rect 12966 3756 13000 3790
rect 13158 3756 13192 3790
rect 13350 3756 13384 3790
rect 13542 3756 13576 3790
rect 13734 3756 13768 3790
rect 13926 3756 13960 3790
rect 14118 3756 14152 3790
rect 14310 3756 14344 3790
rect 14502 3756 14536 3790
rect 14694 3756 14728 3790
rect 14886 3756 14920 3790
rect 12198 3648 12232 3682
rect 12390 3648 12424 3682
rect 12582 3648 12616 3682
rect 12774 3648 12808 3682
rect 12966 3648 13000 3682
rect 13158 3648 13192 3682
rect 13350 3648 13384 3682
rect 13542 3648 13576 3682
rect 13734 3648 13768 3682
rect 13926 3648 13960 3682
rect 14118 3648 14152 3682
rect 14310 3648 14344 3682
rect 14502 3648 14536 3682
rect 14694 3648 14728 3682
rect 14886 3648 14920 3682
rect 12054 3222 12088 3598
rect 12150 3222 12184 3598
rect 12246 3222 12280 3598
rect 12342 3222 12376 3598
rect 12438 3222 12472 3598
rect 12534 3222 12568 3598
rect 12630 3222 12664 3598
rect 12726 3222 12760 3598
rect 12822 3222 12856 3598
rect 12918 3222 12952 3598
rect 13014 3222 13048 3598
rect 13110 3222 13144 3598
rect 13206 3222 13240 3598
rect 13302 3222 13336 3598
rect 13398 3222 13432 3598
rect 13494 3222 13528 3598
rect 13590 3222 13624 3598
rect 13686 3222 13720 3598
rect 13782 3222 13816 3598
rect 13878 3222 13912 3598
rect 13974 3222 14008 3598
rect 14070 3222 14104 3598
rect 14166 3222 14200 3598
rect 14262 3222 14296 3598
rect 14358 3222 14392 3598
rect 14454 3222 14488 3598
rect 14550 3222 14584 3598
rect 14646 3222 14680 3598
rect 14742 3222 14776 3598
rect 14838 3222 14872 3598
rect 14934 3222 14968 3598
rect 12102 3138 12136 3172
rect 12294 3138 12328 3172
rect 12486 3138 12520 3172
rect 12678 3138 12712 3172
rect 12870 3138 12904 3172
rect 13062 3138 13096 3172
rect 13254 3138 13288 3172
rect 13446 3138 13480 3172
rect 13638 3138 13672 3172
rect 13830 3138 13864 3172
rect 14022 3138 14056 3172
rect 14214 3138 14248 3172
rect 14406 3138 14440 3172
rect 14598 3138 14632 3172
rect 14790 3138 14824 3172
rect 15742 5502 15776 5536
rect 15934 5502 15968 5536
rect 16126 5502 16160 5536
rect 16318 5502 16352 5536
rect 16510 5502 16544 5536
rect 16702 5502 16736 5536
rect 16894 5502 16928 5536
rect 17086 5502 17120 5536
rect 17278 5502 17312 5536
rect 17470 5502 17504 5536
rect 17662 5502 17696 5536
rect 17854 5502 17888 5536
rect 18046 5502 18080 5536
rect 18238 5502 18272 5536
rect 18430 5502 18464 5536
rect 15694 5076 15728 5452
rect 15790 5076 15824 5452
rect 15886 5076 15920 5452
rect 15982 5076 16016 5452
rect 16078 5076 16112 5452
rect 16174 5076 16208 5452
rect 16270 5076 16304 5452
rect 16366 5076 16400 5452
rect 16462 5076 16496 5452
rect 16558 5076 16592 5452
rect 16654 5076 16688 5452
rect 16750 5076 16784 5452
rect 16846 5076 16880 5452
rect 16942 5076 16976 5452
rect 17038 5076 17072 5452
rect 17134 5076 17168 5452
rect 17230 5076 17264 5452
rect 17326 5076 17360 5452
rect 17422 5076 17456 5452
rect 17518 5076 17552 5452
rect 17614 5076 17648 5452
rect 17710 5076 17744 5452
rect 17806 5076 17840 5452
rect 17902 5076 17936 5452
rect 17998 5076 18032 5452
rect 18094 5076 18128 5452
rect 18190 5076 18224 5452
rect 18286 5076 18320 5452
rect 18382 5076 18416 5452
rect 18478 5076 18512 5452
rect 18574 5076 18608 5452
rect 15838 4992 15872 5026
rect 16030 4992 16064 5026
rect 16222 4992 16256 5026
rect 16414 4992 16448 5026
rect 16606 4992 16640 5026
rect 16798 4992 16832 5026
rect 16990 4992 17024 5026
rect 17182 4992 17216 5026
rect 17374 4992 17408 5026
rect 17566 4992 17600 5026
rect 17758 4992 17792 5026
rect 17950 4992 17984 5026
rect 18142 4992 18176 5026
rect 18334 4992 18368 5026
rect 18526 4992 18560 5026
rect 15838 4884 15872 4918
rect 16030 4884 16064 4918
rect 16222 4884 16256 4918
rect 16414 4884 16448 4918
rect 16606 4884 16640 4918
rect 16798 4884 16832 4918
rect 16990 4884 17024 4918
rect 17182 4884 17216 4918
rect 17374 4884 17408 4918
rect 17566 4884 17600 4918
rect 17758 4884 17792 4918
rect 17950 4884 17984 4918
rect 18142 4884 18176 4918
rect 18334 4884 18368 4918
rect 18526 4884 18560 4918
rect 15694 4458 15728 4834
rect 15790 4458 15824 4834
rect 15886 4458 15920 4834
rect 15982 4458 16016 4834
rect 16078 4458 16112 4834
rect 16174 4458 16208 4834
rect 16270 4458 16304 4834
rect 16366 4458 16400 4834
rect 16462 4458 16496 4834
rect 16558 4458 16592 4834
rect 16654 4458 16688 4834
rect 16750 4458 16784 4834
rect 16846 4458 16880 4834
rect 16942 4458 16976 4834
rect 17038 4458 17072 4834
rect 17134 4458 17168 4834
rect 17230 4458 17264 4834
rect 17326 4458 17360 4834
rect 17422 4458 17456 4834
rect 17518 4458 17552 4834
rect 17614 4458 17648 4834
rect 17710 4458 17744 4834
rect 17806 4458 17840 4834
rect 17902 4458 17936 4834
rect 17998 4458 18032 4834
rect 18094 4458 18128 4834
rect 18190 4458 18224 4834
rect 18286 4458 18320 4834
rect 18382 4458 18416 4834
rect 18478 4458 18512 4834
rect 18574 4458 18608 4834
rect 15742 4374 15776 4408
rect 15934 4374 15968 4408
rect 16126 4374 16160 4408
rect 16318 4374 16352 4408
rect 16510 4374 16544 4408
rect 16702 4374 16736 4408
rect 16894 4374 16928 4408
rect 17086 4374 17120 4408
rect 17278 4374 17312 4408
rect 17470 4374 17504 4408
rect 17662 4374 17696 4408
rect 17854 4374 17888 4408
rect 18046 4374 18080 4408
rect 18238 4374 18272 4408
rect 18430 4374 18464 4408
rect 15742 4266 15776 4300
rect 15934 4266 15968 4300
rect 16126 4266 16160 4300
rect 16318 4266 16352 4300
rect 16510 4266 16544 4300
rect 16702 4266 16736 4300
rect 16894 4266 16928 4300
rect 17086 4266 17120 4300
rect 17278 4266 17312 4300
rect 17470 4266 17504 4300
rect 17662 4266 17696 4300
rect 17854 4266 17888 4300
rect 18046 4266 18080 4300
rect 18238 4266 18272 4300
rect 18430 4266 18464 4300
rect 15694 3840 15728 4216
rect 15790 3840 15824 4216
rect 15886 3840 15920 4216
rect 15982 3840 16016 4216
rect 16078 3840 16112 4216
rect 16174 3840 16208 4216
rect 16270 3840 16304 4216
rect 16366 3840 16400 4216
rect 16462 3840 16496 4216
rect 16558 3840 16592 4216
rect 16654 3840 16688 4216
rect 16750 3840 16784 4216
rect 16846 3840 16880 4216
rect 16942 3840 16976 4216
rect 17038 3840 17072 4216
rect 17134 3840 17168 4216
rect 17230 3840 17264 4216
rect 17326 3840 17360 4216
rect 17422 3840 17456 4216
rect 17518 3840 17552 4216
rect 17614 3840 17648 4216
rect 17710 3840 17744 4216
rect 17806 3840 17840 4216
rect 17902 3840 17936 4216
rect 17998 3840 18032 4216
rect 18094 3840 18128 4216
rect 18190 3840 18224 4216
rect 18286 3840 18320 4216
rect 18382 3840 18416 4216
rect 18478 3840 18512 4216
rect 18574 3840 18608 4216
rect 15838 3756 15872 3790
rect 16030 3756 16064 3790
rect 16222 3756 16256 3790
rect 16414 3756 16448 3790
rect 16606 3756 16640 3790
rect 16798 3756 16832 3790
rect 16990 3756 17024 3790
rect 17182 3756 17216 3790
rect 17374 3756 17408 3790
rect 17566 3756 17600 3790
rect 17758 3756 17792 3790
rect 17950 3756 17984 3790
rect 18142 3756 18176 3790
rect 18334 3756 18368 3790
rect 18526 3756 18560 3790
rect 15838 3648 15872 3682
rect 16030 3648 16064 3682
rect 16222 3648 16256 3682
rect 16414 3648 16448 3682
rect 16606 3648 16640 3682
rect 16798 3648 16832 3682
rect 16990 3648 17024 3682
rect 17182 3648 17216 3682
rect 17374 3648 17408 3682
rect 17566 3648 17600 3682
rect 17758 3648 17792 3682
rect 17950 3648 17984 3682
rect 18142 3648 18176 3682
rect 18334 3648 18368 3682
rect 18526 3648 18560 3682
rect 15694 3222 15728 3598
rect 15790 3222 15824 3598
rect 15886 3222 15920 3598
rect 15982 3222 16016 3598
rect 16078 3222 16112 3598
rect 16174 3222 16208 3598
rect 16270 3222 16304 3598
rect 16366 3222 16400 3598
rect 16462 3222 16496 3598
rect 16558 3222 16592 3598
rect 16654 3222 16688 3598
rect 16750 3222 16784 3598
rect 16846 3222 16880 3598
rect 16942 3222 16976 3598
rect 17038 3222 17072 3598
rect 17134 3222 17168 3598
rect 17230 3222 17264 3598
rect 17326 3222 17360 3598
rect 17422 3222 17456 3598
rect 17518 3222 17552 3598
rect 17614 3222 17648 3598
rect 17710 3222 17744 3598
rect 17806 3222 17840 3598
rect 17902 3222 17936 3598
rect 17998 3222 18032 3598
rect 18094 3222 18128 3598
rect 18190 3222 18224 3598
rect 18286 3222 18320 3598
rect 18382 3222 18416 3598
rect 18478 3222 18512 3598
rect 18574 3222 18608 3598
rect 15742 3138 15776 3172
rect 15934 3138 15968 3172
rect 16126 3138 16160 3172
rect 16318 3138 16352 3172
rect 16510 3138 16544 3172
rect 16702 3138 16736 3172
rect 16894 3138 16928 3172
rect 17086 3138 17120 3172
rect 17278 3138 17312 3172
rect 17470 3138 17504 3172
rect 17662 3138 17696 3172
rect 17854 3138 17888 3172
rect 18046 3138 18080 3172
rect 18238 3138 18272 3172
rect 18430 3138 18464 3172
rect -1522 2670 -1488 2704
rect -1330 2670 -1296 2704
rect -1138 2670 -1104 2704
rect -1570 2244 -1536 2620
rect -1474 2244 -1440 2620
rect -1378 2244 -1344 2620
rect -1282 2244 -1248 2620
rect -1186 2244 -1152 2620
rect -1090 2244 -1056 2620
rect -994 2244 -960 2620
rect -1426 2160 -1392 2194
rect -1234 2160 -1200 2194
rect -1042 2160 -1008 2194
rect -1426 2052 -1392 2086
rect -1234 2052 -1200 2086
rect -1042 2052 -1008 2086
rect -1570 1626 -1536 2002
rect -1474 1626 -1440 2002
rect -1378 1626 -1344 2002
rect -1282 1626 -1248 2002
rect -1186 1626 -1152 2002
rect -1090 1626 -1056 2002
rect -994 1626 -960 2002
rect -1522 1542 -1488 1576
rect -1330 1542 -1296 1576
rect -1138 1542 -1104 1576
rect -482 2670 -448 2704
rect -290 2670 -256 2704
rect -98 2670 -64 2704
rect -530 2244 -496 2620
rect -434 2244 -400 2620
rect -338 2244 -304 2620
rect -242 2244 -208 2620
rect -146 2244 -112 2620
rect -50 2244 -16 2620
rect 46 2244 80 2620
rect -386 2160 -352 2194
rect -194 2160 -160 2194
rect -2 2160 32 2194
rect -386 2052 -352 2086
rect -194 2052 -160 2086
rect -2 2052 32 2086
rect -530 1626 -496 2002
rect -434 1626 -400 2002
rect -338 1626 -304 2002
rect -242 1626 -208 2002
rect -146 1626 -112 2002
rect -50 1626 -16 2002
rect 46 1626 80 2002
rect -482 1542 -448 1576
rect -290 1542 -256 1576
rect -98 1542 -64 1576
rect 558 2670 592 2704
rect 750 2670 784 2704
rect 942 2670 976 2704
rect 510 2244 544 2620
rect 606 2244 640 2620
rect 702 2244 736 2620
rect 798 2244 832 2620
rect 894 2244 928 2620
rect 990 2244 1024 2620
rect 1086 2244 1120 2620
rect 654 2160 688 2194
rect 846 2160 880 2194
rect 1038 2160 1072 2194
rect 654 2052 688 2086
rect 846 2052 880 2086
rect 1038 2052 1072 2086
rect 510 1626 544 2002
rect 606 1626 640 2002
rect 702 1626 736 2002
rect 798 1626 832 2002
rect 894 1626 928 2002
rect 990 1626 1024 2002
rect 1086 1626 1120 2002
rect 558 1542 592 1576
rect 750 1542 784 1576
rect 942 1542 976 1576
rect 1598 2670 1632 2704
rect 1790 2670 1824 2704
rect 1982 2670 2016 2704
rect 1550 2244 1584 2620
rect 1646 2244 1680 2620
rect 1742 2244 1776 2620
rect 1838 2244 1872 2620
rect 1934 2244 1968 2620
rect 2030 2244 2064 2620
rect 2126 2244 2160 2620
rect 1694 2160 1728 2194
rect 1886 2160 1920 2194
rect 2078 2160 2112 2194
rect 1694 2052 1728 2086
rect 1886 2052 1920 2086
rect 2078 2052 2112 2086
rect 1550 1626 1584 2002
rect 1646 1626 1680 2002
rect 1742 1626 1776 2002
rect 1838 1626 1872 2002
rect 1934 1626 1968 2002
rect 2030 1626 2064 2002
rect 2126 1626 2160 2002
rect 1598 1542 1632 1576
rect 1790 1542 1824 1576
rect 1982 1542 2016 1576
rect 2638 2670 2672 2704
rect 2830 2670 2864 2704
rect 3022 2670 3056 2704
rect 2590 2244 2624 2620
rect 2686 2244 2720 2620
rect 2782 2244 2816 2620
rect 2878 2244 2912 2620
rect 2974 2244 3008 2620
rect 3070 2244 3104 2620
rect 3166 2244 3200 2620
rect 2734 2160 2768 2194
rect 2926 2160 2960 2194
rect 3118 2160 3152 2194
rect 2734 2052 2768 2086
rect 2926 2052 2960 2086
rect 3118 2052 3152 2086
rect 2590 1626 2624 2002
rect 2686 1626 2720 2002
rect 2782 1626 2816 2002
rect 2878 1626 2912 2002
rect 2974 1626 3008 2002
rect 3070 1626 3104 2002
rect 3166 1626 3200 2002
rect 2638 1542 2672 1576
rect 2830 1542 2864 1576
rect 3022 1542 3056 1576
rect 4282 2830 4316 2864
rect 4474 2830 4508 2864
rect 4666 2830 4700 2864
rect 4234 2404 4268 2780
rect 4330 2404 4364 2780
rect 4426 2404 4460 2780
rect 4522 2404 4556 2780
rect 4618 2404 4652 2780
rect 4714 2404 4748 2780
rect 4810 2404 4844 2780
rect 4378 2320 4412 2354
rect 4570 2320 4604 2354
rect 4762 2320 4796 2354
rect 4378 2212 4412 2246
rect 4570 2212 4604 2246
rect 4762 2212 4796 2246
rect 4234 1786 4268 2162
rect 4330 1786 4364 2162
rect 4426 1786 4460 2162
rect 4522 1786 4556 2162
rect 4618 1786 4652 2162
rect 4714 1786 4748 2162
rect 4810 1786 4844 2162
rect 4282 1702 4316 1736
rect 4474 1702 4508 1736
rect 4666 1702 4700 1736
rect 5322 2830 5356 2864
rect 5514 2830 5548 2864
rect 5706 2830 5740 2864
rect 5274 2404 5308 2780
rect 5370 2404 5404 2780
rect 5466 2404 5500 2780
rect 5562 2404 5596 2780
rect 5658 2404 5692 2780
rect 5754 2404 5788 2780
rect 5850 2404 5884 2780
rect 5418 2320 5452 2354
rect 5610 2320 5644 2354
rect 5802 2320 5836 2354
rect 5418 2212 5452 2246
rect 5610 2212 5644 2246
rect 5802 2212 5836 2246
rect 5274 1786 5308 2162
rect 5370 1786 5404 2162
rect 5466 1786 5500 2162
rect 5562 1786 5596 2162
rect 5658 1786 5692 2162
rect 5754 1786 5788 2162
rect 5850 1786 5884 2162
rect 5322 1702 5356 1736
rect 5514 1702 5548 1736
rect 5706 1702 5740 1736
rect 6362 2830 6396 2864
rect 6554 2830 6588 2864
rect 6746 2830 6780 2864
rect 6314 2404 6348 2780
rect 6410 2404 6444 2780
rect 6506 2404 6540 2780
rect 6602 2404 6636 2780
rect 6698 2404 6732 2780
rect 6794 2404 6828 2780
rect 6890 2404 6924 2780
rect 6458 2320 6492 2354
rect 6650 2320 6684 2354
rect 6842 2320 6876 2354
rect 6458 2212 6492 2246
rect 6650 2212 6684 2246
rect 6842 2212 6876 2246
rect 6314 1786 6348 2162
rect 6410 1786 6444 2162
rect 6506 1786 6540 2162
rect 6602 1786 6636 2162
rect 6698 1786 6732 2162
rect 6794 1786 6828 2162
rect 6890 1786 6924 2162
rect 6362 1702 6396 1736
rect 6554 1702 6588 1736
rect 6746 1702 6780 1736
rect 7402 2830 7436 2864
rect 7594 2830 7628 2864
rect 7786 2830 7820 2864
rect 7354 2404 7388 2780
rect 7450 2404 7484 2780
rect 7546 2404 7580 2780
rect 7642 2404 7676 2780
rect 7738 2404 7772 2780
rect 7834 2404 7868 2780
rect 7930 2404 7964 2780
rect 7498 2320 7532 2354
rect 7690 2320 7724 2354
rect 7882 2320 7916 2354
rect 7498 2212 7532 2246
rect 7690 2212 7724 2246
rect 7882 2212 7916 2246
rect 7354 1786 7388 2162
rect 7450 1786 7484 2162
rect 7546 1786 7580 2162
rect 7642 1786 7676 2162
rect 7738 1786 7772 2162
rect 7834 1786 7868 2162
rect 7930 1786 7964 2162
rect 7402 1702 7436 1736
rect 7594 1702 7628 1736
rect 7786 1702 7820 1736
rect 8442 2830 8476 2864
rect 8634 2830 8668 2864
rect 8826 2830 8860 2864
rect 8394 2404 8428 2780
rect 8490 2404 8524 2780
rect 8586 2404 8620 2780
rect 8682 2404 8716 2780
rect 8778 2404 8812 2780
rect 8874 2404 8908 2780
rect 8970 2404 9004 2780
rect 8538 2320 8572 2354
rect 8730 2320 8764 2354
rect 8922 2320 8956 2354
rect 8538 2212 8572 2246
rect 8730 2212 8764 2246
rect 8922 2212 8956 2246
rect 8394 1786 8428 2162
rect 8490 1786 8524 2162
rect 8586 1786 8620 2162
rect 8682 1786 8716 2162
rect 8778 1786 8812 2162
rect 8874 1786 8908 2162
rect 8970 1786 9004 2162
rect 8442 1702 8476 1736
rect 8634 1702 8668 1736
rect 8826 1702 8860 1736
rect 9482 2830 9516 2864
rect 9674 2830 9708 2864
rect 9866 2830 9900 2864
rect 9434 2404 9468 2780
rect 9530 2404 9564 2780
rect 9626 2404 9660 2780
rect 9722 2404 9756 2780
rect 9818 2404 9852 2780
rect 9914 2404 9948 2780
rect 10010 2404 10044 2780
rect 9578 2320 9612 2354
rect 9770 2320 9804 2354
rect 9962 2320 9996 2354
rect 9578 2212 9612 2246
rect 9770 2212 9804 2246
rect 9962 2212 9996 2246
rect 9434 1786 9468 2162
rect 9530 1786 9564 2162
rect 9626 1786 9660 2162
rect 9722 1786 9756 2162
rect 9818 1786 9852 2162
rect 9914 1786 9948 2162
rect 10010 1786 10044 2162
rect 9482 1702 9516 1736
rect 9674 1702 9708 1736
rect 9866 1702 9900 1736
rect 10522 2830 10556 2864
rect 10714 2830 10748 2864
rect 10906 2830 10940 2864
rect 10474 2404 10508 2780
rect 10570 2404 10604 2780
rect 10666 2404 10700 2780
rect 10762 2404 10796 2780
rect 10858 2404 10892 2780
rect 10954 2404 10988 2780
rect 11050 2404 11084 2780
rect 10618 2320 10652 2354
rect 10810 2320 10844 2354
rect 11002 2320 11036 2354
rect 10618 2212 10652 2246
rect 10810 2212 10844 2246
rect 11002 2212 11036 2246
rect 10474 1786 10508 2162
rect 10570 1786 10604 2162
rect 10666 1786 10700 2162
rect 10762 1786 10796 2162
rect 10858 1786 10892 2162
rect 10954 1786 10988 2162
rect 11050 1786 11084 2162
rect 10522 1702 10556 1736
rect 10714 1702 10748 1736
rect 10906 1702 10940 1736
rect 11902 2830 11936 2864
rect 12094 2830 12128 2864
rect 12286 2830 12320 2864
rect 11854 2404 11888 2780
rect 11950 2404 11984 2780
rect 12046 2404 12080 2780
rect 12142 2404 12176 2780
rect 12238 2404 12272 2780
rect 12334 2404 12368 2780
rect 12430 2404 12464 2780
rect 11998 2320 12032 2354
rect 12190 2320 12224 2354
rect 12382 2320 12416 2354
rect 11998 2212 12032 2246
rect 12190 2212 12224 2246
rect 12382 2212 12416 2246
rect 11854 1786 11888 2162
rect 11950 1786 11984 2162
rect 12046 1786 12080 2162
rect 12142 1786 12176 2162
rect 12238 1786 12272 2162
rect 12334 1786 12368 2162
rect 12430 1786 12464 2162
rect 11902 1702 11936 1736
rect 12094 1702 12128 1736
rect 12286 1702 12320 1736
rect 12942 2830 12976 2864
rect 13134 2830 13168 2864
rect 13326 2830 13360 2864
rect 12894 2404 12928 2780
rect 12990 2404 13024 2780
rect 13086 2404 13120 2780
rect 13182 2404 13216 2780
rect 13278 2404 13312 2780
rect 13374 2404 13408 2780
rect 13470 2404 13504 2780
rect 13038 2320 13072 2354
rect 13230 2320 13264 2354
rect 13422 2320 13456 2354
rect 13038 2212 13072 2246
rect 13230 2212 13264 2246
rect 13422 2212 13456 2246
rect 12894 1786 12928 2162
rect 12990 1786 13024 2162
rect 13086 1786 13120 2162
rect 13182 1786 13216 2162
rect 13278 1786 13312 2162
rect 13374 1786 13408 2162
rect 13470 1786 13504 2162
rect 12942 1702 12976 1736
rect 13134 1702 13168 1736
rect 13326 1702 13360 1736
rect 13982 2830 14016 2864
rect 14174 2830 14208 2864
rect 14366 2830 14400 2864
rect 13934 2404 13968 2780
rect 14030 2404 14064 2780
rect 14126 2404 14160 2780
rect 14222 2404 14256 2780
rect 14318 2404 14352 2780
rect 14414 2404 14448 2780
rect 14510 2404 14544 2780
rect 14078 2320 14112 2354
rect 14270 2320 14304 2354
rect 14462 2320 14496 2354
rect 14078 2212 14112 2246
rect 14270 2212 14304 2246
rect 14462 2212 14496 2246
rect 13934 1786 13968 2162
rect 14030 1786 14064 2162
rect 14126 1786 14160 2162
rect 14222 1786 14256 2162
rect 14318 1786 14352 2162
rect 14414 1786 14448 2162
rect 14510 1786 14544 2162
rect 13982 1702 14016 1736
rect 14174 1702 14208 1736
rect 14366 1702 14400 1736
rect 15022 2830 15056 2864
rect 15214 2830 15248 2864
rect 15406 2830 15440 2864
rect 14974 2404 15008 2780
rect 15070 2404 15104 2780
rect 15166 2404 15200 2780
rect 15262 2404 15296 2780
rect 15358 2404 15392 2780
rect 15454 2404 15488 2780
rect 15550 2404 15584 2780
rect 15118 2320 15152 2354
rect 15310 2320 15344 2354
rect 15502 2320 15536 2354
rect 15118 2212 15152 2246
rect 15310 2212 15344 2246
rect 15502 2212 15536 2246
rect 14974 1786 15008 2162
rect 15070 1786 15104 2162
rect 15166 1786 15200 2162
rect 15262 1786 15296 2162
rect 15358 1786 15392 2162
rect 15454 1786 15488 2162
rect 15550 1786 15584 2162
rect 15022 1702 15056 1736
rect 15214 1702 15248 1736
rect 15406 1702 15440 1736
rect 16062 2830 16096 2864
rect 16254 2830 16288 2864
rect 16446 2830 16480 2864
rect 16014 2404 16048 2780
rect 16110 2404 16144 2780
rect 16206 2404 16240 2780
rect 16302 2404 16336 2780
rect 16398 2404 16432 2780
rect 16494 2404 16528 2780
rect 16590 2404 16624 2780
rect 16158 2320 16192 2354
rect 16350 2320 16384 2354
rect 16542 2320 16576 2354
rect 16158 2212 16192 2246
rect 16350 2212 16384 2246
rect 16542 2212 16576 2246
rect 16014 1786 16048 2162
rect 16110 1786 16144 2162
rect 16206 1786 16240 2162
rect 16302 1786 16336 2162
rect 16398 1786 16432 2162
rect 16494 1786 16528 2162
rect 16590 1786 16624 2162
rect 16062 1702 16096 1736
rect 16254 1702 16288 1736
rect 16446 1702 16480 1736
rect 17102 2830 17136 2864
rect 17294 2830 17328 2864
rect 17486 2830 17520 2864
rect 17054 2404 17088 2780
rect 17150 2404 17184 2780
rect 17246 2404 17280 2780
rect 17342 2404 17376 2780
rect 17438 2404 17472 2780
rect 17534 2404 17568 2780
rect 17630 2404 17664 2780
rect 17198 2320 17232 2354
rect 17390 2320 17424 2354
rect 17582 2320 17616 2354
rect 17198 2212 17232 2246
rect 17390 2212 17424 2246
rect 17582 2212 17616 2246
rect 17054 1786 17088 2162
rect 17150 1786 17184 2162
rect 17246 1786 17280 2162
rect 17342 1786 17376 2162
rect 17438 1786 17472 2162
rect 17534 1786 17568 2162
rect 17630 1786 17664 2162
rect 17102 1702 17136 1736
rect 17294 1702 17328 1736
rect 17486 1702 17520 1736
rect 18142 2830 18176 2864
rect 18334 2830 18368 2864
rect 18526 2830 18560 2864
rect 18094 2404 18128 2780
rect 18190 2404 18224 2780
rect 18286 2404 18320 2780
rect 18382 2404 18416 2780
rect 18478 2404 18512 2780
rect 18574 2404 18608 2780
rect 18670 2404 18704 2780
rect 18238 2320 18272 2354
rect 18430 2320 18464 2354
rect 18622 2320 18656 2354
rect 18238 2212 18272 2246
rect 18430 2212 18464 2246
rect 18622 2212 18656 2246
rect 18094 1786 18128 2162
rect 18190 1786 18224 2162
rect 18286 1786 18320 2162
rect 18382 1786 18416 2162
rect 18478 1786 18512 2162
rect 18574 1786 18608 2162
rect 18670 1786 18704 2162
rect 18142 1702 18176 1736
rect 18334 1702 18368 1736
rect 18526 1702 18560 1736
rect -1511 1248 -1477 1282
rect -1393 1248 -1359 1282
rect -1275 1248 -1241 1282
rect -1157 1248 -1123 1282
rect -1039 1248 -1005 1282
rect -921 1248 -887 1282
rect -1570 822 -1536 1198
rect -1452 822 -1418 1198
rect -1334 822 -1300 1198
rect -1216 822 -1182 1198
rect -1098 822 -1064 1198
rect -980 822 -946 1198
rect -862 822 -828 1198
rect -1511 738 -1477 772
rect -1393 738 -1359 772
rect -1275 738 -1241 772
rect -1157 738 -1123 772
rect -1039 738 -1005 772
rect -921 738 -887 772
rect -471 1248 -437 1282
rect -353 1248 -319 1282
rect -235 1248 -201 1282
rect -117 1248 -83 1282
rect 1 1248 35 1282
rect 119 1248 153 1282
rect -530 822 -496 1198
rect -412 822 -378 1198
rect -294 822 -260 1198
rect -176 822 -142 1198
rect -58 822 -24 1198
rect 60 822 94 1198
rect 178 822 212 1198
rect -471 738 -437 772
rect -353 738 -319 772
rect -235 738 -201 772
rect -117 738 -83 772
rect 1 738 35 772
rect 119 738 153 772
rect 569 1248 603 1282
rect 687 1248 721 1282
rect 805 1248 839 1282
rect 923 1248 957 1282
rect 1041 1248 1075 1282
rect 1159 1248 1193 1282
rect 510 822 544 1198
rect 628 822 662 1198
rect 746 822 780 1198
rect 864 822 898 1198
rect 982 822 1016 1198
rect 1100 822 1134 1198
rect 1218 822 1252 1198
rect 569 738 603 772
rect 687 738 721 772
rect 805 738 839 772
rect 923 738 957 772
rect 1041 738 1075 772
rect 1159 738 1193 772
rect 1609 1248 1643 1282
rect 1727 1248 1761 1282
rect 1845 1248 1879 1282
rect 1963 1248 1997 1282
rect 2081 1248 2115 1282
rect 2199 1248 2233 1282
rect 1550 822 1584 1198
rect 1668 822 1702 1198
rect 1786 822 1820 1198
rect 1904 822 1938 1198
rect 2022 822 2056 1198
rect 2140 822 2174 1198
rect 2258 822 2292 1198
rect 1609 738 1643 772
rect 1727 738 1761 772
rect 1845 738 1879 772
rect 1963 738 1997 772
rect 2081 738 2115 772
rect 2199 738 2233 772
rect 2649 1248 2683 1282
rect 2767 1248 2801 1282
rect 2885 1248 2919 1282
rect 3003 1248 3037 1282
rect 3121 1248 3155 1282
rect 3239 1248 3273 1282
rect 2590 822 2624 1198
rect 2708 822 2742 1198
rect 2826 822 2860 1198
rect 2944 822 2978 1198
rect 3062 822 3096 1198
rect 3180 822 3214 1198
rect 3298 822 3332 1198
rect 2649 738 2683 772
rect 2767 738 2801 772
rect 2885 738 2919 772
rect 3003 738 3037 772
rect 3121 738 3155 772
rect 3239 738 3273 772
rect 4293 1408 4327 1442
rect 4411 1408 4445 1442
rect 4529 1408 4563 1442
rect 4647 1408 4681 1442
rect 4765 1408 4799 1442
rect 4883 1408 4917 1442
rect 4234 982 4268 1358
rect 4352 982 4386 1358
rect 4470 982 4504 1358
rect 4588 982 4622 1358
rect 4706 982 4740 1358
rect 4824 982 4858 1358
rect 4942 982 4976 1358
rect 4293 898 4327 932
rect 4411 898 4445 932
rect 4529 898 4563 932
rect 4647 898 4681 932
rect 4765 898 4799 932
rect 4883 898 4917 932
rect 5333 1408 5367 1442
rect 5451 1408 5485 1442
rect 5569 1408 5603 1442
rect 5687 1408 5721 1442
rect 5805 1408 5839 1442
rect 5923 1408 5957 1442
rect 5274 982 5308 1358
rect 5392 982 5426 1358
rect 5510 982 5544 1358
rect 5628 982 5662 1358
rect 5746 982 5780 1358
rect 5864 982 5898 1358
rect 5982 982 6016 1358
rect 5333 898 5367 932
rect 5451 898 5485 932
rect 5569 898 5603 932
rect 5687 898 5721 932
rect 5805 898 5839 932
rect 5923 898 5957 932
rect 6373 1408 6407 1442
rect 6491 1408 6525 1442
rect 6609 1408 6643 1442
rect 6727 1408 6761 1442
rect 6845 1408 6879 1442
rect 6963 1408 6997 1442
rect 6314 982 6348 1358
rect 6432 982 6466 1358
rect 6550 982 6584 1358
rect 6668 982 6702 1358
rect 6786 982 6820 1358
rect 6904 982 6938 1358
rect 7022 982 7056 1358
rect 6373 898 6407 932
rect 6491 898 6525 932
rect 6609 898 6643 932
rect 6727 898 6761 932
rect 6845 898 6879 932
rect 6963 898 6997 932
rect 7413 1408 7447 1442
rect 7531 1408 7565 1442
rect 7649 1408 7683 1442
rect 7767 1408 7801 1442
rect 7885 1408 7919 1442
rect 8003 1408 8037 1442
rect 7354 982 7388 1358
rect 7472 982 7506 1358
rect 7590 982 7624 1358
rect 7708 982 7742 1358
rect 7826 982 7860 1358
rect 7944 982 7978 1358
rect 8062 982 8096 1358
rect 7413 898 7447 932
rect 7531 898 7565 932
rect 7649 898 7683 932
rect 7767 898 7801 932
rect 7885 898 7919 932
rect 8003 898 8037 932
rect 8453 1408 8487 1442
rect 8571 1408 8605 1442
rect 8689 1408 8723 1442
rect 8807 1408 8841 1442
rect 8925 1408 8959 1442
rect 9043 1408 9077 1442
rect 8394 982 8428 1358
rect 8512 982 8546 1358
rect 8630 982 8664 1358
rect 8748 982 8782 1358
rect 8866 982 8900 1358
rect 8984 982 9018 1358
rect 9102 982 9136 1358
rect 8453 898 8487 932
rect 8571 898 8605 932
rect 8689 898 8723 932
rect 8807 898 8841 932
rect 8925 898 8959 932
rect 9043 898 9077 932
rect 9493 1408 9527 1442
rect 9611 1408 9645 1442
rect 9729 1408 9763 1442
rect 9847 1408 9881 1442
rect 9965 1408 9999 1442
rect 10083 1408 10117 1442
rect 9434 982 9468 1358
rect 9552 982 9586 1358
rect 9670 982 9704 1358
rect 9788 982 9822 1358
rect 9906 982 9940 1358
rect 10024 982 10058 1358
rect 10142 982 10176 1358
rect 9493 898 9527 932
rect 9611 898 9645 932
rect 9729 898 9763 932
rect 9847 898 9881 932
rect 9965 898 9999 932
rect 10083 898 10117 932
rect 10533 1408 10567 1442
rect 10651 1408 10685 1442
rect 10769 1408 10803 1442
rect 10887 1408 10921 1442
rect 11005 1408 11039 1442
rect 11123 1408 11157 1442
rect 10474 982 10508 1358
rect 10592 982 10626 1358
rect 10710 982 10744 1358
rect 10828 982 10862 1358
rect 10946 982 10980 1358
rect 11064 982 11098 1358
rect 11182 982 11216 1358
rect 10533 898 10567 932
rect 10651 898 10685 932
rect 10769 898 10803 932
rect 10887 898 10921 932
rect 11005 898 11039 932
rect 11123 898 11157 932
rect 11913 1408 11947 1442
rect 12031 1408 12065 1442
rect 12149 1408 12183 1442
rect 12267 1408 12301 1442
rect 12385 1408 12419 1442
rect 12503 1408 12537 1442
rect 11854 982 11888 1358
rect 11972 982 12006 1358
rect 12090 982 12124 1358
rect 12208 982 12242 1358
rect 12326 982 12360 1358
rect 12444 982 12478 1358
rect 12562 982 12596 1358
rect 11913 898 11947 932
rect 12031 898 12065 932
rect 12149 898 12183 932
rect 12267 898 12301 932
rect 12385 898 12419 932
rect 12503 898 12537 932
rect 12953 1408 12987 1442
rect 13071 1408 13105 1442
rect 13189 1408 13223 1442
rect 13307 1408 13341 1442
rect 13425 1408 13459 1442
rect 13543 1408 13577 1442
rect 12894 982 12928 1358
rect 13012 982 13046 1358
rect 13130 982 13164 1358
rect 13248 982 13282 1358
rect 13366 982 13400 1358
rect 13484 982 13518 1358
rect 13602 982 13636 1358
rect 12953 898 12987 932
rect 13071 898 13105 932
rect 13189 898 13223 932
rect 13307 898 13341 932
rect 13425 898 13459 932
rect 13543 898 13577 932
rect 13993 1408 14027 1442
rect 14111 1408 14145 1442
rect 14229 1408 14263 1442
rect 14347 1408 14381 1442
rect 14465 1408 14499 1442
rect 14583 1408 14617 1442
rect 13934 982 13968 1358
rect 14052 982 14086 1358
rect 14170 982 14204 1358
rect 14288 982 14322 1358
rect 14406 982 14440 1358
rect 14524 982 14558 1358
rect 14642 982 14676 1358
rect 13993 898 14027 932
rect 14111 898 14145 932
rect 14229 898 14263 932
rect 14347 898 14381 932
rect 14465 898 14499 932
rect 14583 898 14617 932
rect 15033 1408 15067 1442
rect 15151 1408 15185 1442
rect 15269 1408 15303 1442
rect 15387 1408 15421 1442
rect 15505 1408 15539 1442
rect 15623 1408 15657 1442
rect 14974 982 15008 1358
rect 15092 982 15126 1358
rect 15210 982 15244 1358
rect 15328 982 15362 1358
rect 15446 982 15480 1358
rect 15564 982 15598 1358
rect 15682 982 15716 1358
rect 15033 898 15067 932
rect 15151 898 15185 932
rect 15269 898 15303 932
rect 15387 898 15421 932
rect 15505 898 15539 932
rect 15623 898 15657 932
rect 16073 1408 16107 1442
rect 16191 1408 16225 1442
rect 16309 1408 16343 1442
rect 16427 1408 16461 1442
rect 16545 1408 16579 1442
rect 16663 1408 16697 1442
rect 16014 982 16048 1358
rect 16132 982 16166 1358
rect 16250 982 16284 1358
rect 16368 982 16402 1358
rect 16486 982 16520 1358
rect 16604 982 16638 1358
rect 16722 982 16756 1358
rect 16073 898 16107 932
rect 16191 898 16225 932
rect 16309 898 16343 932
rect 16427 898 16461 932
rect 16545 898 16579 932
rect 16663 898 16697 932
rect 17113 1408 17147 1442
rect 17231 1408 17265 1442
rect 17349 1408 17383 1442
rect 17467 1408 17501 1442
rect 17585 1408 17619 1442
rect 17703 1408 17737 1442
rect 17054 982 17088 1358
rect 17172 982 17206 1358
rect 17290 982 17324 1358
rect 17408 982 17442 1358
rect 17526 982 17560 1358
rect 17644 982 17678 1358
rect 17762 982 17796 1358
rect 17113 898 17147 932
rect 17231 898 17265 932
rect 17349 898 17383 932
rect 17467 898 17501 932
rect 17585 898 17619 932
rect 17703 898 17737 932
rect 18153 1408 18187 1442
rect 18271 1408 18305 1442
rect 18389 1408 18423 1442
rect 18507 1408 18541 1442
rect 18625 1408 18659 1442
rect 18743 1408 18777 1442
rect 18094 982 18128 1358
rect 18212 982 18246 1358
rect 18330 982 18364 1358
rect 18448 982 18482 1358
rect 18566 982 18600 1358
rect 18684 982 18718 1358
rect 18802 982 18836 1358
rect 18153 898 18187 932
rect 18271 898 18305 932
rect 18389 898 18423 932
rect 18507 898 18541 932
rect 18625 898 18659 932
rect 18743 898 18777 932
rect -1308 412 -1128 476
rect 2800 408 3068 492
rect -7352 -16 -7318 18
rect -7160 -16 -7126 18
rect -6968 -16 -6934 18
rect -6776 -16 -6742 18
rect -6584 -16 -6550 18
rect -7400 -442 -7366 -66
rect -7304 -442 -7270 -66
rect -7208 -442 -7174 -66
rect -7112 -442 -7078 -66
rect -7016 -442 -6982 -66
rect -6920 -442 -6886 -66
rect -6824 -442 -6790 -66
rect -6728 -442 -6694 -66
rect -6632 -442 -6598 -66
rect -6536 -442 -6502 -66
rect -6440 -442 -6406 -66
rect -7256 -526 -7222 -492
rect -7064 -526 -7030 -492
rect -6872 -526 -6838 -492
rect -6680 -526 -6646 -492
rect -6488 -526 -6454 -492
rect -7256 -634 -7222 -600
rect -7064 -634 -7030 -600
rect -6872 -634 -6838 -600
rect -6680 -634 -6646 -600
rect -6488 -634 -6454 -600
rect -7400 -1060 -7366 -684
rect -7304 -1060 -7270 -684
rect -7208 -1060 -7174 -684
rect -7112 -1060 -7078 -684
rect -7016 -1060 -6982 -684
rect -6920 -1060 -6886 -684
rect -6824 -1060 -6790 -684
rect -6728 -1060 -6694 -684
rect -6632 -1060 -6598 -684
rect -6536 -1060 -6502 -684
rect -6440 -1060 -6406 -684
rect -7352 -1144 -7318 -1110
rect -7160 -1144 -7126 -1110
rect -6968 -1144 -6934 -1110
rect -6776 -1144 -6742 -1110
rect -6584 -1144 -6550 -1110
rect -7352 -1852 -7318 -1818
rect -7160 -1852 -7126 -1818
rect -6968 -1852 -6934 -1818
rect -7400 -2278 -7366 -1902
rect -7304 -2278 -7270 -1902
rect -7208 -2278 -7174 -1902
rect -7112 -2278 -7078 -1902
rect -7016 -2278 -6982 -1902
rect -6920 -2278 -6886 -1902
rect -6824 -2278 -6790 -1902
rect -7256 -2362 -7222 -2328
rect -7064 -2362 -7030 -2328
rect -6872 -2362 -6838 -2328
rect -7256 -2470 -7222 -2436
rect -7064 -2470 -7030 -2436
rect -6872 -2470 -6838 -2436
rect -7400 -2896 -7366 -2520
rect -7304 -2896 -7270 -2520
rect -7208 -2896 -7174 -2520
rect -7112 -2896 -7078 -2520
rect -7016 -2896 -6982 -2520
rect -6920 -2896 -6886 -2520
rect -6824 -2896 -6790 -2520
rect -7352 -2980 -7318 -2946
rect -7160 -2980 -7126 -2946
rect -6968 -2980 -6934 -2946
rect -5988 -42 -5812 -8
rect -6072 -1638 -6038 -70
rect -5762 -1638 -5728 -70
rect -5988 -1700 -5812 -1666
rect 4282 590 4316 624
rect 4474 590 4508 624
rect 4666 590 4700 624
rect 4234 164 4268 540
rect 4330 164 4364 540
rect 4426 164 4460 540
rect 4522 164 4556 540
rect 4618 164 4652 540
rect 4714 164 4748 540
rect 4810 164 4844 540
rect 4378 80 4412 114
rect 4570 80 4604 114
rect 4762 80 4796 114
rect 4378 -28 4412 6
rect 4570 -28 4604 6
rect 4762 -28 4796 6
rect 4234 -454 4268 -78
rect 4330 -454 4364 -78
rect 4426 -454 4460 -78
rect 4522 -454 4556 -78
rect 4618 -454 4652 -78
rect 4714 -454 4748 -78
rect 4810 -454 4844 -78
rect 4282 -538 4316 -504
rect 4474 -538 4508 -504
rect 4666 -538 4700 -504
rect 5322 590 5356 624
rect 5514 590 5548 624
rect 5706 590 5740 624
rect 5274 164 5308 540
rect 5370 164 5404 540
rect 5466 164 5500 540
rect 5562 164 5596 540
rect 5658 164 5692 540
rect 5754 164 5788 540
rect 5850 164 5884 540
rect 5418 80 5452 114
rect 5610 80 5644 114
rect 5802 80 5836 114
rect 5418 -28 5452 6
rect 5610 -28 5644 6
rect 5802 -28 5836 6
rect 5274 -454 5308 -78
rect 5370 -454 5404 -78
rect 5466 -454 5500 -78
rect 5562 -454 5596 -78
rect 5658 -454 5692 -78
rect 5754 -454 5788 -78
rect 5850 -454 5884 -78
rect 5322 -538 5356 -504
rect 5514 -538 5548 -504
rect 5706 -538 5740 -504
rect 6362 590 6396 624
rect 6554 590 6588 624
rect 6746 590 6780 624
rect 6314 164 6348 540
rect 6410 164 6444 540
rect 6506 164 6540 540
rect 6602 164 6636 540
rect 6698 164 6732 540
rect 6794 164 6828 540
rect 6890 164 6924 540
rect 6458 80 6492 114
rect 6650 80 6684 114
rect 6842 80 6876 114
rect 6458 -28 6492 6
rect 6650 -28 6684 6
rect 6842 -28 6876 6
rect 6314 -454 6348 -78
rect 6410 -454 6444 -78
rect 6506 -454 6540 -78
rect 6602 -454 6636 -78
rect 6698 -454 6732 -78
rect 6794 -454 6828 -78
rect 6890 -454 6924 -78
rect 6362 -538 6396 -504
rect 6554 -538 6588 -504
rect 6746 -538 6780 -504
rect 7402 590 7436 624
rect 7594 590 7628 624
rect 7786 590 7820 624
rect 7354 164 7388 540
rect 7450 164 7484 540
rect 7546 164 7580 540
rect 7642 164 7676 540
rect 7738 164 7772 540
rect 7834 164 7868 540
rect 7930 164 7964 540
rect 7498 80 7532 114
rect 7690 80 7724 114
rect 7882 80 7916 114
rect 7498 -28 7532 6
rect 7690 -28 7724 6
rect 7882 -28 7916 6
rect 7354 -454 7388 -78
rect 7450 -454 7484 -78
rect 7546 -454 7580 -78
rect 7642 -454 7676 -78
rect 7738 -454 7772 -78
rect 7834 -454 7868 -78
rect 7930 -454 7964 -78
rect 7402 -538 7436 -504
rect 7594 -538 7628 -504
rect 7786 -538 7820 -504
rect 8442 590 8476 624
rect 8634 590 8668 624
rect 8826 590 8860 624
rect 8394 164 8428 540
rect 8490 164 8524 540
rect 8586 164 8620 540
rect 8682 164 8716 540
rect 8778 164 8812 540
rect 8874 164 8908 540
rect 8970 164 9004 540
rect 8538 80 8572 114
rect 8730 80 8764 114
rect 8922 80 8956 114
rect 8538 -28 8572 6
rect 8730 -28 8764 6
rect 8922 -28 8956 6
rect 8394 -454 8428 -78
rect 8490 -454 8524 -78
rect 8586 -454 8620 -78
rect 8682 -454 8716 -78
rect 8778 -454 8812 -78
rect 8874 -454 8908 -78
rect 8970 -454 9004 -78
rect 8442 -538 8476 -504
rect 8634 -538 8668 -504
rect 8826 -538 8860 -504
rect 9482 590 9516 624
rect 9674 590 9708 624
rect 9866 590 9900 624
rect 9434 164 9468 540
rect 9530 164 9564 540
rect 9626 164 9660 540
rect 9722 164 9756 540
rect 9818 164 9852 540
rect 9914 164 9948 540
rect 10010 164 10044 540
rect 9578 80 9612 114
rect 9770 80 9804 114
rect 9962 80 9996 114
rect 9578 -28 9612 6
rect 9770 -28 9804 6
rect 9962 -28 9996 6
rect 9434 -454 9468 -78
rect 9530 -454 9564 -78
rect 9626 -454 9660 -78
rect 9722 -454 9756 -78
rect 9818 -454 9852 -78
rect 9914 -454 9948 -78
rect 10010 -454 10044 -78
rect 9482 -538 9516 -504
rect 9674 -538 9708 -504
rect 9866 -538 9900 -504
rect 10522 590 10556 624
rect 10714 590 10748 624
rect 10906 590 10940 624
rect 10474 164 10508 540
rect 10570 164 10604 540
rect 10666 164 10700 540
rect 10762 164 10796 540
rect 10858 164 10892 540
rect 10954 164 10988 540
rect 11050 164 11084 540
rect 10618 80 10652 114
rect 10810 80 10844 114
rect 11002 80 11036 114
rect 10618 -28 10652 6
rect 10810 -28 10844 6
rect 11002 -28 11036 6
rect 10474 -454 10508 -78
rect 10570 -454 10604 -78
rect 10666 -454 10700 -78
rect 10762 -454 10796 -78
rect 10858 -454 10892 -78
rect 10954 -454 10988 -78
rect 11050 -454 11084 -78
rect 10522 -538 10556 -504
rect 10714 -538 10748 -504
rect 10906 -538 10940 -504
rect 11902 590 11936 624
rect 12094 590 12128 624
rect 12286 590 12320 624
rect 11854 164 11888 540
rect 11950 164 11984 540
rect 12046 164 12080 540
rect 12142 164 12176 540
rect 12238 164 12272 540
rect 12334 164 12368 540
rect 12430 164 12464 540
rect 11998 80 12032 114
rect 12190 80 12224 114
rect 12382 80 12416 114
rect 11998 -28 12032 6
rect 12190 -28 12224 6
rect 12382 -28 12416 6
rect 11854 -454 11888 -78
rect 11950 -454 11984 -78
rect 12046 -454 12080 -78
rect 12142 -454 12176 -78
rect 12238 -454 12272 -78
rect 12334 -454 12368 -78
rect 12430 -454 12464 -78
rect 11902 -538 11936 -504
rect 12094 -538 12128 -504
rect 12286 -538 12320 -504
rect 12942 590 12976 624
rect 13134 590 13168 624
rect 13326 590 13360 624
rect 12894 164 12928 540
rect 12990 164 13024 540
rect 13086 164 13120 540
rect 13182 164 13216 540
rect 13278 164 13312 540
rect 13374 164 13408 540
rect 13470 164 13504 540
rect 13038 80 13072 114
rect 13230 80 13264 114
rect 13422 80 13456 114
rect 13038 -28 13072 6
rect 13230 -28 13264 6
rect 13422 -28 13456 6
rect 12894 -454 12928 -78
rect 12990 -454 13024 -78
rect 13086 -454 13120 -78
rect 13182 -454 13216 -78
rect 13278 -454 13312 -78
rect 13374 -454 13408 -78
rect 13470 -454 13504 -78
rect 12942 -538 12976 -504
rect 13134 -538 13168 -504
rect 13326 -538 13360 -504
rect 13982 590 14016 624
rect 14174 590 14208 624
rect 14366 590 14400 624
rect 13934 164 13968 540
rect 14030 164 14064 540
rect 14126 164 14160 540
rect 14222 164 14256 540
rect 14318 164 14352 540
rect 14414 164 14448 540
rect 14510 164 14544 540
rect 14078 80 14112 114
rect 14270 80 14304 114
rect 14462 80 14496 114
rect 14078 -28 14112 6
rect 14270 -28 14304 6
rect 14462 -28 14496 6
rect 13934 -454 13968 -78
rect 14030 -454 14064 -78
rect 14126 -454 14160 -78
rect 14222 -454 14256 -78
rect 14318 -454 14352 -78
rect 14414 -454 14448 -78
rect 14510 -454 14544 -78
rect 13982 -538 14016 -504
rect 14174 -538 14208 -504
rect 14366 -538 14400 -504
rect 15022 590 15056 624
rect 15214 590 15248 624
rect 15406 590 15440 624
rect 14974 164 15008 540
rect 15070 164 15104 540
rect 15166 164 15200 540
rect 15262 164 15296 540
rect 15358 164 15392 540
rect 15454 164 15488 540
rect 15550 164 15584 540
rect 15118 80 15152 114
rect 15310 80 15344 114
rect 15502 80 15536 114
rect 15118 -28 15152 6
rect 15310 -28 15344 6
rect 15502 -28 15536 6
rect 14974 -454 15008 -78
rect 15070 -454 15104 -78
rect 15166 -454 15200 -78
rect 15262 -454 15296 -78
rect 15358 -454 15392 -78
rect 15454 -454 15488 -78
rect 15550 -454 15584 -78
rect 15022 -538 15056 -504
rect 15214 -538 15248 -504
rect 15406 -538 15440 -504
rect 16062 590 16096 624
rect 16254 590 16288 624
rect 16446 590 16480 624
rect 16014 164 16048 540
rect 16110 164 16144 540
rect 16206 164 16240 540
rect 16302 164 16336 540
rect 16398 164 16432 540
rect 16494 164 16528 540
rect 16590 164 16624 540
rect 16158 80 16192 114
rect 16350 80 16384 114
rect 16542 80 16576 114
rect 16158 -28 16192 6
rect 16350 -28 16384 6
rect 16542 -28 16576 6
rect 16014 -454 16048 -78
rect 16110 -454 16144 -78
rect 16206 -454 16240 -78
rect 16302 -454 16336 -78
rect 16398 -454 16432 -78
rect 16494 -454 16528 -78
rect 16590 -454 16624 -78
rect 16062 -538 16096 -504
rect 16254 -538 16288 -504
rect 16446 -538 16480 -504
rect 17102 590 17136 624
rect 17294 590 17328 624
rect 17486 590 17520 624
rect 17054 164 17088 540
rect 17150 164 17184 540
rect 17246 164 17280 540
rect 17342 164 17376 540
rect 17438 164 17472 540
rect 17534 164 17568 540
rect 17630 164 17664 540
rect 17198 80 17232 114
rect 17390 80 17424 114
rect 17582 80 17616 114
rect 17198 -28 17232 6
rect 17390 -28 17424 6
rect 17582 -28 17616 6
rect 17054 -454 17088 -78
rect 17150 -454 17184 -78
rect 17246 -454 17280 -78
rect 17342 -454 17376 -78
rect 17438 -454 17472 -78
rect 17534 -454 17568 -78
rect 17630 -454 17664 -78
rect 17102 -538 17136 -504
rect 17294 -538 17328 -504
rect 17486 -538 17520 -504
rect 18142 590 18176 624
rect 18334 590 18368 624
rect 18526 590 18560 624
rect 18094 164 18128 540
rect 18190 164 18224 540
rect 18286 164 18320 540
rect 18382 164 18416 540
rect 18478 164 18512 540
rect 18574 164 18608 540
rect 18670 164 18704 540
rect 18238 80 18272 114
rect 18430 80 18464 114
rect 18622 80 18656 114
rect 18238 -28 18272 6
rect 18430 -28 18464 6
rect 18622 -28 18656 6
rect 18094 -454 18128 -78
rect 18190 -454 18224 -78
rect 18286 -454 18320 -78
rect 18382 -454 18416 -78
rect 18478 -454 18512 -78
rect 18574 -454 18608 -78
rect 18670 -454 18704 -78
rect 18142 -538 18176 -504
rect 18334 -538 18368 -504
rect 18526 -538 18560 -504
rect 4293 -832 4327 -798
rect 4411 -832 4445 -798
rect 4529 -832 4563 -798
rect 4647 -832 4681 -798
rect 4765 -832 4799 -798
rect 4883 -832 4917 -798
rect 4234 -1258 4268 -882
rect 4352 -1258 4386 -882
rect 4470 -1258 4504 -882
rect 4588 -1258 4622 -882
rect 4706 -1258 4740 -882
rect 4824 -1258 4858 -882
rect 4942 -1258 4976 -882
rect 4293 -1342 4327 -1308
rect 4411 -1342 4445 -1308
rect 4529 -1342 4563 -1308
rect 4647 -1342 4681 -1308
rect 4765 -1342 4799 -1308
rect 4883 -1342 4917 -1308
rect 5333 -832 5367 -798
rect 5451 -832 5485 -798
rect 5569 -832 5603 -798
rect 5687 -832 5721 -798
rect 5805 -832 5839 -798
rect 5923 -832 5957 -798
rect 5274 -1258 5308 -882
rect 5392 -1258 5426 -882
rect 5510 -1258 5544 -882
rect 5628 -1258 5662 -882
rect 5746 -1258 5780 -882
rect 5864 -1258 5898 -882
rect 5982 -1258 6016 -882
rect 5333 -1342 5367 -1308
rect 5451 -1342 5485 -1308
rect 5569 -1342 5603 -1308
rect 5687 -1342 5721 -1308
rect 5805 -1342 5839 -1308
rect 5923 -1342 5957 -1308
rect 6373 -832 6407 -798
rect 6491 -832 6525 -798
rect 6609 -832 6643 -798
rect 6727 -832 6761 -798
rect 6845 -832 6879 -798
rect 6963 -832 6997 -798
rect 6314 -1258 6348 -882
rect 6432 -1258 6466 -882
rect 6550 -1258 6584 -882
rect 6668 -1258 6702 -882
rect 6786 -1258 6820 -882
rect 6904 -1258 6938 -882
rect 7022 -1258 7056 -882
rect 6373 -1342 6407 -1308
rect 6491 -1342 6525 -1308
rect 6609 -1342 6643 -1308
rect 6727 -1342 6761 -1308
rect 6845 -1342 6879 -1308
rect 6963 -1342 6997 -1308
rect 7413 -832 7447 -798
rect 7531 -832 7565 -798
rect 7649 -832 7683 -798
rect 7767 -832 7801 -798
rect 7885 -832 7919 -798
rect 8003 -832 8037 -798
rect 7354 -1258 7388 -882
rect 7472 -1258 7506 -882
rect 7590 -1258 7624 -882
rect 7708 -1258 7742 -882
rect 7826 -1258 7860 -882
rect 7944 -1258 7978 -882
rect 8062 -1258 8096 -882
rect 7413 -1342 7447 -1308
rect 7531 -1342 7565 -1308
rect 7649 -1342 7683 -1308
rect 7767 -1342 7801 -1308
rect 7885 -1342 7919 -1308
rect 8003 -1342 8037 -1308
rect 8453 -832 8487 -798
rect 8571 -832 8605 -798
rect 8689 -832 8723 -798
rect 8807 -832 8841 -798
rect 8925 -832 8959 -798
rect 9043 -832 9077 -798
rect 8394 -1258 8428 -882
rect 8512 -1258 8546 -882
rect 8630 -1258 8664 -882
rect 8748 -1258 8782 -882
rect 8866 -1258 8900 -882
rect 8984 -1258 9018 -882
rect 9102 -1258 9136 -882
rect 8453 -1342 8487 -1308
rect 8571 -1342 8605 -1308
rect 8689 -1342 8723 -1308
rect 8807 -1342 8841 -1308
rect 8925 -1342 8959 -1308
rect 9043 -1342 9077 -1308
rect 9493 -832 9527 -798
rect 9611 -832 9645 -798
rect 9729 -832 9763 -798
rect 9847 -832 9881 -798
rect 9965 -832 9999 -798
rect 10083 -832 10117 -798
rect 9434 -1258 9468 -882
rect 9552 -1258 9586 -882
rect 9670 -1258 9704 -882
rect 9788 -1258 9822 -882
rect 9906 -1258 9940 -882
rect 10024 -1258 10058 -882
rect 10142 -1258 10176 -882
rect 9493 -1342 9527 -1308
rect 9611 -1342 9645 -1308
rect 9729 -1342 9763 -1308
rect 9847 -1342 9881 -1308
rect 9965 -1342 9999 -1308
rect 10083 -1342 10117 -1308
rect 10533 -832 10567 -798
rect 10651 -832 10685 -798
rect 10769 -832 10803 -798
rect 10887 -832 10921 -798
rect 11005 -832 11039 -798
rect 11123 -832 11157 -798
rect 10474 -1258 10508 -882
rect 10592 -1258 10626 -882
rect 10710 -1258 10744 -882
rect 10828 -1258 10862 -882
rect 10946 -1258 10980 -882
rect 11064 -1258 11098 -882
rect 11182 -1258 11216 -882
rect 10533 -1342 10567 -1308
rect 10651 -1342 10685 -1308
rect 10769 -1342 10803 -1308
rect 10887 -1342 10921 -1308
rect 11005 -1342 11039 -1308
rect 11123 -1342 11157 -1308
rect 11913 -832 11947 -798
rect 12031 -832 12065 -798
rect 12149 -832 12183 -798
rect 12267 -832 12301 -798
rect 12385 -832 12419 -798
rect 12503 -832 12537 -798
rect 11854 -1258 11888 -882
rect 11972 -1258 12006 -882
rect 12090 -1258 12124 -882
rect 12208 -1258 12242 -882
rect 12326 -1258 12360 -882
rect 12444 -1258 12478 -882
rect 12562 -1258 12596 -882
rect 11913 -1342 11947 -1308
rect 12031 -1342 12065 -1308
rect 12149 -1342 12183 -1308
rect 12267 -1342 12301 -1308
rect 12385 -1342 12419 -1308
rect 12503 -1342 12537 -1308
rect 12953 -832 12987 -798
rect 13071 -832 13105 -798
rect 13189 -832 13223 -798
rect 13307 -832 13341 -798
rect 13425 -832 13459 -798
rect 13543 -832 13577 -798
rect 12894 -1258 12928 -882
rect 13012 -1258 13046 -882
rect 13130 -1258 13164 -882
rect 13248 -1258 13282 -882
rect 13366 -1258 13400 -882
rect 13484 -1258 13518 -882
rect 13602 -1258 13636 -882
rect 12953 -1342 12987 -1308
rect 13071 -1342 13105 -1308
rect 13189 -1342 13223 -1308
rect 13307 -1342 13341 -1308
rect 13425 -1342 13459 -1308
rect 13543 -1342 13577 -1308
rect 13993 -832 14027 -798
rect 14111 -832 14145 -798
rect 14229 -832 14263 -798
rect 14347 -832 14381 -798
rect 14465 -832 14499 -798
rect 14583 -832 14617 -798
rect 13934 -1258 13968 -882
rect 14052 -1258 14086 -882
rect 14170 -1258 14204 -882
rect 14288 -1258 14322 -882
rect 14406 -1258 14440 -882
rect 14524 -1258 14558 -882
rect 14642 -1258 14676 -882
rect 13993 -1342 14027 -1308
rect 14111 -1342 14145 -1308
rect 14229 -1342 14263 -1308
rect 14347 -1342 14381 -1308
rect 14465 -1342 14499 -1308
rect 14583 -1342 14617 -1308
rect 15033 -832 15067 -798
rect 15151 -832 15185 -798
rect 15269 -832 15303 -798
rect 15387 -832 15421 -798
rect 15505 -832 15539 -798
rect 15623 -832 15657 -798
rect 14974 -1258 15008 -882
rect 15092 -1258 15126 -882
rect 15210 -1258 15244 -882
rect 15328 -1258 15362 -882
rect 15446 -1258 15480 -882
rect 15564 -1258 15598 -882
rect 15682 -1258 15716 -882
rect 15033 -1342 15067 -1308
rect 15151 -1342 15185 -1308
rect 15269 -1342 15303 -1308
rect 15387 -1342 15421 -1308
rect 15505 -1342 15539 -1308
rect 15623 -1342 15657 -1308
rect 16073 -832 16107 -798
rect 16191 -832 16225 -798
rect 16309 -832 16343 -798
rect 16427 -832 16461 -798
rect 16545 -832 16579 -798
rect 16663 -832 16697 -798
rect 16014 -1258 16048 -882
rect 16132 -1258 16166 -882
rect 16250 -1258 16284 -882
rect 16368 -1258 16402 -882
rect 16486 -1258 16520 -882
rect 16604 -1258 16638 -882
rect 16722 -1258 16756 -882
rect 16073 -1342 16107 -1308
rect 16191 -1342 16225 -1308
rect 16309 -1342 16343 -1308
rect 16427 -1342 16461 -1308
rect 16545 -1342 16579 -1308
rect 16663 -1342 16697 -1308
rect 17113 -832 17147 -798
rect 17231 -832 17265 -798
rect 17349 -832 17383 -798
rect 17467 -832 17501 -798
rect 17585 -832 17619 -798
rect 17703 -832 17737 -798
rect 17054 -1258 17088 -882
rect 17172 -1258 17206 -882
rect 17290 -1258 17324 -882
rect 17408 -1258 17442 -882
rect 17526 -1258 17560 -882
rect 17644 -1258 17678 -882
rect 17762 -1258 17796 -882
rect 17113 -1342 17147 -1308
rect 17231 -1342 17265 -1308
rect 17349 -1342 17383 -1308
rect 17467 -1342 17501 -1308
rect 17585 -1342 17619 -1308
rect 17703 -1342 17737 -1308
rect 18153 -832 18187 -798
rect 18271 -832 18305 -798
rect 18389 -832 18423 -798
rect 18507 -832 18541 -798
rect 18625 -832 18659 -798
rect 18743 -832 18777 -798
rect 18094 -1258 18128 -882
rect 18212 -1258 18246 -882
rect 18330 -1258 18364 -882
rect 18448 -1258 18482 -882
rect 18566 -1258 18600 -882
rect 18684 -1258 18718 -882
rect 18802 -1258 18836 -882
rect 18153 -1342 18187 -1308
rect 18271 -1342 18305 -1308
rect 18389 -1342 18423 -1308
rect 18507 -1342 18541 -1308
rect 18625 -1342 18659 -1308
rect 18743 -1342 18777 -1308
rect -6186 -1780 -5790 -1754
rect -6186 -1814 -6078 -1780
rect -6078 -1814 -5790 -1780
rect -6186 -1834 -5790 -1814
rect 4282 -1650 4316 -1616
rect 4474 -1650 4508 -1616
rect 4666 -1650 4700 -1616
rect 4234 -2076 4268 -1700
rect 4330 -2076 4364 -1700
rect 4426 -2076 4460 -1700
rect 4522 -2076 4556 -1700
rect 4618 -2076 4652 -1700
rect 4714 -2076 4748 -1700
rect 4810 -2076 4844 -1700
rect 4378 -2160 4412 -2126
rect 4570 -2160 4604 -2126
rect 4762 -2160 4796 -2126
rect 4378 -2268 4412 -2234
rect 4570 -2268 4604 -2234
rect 4762 -2268 4796 -2234
rect 4234 -2694 4268 -2318
rect 4330 -2694 4364 -2318
rect 4426 -2694 4460 -2318
rect 4522 -2694 4556 -2318
rect 4618 -2694 4652 -2318
rect 4714 -2694 4748 -2318
rect 4810 -2694 4844 -2318
rect 4282 -2778 4316 -2744
rect 4474 -2778 4508 -2744
rect 4666 -2778 4700 -2744
rect 5322 -1650 5356 -1616
rect 5514 -1650 5548 -1616
rect 5706 -1650 5740 -1616
rect 5274 -2076 5308 -1700
rect 5370 -2076 5404 -1700
rect 5466 -2076 5500 -1700
rect 5562 -2076 5596 -1700
rect 5658 -2076 5692 -1700
rect 5754 -2076 5788 -1700
rect 5850 -2076 5884 -1700
rect 5418 -2160 5452 -2126
rect 5610 -2160 5644 -2126
rect 5802 -2160 5836 -2126
rect 5418 -2268 5452 -2234
rect 5610 -2268 5644 -2234
rect 5802 -2268 5836 -2234
rect 5274 -2694 5308 -2318
rect 5370 -2694 5404 -2318
rect 5466 -2694 5500 -2318
rect 5562 -2694 5596 -2318
rect 5658 -2694 5692 -2318
rect 5754 -2694 5788 -2318
rect 5850 -2694 5884 -2318
rect 5322 -2778 5356 -2744
rect 5514 -2778 5548 -2744
rect 5706 -2778 5740 -2744
rect 6362 -1650 6396 -1616
rect 6554 -1650 6588 -1616
rect 6746 -1650 6780 -1616
rect 6314 -2076 6348 -1700
rect 6410 -2076 6444 -1700
rect 6506 -2076 6540 -1700
rect 6602 -2076 6636 -1700
rect 6698 -2076 6732 -1700
rect 6794 -2076 6828 -1700
rect 6890 -2076 6924 -1700
rect 6458 -2160 6492 -2126
rect 6650 -2160 6684 -2126
rect 6842 -2160 6876 -2126
rect 6458 -2268 6492 -2234
rect 6650 -2268 6684 -2234
rect 6842 -2268 6876 -2234
rect 6314 -2694 6348 -2318
rect 6410 -2694 6444 -2318
rect 6506 -2694 6540 -2318
rect 6602 -2694 6636 -2318
rect 6698 -2694 6732 -2318
rect 6794 -2694 6828 -2318
rect 6890 -2694 6924 -2318
rect 6362 -2778 6396 -2744
rect 6554 -2778 6588 -2744
rect 6746 -2778 6780 -2744
rect 7402 -1650 7436 -1616
rect 7594 -1650 7628 -1616
rect 7786 -1650 7820 -1616
rect 7354 -2076 7388 -1700
rect 7450 -2076 7484 -1700
rect 7546 -2076 7580 -1700
rect 7642 -2076 7676 -1700
rect 7738 -2076 7772 -1700
rect 7834 -2076 7868 -1700
rect 7930 -2076 7964 -1700
rect 7498 -2160 7532 -2126
rect 7690 -2160 7724 -2126
rect 7882 -2160 7916 -2126
rect 7498 -2268 7532 -2234
rect 7690 -2268 7724 -2234
rect 7882 -2268 7916 -2234
rect 7354 -2694 7388 -2318
rect 7450 -2694 7484 -2318
rect 7546 -2694 7580 -2318
rect 7642 -2694 7676 -2318
rect 7738 -2694 7772 -2318
rect 7834 -2694 7868 -2318
rect 7930 -2694 7964 -2318
rect 7402 -2778 7436 -2744
rect 7594 -2778 7628 -2744
rect 7786 -2778 7820 -2744
rect 8442 -1650 8476 -1616
rect 8634 -1650 8668 -1616
rect 8826 -1650 8860 -1616
rect 8394 -2076 8428 -1700
rect 8490 -2076 8524 -1700
rect 8586 -2076 8620 -1700
rect 8682 -2076 8716 -1700
rect 8778 -2076 8812 -1700
rect 8874 -2076 8908 -1700
rect 8970 -2076 9004 -1700
rect 8538 -2160 8572 -2126
rect 8730 -2160 8764 -2126
rect 8922 -2160 8956 -2126
rect 8538 -2268 8572 -2234
rect 8730 -2268 8764 -2234
rect 8922 -2268 8956 -2234
rect 8394 -2694 8428 -2318
rect 8490 -2694 8524 -2318
rect 8586 -2694 8620 -2318
rect 8682 -2694 8716 -2318
rect 8778 -2694 8812 -2318
rect 8874 -2694 8908 -2318
rect 8970 -2694 9004 -2318
rect 8442 -2778 8476 -2744
rect 8634 -2778 8668 -2744
rect 8826 -2778 8860 -2744
rect 11902 -1650 11936 -1616
rect 12094 -1650 12128 -1616
rect 12286 -1650 12320 -1616
rect 11854 -2076 11888 -1700
rect 11950 -2076 11984 -1700
rect 12046 -2076 12080 -1700
rect 12142 -2076 12176 -1700
rect 12238 -2076 12272 -1700
rect 12334 -2076 12368 -1700
rect 12430 -2076 12464 -1700
rect 11998 -2160 12032 -2126
rect 12190 -2160 12224 -2126
rect 12382 -2160 12416 -2126
rect 11998 -2268 12032 -2234
rect 12190 -2268 12224 -2234
rect 12382 -2268 12416 -2234
rect 11854 -2694 11888 -2318
rect 11950 -2694 11984 -2318
rect 12046 -2694 12080 -2318
rect 12142 -2694 12176 -2318
rect 12238 -2694 12272 -2318
rect 12334 -2694 12368 -2318
rect 12430 -2694 12464 -2318
rect 11902 -2778 11936 -2744
rect 12094 -2778 12128 -2744
rect 12286 -2778 12320 -2744
rect 12942 -1650 12976 -1616
rect 13134 -1650 13168 -1616
rect 13326 -1650 13360 -1616
rect 12894 -2076 12928 -1700
rect 12990 -2076 13024 -1700
rect 13086 -2076 13120 -1700
rect 13182 -2076 13216 -1700
rect 13278 -2076 13312 -1700
rect 13374 -2076 13408 -1700
rect 13470 -2076 13504 -1700
rect 13038 -2160 13072 -2126
rect 13230 -2160 13264 -2126
rect 13422 -2160 13456 -2126
rect 13038 -2268 13072 -2234
rect 13230 -2268 13264 -2234
rect 13422 -2268 13456 -2234
rect 12894 -2694 12928 -2318
rect 12990 -2694 13024 -2318
rect 13086 -2694 13120 -2318
rect 13182 -2694 13216 -2318
rect 13278 -2694 13312 -2318
rect 13374 -2694 13408 -2318
rect 13470 -2694 13504 -2318
rect 12942 -2778 12976 -2744
rect 13134 -2778 13168 -2744
rect 13326 -2778 13360 -2744
rect 13982 -1650 14016 -1616
rect 14174 -1650 14208 -1616
rect 14366 -1650 14400 -1616
rect 13934 -2076 13968 -1700
rect 14030 -2076 14064 -1700
rect 14126 -2076 14160 -1700
rect 14222 -2076 14256 -1700
rect 14318 -2076 14352 -1700
rect 14414 -2076 14448 -1700
rect 14510 -2076 14544 -1700
rect 14078 -2160 14112 -2126
rect 14270 -2160 14304 -2126
rect 14462 -2160 14496 -2126
rect 14078 -2268 14112 -2234
rect 14270 -2268 14304 -2234
rect 14462 -2268 14496 -2234
rect 13934 -2694 13968 -2318
rect 14030 -2694 14064 -2318
rect 14126 -2694 14160 -2318
rect 14222 -2694 14256 -2318
rect 14318 -2694 14352 -2318
rect 14414 -2694 14448 -2318
rect 14510 -2694 14544 -2318
rect 13982 -2778 14016 -2744
rect 14174 -2778 14208 -2744
rect 14366 -2778 14400 -2744
rect 15022 -1650 15056 -1616
rect 15214 -1650 15248 -1616
rect 15406 -1650 15440 -1616
rect 14974 -2076 15008 -1700
rect 15070 -2076 15104 -1700
rect 15166 -2076 15200 -1700
rect 15262 -2076 15296 -1700
rect 15358 -2076 15392 -1700
rect 15454 -2076 15488 -1700
rect 15550 -2076 15584 -1700
rect 15118 -2160 15152 -2126
rect 15310 -2160 15344 -2126
rect 15502 -2160 15536 -2126
rect 15118 -2268 15152 -2234
rect 15310 -2268 15344 -2234
rect 15502 -2268 15536 -2234
rect 14974 -2694 15008 -2318
rect 15070 -2694 15104 -2318
rect 15166 -2694 15200 -2318
rect 15262 -2694 15296 -2318
rect 15358 -2694 15392 -2318
rect 15454 -2694 15488 -2318
rect 15550 -2694 15584 -2318
rect 15022 -2778 15056 -2744
rect 15214 -2778 15248 -2744
rect 15406 -2778 15440 -2744
rect 16062 -1650 16096 -1616
rect 16254 -1650 16288 -1616
rect 16446 -1650 16480 -1616
rect 16014 -2076 16048 -1700
rect 16110 -2076 16144 -1700
rect 16206 -2076 16240 -1700
rect 16302 -2076 16336 -1700
rect 16398 -2076 16432 -1700
rect 16494 -2076 16528 -1700
rect 16590 -2076 16624 -1700
rect 16158 -2160 16192 -2126
rect 16350 -2160 16384 -2126
rect 16542 -2160 16576 -2126
rect 16158 -2268 16192 -2234
rect 16350 -2268 16384 -2234
rect 16542 -2268 16576 -2234
rect 16014 -2694 16048 -2318
rect 16110 -2694 16144 -2318
rect 16206 -2694 16240 -2318
rect 16302 -2694 16336 -2318
rect 16398 -2694 16432 -2318
rect 16494 -2694 16528 -2318
rect 16590 -2694 16624 -2318
rect 16062 -2778 16096 -2744
rect 16254 -2778 16288 -2744
rect 16446 -2778 16480 -2744
rect -7341 -3274 -7307 -3240
rect -7223 -3274 -7189 -3240
rect -7105 -3274 -7071 -3240
rect -6987 -3274 -6953 -3240
rect -6869 -3274 -6835 -3240
rect -6751 -3274 -6717 -3240
rect -7400 -3700 -7366 -3324
rect -7282 -3700 -7248 -3324
rect -7164 -3700 -7130 -3324
rect -7046 -3700 -7012 -3324
rect -6928 -3700 -6894 -3324
rect -6810 -3700 -6776 -3324
rect -6692 -3700 -6658 -3324
rect -7341 -3784 -7307 -3750
rect -7223 -3784 -7189 -3750
rect -7105 -3784 -7071 -3750
rect -6987 -3784 -6953 -3750
rect -6869 -3784 -6835 -3750
rect -6751 -3784 -6717 -3750
rect 4293 -3072 4327 -3038
rect 4411 -3072 4445 -3038
rect 4529 -3072 4563 -3038
rect 4647 -3072 4681 -3038
rect 4765 -3072 4799 -3038
rect 4883 -3072 4917 -3038
rect 4234 -3498 4268 -3122
rect 4352 -3498 4386 -3122
rect 4470 -3498 4504 -3122
rect 4588 -3498 4622 -3122
rect 4706 -3498 4740 -3122
rect 4824 -3498 4858 -3122
rect 4942 -3498 4976 -3122
rect 4293 -3582 4327 -3548
rect 4411 -3582 4445 -3548
rect 4529 -3582 4563 -3548
rect 4647 -3582 4681 -3548
rect 4765 -3582 4799 -3548
rect 4883 -3582 4917 -3548
rect 5333 -3072 5367 -3038
rect 5451 -3072 5485 -3038
rect 5569 -3072 5603 -3038
rect 5687 -3072 5721 -3038
rect 5805 -3072 5839 -3038
rect 5923 -3072 5957 -3038
rect 5274 -3498 5308 -3122
rect 5392 -3498 5426 -3122
rect 5510 -3498 5544 -3122
rect 5628 -3498 5662 -3122
rect 5746 -3498 5780 -3122
rect 5864 -3498 5898 -3122
rect 5982 -3498 6016 -3122
rect 5333 -3582 5367 -3548
rect 5451 -3582 5485 -3548
rect 5569 -3582 5603 -3548
rect 5687 -3582 5721 -3548
rect 5805 -3582 5839 -3548
rect 5923 -3582 5957 -3548
rect 6373 -3072 6407 -3038
rect 6491 -3072 6525 -3038
rect 6609 -3072 6643 -3038
rect 6727 -3072 6761 -3038
rect 6845 -3072 6879 -3038
rect 6963 -3072 6997 -3038
rect 6314 -3498 6348 -3122
rect 6432 -3498 6466 -3122
rect 6550 -3498 6584 -3122
rect 6668 -3498 6702 -3122
rect 6786 -3498 6820 -3122
rect 6904 -3498 6938 -3122
rect 7022 -3498 7056 -3122
rect 6373 -3582 6407 -3548
rect 6491 -3582 6525 -3548
rect 6609 -3582 6643 -3548
rect 6727 -3582 6761 -3548
rect 6845 -3582 6879 -3548
rect 6963 -3582 6997 -3548
rect 7413 -3072 7447 -3038
rect 7531 -3072 7565 -3038
rect 7649 -3072 7683 -3038
rect 7767 -3072 7801 -3038
rect 7885 -3072 7919 -3038
rect 8003 -3072 8037 -3038
rect 7354 -3498 7388 -3122
rect 7472 -3498 7506 -3122
rect 7590 -3498 7624 -3122
rect 7708 -3498 7742 -3122
rect 7826 -3498 7860 -3122
rect 7944 -3498 7978 -3122
rect 8062 -3498 8096 -3122
rect 7413 -3582 7447 -3548
rect 7531 -3582 7565 -3548
rect 7649 -3582 7683 -3548
rect 7767 -3582 7801 -3548
rect 7885 -3582 7919 -3548
rect 8003 -3582 8037 -3548
rect 8453 -3072 8487 -3038
rect 8571 -3072 8605 -3038
rect 8689 -3072 8723 -3038
rect 8807 -3072 8841 -3038
rect 8925 -3072 8959 -3038
rect 9043 -3072 9077 -3038
rect 8394 -3498 8428 -3122
rect 8512 -3498 8546 -3122
rect 8630 -3498 8664 -3122
rect 8748 -3498 8782 -3122
rect 8866 -3498 8900 -3122
rect 8984 -3498 9018 -3122
rect 9102 -3498 9136 -3122
rect 8453 -3582 8487 -3548
rect 8571 -3582 8605 -3548
rect 8689 -3582 8723 -3548
rect 8807 -3582 8841 -3548
rect 8925 -3582 8959 -3548
rect 9043 -3582 9077 -3548
rect 11913 -3072 11947 -3038
rect 12031 -3072 12065 -3038
rect 12149 -3072 12183 -3038
rect 12267 -3072 12301 -3038
rect 12385 -3072 12419 -3038
rect 12503 -3072 12537 -3038
rect 11854 -3498 11888 -3122
rect 11972 -3498 12006 -3122
rect 12090 -3498 12124 -3122
rect 12208 -3498 12242 -3122
rect 12326 -3498 12360 -3122
rect 12444 -3498 12478 -3122
rect 12562 -3498 12596 -3122
rect 11913 -3582 11947 -3548
rect 12031 -3582 12065 -3548
rect 12149 -3582 12183 -3548
rect 12267 -3582 12301 -3548
rect 12385 -3582 12419 -3548
rect 12503 -3582 12537 -3548
rect 12953 -3072 12987 -3038
rect 13071 -3072 13105 -3038
rect 13189 -3072 13223 -3038
rect 13307 -3072 13341 -3038
rect 13425 -3072 13459 -3038
rect 13543 -3072 13577 -3038
rect 12894 -3498 12928 -3122
rect 13012 -3498 13046 -3122
rect 13130 -3498 13164 -3122
rect 13248 -3498 13282 -3122
rect 13366 -3498 13400 -3122
rect 13484 -3498 13518 -3122
rect 13602 -3498 13636 -3122
rect 12953 -3582 12987 -3548
rect 13071 -3582 13105 -3548
rect 13189 -3582 13223 -3548
rect 13307 -3582 13341 -3548
rect 13425 -3582 13459 -3548
rect 13543 -3582 13577 -3548
rect 13993 -3072 14027 -3038
rect 14111 -3072 14145 -3038
rect 14229 -3072 14263 -3038
rect 14347 -3072 14381 -3038
rect 14465 -3072 14499 -3038
rect 14583 -3072 14617 -3038
rect 13934 -3498 13968 -3122
rect 14052 -3498 14086 -3122
rect 14170 -3498 14204 -3122
rect 14288 -3498 14322 -3122
rect 14406 -3498 14440 -3122
rect 14524 -3498 14558 -3122
rect 14642 -3498 14676 -3122
rect 13993 -3582 14027 -3548
rect 14111 -3582 14145 -3548
rect 14229 -3582 14263 -3548
rect 14347 -3582 14381 -3548
rect 14465 -3582 14499 -3548
rect 14583 -3582 14617 -3548
rect 15033 -3072 15067 -3038
rect 15151 -3072 15185 -3038
rect 15269 -3072 15303 -3038
rect 15387 -3072 15421 -3038
rect 15505 -3072 15539 -3038
rect 15623 -3072 15657 -3038
rect 14974 -3498 15008 -3122
rect 15092 -3498 15126 -3122
rect 15210 -3498 15244 -3122
rect 15328 -3498 15362 -3122
rect 15446 -3498 15480 -3122
rect 15564 -3498 15598 -3122
rect 15682 -3498 15716 -3122
rect 15033 -3582 15067 -3548
rect 15151 -3582 15185 -3548
rect 15269 -3582 15303 -3548
rect 15387 -3582 15421 -3548
rect 15505 -3582 15539 -3548
rect 15623 -3582 15657 -3548
rect 16073 -3072 16107 -3038
rect 16191 -3072 16225 -3038
rect 16309 -3072 16343 -3038
rect 16427 -3072 16461 -3038
rect 16545 -3072 16579 -3038
rect 16663 -3072 16697 -3038
rect 16014 -3498 16048 -3122
rect 16132 -3498 16166 -3122
rect 16250 -3498 16284 -3122
rect 16368 -3498 16402 -3122
rect 16486 -3498 16520 -3122
rect 16604 -3498 16638 -3122
rect 16722 -3498 16756 -3122
rect 16073 -3582 16107 -3548
rect 16191 -3582 16225 -3548
rect 16309 -3582 16343 -3548
rect 16427 -3582 16461 -3548
rect 16545 -3582 16579 -3548
rect 16663 -3582 16697 -3548
rect 4924 -3840 5224 -3720
rect 8564 -3840 8864 -3720
rect 12544 -3840 12844 -3720
rect 16184 -3840 16484 -3720
rect -7230 -3886 -6950 -3862
rect -7230 -3982 -6950 -3886
<< metal1 >>
rect -1436 6596 -88 6604
rect -52 6596 360 6604
rect -1436 6588 360 6596
rect 1364 6596 2712 6604
rect 2748 6596 3160 6604
rect 1364 6588 3160 6596
rect -1436 6584 -28 6588
rect -1436 6580 -1418 6584
rect -1168 6580 -1040 6584
rect -1466 6184 -1456 6580
rect -1044 6187 -1040 6580
rect -790 6187 -662 6584
rect -412 6187 -284 6584
rect -34 6192 -28 6584
rect 384 6192 394 6588
rect 1364 6584 2772 6588
rect 1364 6580 1382 6584
rect 1632 6580 1760 6584
rect -34 6187 94 6192
rect 344 6187 360 6192
rect -1044 6184 360 6187
rect 1334 6184 1344 6580
rect 1756 6187 1760 6580
rect 2010 6187 2138 6584
rect 2388 6187 2516 6584
rect 2766 6192 2772 6584
rect 3184 6192 3194 6588
rect 2766 6187 2894 6192
rect 3144 6187 3160 6192
rect 1756 6184 3160 6187
rect -1436 6175 360 6184
rect -1436 6172 -88 6175
rect -52 6172 360 6175
rect 1364 6175 3160 6184
rect 1364 6172 2712 6175
rect 2748 6172 3160 6175
rect 2700 5768 4324 5780
rect -1436 5765 -88 5768
rect -52 5765 360 5768
rect -1436 5753 360 5765
rect -1436 5356 -1418 5753
rect -1168 5356 -1040 5753
rect -790 5744 -662 5753
rect -412 5744 -284 5753
rect -790 5356 -662 5368
rect -412 5356 -284 5368
rect -34 5356 94 5753
rect 344 5356 360 5753
rect -1436 5344 360 5356
rect -1436 5336 -88 5344
rect -52 5336 360 5344
rect 1364 5753 4324 5768
rect 1364 5356 1382 5753
rect 1632 5356 1760 5753
rect 2010 5744 2138 5753
rect 2388 5744 2516 5753
rect 2010 5356 2138 5368
rect 2388 5356 2516 5368
rect 2766 5356 2894 5753
rect 3144 5620 4324 5753
rect 15070 5620 15080 5780
rect 3144 5536 10864 5620
rect 3144 5502 4482 5536
rect 4516 5502 4674 5536
rect 4708 5502 4866 5536
rect 4900 5502 5058 5536
rect 5092 5502 5250 5536
rect 5284 5502 5442 5536
rect 5476 5502 5634 5536
rect 5668 5502 5826 5536
rect 5860 5502 6018 5536
rect 6052 5502 6210 5536
rect 6244 5502 6402 5536
rect 6436 5502 6594 5536
rect 6628 5502 6786 5536
rect 6820 5502 6978 5536
rect 7012 5502 7170 5536
rect 7204 5502 8122 5536
rect 8156 5502 8314 5536
rect 8348 5502 8506 5536
rect 8540 5502 8698 5536
rect 8732 5502 8890 5536
rect 8924 5502 9082 5536
rect 9116 5502 9274 5536
rect 9308 5502 9466 5536
rect 9500 5502 9658 5536
rect 9692 5502 9850 5536
rect 9884 5502 10042 5536
rect 10076 5502 10234 5536
rect 10268 5502 10426 5536
rect 10460 5502 10618 5536
rect 10652 5502 10810 5536
rect 10844 5502 10864 5536
rect 3144 5496 10864 5502
rect 12084 5536 15080 5620
rect 12084 5502 12102 5536
rect 12136 5502 12294 5536
rect 12328 5502 12486 5536
rect 12520 5502 12678 5536
rect 12712 5502 12870 5536
rect 12904 5502 13062 5536
rect 13096 5502 13254 5536
rect 13288 5502 13446 5536
rect 13480 5502 13638 5536
rect 13672 5502 13830 5536
rect 13864 5502 14022 5536
rect 14056 5502 14214 5536
rect 14248 5502 14406 5536
rect 14440 5502 14598 5536
rect 14632 5502 14790 5536
rect 14824 5502 15080 5536
rect 12084 5496 15080 5502
rect 3144 5356 4324 5496
rect 1364 5340 4324 5356
rect 1364 5336 2712 5340
rect 2748 5336 3160 5340
rect -1436 5228 -88 5236
rect -52 5228 360 5236
rect -1436 5220 360 5228
rect 1364 5228 2712 5236
rect 2748 5228 3160 5236
rect 1364 5220 3160 5228
rect -1436 5216 -28 5220
rect -1436 5212 -1418 5216
rect -1168 5212 -1040 5216
rect -1466 4816 -1456 5212
rect -1044 4819 -1040 5212
rect -790 4819 -662 5216
rect -412 4819 -284 5216
rect -34 4824 -28 5216
rect 384 4824 394 5220
rect 1364 5216 2772 5220
rect 1364 5212 1382 5216
rect 1632 5212 1760 5216
rect -34 4819 94 4824
rect 344 4819 360 4824
rect -1044 4816 360 4819
rect 1334 4816 1344 5212
rect 1756 4819 1760 5212
rect 2010 4819 2138 5216
rect 2388 4819 2516 5216
rect 2766 4824 2772 5216
rect 3184 4824 3194 5220
rect 4160 5032 4324 5340
rect 4428 5452 4474 5464
rect 4428 5248 4434 5452
rect 4468 5248 4474 5452
rect 4510 5284 4520 5468
rect 4572 5284 4582 5468
rect 4620 5452 4666 5464
rect 4414 5064 4424 5248
rect 4476 5064 4486 5248
rect 4524 5076 4530 5284
rect 4564 5076 4570 5284
rect 4620 5248 4626 5452
rect 4660 5248 4666 5452
rect 4702 5284 4712 5468
rect 4764 5284 4774 5468
rect 4812 5452 4858 5464
rect 4524 5064 4570 5076
rect 4606 5064 4616 5248
rect 4668 5064 4678 5248
rect 4716 5076 4722 5284
rect 4756 5076 4762 5284
rect 4812 5248 4818 5452
rect 4852 5248 4858 5452
rect 4894 5284 4904 5468
rect 4956 5284 4966 5468
rect 5004 5452 5050 5464
rect 4716 5064 4762 5076
rect 4798 5064 4808 5248
rect 4860 5064 4870 5248
rect 4908 5076 4914 5284
rect 4948 5076 4954 5284
rect 5004 5248 5010 5452
rect 5044 5248 5050 5452
rect 5086 5284 5096 5468
rect 5148 5284 5158 5468
rect 5196 5452 5242 5464
rect 4908 5064 4954 5076
rect 4990 5064 5000 5248
rect 5052 5064 5062 5248
rect 5100 5076 5106 5284
rect 5140 5076 5146 5284
rect 5196 5248 5202 5452
rect 5236 5248 5242 5452
rect 5278 5284 5288 5468
rect 5340 5284 5350 5468
rect 5388 5452 5434 5464
rect 5100 5064 5146 5076
rect 5182 5064 5192 5248
rect 5244 5064 5254 5248
rect 5292 5076 5298 5284
rect 5332 5076 5338 5284
rect 5388 5248 5394 5452
rect 5428 5248 5434 5452
rect 5470 5284 5480 5468
rect 5532 5284 5542 5468
rect 5580 5452 5626 5464
rect 5292 5064 5338 5076
rect 5374 5064 5384 5248
rect 5436 5064 5446 5248
rect 5484 5076 5490 5284
rect 5524 5076 5530 5284
rect 5580 5248 5586 5452
rect 5620 5248 5626 5452
rect 5662 5284 5672 5468
rect 5724 5284 5734 5468
rect 5772 5452 5818 5464
rect 5484 5064 5530 5076
rect 5566 5064 5576 5248
rect 5628 5064 5638 5248
rect 5676 5076 5682 5284
rect 5716 5076 5722 5284
rect 5772 5248 5778 5452
rect 5812 5248 5818 5452
rect 5854 5284 5864 5468
rect 5916 5284 5926 5468
rect 5964 5452 6010 5464
rect 5676 5064 5722 5076
rect 5758 5064 5768 5248
rect 5820 5064 5830 5248
rect 5868 5076 5874 5284
rect 5908 5076 5914 5284
rect 5964 5248 5970 5452
rect 6004 5248 6010 5452
rect 6046 5284 6056 5468
rect 6108 5284 6118 5468
rect 6156 5452 6202 5464
rect 5868 5064 5914 5076
rect 5950 5064 5960 5248
rect 6012 5064 6022 5248
rect 6060 5076 6066 5284
rect 6100 5076 6106 5284
rect 6156 5248 6162 5452
rect 6196 5248 6202 5452
rect 6238 5284 6248 5468
rect 6300 5284 6310 5468
rect 6348 5452 6394 5464
rect 6060 5064 6106 5076
rect 6142 5064 6152 5248
rect 6204 5064 6214 5248
rect 6252 5076 6258 5284
rect 6292 5076 6298 5284
rect 6348 5248 6354 5452
rect 6388 5248 6394 5452
rect 6430 5284 6440 5468
rect 6492 5284 6502 5468
rect 6540 5452 6586 5464
rect 6252 5064 6298 5076
rect 6334 5064 6344 5248
rect 6396 5064 6406 5248
rect 6444 5076 6450 5284
rect 6484 5076 6490 5284
rect 6540 5248 6546 5452
rect 6580 5248 6586 5452
rect 6622 5284 6632 5468
rect 6684 5284 6694 5468
rect 6732 5452 6778 5464
rect 6444 5064 6490 5076
rect 6526 5064 6536 5248
rect 6588 5064 6598 5248
rect 6636 5076 6642 5284
rect 6676 5076 6682 5284
rect 6732 5248 6738 5452
rect 6772 5248 6778 5452
rect 6814 5284 6824 5468
rect 6876 5284 6886 5468
rect 6924 5452 6970 5464
rect 6636 5064 6682 5076
rect 6718 5064 6728 5248
rect 6780 5064 6790 5248
rect 6828 5076 6834 5284
rect 6868 5076 6874 5284
rect 6924 5248 6930 5452
rect 6964 5248 6970 5452
rect 7006 5284 7016 5468
rect 7068 5284 7078 5468
rect 7116 5452 7162 5464
rect 6828 5064 6874 5076
rect 6910 5064 6920 5248
rect 6972 5064 6982 5248
rect 7020 5076 7026 5284
rect 7060 5076 7066 5284
rect 7116 5248 7122 5452
rect 7156 5248 7162 5452
rect 7198 5284 7208 5468
rect 7260 5284 7270 5468
rect 7308 5452 7354 5464
rect 7020 5064 7066 5076
rect 7102 5064 7112 5248
rect 7164 5064 7174 5248
rect 7212 5076 7218 5284
rect 7252 5076 7258 5284
rect 7308 5248 7314 5452
rect 7348 5248 7354 5452
rect 7212 5064 7258 5076
rect 7294 5064 7304 5248
rect 7356 5064 7366 5248
rect 7468 5032 7916 5496
rect 8068 5452 8114 5464
rect 8068 5248 8074 5452
rect 8108 5248 8114 5452
rect 8150 5284 8160 5468
rect 8212 5284 8222 5468
rect 8260 5452 8306 5464
rect 8054 5064 8064 5248
rect 8116 5064 8126 5248
rect 8164 5076 8170 5284
rect 8204 5076 8210 5284
rect 8260 5248 8266 5452
rect 8300 5248 8306 5452
rect 8342 5284 8352 5468
rect 8404 5284 8414 5468
rect 8452 5452 8498 5464
rect 8164 5064 8210 5076
rect 8246 5064 8256 5248
rect 8308 5064 8318 5248
rect 8356 5076 8362 5284
rect 8396 5076 8402 5284
rect 8452 5248 8458 5452
rect 8492 5248 8498 5452
rect 8534 5284 8544 5468
rect 8596 5284 8606 5468
rect 8644 5452 8690 5464
rect 8356 5064 8402 5076
rect 8438 5064 8448 5248
rect 8500 5064 8510 5248
rect 8548 5076 8554 5284
rect 8588 5076 8594 5284
rect 8644 5248 8650 5452
rect 8684 5248 8690 5452
rect 8726 5284 8736 5468
rect 8788 5284 8798 5468
rect 8836 5452 8882 5464
rect 8548 5064 8594 5076
rect 8630 5064 8640 5248
rect 8692 5064 8702 5248
rect 8740 5076 8746 5284
rect 8780 5076 8786 5284
rect 8836 5248 8842 5452
rect 8876 5248 8882 5452
rect 8918 5284 8928 5468
rect 8980 5284 8990 5468
rect 9028 5452 9074 5464
rect 8740 5064 8786 5076
rect 8822 5064 8832 5248
rect 8884 5064 8894 5248
rect 8932 5076 8938 5284
rect 8972 5076 8978 5284
rect 9028 5248 9034 5452
rect 9068 5248 9074 5452
rect 9110 5284 9120 5468
rect 9172 5284 9182 5468
rect 9220 5452 9266 5464
rect 8932 5064 8978 5076
rect 9014 5064 9024 5248
rect 9076 5064 9086 5248
rect 9124 5076 9130 5284
rect 9164 5076 9170 5284
rect 9220 5248 9226 5452
rect 9260 5248 9266 5452
rect 9302 5284 9312 5468
rect 9364 5284 9374 5468
rect 9412 5452 9458 5464
rect 9124 5064 9170 5076
rect 9206 5064 9216 5248
rect 9268 5064 9278 5248
rect 9316 5076 9322 5284
rect 9356 5076 9362 5284
rect 9412 5248 9418 5452
rect 9452 5248 9458 5452
rect 9494 5284 9504 5468
rect 9556 5284 9566 5468
rect 9604 5452 9650 5464
rect 9316 5064 9362 5076
rect 9398 5064 9408 5248
rect 9460 5064 9470 5248
rect 9508 5076 9514 5284
rect 9548 5076 9554 5284
rect 9604 5248 9610 5452
rect 9644 5248 9650 5452
rect 9686 5284 9696 5468
rect 9748 5284 9758 5468
rect 9796 5452 9842 5464
rect 9508 5064 9554 5076
rect 9590 5064 9600 5248
rect 9652 5064 9662 5248
rect 9700 5076 9706 5284
rect 9740 5076 9746 5284
rect 9796 5248 9802 5452
rect 9836 5248 9842 5452
rect 9878 5284 9888 5468
rect 9940 5284 9950 5468
rect 9988 5452 10034 5464
rect 9700 5064 9746 5076
rect 9782 5064 9792 5248
rect 9844 5064 9854 5248
rect 9892 5076 9898 5284
rect 9932 5076 9938 5284
rect 9988 5248 9994 5452
rect 10028 5248 10034 5452
rect 10070 5284 10080 5468
rect 10132 5284 10142 5468
rect 10180 5452 10226 5464
rect 9892 5064 9938 5076
rect 9974 5064 9984 5248
rect 10036 5064 10046 5248
rect 10084 5076 10090 5284
rect 10124 5076 10130 5284
rect 10180 5248 10186 5452
rect 10220 5248 10226 5452
rect 10262 5284 10272 5468
rect 10324 5284 10334 5468
rect 10372 5452 10418 5464
rect 10084 5064 10130 5076
rect 10166 5064 10176 5248
rect 10228 5064 10238 5248
rect 10276 5076 10282 5284
rect 10316 5076 10322 5284
rect 10372 5248 10378 5452
rect 10412 5248 10418 5452
rect 10454 5284 10464 5468
rect 10516 5284 10526 5468
rect 10564 5452 10610 5464
rect 10276 5064 10322 5076
rect 10358 5064 10368 5248
rect 10420 5064 10430 5248
rect 10468 5076 10474 5284
rect 10508 5076 10514 5284
rect 10564 5248 10570 5452
rect 10604 5248 10610 5452
rect 10646 5284 10656 5468
rect 10708 5284 10718 5468
rect 10756 5452 10802 5464
rect 10468 5064 10514 5076
rect 10550 5064 10560 5248
rect 10612 5064 10622 5248
rect 10660 5076 10666 5284
rect 10700 5076 10706 5284
rect 10756 5248 10762 5452
rect 10796 5248 10802 5452
rect 10838 5284 10848 5468
rect 10900 5284 10910 5468
rect 10948 5452 10994 5464
rect 10660 5064 10706 5076
rect 10742 5064 10752 5248
rect 10804 5064 10814 5248
rect 10852 5076 10858 5284
rect 10892 5076 10898 5284
rect 10948 5248 10954 5452
rect 10988 5248 10994 5452
rect 12048 5452 12094 5464
rect 12048 5248 12054 5452
rect 12088 5248 12094 5452
rect 12130 5284 12140 5468
rect 12192 5284 12202 5468
rect 12240 5452 12286 5464
rect 10852 5064 10898 5076
rect 10934 5064 10944 5248
rect 10996 5064 11006 5248
rect 12034 5064 12044 5248
rect 12096 5064 12106 5248
rect 12144 5076 12150 5284
rect 12184 5076 12190 5284
rect 12240 5248 12246 5452
rect 12280 5248 12286 5452
rect 12322 5284 12332 5468
rect 12384 5284 12394 5468
rect 12432 5452 12478 5464
rect 12144 5064 12190 5076
rect 12226 5064 12236 5248
rect 12288 5064 12298 5248
rect 12336 5076 12342 5284
rect 12376 5076 12382 5284
rect 12432 5248 12438 5452
rect 12472 5248 12478 5452
rect 12514 5284 12524 5468
rect 12576 5284 12586 5468
rect 12624 5452 12670 5464
rect 12336 5064 12382 5076
rect 12418 5064 12428 5248
rect 12480 5064 12490 5248
rect 12528 5076 12534 5284
rect 12568 5076 12574 5284
rect 12624 5248 12630 5452
rect 12664 5248 12670 5452
rect 12706 5284 12716 5468
rect 12768 5284 12778 5468
rect 12816 5452 12862 5464
rect 12528 5064 12574 5076
rect 12610 5064 12620 5248
rect 12672 5064 12682 5248
rect 12720 5076 12726 5284
rect 12760 5076 12766 5284
rect 12816 5248 12822 5452
rect 12856 5248 12862 5452
rect 12898 5284 12908 5468
rect 12960 5284 12970 5468
rect 13008 5452 13054 5464
rect 12720 5064 12766 5076
rect 12802 5064 12812 5248
rect 12864 5064 12874 5248
rect 12912 5076 12918 5284
rect 12952 5076 12958 5284
rect 13008 5248 13014 5452
rect 13048 5248 13054 5452
rect 13090 5284 13100 5468
rect 13152 5284 13162 5468
rect 13200 5452 13246 5464
rect 12912 5064 12958 5076
rect 12994 5064 13004 5248
rect 13056 5064 13066 5248
rect 13104 5076 13110 5284
rect 13144 5076 13150 5284
rect 13200 5248 13206 5452
rect 13240 5248 13246 5452
rect 13282 5284 13292 5468
rect 13344 5284 13354 5468
rect 13392 5452 13438 5464
rect 13104 5064 13150 5076
rect 13186 5064 13196 5248
rect 13248 5064 13258 5248
rect 13296 5076 13302 5284
rect 13336 5076 13342 5284
rect 13392 5248 13398 5452
rect 13432 5248 13438 5452
rect 13474 5284 13484 5468
rect 13536 5284 13546 5468
rect 13584 5452 13630 5464
rect 13296 5064 13342 5076
rect 13378 5064 13388 5248
rect 13440 5064 13450 5248
rect 13488 5076 13494 5284
rect 13528 5076 13534 5284
rect 13584 5248 13590 5452
rect 13624 5248 13630 5452
rect 13666 5284 13676 5468
rect 13728 5284 13738 5468
rect 13776 5452 13822 5464
rect 13488 5064 13534 5076
rect 13570 5064 13580 5248
rect 13632 5064 13642 5248
rect 13680 5076 13686 5284
rect 13720 5076 13726 5284
rect 13776 5248 13782 5452
rect 13816 5248 13822 5452
rect 13858 5284 13868 5468
rect 13920 5284 13930 5468
rect 13968 5452 14014 5464
rect 13680 5064 13726 5076
rect 13762 5064 13772 5248
rect 13824 5064 13834 5248
rect 13872 5076 13878 5284
rect 13912 5076 13918 5284
rect 13968 5248 13974 5452
rect 14008 5248 14014 5452
rect 14050 5284 14060 5468
rect 14112 5284 14122 5468
rect 14160 5452 14206 5464
rect 13872 5064 13918 5076
rect 13954 5064 13964 5248
rect 14016 5064 14026 5248
rect 14064 5076 14070 5284
rect 14104 5076 14110 5284
rect 14160 5248 14166 5452
rect 14200 5248 14206 5452
rect 14242 5284 14252 5468
rect 14304 5284 14314 5468
rect 14352 5452 14398 5464
rect 14064 5064 14110 5076
rect 14146 5064 14156 5248
rect 14208 5064 14218 5248
rect 14256 5076 14262 5284
rect 14296 5076 14302 5284
rect 14352 5248 14358 5452
rect 14392 5248 14398 5452
rect 14434 5284 14444 5468
rect 14496 5284 14506 5468
rect 14544 5452 14590 5464
rect 14256 5064 14302 5076
rect 14338 5064 14348 5248
rect 14400 5064 14410 5248
rect 14448 5076 14454 5284
rect 14488 5076 14494 5284
rect 14544 5248 14550 5452
rect 14584 5248 14590 5452
rect 14626 5284 14636 5468
rect 14688 5284 14698 5468
rect 14736 5452 14782 5464
rect 14448 5064 14494 5076
rect 14530 5064 14540 5248
rect 14592 5064 14602 5248
rect 14640 5076 14646 5284
rect 14680 5076 14686 5284
rect 14736 5248 14742 5452
rect 14776 5248 14782 5452
rect 14818 5284 14828 5468
rect 14880 5284 14890 5468
rect 14928 5452 14974 5464
rect 14640 5064 14686 5076
rect 14722 5064 14732 5248
rect 14784 5064 14794 5248
rect 14832 5076 14838 5284
rect 14872 5076 14878 5284
rect 14928 5248 14934 5452
rect 14968 5248 14974 5452
rect 15070 5420 15080 5496
rect 15540 5620 15550 5780
rect 15540 5536 18484 5620
rect 15540 5502 15742 5536
rect 15776 5502 15934 5536
rect 15968 5502 16126 5536
rect 16160 5502 16318 5536
rect 16352 5502 16510 5536
rect 16544 5502 16702 5536
rect 16736 5502 16894 5536
rect 16928 5502 17086 5536
rect 17120 5502 17278 5536
rect 17312 5502 17470 5536
rect 17504 5502 17662 5536
rect 17696 5502 17854 5536
rect 17888 5502 18046 5536
rect 18080 5502 18238 5536
rect 18272 5502 18430 5536
rect 18464 5502 18484 5536
rect 15540 5496 18484 5502
rect 15540 5420 15550 5496
rect 15688 5452 15734 5464
rect 14832 5064 14878 5076
rect 14914 5064 14924 5248
rect 14976 5064 14986 5248
rect 15088 5032 15536 5420
rect 15688 5248 15694 5452
rect 15728 5248 15734 5452
rect 15770 5284 15780 5468
rect 15832 5284 15842 5468
rect 15880 5452 15926 5464
rect 15674 5064 15684 5248
rect 15736 5064 15746 5248
rect 15784 5076 15790 5284
rect 15824 5076 15830 5284
rect 15880 5248 15886 5452
rect 15920 5248 15926 5452
rect 15962 5284 15972 5468
rect 16024 5284 16034 5468
rect 16072 5452 16118 5464
rect 15784 5064 15830 5076
rect 15866 5064 15876 5248
rect 15928 5064 15938 5248
rect 15976 5076 15982 5284
rect 16016 5076 16022 5284
rect 16072 5248 16078 5452
rect 16112 5248 16118 5452
rect 16154 5284 16164 5468
rect 16216 5284 16226 5468
rect 16264 5452 16310 5464
rect 15976 5064 16022 5076
rect 16058 5064 16068 5248
rect 16120 5064 16130 5248
rect 16168 5076 16174 5284
rect 16208 5076 16214 5284
rect 16264 5248 16270 5452
rect 16304 5248 16310 5452
rect 16346 5284 16356 5468
rect 16408 5284 16418 5468
rect 16456 5452 16502 5464
rect 16168 5064 16214 5076
rect 16250 5064 16260 5248
rect 16312 5064 16322 5248
rect 16360 5076 16366 5284
rect 16400 5076 16406 5284
rect 16456 5248 16462 5452
rect 16496 5248 16502 5452
rect 16538 5284 16548 5468
rect 16600 5284 16610 5468
rect 16648 5452 16694 5464
rect 16360 5064 16406 5076
rect 16442 5064 16452 5248
rect 16504 5064 16514 5248
rect 16552 5076 16558 5284
rect 16592 5076 16598 5284
rect 16648 5248 16654 5452
rect 16688 5248 16694 5452
rect 16730 5284 16740 5468
rect 16792 5284 16802 5468
rect 16840 5452 16886 5464
rect 16552 5064 16598 5076
rect 16634 5064 16644 5248
rect 16696 5064 16706 5248
rect 16744 5076 16750 5284
rect 16784 5076 16790 5284
rect 16840 5248 16846 5452
rect 16880 5248 16886 5452
rect 16922 5284 16932 5468
rect 16984 5284 16994 5468
rect 17032 5452 17078 5464
rect 16744 5064 16790 5076
rect 16826 5064 16836 5248
rect 16888 5064 16898 5248
rect 16936 5076 16942 5284
rect 16976 5076 16982 5284
rect 17032 5248 17038 5452
rect 17072 5248 17078 5452
rect 17114 5284 17124 5468
rect 17176 5284 17186 5468
rect 17224 5452 17270 5464
rect 16936 5064 16982 5076
rect 17018 5064 17028 5248
rect 17080 5064 17090 5248
rect 17128 5076 17134 5284
rect 17168 5076 17174 5284
rect 17224 5248 17230 5452
rect 17264 5248 17270 5452
rect 17306 5284 17316 5468
rect 17368 5284 17378 5468
rect 17416 5452 17462 5464
rect 17128 5064 17174 5076
rect 17210 5064 17220 5248
rect 17272 5064 17282 5248
rect 17320 5076 17326 5284
rect 17360 5076 17366 5284
rect 17416 5248 17422 5452
rect 17456 5248 17462 5452
rect 17498 5284 17508 5468
rect 17560 5284 17570 5468
rect 17608 5452 17654 5464
rect 17320 5064 17366 5076
rect 17402 5064 17412 5248
rect 17464 5064 17474 5248
rect 17512 5076 17518 5284
rect 17552 5076 17558 5284
rect 17608 5248 17614 5452
rect 17648 5248 17654 5452
rect 17690 5284 17700 5468
rect 17752 5284 17762 5468
rect 17800 5452 17846 5464
rect 17512 5064 17558 5076
rect 17594 5064 17604 5248
rect 17656 5064 17666 5248
rect 17704 5076 17710 5284
rect 17744 5076 17750 5284
rect 17800 5248 17806 5452
rect 17840 5248 17846 5452
rect 17882 5284 17892 5468
rect 17944 5284 17954 5468
rect 17992 5452 18038 5464
rect 17704 5064 17750 5076
rect 17786 5064 17796 5248
rect 17848 5064 17858 5248
rect 17896 5076 17902 5284
rect 17936 5076 17942 5284
rect 17992 5248 17998 5452
rect 18032 5248 18038 5452
rect 18074 5284 18084 5468
rect 18136 5284 18146 5468
rect 18184 5452 18230 5464
rect 17896 5064 17942 5076
rect 17978 5064 17988 5248
rect 18040 5064 18050 5248
rect 18088 5076 18094 5284
rect 18128 5076 18134 5284
rect 18184 5248 18190 5452
rect 18224 5248 18230 5452
rect 18266 5284 18276 5468
rect 18328 5284 18338 5468
rect 18376 5452 18422 5464
rect 18088 5064 18134 5076
rect 18170 5064 18180 5248
rect 18232 5064 18242 5248
rect 18280 5076 18286 5284
rect 18320 5076 18326 5284
rect 18376 5248 18382 5452
rect 18416 5248 18422 5452
rect 18458 5284 18468 5468
rect 18520 5284 18530 5468
rect 18568 5452 18614 5464
rect 18280 5064 18326 5076
rect 18362 5064 18372 5248
rect 18424 5064 18434 5248
rect 18472 5076 18478 5284
rect 18512 5076 18518 5284
rect 18568 5248 18574 5452
rect 18608 5248 18614 5452
rect 18472 5064 18518 5076
rect 18554 5064 18564 5248
rect 18616 5064 18626 5248
rect 4160 5026 10960 5032
rect 4160 4992 4578 5026
rect 4612 4992 4770 5026
rect 4804 4992 4962 5026
rect 4996 4992 5154 5026
rect 5188 4992 5346 5026
rect 5380 4992 5538 5026
rect 5572 4992 5730 5026
rect 5764 4992 5922 5026
rect 5956 4992 6114 5026
rect 6148 4992 6306 5026
rect 6340 4992 6498 5026
rect 6532 4992 6690 5026
rect 6724 4992 6882 5026
rect 6916 4992 7074 5026
rect 7108 4992 7266 5026
rect 7300 4992 8218 5026
rect 8252 4992 8410 5026
rect 8444 4992 8602 5026
rect 8636 4992 8794 5026
rect 8828 4992 8986 5026
rect 9020 4992 9178 5026
rect 9212 4992 9370 5026
rect 9404 4992 9562 5026
rect 9596 4992 9754 5026
rect 9788 4992 9946 5026
rect 9980 4992 10138 5026
rect 10172 4992 10330 5026
rect 10364 4992 10522 5026
rect 10556 4992 10714 5026
rect 10748 4992 10906 5026
rect 10940 4992 10960 5026
rect 4160 4918 10960 4992
rect 4160 4884 4578 4918
rect 4612 4884 4770 4918
rect 4804 4884 4962 4918
rect 4996 4884 5154 4918
rect 5188 4884 5346 4918
rect 5380 4884 5538 4918
rect 5572 4884 5730 4918
rect 5764 4884 5922 4918
rect 5956 4884 6114 4918
rect 6148 4884 6306 4918
rect 6340 4884 6498 4918
rect 6532 4884 6690 4918
rect 6724 4884 6882 4918
rect 6916 4884 7074 4918
rect 7108 4884 7266 4918
rect 7300 4884 8218 4918
rect 8252 4884 8410 4918
rect 8444 4884 8602 4918
rect 8636 4884 8794 4918
rect 8828 4884 8986 4918
rect 9020 4884 9178 4918
rect 9212 4884 9370 4918
rect 9404 4884 9562 4918
rect 9596 4884 9754 4918
rect 9788 4884 9946 4918
rect 9980 4884 10138 4918
rect 10172 4884 10330 4918
rect 10364 4884 10522 4918
rect 10556 4884 10714 4918
rect 10748 4884 10906 4918
rect 10940 4884 10960 4918
rect 4160 4876 10960 4884
rect 12180 5026 18580 5032
rect 12180 4992 12198 5026
rect 12232 4992 12390 5026
rect 12424 4992 12582 5026
rect 12616 4992 12774 5026
rect 12808 4992 12966 5026
rect 13000 4992 13158 5026
rect 13192 4992 13350 5026
rect 13384 4992 13542 5026
rect 13576 4992 13734 5026
rect 13768 4992 13926 5026
rect 13960 4992 14118 5026
rect 14152 4992 14310 5026
rect 14344 4992 14502 5026
rect 14536 4992 14694 5026
rect 14728 4992 14886 5026
rect 14920 4992 15838 5026
rect 15872 4992 16030 5026
rect 16064 4992 16222 5026
rect 16256 4992 16414 5026
rect 16448 4992 16606 5026
rect 16640 4992 16798 5026
rect 16832 4992 16990 5026
rect 17024 4992 17182 5026
rect 17216 4992 17374 5026
rect 17408 4992 17566 5026
rect 17600 4992 17758 5026
rect 17792 4992 17950 5026
rect 17984 4992 18142 5026
rect 18176 4992 18334 5026
rect 18368 4992 18526 5026
rect 18560 4992 18580 5026
rect 12180 4918 18580 4992
rect 12180 4884 12198 4918
rect 12232 4884 12390 4918
rect 12424 4884 12582 4918
rect 12616 4884 12774 4918
rect 12808 4884 12966 4918
rect 13000 4884 13158 4918
rect 13192 4884 13350 4918
rect 13384 4884 13542 4918
rect 13576 4884 13734 4918
rect 13768 4884 13926 4918
rect 13960 4884 14118 4918
rect 14152 4884 14310 4918
rect 14344 4884 14502 4918
rect 14536 4884 14694 4918
rect 14728 4884 14886 4918
rect 14920 4884 15838 4918
rect 15872 4884 16030 4918
rect 16064 4884 16222 4918
rect 16256 4884 16414 4918
rect 16448 4884 16606 4918
rect 16640 4884 16798 4918
rect 16832 4884 16990 4918
rect 17024 4884 17182 4918
rect 17216 4884 17374 4918
rect 17408 4884 17566 4918
rect 17600 4884 17758 4918
rect 17792 4884 17950 4918
rect 17984 4884 18142 4918
rect 18176 4884 18334 4918
rect 18368 4884 18526 4918
rect 18560 4884 18580 4918
rect 12180 4876 18580 4884
rect 2766 4819 2894 4824
rect 3144 4819 3160 4824
rect 1756 4816 3160 4819
rect -1436 4807 360 4816
rect -1436 4804 -88 4807
rect -52 4804 360 4807
rect 1364 4807 3160 4816
rect 1364 4804 2712 4807
rect 2748 4804 3160 4807
rect 4160 4416 4324 4876
rect 4428 4834 4474 4846
rect 4428 4628 4434 4834
rect 4468 4628 4474 4834
rect 4510 4664 4520 4848
rect 4572 4664 4582 4848
rect 4620 4834 4666 4846
rect 4414 4444 4424 4628
rect 4476 4444 4486 4628
rect 4524 4458 4530 4664
rect 4564 4458 4570 4664
rect 4620 4628 4626 4834
rect 4660 4628 4666 4834
rect 4702 4664 4712 4848
rect 4764 4664 4774 4848
rect 4812 4834 4858 4846
rect 4524 4446 4570 4458
rect 4606 4444 4616 4628
rect 4668 4444 4678 4628
rect 4716 4458 4722 4664
rect 4756 4458 4762 4664
rect 4812 4628 4818 4834
rect 4852 4628 4858 4834
rect 4894 4664 4904 4848
rect 4956 4664 4966 4848
rect 5004 4834 5050 4846
rect 4716 4446 4762 4458
rect 4798 4444 4808 4628
rect 4860 4444 4870 4628
rect 4908 4458 4914 4664
rect 4948 4458 4954 4664
rect 5004 4628 5010 4834
rect 5044 4628 5050 4834
rect 5086 4664 5096 4848
rect 5148 4664 5158 4848
rect 5196 4834 5242 4846
rect 4908 4446 4954 4458
rect 4990 4444 5000 4628
rect 5052 4444 5062 4628
rect 5100 4458 5106 4664
rect 5140 4458 5146 4664
rect 5196 4628 5202 4834
rect 5236 4628 5242 4834
rect 5278 4664 5288 4848
rect 5340 4664 5350 4848
rect 5388 4834 5434 4846
rect 5100 4446 5146 4458
rect 5182 4444 5192 4628
rect 5244 4444 5254 4628
rect 5292 4458 5298 4664
rect 5332 4458 5338 4664
rect 5388 4628 5394 4834
rect 5428 4628 5434 4834
rect 5470 4664 5480 4848
rect 5532 4664 5542 4848
rect 5580 4834 5626 4846
rect 5292 4446 5338 4458
rect 5374 4444 5384 4628
rect 5436 4444 5446 4628
rect 5484 4458 5490 4664
rect 5524 4458 5530 4664
rect 5580 4628 5586 4834
rect 5620 4628 5626 4834
rect 5662 4664 5672 4848
rect 5724 4664 5734 4848
rect 5772 4834 5818 4846
rect 5484 4446 5530 4458
rect 5566 4444 5576 4628
rect 5628 4444 5638 4628
rect 5676 4458 5682 4664
rect 5716 4458 5722 4664
rect 5772 4628 5778 4834
rect 5812 4628 5818 4834
rect 5854 4664 5864 4848
rect 5916 4664 5926 4848
rect 5964 4834 6010 4846
rect 5676 4446 5722 4458
rect 5758 4444 5768 4628
rect 5820 4444 5830 4628
rect 5868 4458 5874 4664
rect 5908 4458 5914 4664
rect 5964 4628 5970 4834
rect 6004 4628 6010 4834
rect 6046 4664 6056 4848
rect 6108 4664 6118 4848
rect 6156 4834 6202 4846
rect 5868 4446 5914 4458
rect 5950 4444 5960 4628
rect 6012 4444 6022 4628
rect 6060 4458 6066 4664
rect 6100 4458 6106 4664
rect 6156 4628 6162 4834
rect 6196 4628 6202 4834
rect 6238 4664 6248 4848
rect 6300 4664 6310 4848
rect 6348 4834 6394 4846
rect 6060 4446 6106 4458
rect 6142 4444 6152 4628
rect 6204 4444 6214 4628
rect 6252 4458 6258 4664
rect 6292 4458 6298 4664
rect 6348 4628 6354 4834
rect 6388 4628 6394 4834
rect 6430 4664 6440 4848
rect 6492 4664 6502 4848
rect 6540 4834 6586 4846
rect 6252 4446 6298 4458
rect 6334 4444 6344 4628
rect 6396 4444 6406 4628
rect 6444 4458 6450 4664
rect 6484 4458 6490 4664
rect 6540 4628 6546 4834
rect 6580 4628 6586 4834
rect 6622 4664 6632 4848
rect 6684 4664 6694 4848
rect 6732 4834 6778 4846
rect 6444 4446 6490 4458
rect 6526 4444 6536 4628
rect 6588 4444 6598 4628
rect 6636 4458 6642 4664
rect 6676 4458 6682 4664
rect 6732 4628 6738 4834
rect 6772 4628 6778 4834
rect 6814 4664 6824 4848
rect 6876 4664 6886 4848
rect 6924 4834 6970 4846
rect 6636 4446 6682 4458
rect 6718 4444 6728 4628
rect 6780 4444 6790 4628
rect 6828 4458 6834 4664
rect 6868 4458 6874 4664
rect 6924 4628 6930 4834
rect 6964 4628 6970 4834
rect 7006 4664 7016 4848
rect 7068 4664 7078 4848
rect 7116 4834 7162 4846
rect 6828 4446 6874 4458
rect 6910 4444 6920 4628
rect 6972 4444 6982 4628
rect 7020 4458 7026 4664
rect 7060 4458 7066 4664
rect 7116 4628 7122 4834
rect 7156 4628 7162 4834
rect 7198 4664 7208 4848
rect 7260 4664 7270 4848
rect 7308 4834 7354 4846
rect 7020 4446 7066 4458
rect 7102 4444 7112 4628
rect 7164 4444 7174 4628
rect 7212 4458 7218 4664
rect 7252 4458 7258 4664
rect 7308 4628 7314 4834
rect 7348 4628 7354 4834
rect 7212 4446 7258 4458
rect 7294 4444 7304 4628
rect 7356 4444 7366 4628
rect 7468 4416 7916 4876
rect 8068 4834 8114 4846
rect 8068 4628 8074 4834
rect 8108 4628 8114 4834
rect 8150 4664 8160 4848
rect 8212 4664 8222 4848
rect 8260 4834 8306 4846
rect 8054 4444 8064 4628
rect 8116 4444 8126 4628
rect 8164 4458 8170 4664
rect 8204 4458 8210 4664
rect 8260 4628 8266 4834
rect 8300 4628 8306 4834
rect 8342 4664 8352 4848
rect 8404 4664 8414 4848
rect 8452 4834 8498 4846
rect 8164 4446 8210 4458
rect 8246 4444 8256 4628
rect 8308 4444 8318 4628
rect 8356 4458 8362 4664
rect 8396 4458 8402 4664
rect 8452 4628 8458 4834
rect 8492 4628 8498 4834
rect 8534 4664 8544 4848
rect 8596 4664 8606 4848
rect 8644 4834 8690 4846
rect 8356 4446 8402 4458
rect 8438 4444 8448 4628
rect 8500 4444 8510 4628
rect 8548 4458 8554 4664
rect 8588 4458 8594 4664
rect 8644 4628 8650 4834
rect 8684 4628 8690 4834
rect 8726 4664 8736 4848
rect 8788 4664 8798 4848
rect 8836 4834 8882 4846
rect 8548 4446 8594 4458
rect 8630 4444 8640 4628
rect 8692 4444 8702 4628
rect 8740 4458 8746 4664
rect 8780 4458 8786 4664
rect 8836 4628 8842 4834
rect 8876 4628 8882 4834
rect 8918 4664 8928 4848
rect 8980 4664 8990 4848
rect 9028 4834 9074 4846
rect 8740 4446 8786 4458
rect 8822 4444 8832 4628
rect 8884 4444 8894 4628
rect 8932 4458 8938 4664
rect 8972 4458 8978 4664
rect 9028 4628 9034 4834
rect 9068 4628 9074 4834
rect 9110 4664 9120 4848
rect 9172 4664 9182 4848
rect 9220 4834 9266 4846
rect 8932 4446 8978 4458
rect 9014 4444 9024 4628
rect 9076 4444 9086 4628
rect 9124 4458 9130 4664
rect 9164 4458 9170 4664
rect 9220 4628 9226 4834
rect 9260 4628 9266 4834
rect 9302 4664 9312 4848
rect 9364 4664 9374 4848
rect 9412 4834 9458 4846
rect 9124 4446 9170 4458
rect 9206 4444 9216 4628
rect 9268 4444 9278 4628
rect 9316 4458 9322 4664
rect 9356 4458 9362 4664
rect 9412 4628 9418 4834
rect 9452 4628 9458 4834
rect 9494 4664 9504 4848
rect 9556 4664 9566 4848
rect 9604 4834 9650 4846
rect 9316 4446 9362 4458
rect 9398 4444 9408 4628
rect 9460 4444 9470 4628
rect 9508 4458 9514 4664
rect 9548 4458 9554 4664
rect 9604 4628 9610 4834
rect 9644 4628 9650 4834
rect 9686 4664 9696 4848
rect 9748 4664 9758 4848
rect 9796 4834 9842 4846
rect 9508 4446 9554 4458
rect 9590 4444 9600 4628
rect 9652 4444 9662 4628
rect 9700 4458 9706 4664
rect 9740 4458 9746 4664
rect 9796 4628 9802 4834
rect 9836 4628 9842 4834
rect 9878 4664 9888 4848
rect 9940 4664 9950 4848
rect 9988 4834 10034 4846
rect 9700 4446 9746 4458
rect 9782 4444 9792 4628
rect 9844 4444 9854 4628
rect 9892 4458 9898 4664
rect 9932 4458 9938 4664
rect 9988 4628 9994 4834
rect 10028 4628 10034 4834
rect 10070 4664 10080 4848
rect 10132 4664 10142 4848
rect 10180 4834 10226 4846
rect 9892 4446 9938 4458
rect 9974 4444 9984 4628
rect 10036 4444 10046 4628
rect 10084 4458 10090 4664
rect 10124 4458 10130 4664
rect 10180 4628 10186 4834
rect 10220 4628 10226 4834
rect 10262 4664 10272 4848
rect 10324 4664 10334 4848
rect 10372 4834 10418 4846
rect 10084 4446 10130 4458
rect 10166 4444 10176 4628
rect 10228 4444 10238 4628
rect 10276 4458 10282 4664
rect 10316 4458 10322 4664
rect 10372 4628 10378 4834
rect 10412 4628 10418 4834
rect 10454 4664 10464 4848
rect 10516 4664 10526 4848
rect 10564 4834 10610 4846
rect 10276 4446 10322 4458
rect 10358 4444 10368 4628
rect 10420 4444 10430 4628
rect 10468 4458 10474 4664
rect 10508 4458 10514 4664
rect 10564 4628 10570 4834
rect 10604 4628 10610 4834
rect 10646 4664 10656 4848
rect 10708 4664 10718 4848
rect 10756 4834 10802 4846
rect 10468 4446 10514 4458
rect 10550 4444 10560 4628
rect 10612 4444 10622 4628
rect 10660 4458 10666 4664
rect 10700 4458 10706 4664
rect 10756 4628 10762 4834
rect 10796 4628 10802 4834
rect 10838 4664 10848 4848
rect 10900 4664 10910 4848
rect 10948 4834 10994 4846
rect 10660 4446 10706 4458
rect 10742 4444 10752 4628
rect 10804 4444 10814 4628
rect 10852 4458 10858 4664
rect 10892 4458 10898 4664
rect 10948 4628 10954 4834
rect 10988 4628 10994 4834
rect 12048 4834 12094 4846
rect 12048 4628 12054 4834
rect 12088 4628 12094 4834
rect 12130 4664 12140 4848
rect 12192 4664 12202 4848
rect 12240 4834 12286 4846
rect 10852 4446 10898 4458
rect 10934 4444 10944 4628
rect 10996 4444 11006 4628
rect 12034 4444 12044 4628
rect 12096 4444 12106 4628
rect 12144 4458 12150 4664
rect 12184 4458 12190 4664
rect 12240 4628 12246 4834
rect 12280 4628 12286 4834
rect 12322 4664 12332 4848
rect 12384 4664 12394 4848
rect 12432 4834 12478 4846
rect 12144 4446 12190 4458
rect 12226 4444 12236 4628
rect 12288 4444 12298 4628
rect 12336 4458 12342 4664
rect 12376 4458 12382 4664
rect 12432 4628 12438 4834
rect 12472 4628 12478 4834
rect 12514 4664 12524 4848
rect 12576 4664 12586 4848
rect 12624 4834 12670 4846
rect 12336 4446 12382 4458
rect 12418 4444 12428 4628
rect 12480 4444 12490 4628
rect 12528 4458 12534 4664
rect 12568 4458 12574 4664
rect 12624 4628 12630 4834
rect 12664 4628 12670 4834
rect 12706 4664 12716 4848
rect 12768 4664 12778 4848
rect 12816 4834 12862 4846
rect 12528 4446 12574 4458
rect 12610 4444 12620 4628
rect 12672 4444 12682 4628
rect 12720 4458 12726 4664
rect 12760 4458 12766 4664
rect 12816 4628 12822 4834
rect 12856 4628 12862 4834
rect 12898 4664 12908 4848
rect 12960 4664 12970 4848
rect 13008 4834 13054 4846
rect 12720 4446 12766 4458
rect 12802 4444 12812 4628
rect 12864 4444 12874 4628
rect 12912 4458 12918 4664
rect 12952 4458 12958 4664
rect 13008 4628 13014 4834
rect 13048 4628 13054 4834
rect 13090 4664 13100 4848
rect 13152 4664 13162 4848
rect 13200 4834 13246 4846
rect 12912 4446 12958 4458
rect 12994 4444 13004 4628
rect 13056 4444 13066 4628
rect 13104 4458 13110 4664
rect 13144 4458 13150 4664
rect 13200 4628 13206 4834
rect 13240 4628 13246 4834
rect 13282 4664 13292 4848
rect 13344 4664 13354 4848
rect 13392 4834 13438 4846
rect 13104 4446 13150 4458
rect 13186 4444 13196 4628
rect 13248 4444 13258 4628
rect 13296 4458 13302 4664
rect 13336 4458 13342 4664
rect 13392 4628 13398 4834
rect 13432 4628 13438 4834
rect 13474 4664 13484 4848
rect 13536 4664 13546 4848
rect 13584 4834 13630 4846
rect 13296 4446 13342 4458
rect 13378 4444 13388 4628
rect 13440 4444 13450 4628
rect 13488 4458 13494 4664
rect 13528 4458 13534 4664
rect 13584 4628 13590 4834
rect 13624 4628 13630 4834
rect 13666 4664 13676 4848
rect 13728 4664 13738 4848
rect 13776 4834 13822 4846
rect 13488 4446 13534 4458
rect 13570 4444 13580 4628
rect 13632 4444 13642 4628
rect 13680 4458 13686 4664
rect 13720 4458 13726 4664
rect 13776 4628 13782 4834
rect 13816 4628 13822 4834
rect 13858 4664 13868 4848
rect 13920 4664 13930 4848
rect 13968 4834 14014 4846
rect 13680 4446 13726 4458
rect 13762 4444 13772 4628
rect 13824 4444 13834 4628
rect 13872 4458 13878 4664
rect 13912 4458 13918 4664
rect 13968 4628 13974 4834
rect 14008 4628 14014 4834
rect 14050 4664 14060 4848
rect 14112 4664 14122 4848
rect 14160 4834 14206 4846
rect 13872 4446 13918 4458
rect 13954 4444 13964 4628
rect 14016 4444 14026 4628
rect 14064 4458 14070 4664
rect 14104 4458 14110 4664
rect 14160 4628 14166 4834
rect 14200 4628 14206 4834
rect 14242 4664 14252 4848
rect 14304 4664 14314 4848
rect 14352 4834 14398 4846
rect 14064 4446 14110 4458
rect 14146 4444 14156 4628
rect 14208 4444 14218 4628
rect 14256 4458 14262 4664
rect 14296 4458 14302 4664
rect 14352 4628 14358 4834
rect 14392 4628 14398 4834
rect 14434 4664 14444 4848
rect 14496 4664 14506 4848
rect 14544 4834 14590 4846
rect 14256 4446 14302 4458
rect 14338 4444 14348 4628
rect 14400 4444 14410 4628
rect 14448 4458 14454 4664
rect 14488 4458 14494 4664
rect 14544 4628 14550 4834
rect 14584 4628 14590 4834
rect 14626 4664 14636 4848
rect 14688 4664 14698 4848
rect 14736 4834 14782 4846
rect 14448 4446 14494 4458
rect 14530 4444 14540 4628
rect 14592 4444 14602 4628
rect 14640 4458 14646 4664
rect 14680 4458 14686 4664
rect 14736 4628 14742 4834
rect 14776 4628 14782 4834
rect 14818 4664 14828 4848
rect 14880 4664 14890 4848
rect 14928 4834 14974 4846
rect 14640 4446 14686 4458
rect 14722 4444 14732 4628
rect 14784 4444 14794 4628
rect 14832 4458 14838 4664
rect 14872 4458 14878 4664
rect 14928 4628 14934 4834
rect 14968 4628 14974 4834
rect 14832 4446 14878 4458
rect 14914 4444 14924 4628
rect 14976 4444 14986 4628
rect 15088 4416 15536 4876
rect 15688 4834 15734 4846
rect 15688 4628 15694 4834
rect 15728 4628 15734 4834
rect 15770 4664 15780 4848
rect 15832 4664 15842 4848
rect 15880 4834 15926 4846
rect 15674 4444 15684 4628
rect 15736 4444 15746 4628
rect 15784 4458 15790 4664
rect 15824 4458 15830 4664
rect 15880 4628 15886 4834
rect 15920 4628 15926 4834
rect 15962 4664 15972 4848
rect 16024 4664 16034 4848
rect 16072 4834 16118 4846
rect 15784 4446 15830 4458
rect 15866 4444 15876 4628
rect 15928 4444 15938 4628
rect 15976 4458 15982 4664
rect 16016 4458 16022 4664
rect 16072 4628 16078 4834
rect 16112 4628 16118 4834
rect 16154 4664 16164 4848
rect 16216 4664 16226 4848
rect 16264 4834 16310 4846
rect 15976 4446 16022 4458
rect 16058 4444 16068 4628
rect 16120 4444 16130 4628
rect 16168 4458 16174 4664
rect 16208 4458 16214 4664
rect 16264 4628 16270 4834
rect 16304 4628 16310 4834
rect 16346 4664 16356 4848
rect 16408 4664 16418 4848
rect 16456 4834 16502 4846
rect 16168 4446 16214 4458
rect 16250 4444 16260 4628
rect 16312 4444 16322 4628
rect 16360 4458 16366 4664
rect 16400 4458 16406 4664
rect 16456 4628 16462 4834
rect 16496 4628 16502 4834
rect 16538 4664 16548 4848
rect 16600 4664 16610 4848
rect 16648 4834 16694 4846
rect 16360 4446 16406 4458
rect 16442 4444 16452 4628
rect 16504 4444 16514 4628
rect 16552 4458 16558 4664
rect 16592 4458 16598 4664
rect 16648 4628 16654 4834
rect 16688 4628 16694 4834
rect 16730 4664 16740 4848
rect 16792 4664 16802 4848
rect 16840 4834 16886 4846
rect 16552 4446 16598 4458
rect 16634 4444 16644 4628
rect 16696 4444 16706 4628
rect 16744 4458 16750 4664
rect 16784 4458 16790 4664
rect 16840 4628 16846 4834
rect 16880 4628 16886 4834
rect 16922 4664 16932 4848
rect 16984 4664 16994 4848
rect 17032 4834 17078 4846
rect 16744 4446 16790 4458
rect 16826 4444 16836 4628
rect 16888 4444 16898 4628
rect 16936 4458 16942 4664
rect 16976 4458 16982 4664
rect 17032 4628 17038 4834
rect 17072 4628 17078 4834
rect 17114 4664 17124 4848
rect 17176 4664 17186 4848
rect 17224 4834 17270 4846
rect 16936 4446 16982 4458
rect 17018 4444 17028 4628
rect 17080 4444 17090 4628
rect 17128 4458 17134 4664
rect 17168 4458 17174 4664
rect 17224 4628 17230 4834
rect 17264 4628 17270 4834
rect 17306 4664 17316 4848
rect 17368 4664 17378 4848
rect 17416 4834 17462 4846
rect 17128 4446 17174 4458
rect 17210 4444 17220 4628
rect 17272 4444 17282 4628
rect 17320 4458 17326 4664
rect 17360 4458 17366 4664
rect 17416 4628 17422 4834
rect 17456 4628 17462 4834
rect 17498 4664 17508 4848
rect 17560 4664 17570 4848
rect 17608 4834 17654 4846
rect 17320 4446 17366 4458
rect 17402 4444 17412 4628
rect 17464 4444 17474 4628
rect 17512 4458 17518 4664
rect 17552 4458 17558 4664
rect 17608 4628 17614 4834
rect 17648 4628 17654 4834
rect 17690 4664 17700 4848
rect 17752 4664 17762 4848
rect 17800 4834 17846 4846
rect 17512 4446 17558 4458
rect 17594 4444 17604 4628
rect 17656 4444 17666 4628
rect 17704 4458 17710 4664
rect 17744 4458 17750 4664
rect 17800 4628 17806 4834
rect 17840 4628 17846 4834
rect 17882 4664 17892 4848
rect 17944 4664 17954 4848
rect 17992 4834 18038 4846
rect 17704 4446 17750 4458
rect 17786 4444 17796 4628
rect 17848 4444 17858 4628
rect 17896 4458 17902 4664
rect 17936 4458 17942 4664
rect 17992 4628 17998 4834
rect 18032 4628 18038 4834
rect 18074 4664 18084 4848
rect 18136 4664 18146 4848
rect 18184 4834 18230 4846
rect 17896 4446 17942 4458
rect 17978 4444 17988 4628
rect 18040 4444 18050 4628
rect 18088 4458 18094 4664
rect 18128 4458 18134 4664
rect 18184 4628 18190 4834
rect 18224 4628 18230 4834
rect 18266 4664 18276 4848
rect 18328 4664 18338 4848
rect 18376 4834 18422 4846
rect 18088 4446 18134 4458
rect 18170 4444 18180 4628
rect 18232 4444 18242 4628
rect 18280 4458 18286 4664
rect 18320 4458 18326 4664
rect 18376 4628 18382 4834
rect 18416 4628 18422 4834
rect 18458 4664 18468 4848
rect 18520 4664 18530 4848
rect 18568 4834 18614 4846
rect 18280 4446 18326 4458
rect 18362 4444 18372 4628
rect 18424 4444 18434 4628
rect 18472 4458 18478 4664
rect 18512 4458 18518 4664
rect 18568 4628 18574 4834
rect 18608 4628 18614 4834
rect 18472 4446 18518 4458
rect 18554 4444 18564 4628
rect 18616 4444 18626 4628
rect 4160 4408 10864 4416
rect -1436 4385 360 4404
rect -1436 3988 -1418 4385
rect -1168 3988 -1040 4385
rect -790 4372 -662 4385
rect -412 4372 -284 4385
rect -790 3988 -662 3996
rect -412 3988 -284 3996
rect -34 3988 94 4385
rect 344 3988 360 4385
rect -1436 3972 360 3988
rect 1364 4400 3160 4404
rect 4160 4400 4482 4408
rect 1364 4385 4482 4400
rect 1364 3988 1382 4385
rect 1632 3988 1760 4385
rect 2010 4372 2138 4385
rect 2388 4372 2516 4385
rect 2010 3988 2138 3996
rect 2388 3988 2516 3996
rect 2766 3988 2894 4385
rect 3144 4374 4482 4385
rect 4516 4374 4674 4408
rect 4708 4374 4866 4408
rect 4900 4374 5058 4408
rect 5092 4374 5250 4408
rect 5284 4374 5442 4408
rect 5476 4374 5634 4408
rect 5668 4374 5826 4408
rect 5860 4374 6018 4408
rect 6052 4374 6210 4408
rect 6244 4374 6402 4408
rect 6436 4374 6594 4408
rect 6628 4374 6786 4408
rect 6820 4374 6978 4408
rect 7012 4374 7170 4408
rect 7204 4374 8122 4408
rect 8156 4374 8314 4408
rect 8348 4374 8506 4408
rect 8540 4374 8698 4408
rect 8732 4374 8890 4408
rect 8924 4374 9082 4408
rect 9116 4374 9274 4408
rect 9308 4374 9466 4408
rect 9500 4374 9658 4408
rect 9692 4374 9850 4408
rect 9884 4374 10042 4408
rect 10076 4374 10234 4408
rect 10268 4374 10426 4408
rect 10460 4374 10618 4408
rect 10652 4374 10810 4408
rect 10844 4374 10864 4408
rect 3144 4300 10864 4374
rect 3144 4266 4482 4300
rect 4516 4266 4674 4300
rect 4708 4266 4866 4300
rect 4900 4266 5058 4300
rect 5092 4266 5250 4300
rect 5284 4266 5442 4300
rect 5476 4266 5634 4300
rect 5668 4266 5826 4300
rect 5860 4266 6018 4300
rect 6052 4266 6210 4300
rect 6244 4266 6402 4300
rect 6436 4266 6594 4300
rect 6628 4266 6786 4300
rect 6820 4266 6978 4300
rect 7012 4266 7170 4300
rect 7204 4266 8122 4300
rect 8156 4266 8314 4300
rect 8348 4266 8506 4300
rect 8540 4266 8698 4300
rect 8732 4266 8890 4300
rect 8924 4266 9082 4300
rect 9116 4266 9274 4300
rect 9308 4266 9466 4300
rect 9500 4266 9658 4300
rect 9692 4266 9850 4300
rect 9884 4266 10042 4300
rect 10076 4266 10234 4300
rect 10268 4266 10426 4300
rect 10460 4266 10618 4300
rect 10652 4266 10810 4300
rect 10844 4266 10864 4300
rect 3144 4260 10864 4266
rect 12084 4408 18484 4416
rect 12084 4374 12102 4408
rect 12136 4374 12294 4408
rect 12328 4374 12486 4408
rect 12520 4374 12678 4408
rect 12712 4374 12870 4408
rect 12904 4374 13062 4408
rect 13096 4374 13254 4408
rect 13288 4374 13446 4408
rect 13480 4374 13638 4408
rect 13672 4374 13830 4408
rect 13864 4374 14022 4408
rect 14056 4374 14214 4408
rect 14248 4374 14406 4408
rect 14440 4374 14598 4408
rect 14632 4374 14790 4408
rect 14824 4374 15742 4408
rect 15776 4374 15934 4408
rect 15968 4374 16126 4408
rect 16160 4374 16318 4408
rect 16352 4374 16510 4408
rect 16544 4374 16702 4408
rect 16736 4374 16894 4408
rect 16928 4374 17086 4408
rect 17120 4374 17278 4408
rect 17312 4374 17470 4408
rect 17504 4374 17662 4408
rect 17696 4374 17854 4408
rect 17888 4374 18046 4408
rect 18080 4374 18238 4408
rect 18272 4374 18430 4408
rect 18464 4374 18484 4408
rect 12084 4300 18484 4374
rect 12084 4266 12102 4300
rect 12136 4266 12294 4300
rect 12328 4266 12486 4300
rect 12520 4266 12678 4300
rect 12712 4266 12870 4300
rect 12904 4266 13062 4300
rect 13096 4266 13254 4300
rect 13288 4266 13446 4300
rect 13480 4266 13638 4300
rect 13672 4266 13830 4300
rect 13864 4266 14022 4300
rect 14056 4266 14214 4300
rect 14248 4266 14406 4300
rect 14440 4266 14598 4300
rect 14632 4266 14790 4300
rect 14824 4266 15742 4300
rect 15776 4266 15934 4300
rect 15968 4266 16126 4300
rect 16160 4266 16318 4300
rect 16352 4266 16510 4300
rect 16544 4266 16702 4300
rect 16736 4266 16894 4300
rect 16928 4266 17086 4300
rect 17120 4266 17278 4300
rect 17312 4266 17470 4300
rect 17504 4266 17662 4300
rect 17696 4266 17854 4300
rect 17888 4266 18046 4300
rect 18080 4266 18238 4300
rect 18272 4266 18430 4300
rect 18464 4266 18484 4300
rect 12084 4260 18484 4266
rect 3144 3988 4324 4260
rect 4428 4216 4474 4228
rect 4428 4012 4434 4216
rect 4468 4012 4474 4216
rect 4510 4048 4520 4232
rect 4572 4048 4582 4232
rect 4620 4216 4666 4228
rect 1364 3972 4324 3988
rect 2960 3960 4324 3972
rect 4160 3796 4324 3960
rect 4414 3828 4424 4012
rect 4476 3828 4486 4012
rect 4524 3840 4530 4048
rect 4564 3840 4570 4048
rect 4620 4012 4626 4216
rect 4660 4012 4666 4216
rect 4702 4048 4712 4232
rect 4764 4048 4774 4232
rect 4812 4216 4858 4228
rect 4524 3828 4570 3840
rect 4606 3828 4616 4012
rect 4668 3828 4678 4012
rect 4716 3840 4722 4048
rect 4756 3840 4762 4048
rect 4812 4012 4818 4216
rect 4852 4012 4858 4216
rect 4894 4048 4904 4232
rect 4956 4048 4966 4232
rect 5004 4216 5050 4228
rect 4716 3828 4762 3840
rect 4798 3828 4808 4012
rect 4860 3828 4870 4012
rect 4908 3840 4914 4048
rect 4948 3840 4954 4048
rect 5004 4012 5010 4216
rect 5044 4012 5050 4216
rect 5086 4048 5096 4232
rect 5148 4048 5158 4232
rect 5196 4216 5242 4228
rect 4908 3828 4954 3840
rect 4990 3828 5000 4012
rect 5052 3828 5062 4012
rect 5100 3840 5106 4048
rect 5140 3840 5146 4048
rect 5196 4012 5202 4216
rect 5236 4012 5242 4216
rect 5278 4048 5288 4232
rect 5340 4048 5350 4232
rect 5388 4216 5434 4228
rect 5100 3828 5146 3840
rect 5182 3828 5192 4012
rect 5244 3828 5254 4012
rect 5292 3840 5298 4048
rect 5332 3840 5338 4048
rect 5388 4012 5394 4216
rect 5428 4012 5434 4216
rect 5470 4048 5480 4232
rect 5532 4048 5542 4232
rect 5580 4216 5626 4228
rect 5292 3828 5338 3840
rect 5374 3828 5384 4012
rect 5436 3828 5446 4012
rect 5484 3840 5490 4048
rect 5524 3840 5530 4048
rect 5580 4012 5586 4216
rect 5620 4012 5626 4216
rect 5662 4048 5672 4232
rect 5724 4048 5734 4232
rect 5772 4216 5818 4228
rect 5484 3828 5530 3840
rect 5566 3828 5576 4012
rect 5628 3828 5638 4012
rect 5676 3840 5682 4048
rect 5716 3840 5722 4048
rect 5772 4012 5778 4216
rect 5812 4012 5818 4216
rect 5854 4048 5864 4232
rect 5916 4048 5926 4232
rect 5964 4216 6010 4228
rect 5676 3828 5722 3840
rect 5758 3828 5768 4012
rect 5820 3828 5830 4012
rect 5868 3840 5874 4048
rect 5908 3840 5914 4048
rect 5964 4012 5970 4216
rect 6004 4012 6010 4216
rect 6046 4048 6056 4232
rect 6108 4048 6118 4232
rect 6156 4216 6202 4228
rect 5868 3828 5914 3840
rect 5950 3828 5960 4012
rect 6012 3828 6022 4012
rect 6060 3840 6066 4048
rect 6100 3840 6106 4048
rect 6156 4012 6162 4216
rect 6196 4012 6202 4216
rect 6238 4048 6248 4232
rect 6300 4048 6310 4232
rect 6348 4216 6394 4228
rect 6060 3828 6106 3840
rect 6142 3828 6152 4012
rect 6204 3828 6214 4012
rect 6252 3840 6258 4048
rect 6292 3840 6298 4048
rect 6348 4012 6354 4216
rect 6388 4012 6394 4216
rect 6430 4048 6440 4232
rect 6492 4048 6502 4232
rect 6540 4216 6586 4228
rect 6252 3828 6298 3840
rect 6334 3828 6344 4012
rect 6396 3828 6406 4012
rect 6444 3840 6450 4048
rect 6484 3840 6490 4048
rect 6540 4012 6546 4216
rect 6580 4012 6586 4216
rect 6622 4048 6632 4232
rect 6684 4048 6694 4232
rect 6732 4216 6778 4228
rect 6444 3828 6490 3840
rect 6526 3828 6536 4012
rect 6588 3828 6598 4012
rect 6636 3840 6642 4048
rect 6676 3840 6682 4048
rect 6732 4012 6738 4216
rect 6772 4012 6778 4216
rect 6814 4048 6824 4232
rect 6876 4048 6886 4232
rect 6924 4216 6970 4228
rect 6636 3828 6682 3840
rect 6718 3828 6728 4012
rect 6780 3828 6790 4012
rect 6828 3840 6834 4048
rect 6868 3840 6874 4048
rect 6924 4012 6930 4216
rect 6964 4012 6970 4216
rect 7006 4048 7016 4232
rect 7068 4048 7078 4232
rect 7116 4216 7162 4228
rect 6828 3828 6874 3840
rect 6910 3828 6920 4012
rect 6972 3828 6982 4012
rect 7020 3840 7026 4048
rect 7060 3840 7066 4048
rect 7116 4012 7122 4216
rect 7156 4012 7162 4216
rect 7198 4048 7208 4232
rect 7260 4048 7270 4232
rect 7308 4216 7354 4228
rect 7020 3828 7066 3840
rect 7102 3828 7112 4012
rect 7164 3828 7174 4012
rect 7212 3840 7218 4048
rect 7252 3840 7258 4048
rect 7308 4012 7314 4216
rect 7348 4012 7354 4216
rect 7212 3828 7258 3840
rect 7294 3828 7304 4012
rect 7356 3828 7366 4012
rect 7468 3796 7916 4260
rect 8068 4216 8114 4228
rect 8068 4012 8074 4216
rect 8108 4012 8114 4216
rect 8150 4048 8160 4232
rect 8212 4048 8222 4232
rect 8260 4216 8306 4228
rect 8054 3828 8064 4012
rect 8116 3828 8126 4012
rect 8164 3840 8170 4048
rect 8204 3840 8210 4048
rect 8260 4012 8266 4216
rect 8300 4012 8306 4216
rect 8342 4048 8352 4232
rect 8404 4048 8414 4232
rect 8452 4216 8498 4228
rect 8164 3828 8210 3840
rect 8246 3828 8256 4012
rect 8308 3828 8318 4012
rect 8356 3840 8362 4048
rect 8396 3840 8402 4048
rect 8452 4012 8458 4216
rect 8492 4012 8498 4216
rect 8534 4048 8544 4232
rect 8596 4048 8606 4232
rect 8644 4216 8690 4228
rect 8356 3828 8402 3840
rect 8438 3828 8448 4012
rect 8500 3828 8510 4012
rect 8548 3840 8554 4048
rect 8588 3840 8594 4048
rect 8644 4012 8650 4216
rect 8684 4012 8690 4216
rect 8726 4048 8736 4232
rect 8788 4048 8798 4232
rect 8836 4216 8882 4228
rect 8548 3828 8594 3840
rect 8630 3828 8640 4012
rect 8692 3828 8702 4012
rect 8740 3840 8746 4048
rect 8780 3840 8786 4048
rect 8836 4012 8842 4216
rect 8876 4012 8882 4216
rect 8918 4048 8928 4232
rect 8980 4048 8990 4232
rect 9028 4216 9074 4228
rect 8740 3828 8786 3840
rect 8822 3828 8832 4012
rect 8884 3828 8894 4012
rect 8932 3840 8938 4048
rect 8972 3840 8978 4048
rect 9028 4012 9034 4216
rect 9068 4012 9074 4216
rect 9110 4048 9120 4232
rect 9172 4048 9182 4232
rect 9220 4216 9266 4228
rect 8932 3828 8978 3840
rect 9014 3828 9024 4012
rect 9076 3828 9086 4012
rect 9124 3840 9130 4048
rect 9164 3840 9170 4048
rect 9220 4012 9226 4216
rect 9260 4012 9266 4216
rect 9302 4048 9312 4232
rect 9364 4048 9374 4232
rect 9412 4216 9458 4228
rect 9124 3828 9170 3840
rect 9206 3828 9216 4012
rect 9268 3828 9278 4012
rect 9316 3840 9322 4048
rect 9356 3840 9362 4048
rect 9412 4012 9418 4216
rect 9452 4012 9458 4216
rect 9494 4048 9504 4232
rect 9556 4048 9566 4232
rect 9604 4216 9650 4228
rect 9316 3828 9362 3840
rect 9398 3828 9408 4012
rect 9460 3828 9470 4012
rect 9508 3840 9514 4048
rect 9548 3840 9554 4048
rect 9604 4012 9610 4216
rect 9644 4012 9650 4216
rect 9686 4048 9696 4232
rect 9748 4048 9758 4232
rect 9796 4216 9842 4228
rect 9508 3828 9554 3840
rect 9590 3828 9600 4012
rect 9652 3828 9662 4012
rect 9700 3840 9706 4048
rect 9740 3840 9746 4048
rect 9796 4012 9802 4216
rect 9836 4012 9842 4216
rect 9878 4048 9888 4232
rect 9940 4048 9950 4232
rect 9988 4216 10034 4228
rect 9700 3828 9746 3840
rect 9782 3828 9792 4012
rect 9844 3828 9854 4012
rect 9892 3840 9898 4048
rect 9932 3840 9938 4048
rect 9988 4012 9994 4216
rect 10028 4012 10034 4216
rect 10070 4048 10080 4232
rect 10132 4048 10142 4232
rect 10180 4216 10226 4228
rect 9892 3828 9938 3840
rect 9974 3828 9984 4012
rect 10036 3828 10046 4012
rect 10084 3840 10090 4048
rect 10124 3840 10130 4048
rect 10180 4012 10186 4216
rect 10220 4012 10226 4216
rect 10262 4048 10272 4232
rect 10324 4048 10334 4232
rect 10372 4216 10418 4228
rect 10084 3828 10130 3840
rect 10166 3828 10176 4012
rect 10228 3828 10238 4012
rect 10276 3840 10282 4048
rect 10316 3840 10322 4048
rect 10372 4012 10378 4216
rect 10412 4012 10418 4216
rect 10454 4048 10464 4232
rect 10516 4048 10526 4232
rect 10564 4216 10610 4228
rect 10276 3828 10322 3840
rect 10358 3828 10368 4012
rect 10420 3828 10430 4012
rect 10468 3840 10474 4048
rect 10508 3840 10514 4048
rect 10564 4012 10570 4216
rect 10604 4012 10610 4216
rect 10646 4048 10656 4232
rect 10708 4048 10718 4232
rect 10756 4216 10802 4228
rect 10468 3828 10514 3840
rect 10550 3828 10560 4012
rect 10612 3828 10622 4012
rect 10660 3840 10666 4048
rect 10700 3840 10706 4048
rect 10756 4012 10762 4216
rect 10796 4012 10802 4216
rect 10838 4048 10848 4232
rect 10900 4048 10910 4232
rect 10948 4216 10994 4228
rect 10660 3828 10706 3840
rect 10742 3828 10752 4012
rect 10804 3828 10814 4012
rect 10852 3840 10858 4048
rect 10892 3840 10898 4048
rect 10948 4012 10954 4216
rect 10988 4012 10994 4216
rect 12048 4216 12094 4228
rect 12048 4012 12054 4216
rect 12088 4012 12094 4216
rect 12130 4048 12140 4232
rect 12192 4048 12202 4232
rect 12240 4216 12286 4228
rect 10852 3828 10898 3840
rect 10934 3828 10944 4012
rect 10996 3828 11006 4012
rect 12034 3828 12044 4012
rect 12096 3828 12106 4012
rect 12144 3840 12150 4048
rect 12184 3840 12190 4048
rect 12240 4012 12246 4216
rect 12280 4012 12286 4216
rect 12322 4048 12332 4232
rect 12384 4048 12394 4232
rect 12432 4216 12478 4228
rect 12144 3828 12190 3840
rect 12226 3828 12236 4012
rect 12288 3828 12298 4012
rect 12336 3840 12342 4048
rect 12376 3840 12382 4048
rect 12432 4012 12438 4216
rect 12472 4012 12478 4216
rect 12514 4048 12524 4232
rect 12576 4048 12586 4232
rect 12624 4216 12670 4228
rect 12336 3828 12382 3840
rect 12418 3828 12428 4012
rect 12480 3828 12490 4012
rect 12528 3840 12534 4048
rect 12568 3840 12574 4048
rect 12624 4012 12630 4216
rect 12664 4012 12670 4216
rect 12706 4048 12716 4232
rect 12768 4048 12778 4232
rect 12816 4216 12862 4228
rect 12528 3828 12574 3840
rect 12610 3828 12620 4012
rect 12672 3828 12682 4012
rect 12720 3840 12726 4048
rect 12760 3840 12766 4048
rect 12816 4012 12822 4216
rect 12856 4012 12862 4216
rect 12898 4048 12908 4232
rect 12960 4048 12970 4232
rect 13008 4216 13054 4228
rect 12720 3828 12766 3840
rect 12802 3828 12812 4012
rect 12864 3828 12874 4012
rect 12912 3840 12918 4048
rect 12952 3840 12958 4048
rect 13008 4012 13014 4216
rect 13048 4012 13054 4216
rect 13090 4048 13100 4232
rect 13152 4048 13162 4232
rect 13200 4216 13246 4228
rect 12912 3828 12958 3840
rect 12994 3828 13004 4012
rect 13056 3828 13066 4012
rect 13104 3840 13110 4048
rect 13144 3840 13150 4048
rect 13200 4012 13206 4216
rect 13240 4012 13246 4216
rect 13282 4048 13292 4232
rect 13344 4048 13354 4232
rect 13392 4216 13438 4228
rect 13104 3828 13150 3840
rect 13186 3828 13196 4012
rect 13248 3828 13258 4012
rect 13296 3840 13302 4048
rect 13336 3840 13342 4048
rect 13392 4012 13398 4216
rect 13432 4012 13438 4216
rect 13474 4048 13484 4232
rect 13536 4048 13546 4232
rect 13584 4216 13630 4228
rect 13296 3828 13342 3840
rect 13378 3828 13388 4012
rect 13440 3828 13450 4012
rect 13488 3840 13494 4048
rect 13528 3840 13534 4048
rect 13584 4012 13590 4216
rect 13624 4012 13630 4216
rect 13666 4048 13676 4232
rect 13728 4048 13738 4232
rect 13776 4216 13822 4228
rect 13488 3828 13534 3840
rect 13570 3828 13580 4012
rect 13632 3828 13642 4012
rect 13680 3840 13686 4048
rect 13720 3840 13726 4048
rect 13776 4012 13782 4216
rect 13816 4012 13822 4216
rect 13858 4048 13868 4232
rect 13920 4048 13930 4232
rect 13968 4216 14014 4228
rect 13680 3828 13726 3840
rect 13762 3828 13772 4012
rect 13824 3828 13834 4012
rect 13872 3840 13878 4048
rect 13912 3840 13918 4048
rect 13968 4012 13974 4216
rect 14008 4012 14014 4216
rect 14050 4048 14060 4232
rect 14112 4048 14122 4232
rect 14160 4216 14206 4228
rect 13872 3828 13918 3840
rect 13954 3828 13964 4012
rect 14016 3828 14026 4012
rect 14064 3840 14070 4048
rect 14104 3840 14110 4048
rect 14160 4012 14166 4216
rect 14200 4012 14206 4216
rect 14242 4048 14252 4232
rect 14304 4048 14314 4232
rect 14352 4216 14398 4228
rect 14064 3828 14110 3840
rect 14146 3828 14156 4012
rect 14208 3828 14218 4012
rect 14256 3840 14262 4048
rect 14296 3840 14302 4048
rect 14352 4012 14358 4216
rect 14392 4012 14398 4216
rect 14434 4048 14444 4232
rect 14496 4048 14506 4232
rect 14544 4216 14590 4228
rect 14256 3828 14302 3840
rect 14338 3828 14348 4012
rect 14400 3828 14410 4012
rect 14448 3840 14454 4048
rect 14488 3840 14494 4048
rect 14544 4012 14550 4216
rect 14584 4012 14590 4216
rect 14626 4048 14636 4232
rect 14688 4048 14698 4232
rect 14736 4216 14782 4228
rect 14448 3828 14494 3840
rect 14530 3828 14540 4012
rect 14592 3828 14602 4012
rect 14640 3840 14646 4048
rect 14680 3840 14686 4048
rect 14736 4012 14742 4216
rect 14776 4012 14782 4216
rect 14818 4048 14828 4232
rect 14880 4048 14890 4232
rect 14928 4216 14974 4228
rect 14640 3828 14686 3840
rect 14722 3828 14732 4012
rect 14784 3828 14794 4012
rect 14832 3840 14838 4048
rect 14872 3840 14878 4048
rect 14928 4012 14934 4216
rect 14968 4012 14974 4216
rect 14832 3828 14878 3840
rect 14914 3828 14924 4012
rect 14976 3828 14986 4012
rect 15088 3796 15536 4260
rect 15688 4216 15734 4228
rect 15688 4012 15694 4216
rect 15728 4012 15734 4216
rect 15770 4048 15780 4232
rect 15832 4048 15842 4232
rect 15880 4216 15926 4228
rect 15674 3828 15684 4012
rect 15736 3828 15746 4012
rect 15784 3840 15790 4048
rect 15824 3840 15830 4048
rect 15880 4012 15886 4216
rect 15920 4012 15926 4216
rect 15962 4048 15972 4232
rect 16024 4048 16034 4232
rect 16072 4216 16118 4228
rect 15784 3828 15830 3840
rect 15866 3828 15876 4012
rect 15928 3828 15938 4012
rect 15976 3840 15982 4048
rect 16016 3840 16022 4048
rect 16072 4012 16078 4216
rect 16112 4012 16118 4216
rect 16154 4048 16164 4232
rect 16216 4048 16226 4232
rect 16264 4216 16310 4228
rect 15976 3828 16022 3840
rect 16058 3828 16068 4012
rect 16120 3828 16130 4012
rect 16168 3840 16174 4048
rect 16208 3840 16214 4048
rect 16264 4012 16270 4216
rect 16304 4012 16310 4216
rect 16346 4048 16356 4232
rect 16408 4048 16418 4232
rect 16456 4216 16502 4228
rect 16168 3828 16214 3840
rect 16250 3828 16260 4012
rect 16312 3828 16322 4012
rect 16360 3840 16366 4048
rect 16400 3840 16406 4048
rect 16456 4012 16462 4216
rect 16496 4012 16502 4216
rect 16538 4048 16548 4232
rect 16600 4048 16610 4232
rect 16648 4216 16694 4228
rect 16360 3828 16406 3840
rect 16442 3828 16452 4012
rect 16504 3828 16514 4012
rect 16552 3840 16558 4048
rect 16592 3840 16598 4048
rect 16648 4012 16654 4216
rect 16688 4012 16694 4216
rect 16730 4048 16740 4232
rect 16792 4048 16802 4232
rect 16840 4216 16886 4228
rect 16552 3828 16598 3840
rect 16634 3828 16644 4012
rect 16696 3828 16706 4012
rect 16744 3840 16750 4048
rect 16784 3840 16790 4048
rect 16840 4012 16846 4216
rect 16880 4012 16886 4216
rect 16922 4048 16932 4232
rect 16984 4048 16994 4232
rect 17032 4216 17078 4228
rect 16744 3828 16790 3840
rect 16826 3828 16836 4012
rect 16888 3828 16898 4012
rect 16936 3840 16942 4048
rect 16976 3840 16982 4048
rect 17032 4012 17038 4216
rect 17072 4012 17078 4216
rect 17114 4048 17124 4232
rect 17176 4048 17186 4232
rect 17224 4216 17270 4228
rect 16936 3828 16982 3840
rect 17018 3828 17028 4012
rect 17080 3828 17090 4012
rect 17128 3840 17134 4048
rect 17168 3840 17174 4048
rect 17224 4012 17230 4216
rect 17264 4012 17270 4216
rect 17306 4048 17316 4232
rect 17368 4048 17378 4232
rect 17416 4216 17462 4228
rect 17128 3828 17174 3840
rect 17210 3828 17220 4012
rect 17272 3828 17282 4012
rect 17320 3840 17326 4048
rect 17360 3840 17366 4048
rect 17416 4012 17422 4216
rect 17456 4012 17462 4216
rect 17498 4048 17508 4232
rect 17560 4048 17570 4232
rect 17608 4216 17654 4228
rect 17320 3828 17366 3840
rect 17402 3828 17412 4012
rect 17464 3828 17474 4012
rect 17512 3840 17518 4048
rect 17552 3840 17558 4048
rect 17608 4012 17614 4216
rect 17648 4012 17654 4216
rect 17690 4048 17700 4232
rect 17752 4048 17762 4232
rect 17800 4216 17846 4228
rect 17512 3828 17558 3840
rect 17594 3828 17604 4012
rect 17656 3828 17666 4012
rect 17704 3840 17710 4048
rect 17744 3840 17750 4048
rect 17800 4012 17806 4216
rect 17840 4012 17846 4216
rect 17882 4048 17892 4232
rect 17944 4048 17954 4232
rect 17992 4216 18038 4228
rect 17704 3828 17750 3840
rect 17786 3828 17796 4012
rect 17848 3828 17858 4012
rect 17896 3840 17902 4048
rect 17936 3840 17942 4048
rect 17992 4012 17998 4216
rect 18032 4012 18038 4216
rect 18074 4048 18084 4232
rect 18136 4048 18146 4232
rect 18184 4216 18230 4228
rect 17896 3828 17942 3840
rect 17978 3828 17988 4012
rect 18040 3828 18050 4012
rect 18088 3840 18094 4048
rect 18128 3840 18134 4048
rect 18184 4012 18190 4216
rect 18224 4012 18230 4216
rect 18266 4048 18276 4232
rect 18328 4048 18338 4232
rect 18376 4216 18422 4228
rect 18088 3828 18134 3840
rect 18170 3828 18180 4012
rect 18232 3828 18242 4012
rect 18280 3840 18286 4048
rect 18320 3840 18326 4048
rect 18376 4012 18382 4216
rect 18416 4012 18422 4216
rect 18458 4048 18468 4232
rect 18520 4048 18530 4232
rect 18568 4216 18614 4228
rect 18280 3828 18326 3840
rect 18362 3828 18372 4012
rect 18424 3828 18434 4012
rect 18472 3840 18478 4048
rect 18512 3840 18518 4048
rect 18568 4012 18574 4216
rect 18608 4012 18614 4216
rect 18472 3828 18518 3840
rect 18554 3828 18564 4012
rect 18616 3828 18626 4012
rect 4160 3790 10972 3796
rect 4160 3756 4578 3790
rect 4612 3756 4770 3790
rect 4804 3756 4962 3790
rect 4996 3756 5154 3790
rect 5188 3756 5346 3790
rect 5380 3756 5538 3790
rect 5572 3756 5730 3790
rect 5764 3756 5922 3790
rect 5956 3756 6114 3790
rect 6148 3756 6306 3790
rect 6340 3756 6498 3790
rect 6532 3756 6690 3790
rect 6724 3756 6882 3790
rect 6916 3756 7074 3790
rect 7108 3756 7266 3790
rect 7300 3756 8218 3790
rect 8252 3756 8410 3790
rect 8444 3756 8602 3790
rect 8636 3756 8794 3790
rect 8828 3756 8986 3790
rect 9020 3756 9178 3790
rect 9212 3756 9370 3790
rect 9404 3756 9562 3790
rect 9596 3756 9754 3790
rect 9788 3756 9946 3790
rect 9980 3756 10138 3790
rect 10172 3756 10330 3790
rect 10364 3756 10522 3790
rect 10556 3756 10714 3790
rect 10748 3756 10906 3790
rect 10940 3756 10972 3790
rect -1180 3740 116 3748
rect 1620 3740 2916 3748
rect -1180 3682 320 3740
rect -1180 3648 -886 3682
rect -852 3648 -694 3682
rect -660 3648 -502 3682
rect -468 3648 -310 3682
rect -276 3648 -118 3682
rect -84 3648 320 3682
rect -1180 3640 320 3648
rect -1180 3180 -1080 3640
rect -1036 3598 -990 3610
rect -940 3608 -894 3610
rect -1036 3392 -1030 3598
rect -996 3392 -990 3598
rect -954 3428 -944 3608
rect -892 3428 -882 3608
rect -844 3598 -798 3610
rect -748 3608 -702 3610
rect -1050 3212 -1040 3392
rect -988 3212 -978 3392
rect -940 3222 -934 3428
rect -900 3222 -894 3428
rect -844 3392 -838 3598
rect -804 3392 -798 3598
rect -762 3428 -752 3608
rect -700 3428 -690 3608
rect -652 3598 -606 3610
rect -556 3608 -510 3610
rect -1036 3210 -990 3212
rect -940 3210 -894 3222
rect -858 3212 -848 3392
rect -796 3212 -786 3392
rect -748 3222 -742 3428
rect -708 3222 -702 3428
rect -652 3392 -646 3598
rect -612 3392 -606 3598
rect -570 3428 -560 3608
rect -508 3428 -498 3608
rect -460 3598 -414 3610
rect -364 3608 -318 3610
rect -844 3210 -798 3212
rect -748 3210 -702 3222
rect -666 3212 -656 3392
rect -604 3212 -594 3392
rect -556 3222 -550 3428
rect -516 3222 -510 3428
rect -460 3392 -454 3598
rect -420 3392 -414 3598
rect -378 3428 -368 3608
rect -316 3428 -306 3608
rect -268 3598 -222 3610
rect -172 3608 -126 3610
rect -652 3210 -606 3212
rect -556 3210 -510 3222
rect -474 3212 -464 3392
rect -412 3212 -402 3392
rect -364 3222 -358 3428
rect -324 3222 -318 3428
rect -268 3392 -262 3598
rect -228 3392 -222 3598
rect -186 3428 -176 3608
rect -124 3428 -114 3608
rect -76 3598 -30 3610
rect -460 3210 -414 3212
rect -364 3210 -318 3222
rect -282 3212 -272 3392
rect -220 3212 -210 3392
rect -172 3222 -166 3428
rect -132 3222 -126 3428
rect -76 3392 -70 3598
rect -36 3392 -30 3598
rect 16 3460 320 3640
rect 1380 3682 2916 3740
rect 1380 3648 1914 3682
rect 1948 3648 2106 3682
rect 2140 3648 2298 3682
rect 2332 3648 2490 3682
rect 2524 3648 2682 3682
rect 2716 3648 2916 3682
rect 1380 3640 2916 3648
rect 1380 3460 1720 3640
rect -268 3210 -222 3212
rect -172 3210 -126 3222
rect -90 3212 -80 3392
rect -28 3212 -18 3392
rect -76 3210 -30 3212
rect 16 3180 116 3460
rect -1180 3172 116 3180
rect -1180 3138 -982 3172
rect -948 3138 -790 3172
rect -756 3138 -598 3172
rect -564 3138 -406 3172
rect -372 3138 -214 3172
rect -180 3138 116 3172
rect -1180 3072 116 3138
rect 1620 3180 1720 3460
rect 1764 3598 1810 3610
rect 1860 3608 1906 3610
rect 1764 3392 1770 3598
rect 1804 3392 1810 3598
rect 1846 3428 1856 3608
rect 1908 3428 1918 3608
rect 1956 3598 2002 3610
rect 2052 3608 2098 3610
rect 1750 3212 1760 3392
rect 1812 3212 1822 3392
rect 1860 3222 1866 3428
rect 1900 3222 1906 3428
rect 1956 3392 1962 3598
rect 1996 3392 2002 3598
rect 2038 3428 2048 3608
rect 2100 3428 2110 3608
rect 2148 3598 2194 3610
rect 2244 3608 2290 3610
rect 1764 3210 1810 3212
rect 1860 3210 1906 3222
rect 1942 3212 1952 3392
rect 2004 3212 2014 3392
rect 2052 3222 2058 3428
rect 2092 3222 2098 3428
rect 2148 3392 2154 3598
rect 2188 3392 2194 3598
rect 2230 3428 2240 3608
rect 2292 3428 2302 3608
rect 2340 3598 2386 3610
rect 2436 3608 2482 3610
rect 1956 3210 2002 3212
rect 2052 3210 2098 3222
rect 2134 3212 2144 3392
rect 2196 3212 2206 3392
rect 2244 3222 2250 3428
rect 2284 3222 2290 3428
rect 2340 3392 2346 3598
rect 2380 3392 2386 3598
rect 2422 3428 2432 3608
rect 2484 3428 2494 3608
rect 2532 3598 2578 3610
rect 2628 3608 2674 3610
rect 2148 3210 2194 3212
rect 2244 3210 2290 3222
rect 2326 3212 2336 3392
rect 2388 3212 2398 3392
rect 2436 3222 2442 3428
rect 2476 3222 2482 3428
rect 2532 3392 2538 3598
rect 2572 3392 2578 3598
rect 2614 3428 2624 3608
rect 2676 3428 2686 3608
rect 2724 3598 2770 3610
rect 2340 3210 2386 3212
rect 2436 3210 2482 3222
rect 2518 3212 2528 3392
rect 2580 3212 2590 3392
rect 2628 3222 2634 3428
rect 2668 3222 2674 3428
rect 2724 3392 2730 3598
rect 2764 3392 2770 3598
rect 2532 3210 2578 3212
rect 2628 3210 2674 3222
rect 2710 3212 2720 3392
rect 2772 3212 2782 3392
rect 2724 3210 2770 3212
rect 2816 3180 2916 3640
rect 1620 3172 2916 3180
rect 1620 3138 1818 3172
rect 1852 3138 2010 3172
rect 2044 3138 2202 3172
rect 2236 3138 2394 3172
rect 2428 3138 2586 3172
rect 2620 3138 2916 3172
rect 1620 3072 2916 3138
rect 4160 3682 10972 3756
rect 4160 3648 4578 3682
rect 4612 3648 4770 3682
rect 4804 3648 4962 3682
rect 4996 3648 5154 3682
rect 5188 3648 5346 3682
rect 5380 3648 5538 3682
rect 5572 3648 5730 3682
rect 5764 3648 5922 3682
rect 5956 3648 6114 3682
rect 6148 3648 6306 3682
rect 6340 3648 6498 3682
rect 6532 3648 6690 3682
rect 6724 3648 6882 3682
rect 6916 3648 7074 3682
rect 7108 3648 7266 3682
rect 7300 3648 8218 3682
rect 8252 3648 8410 3682
rect 8444 3648 8602 3682
rect 8636 3648 8794 3682
rect 8828 3648 8986 3682
rect 9020 3648 9178 3682
rect 9212 3648 9370 3682
rect 9404 3648 9562 3682
rect 9596 3648 9754 3682
rect 9788 3648 9946 3682
rect 9980 3648 10138 3682
rect 10172 3648 10330 3682
rect 10364 3648 10522 3682
rect 10556 3648 10714 3682
rect 10748 3648 10906 3682
rect 10940 3648 10972 3682
rect 4160 3640 10972 3648
rect 12176 3790 18592 3796
rect 12176 3756 12198 3790
rect 12232 3756 12390 3790
rect 12424 3756 12582 3790
rect 12616 3756 12774 3790
rect 12808 3756 12966 3790
rect 13000 3756 13158 3790
rect 13192 3756 13350 3790
rect 13384 3756 13542 3790
rect 13576 3756 13734 3790
rect 13768 3756 13926 3790
rect 13960 3756 14118 3790
rect 14152 3756 14310 3790
rect 14344 3756 14502 3790
rect 14536 3756 14694 3790
rect 14728 3756 14886 3790
rect 14920 3756 15838 3790
rect 15872 3756 16030 3790
rect 16064 3756 16222 3790
rect 16256 3756 16414 3790
rect 16448 3756 16606 3790
rect 16640 3756 16798 3790
rect 16832 3756 16990 3790
rect 17024 3756 17182 3790
rect 17216 3756 17374 3790
rect 17408 3756 17566 3790
rect 17600 3756 17758 3790
rect 17792 3756 17950 3790
rect 17984 3756 18142 3790
rect 18176 3756 18334 3790
rect 18368 3756 18526 3790
rect 18560 3756 18592 3790
rect 12176 3682 18592 3756
rect 12176 3648 12198 3682
rect 12232 3648 12390 3682
rect 12424 3648 12582 3682
rect 12616 3648 12774 3682
rect 12808 3648 12966 3682
rect 13000 3648 13158 3682
rect 13192 3648 13350 3682
rect 13384 3648 13542 3682
rect 13576 3648 13734 3682
rect 13768 3648 13926 3682
rect 13960 3648 14118 3682
rect 14152 3648 14310 3682
rect 14344 3648 14502 3682
rect 14536 3648 14694 3682
rect 14728 3648 14886 3682
rect 14920 3648 15838 3682
rect 15872 3648 16030 3682
rect 16064 3648 16222 3682
rect 16256 3648 16414 3682
rect 16448 3648 16606 3682
rect 16640 3648 16798 3682
rect 16832 3648 16990 3682
rect 17024 3648 17182 3682
rect 17216 3648 17374 3682
rect 17408 3648 17566 3682
rect 17600 3648 17758 3682
rect 17792 3648 17950 3682
rect 17984 3648 18142 3682
rect 18176 3648 18334 3682
rect 18368 3648 18526 3682
rect 18560 3648 18592 3682
rect 12176 3640 18592 3648
rect 4160 3180 4324 3640
rect 4428 3598 4474 3610
rect 4428 3392 4434 3598
rect 4468 3392 4474 3598
rect 4510 3428 4520 3612
rect 4572 3428 4582 3612
rect 4620 3598 4666 3610
rect 4414 3208 4424 3392
rect 4476 3208 4486 3392
rect 4524 3222 4530 3428
rect 4564 3222 4570 3428
rect 4620 3392 4626 3598
rect 4660 3392 4666 3598
rect 4702 3428 4712 3612
rect 4764 3428 4774 3612
rect 4812 3598 4858 3610
rect 4524 3210 4570 3222
rect 4606 3208 4616 3392
rect 4668 3208 4678 3392
rect 4716 3222 4722 3428
rect 4756 3222 4762 3428
rect 4812 3392 4818 3598
rect 4852 3392 4858 3598
rect 4894 3428 4904 3612
rect 4956 3428 4966 3612
rect 5004 3598 5050 3610
rect 4716 3210 4762 3222
rect 4798 3208 4808 3392
rect 4860 3208 4870 3392
rect 4908 3222 4914 3428
rect 4948 3222 4954 3428
rect 5004 3392 5010 3598
rect 5044 3392 5050 3598
rect 5086 3428 5096 3612
rect 5148 3428 5158 3612
rect 5196 3598 5242 3610
rect 4908 3210 4954 3222
rect 4990 3208 5000 3392
rect 5052 3208 5062 3392
rect 5100 3222 5106 3428
rect 5140 3222 5146 3428
rect 5196 3392 5202 3598
rect 5236 3392 5242 3598
rect 5278 3428 5288 3612
rect 5340 3428 5350 3612
rect 5388 3598 5434 3610
rect 5100 3210 5146 3222
rect 5182 3208 5192 3392
rect 5244 3208 5254 3392
rect 5292 3222 5298 3428
rect 5332 3222 5338 3428
rect 5388 3392 5394 3598
rect 5428 3392 5434 3598
rect 5470 3428 5480 3612
rect 5532 3428 5542 3612
rect 5580 3598 5626 3610
rect 5292 3210 5338 3222
rect 5374 3208 5384 3392
rect 5436 3208 5446 3392
rect 5484 3222 5490 3428
rect 5524 3222 5530 3428
rect 5580 3392 5586 3598
rect 5620 3392 5626 3598
rect 5662 3428 5672 3612
rect 5724 3428 5734 3612
rect 5772 3598 5818 3610
rect 5484 3210 5530 3222
rect 5566 3208 5576 3392
rect 5628 3208 5638 3392
rect 5676 3222 5682 3428
rect 5716 3222 5722 3428
rect 5772 3392 5778 3598
rect 5812 3392 5818 3598
rect 5854 3428 5864 3612
rect 5916 3428 5926 3612
rect 5964 3598 6010 3610
rect 5676 3210 5722 3222
rect 5758 3208 5768 3392
rect 5820 3208 5830 3392
rect 5868 3222 5874 3428
rect 5908 3222 5914 3428
rect 5964 3392 5970 3598
rect 6004 3392 6010 3598
rect 6046 3428 6056 3612
rect 6108 3428 6118 3612
rect 6156 3598 6202 3610
rect 5868 3210 5914 3222
rect 5950 3208 5960 3392
rect 6012 3208 6022 3392
rect 6060 3222 6066 3428
rect 6100 3222 6106 3428
rect 6156 3392 6162 3598
rect 6196 3392 6202 3598
rect 6238 3428 6248 3612
rect 6300 3428 6310 3612
rect 6348 3598 6394 3610
rect 6060 3210 6106 3222
rect 6142 3208 6152 3392
rect 6204 3208 6214 3392
rect 6252 3222 6258 3428
rect 6292 3222 6298 3428
rect 6348 3392 6354 3598
rect 6388 3392 6394 3598
rect 6430 3428 6440 3612
rect 6492 3428 6502 3612
rect 6540 3598 6586 3610
rect 6252 3210 6298 3222
rect 6334 3208 6344 3392
rect 6396 3208 6406 3392
rect 6444 3222 6450 3428
rect 6484 3222 6490 3428
rect 6540 3392 6546 3598
rect 6580 3392 6586 3598
rect 6622 3428 6632 3612
rect 6684 3428 6694 3612
rect 6732 3598 6778 3610
rect 6444 3210 6490 3222
rect 6526 3208 6536 3392
rect 6588 3208 6598 3392
rect 6636 3222 6642 3428
rect 6676 3222 6682 3428
rect 6732 3392 6738 3598
rect 6772 3392 6778 3598
rect 6814 3428 6824 3612
rect 6876 3428 6886 3612
rect 6924 3598 6970 3610
rect 6636 3210 6682 3222
rect 6718 3208 6728 3392
rect 6780 3208 6790 3392
rect 6828 3222 6834 3428
rect 6868 3222 6874 3428
rect 6924 3392 6930 3598
rect 6964 3392 6970 3598
rect 7006 3428 7016 3612
rect 7068 3428 7078 3612
rect 7116 3598 7162 3610
rect 6828 3210 6874 3222
rect 6910 3208 6920 3392
rect 6972 3208 6982 3392
rect 7020 3222 7026 3428
rect 7060 3222 7066 3428
rect 7116 3392 7122 3598
rect 7156 3392 7162 3598
rect 7198 3428 7208 3612
rect 7260 3428 7270 3612
rect 7308 3598 7354 3610
rect 7020 3210 7066 3222
rect 7102 3208 7112 3392
rect 7164 3208 7174 3392
rect 7212 3222 7218 3428
rect 7252 3222 7258 3428
rect 7308 3392 7314 3598
rect 7348 3392 7354 3598
rect 7212 3210 7258 3222
rect 7294 3208 7304 3392
rect 7356 3208 7366 3392
rect 7468 3180 7916 3640
rect 8068 3598 8114 3610
rect 8068 3392 8074 3598
rect 8108 3392 8114 3598
rect 8150 3428 8160 3612
rect 8212 3428 8222 3612
rect 8260 3598 8306 3610
rect 8054 3208 8064 3392
rect 8116 3208 8126 3392
rect 8164 3222 8170 3428
rect 8204 3222 8210 3428
rect 8260 3392 8266 3598
rect 8300 3392 8306 3598
rect 8342 3428 8352 3612
rect 8404 3428 8414 3612
rect 8452 3598 8498 3610
rect 8164 3210 8210 3222
rect 8246 3208 8256 3392
rect 8308 3208 8318 3392
rect 8356 3222 8362 3428
rect 8396 3222 8402 3428
rect 8452 3392 8458 3598
rect 8492 3392 8498 3598
rect 8534 3428 8544 3612
rect 8596 3428 8606 3612
rect 8644 3598 8690 3610
rect 8356 3210 8402 3222
rect 8438 3208 8448 3392
rect 8500 3208 8510 3392
rect 8548 3222 8554 3428
rect 8588 3222 8594 3428
rect 8644 3392 8650 3598
rect 8684 3392 8690 3598
rect 8726 3428 8736 3612
rect 8788 3428 8798 3612
rect 8836 3598 8882 3610
rect 8548 3210 8594 3222
rect 8630 3208 8640 3392
rect 8692 3208 8702 3392
rect 8740 3222 8746 3428
rect 8780 3222 8786 3428
rect 8836 3392 8842 3598
rect 8876 3392 8882 3598
rect 8918 3428 8928 3612
rect 8980 3428 8990 3612
rect 9028 3598 9074 3610
rect 8740 3210 8786 3222
rect 8822 3208 8832 3392
rect 8884 3208 8894 3392
rect 8932 3222 8938 3428
rect 8972 3222 8978 3428
rect 9028 3392 9034 3598
rect 9068 3392 9074 3598
rect 9110 3428 9120 3612
rect 9172 3428 9182 3612
rect 9220 3598 9266 3610
rect 8932 3210 8978 3222
rect 9014 3208 9024 3392
rect 9076 3208 9086 3392
rect 9124 3222 9130 3428
rect 9164 3222 9170 3428
rect 9220 3392 9226 3598
rect 9260 3392 9266 3598
rect 9302 3428 9312 3612
rect 9364 3428 9374 3612
rect 9412 3598 9458 3610
rect 9124 3210 9170 3222
rect 9206 3208 9216 3392
rect 9268 3208 9278 3392
rect 9316 3222 9322 3428
rect 9356 3222 9362 3428
rect 9412 3392 9418 3598
rect 9452 3392 9458 3598
rect 9494 3428 9504 3612
rect 9556 3428 9566 3612
rect 9604 3598 9650 3610
rect 9316 3210 9362 3222
rect 9398 3208 9408 3392
rect 9460 3208 9470 3392
rect 9508 3222 9514 3428
rect 9548 3222 9554 3428
rect 9604 3392 9610 3598
rect 9644 3392 9650 3598
rect 9686 3428 9696 3612
rect 9748 3428 9758 3612
rect 9796 3598 9842 3610
rect 9508 3210 9554 3222
rect 9590 3208 9600 3392
rect 9652 3208 9662 3392
rect 9700 3222 9706 3428
rect 9740 3222 9746 3428
rect 9796 3392 9802 3598
rect 9836 3392 9842 3598
rect 9878 3428 9888 3612
rect 9940 3428 9950 3612
rect 9988 3598 10034 3610
rect 9700 3210 9746 3222
rect 9782 3208 9792 3392
rect 9844 3208 9854 3392
rect 9892 3222 9898 3428
rect 9932 3222 9938 3428
rect 9988 3392 9994 3598
rect 10028 3392 10034 3598
rect 10070 3428 10080 3612
rect 10132 3428 10142 3612
rect 10180 3598 10226 3610
rect 9892 3210 9938 3222
rect 9974 3208 9984 3392
rect 10036 3208 10046 3392
rect 10084 3222 10090 3428
rect 10124 3222 10130 3428
rect 10180 3392 10186 3598
rect 10220 3392 10226 3598
rect 10262 3428 10272 3612
rect 10324 3428 10334 3612
rect 10372 3598 10418 3610
rect 10084 3210 10130 3222
rect 10166 3208 10176 3392
rect 10228 3208 10238 3392
rect 10276 3222 10282 3428
rect 10316 3222 10322 3428
rect 10372 3392 10378 3598
rect 10412 3392 10418 3598
rect 10454 3428 10464 3612
rect 10516 3428 10526 3612
rect 10564 3598 10610 3610
rect 10276 3210 10322 3222
rect 10358 3208 10368 3392
rect 10420 3208 10430 3392
rect 10468 3222 10474 3428
rect 10508 3222 10514 3428
rect 10564 3392 10570 3598
rect 10604 3392 10610 3598
rect 10646 3428 10656 3612
rect 10708 3428 10718 3612
rect 10756 3598 10802 3610
rect 10468 3210 10514 3222
rect 10550 3208 10560 3392
rect 10612 3208 10622 3392
rect 10660 3222 10666 3428
rect 10700 3222 10706 3428
rect 10756 3392 10762 3598
rect 10796 3392 10802 3598
rect 10838 3428 10848 3612
rect 10900 3428 10910 3612
rect 10948 3598 10994 3610
rect 10660 3210 10706 3222
rect 10742 3208 10752 3392
rect 10804 3208 10814 3392
rect 10852 3222 10858 3428
rect 10892 3222 10898 3428
rect 10948 3392 10954 3598
rect 10988 3392 10994 3598
rect 12048 3598 12094 3610
rect 12048 3392 12054 3598
rect 12088 3392 12094 3598
rect 12130 3428 12140 3612
rect 12192 3428 12202 3612
rect 12240 3598 12286 3610
rect 10852 3210 10898 3222
rect 10934 3208 10944 3392
rect 10996 3208 11006 3392
rect 12034 3208 12044 3392
rect 12096 3208 12106 3392
rect 12144 3222 12150 3428
rect 12184 3222 12190 3428
rect 12240 3392 12246 3598
rect 12280 3392 12286 3598
rect 12322 3428 12332 3612
rect 12384 3428 12394 3612
rect 12432 3598 12478 3610
rect 12144 3210 12190 3222
rect 12226 3208 12236 3392
rect 12288 3208 12298 3392
rect 12336 3222 12342 3428
rect 12376 3222 12382 3428
rect 12432 3392 12438 3598
rect 12472 3392 12478 3598
rect 12514 3428 12524 3612
rect 12576 3428 12586 3612
rect 12624 3598 12670 3610
rect 12336 3210 12382 3222
rect 12418 3208 12428 3392
rect 12480 3208 12490 3392
rect 12528 3222 12534 3428
rect 12568 3222 12574 3428
rect 12624 3392 12630 3598
rect 12664 3392 12670 3598
rect 12706 3428 12716 3612
rect 12768 3428 12778 3612
rect 12816 3598 12862 3610
rect 12528 3210 12574 3222
rect 12610 3208 12620 3392
rect 12672 3208 12682 3392
rect 12720 3222 12726 3428
rect 12760 3222 12766 3428
rect 12816 3392 12822 3598
rect 12856 3392 12862 3598
rect 12898 3428 12908 3612
rect 12960 3428 12970 3612
rect 13008 3598 13054 3610
rect 12720 3210 12766 3222
rect 12802 3208 12812 3392
rect 12864 3208 12874 3392
rect 12912 3222 12918 3428
rect 12952 3222 12958 3428
rect 13008 3392 13014 3598
rect 13048 3392 13054 3598
rect 13090 3428 13100 3612
rect 13152 3428 13162 3612
rect 13200 3598 13246 3610
rect 12912 3210 12958 3222
rect 12994 3208 13004 3392
rect 13056 3208 13066 3392
rect 13104 3222 13110 3428
rect 13144 3222 13150 3428
rect 13200 3392 13206 3598
rect 13240 3392 13246 3598
rect 13282 3428 13292 3612
rect 13344 3428 13354 3612
rect 13392 3598 13438 3610
rect 13104 3210 13150 3222
rect 13186 3208 13196 3392
rect 13248 3208 13258 3392
rect 13296 3222 13302 3428
rect 13336 3222 13342 3428
rect 13392 3392 13398 3598
rect 13432 3392 13438 3598
rect 13474 3428 13484 3612
rect 13536 3428 13546 3612
rect 13584 3598 13630 3610
rect 13296 3210 13342 3222
rect 13378 3208 13388 3392
rect 13440 3208 13450 3392
rect 13488 3222 13494 3428
rect 13528 3222 13534 3428
rect 13584 3392 13590 3598
rect 13624 3392 13630 3598
rect 13666 3428 13676 3612
rect 13728 3428 13738 3612
rect 13776 3598 13822 3610
rect 13488 3210 13534 3222
rect 13570 3208 13580 3392
rect 13632 3208 13642 3392
rect 13680 3222 13686 3428
rect 13720 3222 13726 3428
rect 13776 3392 13782 3598
rect 13816 3392 13822 3598
rect 13858 3428 13868 3612
rect 13920 3428 13930 3612
rect 13968 3598 14014 3610
rect 13680 3210 13726 3222
rect 13762 3208 13772 3392
rect 13824 3208 13834 3392
rect 13872 3222 13878 3428
rect 13912 3222 13918 3428
rect 13968 3392 13974 3598
rect 14008 3392 14014 3598
rect 14050 3428 14060 3612
rect 14112 3428 14122 3612
rect 14160 3598 14206 3610
rect 13872 3210 13918 3222
rect 13954 3208 13964 3392
rect 14016 3208 14026 3392
rect 14064 3222 14070 3428
rect 14104 3222 14110 3428
rect 14160 3392 14166 3598
rect 14200 3392 14206 3598
rect 14242 3428 14252 3612
rect 14304 3428 14314 3612
rect 14352 3598 14398 3610
rect 14064 3210 14110 3222
rect 14146 3208 14156 3392
rect 14208 3208 14218 3392
rect 14256 3222 14262 3428
rect 14296 3222 14302 3428
rect 14352 3392 14358 3598
rect 14392 3392 14398 3598
rect 14434 3428 14444 3612
rect 14496 3428 14506 3612
rect 14544 3598 14590 3610
rect 14256 3210 14302 3222
rect 14338 3208 14348 3392
rect 14400 3208 14410 3392
rect 14448 3222 14454 3428
rect 14488 3222 14494 3428
rect 14544 3392 14550 3598
rect 14584 3392 14590 3598
rect 14626 3428 14636 3612
rect 14688 3428 14698 3612
rect 14736 3598 14782 3610
rect 14448 3210 14494 3222
rect 14530 3208 14540 3392
rect 14592 3208 14602 3392
rect 14640 3222 14646 3428
rect 14680 3222 14686 3428
rect 14736 3392 14742 3598
rect 14776 3392 14782 3598
rect 14818 3428 14828 3612
rect 14880 3428 14890 3612
rect 14928 3598 14974 3610
rect 14640 3210 14686 3222
rect 14722 3208 14732 3392
rect 14784 3208 14794 3392
rect 14832 3222 14838 3428
rect 14872 3222 14878 3428
rect 14928 3392 14934 3598
rect 14968 3392 14974 3598
rect 14832 3210 14878 3222
rect 14914 3208 14924 3392
rect 14976 3208 14986 3392
rect 15088 3180 15536 3640
rect 15688 3598 15734 3610
rect 15688 3392 15694 3598
rect 15728 3392 15734 3598
rect 15770 3428 15780 3612
rect 15832 3428 15842 3612
rect 15880 3598 15926 3610
rect 15674 3208 15684 3392
rect 15736 3208 15746 3392
rect 15784 3222 15790 3428
rect 15824 3222 15830 3428
rect 15880 3392 15886 3598
rect 15920 3392 15926 3598
rect 15962 3428 15972 3612
rect 16024 3428 16034 3612
rect 16072 3598 16118 3610
rect 15784 3210 15830 3222
rect 15866 3208 15876 3392
rect 15928 3208 15938 3392
rect 15976 3222 15982 3428
rect 16016 3222 16022 3428
rect 16072 3392 16078 3598
rect 16112 3392 16118 3598
rect 16154 3428 16164 3612
rect 16216 3428 16226 3612
rect 16264 3598 16310 3610
rect 15976 3210 16022 3222
rect 16058 3208 16068 3392
rect 16120 3208 16130 3392
rect 16168 3222 16174 3428
rect 16208 3222 16214 3428
rect 16264 3392 16270 3598
rect 16304 3392 16310 3598
rect 16346 3428 16356 3612
rect 16408 3428 16418 3612
rect 16456 3598 16502 3610
rect 16168 3210 16214 3222
rect 16250 3208 16260 3392
rect 16312 3208 16322 3392
rect 16360 3222 16366 3428
rect 16400 3222 16406 3428
rect 16456 3392 16462 3598
rect 16496 3392 16502 3598
rect 16538 3428 16548 3612
rect 16600 3428 16610 3612
rect 16648 3598 16694 3610
rect 16360 3210 16406 3222
rect 16442 3208 16452 3392
rect 16504 3208 16514 3392
rect 16552 3222 16558 3428
rect 16592 3222 16598 3428
rect 16648 3392 16654 3598
rect 16688 3392 16694 3598
rect 16730 3428 16740 3612
rect 16792 3428 16802 3612
rect 16840 3598 16886 3610
rect 16552 3210 16598 3222
rect 16634 3208 16644 3392
rect 16696 3208 16706 3392
rect 16744 3222 16750 3428
rect 16784 3222 16790 3428
rect 16840 3392 16846 3598
rect 16880 3392 16886 3598
rect 16922 3428 16932 3612
rect 16984 3428 16994 3612
rect 17032 3598 17078 3610
rect 16744 3210 16790 3222
rect 16826 3208 16836 3392
rect 16888 3208 16898 3392
rect 16936 3222 16942 3428
rect 16976 3222 16982 3428
rect 17032 3392 17038 3598
rect 17072 3392 17078 3598
rect 17114 3428 17124 3612
rect 17176 3428 17186 3612
rect 17224 3598 17270 3610
rect 16936 3210 16982 3222
rect 17018 3208 17028 3392
rect 17080 3208 17090 3392
rect 17128 3222 17134 3428
rect 17168 3222 17174 3428
rect 17224 3392 17230 3598
rect 17264 3392 17270 3598
rect 17306 3428 17316 3612
rect 17368 3428 17378 3612
rect 17416 3598 17462 3610
rect 17128 3210 17174 3222
rect 17210 3208 17220 3392
rect 17272 3208 17282 3392
rect 17320 3222 17326 3428
rect 17360 3222 17366 3428
rect 17416 3392 17422 3598
rect 17456 3392 17462 3598
rect 17498 3428 17508 3612
rect 17560 3428 17570 3612
rect 17608 3598 17654 3610
rect 17320 3210 17366 3222
rect 17402 3208 17412 3392
rect 17464 3208 17474 3392
rect 17512 3222 17518 3428
rect 17552 3222 17558 3428
rect 17608 3392 17614 3598
rect 17648 3392 17654 3598
rect 17690 3428 17700 3612
rect 17752 3428 17762 3612
rect 17800 3598 17846 3610
rect 17512 3210 17558 3222
rect 17594 3208 17604 3392
rect 17656 3208 17666 3392
rect 17704 3222 17710 3428
rect 17744 3222 17750 3428
rect 17800 3392 17806 3598
rect 17840 3392 17846 3598
rect 17882 3428 17892 3612
rect 17944 3428 17954 3612
rect 17992 3598 18038 3610
rect 17704 3210 17750 3222
rect 17786 3208 17796 3392
rect 17848 3208 17858 3392
rect 17896 3222 17902 3428
rect 17936 3222 17942 3428
rect 17992 3392 17998 3598
rect 18032 3392 18038 3598
rect 18074 3428 18084 3612
rect 18136 3428 18146 3612
rect 18184 3598 18230 3610
rect 17896 3210 17942 3222
rect 17978 3208 17988 3392
rect 18040 3208 18050 3392
rect 18088 3222 18094 3428
rect 18128 3222 18134 3428
rect 18184 3392 18190 3598
rect 18224 3392 18230 3598
rect 18266 3428 18276 3612
rect 18328 3428 18338 3612
rect 18376 3598 18422 3610
rect 18088 3210 18134 3222
rect 18170 3208 18180 3392
rect 18232 3208 18242 3392
rect 18280 3222 18286 3428
rect 18320 3222 18326 3428
rect 18376 3392 18382 3598
rect 18416 3392 18422 3598
rect 18458 3428 18468 3612
rect 18520 3428 18530 3612
rect 18568 3598 18614 3610
rect 18280 3210 18326 3222
rect 18362 3208 18372 3392
rect 18424 3208 18434 3392
rect 18472 3222 18478 3428
rect 18512 3222 18518 3428
rect 18568 3392 18574 3598
rect 18608 3392 18614 3598
rect 18472 3210 18518 3222
rect 18554 3208 18564 3392
rect 18616 3208 18626 3392
rect 4160 3172 10924 3180
rect 4160 3138 4482 3172
rect 4516 3138 4674 3172
rect 4708 3138 4866 3172
rect 4900 3138 5058 3172
rect 5092 3138 5250 3172
rect 5284 3138 5442 3172
rect 5476 3138 5634 3172
rect 5668 3138 5826 3172
rect 5860 3138 6018 3172
rect 6052 3138 6210 3172
rect 6244 3138 6402 3172
rect 6436 3138 6594 3172
rect 6628 3138 6786 3172
rect 6820 3138 6978 3172
rect 7012 3138 7170 3172
rect 7204 3138 8122 3172
rect 8156 3138 8314 3172
rect 8348 3138 8506 3172
rect 8540 3138 8698 3172
rect 8732 3138 8890 3172
rect 8924 3138 9082 3172
rect 9116 3138 9274 3172
rect 9308 3138 9466 3172
rect 9500 3138 9658 3172
rect 9692 3138 9850 3172
rect 9884 3138 10042 3172
rect 10076 3138 10234 3172
rect 10268 3138 10426 3172
rect 10460 3138 10618 3172
rect 10652 3138 10810 3172
rect 10844 3138 10924 3172
rect 4160 3040 10924 3138
rect 12064 3172 18544 3180
rect 12064 3138 12102 3172
rect 12136 3138 12294 3172
rect 12328 3138 12486 3172
rect 12520 3138 12678 3172
rect 12712 3138 12870 3172
rect 12904 3138 13062 3172
rect 13096 3138 13254 3172
rect 13288 3138 13446 3172
rect 13480 3138 13638 3172
rect 13672 3138 13830 3172
rect 13864 3138 14022 3172
rect 14056 3138 14214 3172
rect 14248 3138 14406 3172
rect 14440 3138 14598 3172
rect 14632 3138 14790 3172
rect 14824 3138 15742 3172
rect 15776 3138 15934 3172
rect 15968 3138 16126 3172
rect 16160 3138 16318 3172
rect 16352 3138 16510 3172
rect 16544 3138 16702 3172
rect 16736 3138 16894 3172
rect 16928 3138 17086 3172
rect 17120 3138 17278 3172
rect 17312 3138 17470 3172
rect 17504 3138 17662 3172
rect 17696 3138 17854 3172
rect 17888 3138 18046 3172
rect 18080 3138 18238 3172
rect 18272 3138 18430 3172
rect 18464 3138 18544 3172
rect 12064 3040 18544 3138
rect 4260 2864 4972 2908
rect 4260 2830 4282 2864
rect 4316 2830 4474 2864
rect 4508 2830 4666 2864
rect 4700 2830 4972 2864
rect 4260 2824 4972 2830
rect 5300 2864 6012 2908
rect 5300 2830 5322 2864
rect 5356 2830 5514 2864
rect 5548 2830 5706 2864
rect 5740 2830 6012 2864
rect 5300 2824 6012 2830
rect 6340 2864 7052 2908
rect 6340 2830 6362 2864
rect 6396 2830 6554 2864
rect 6588 2830 6746 2864
rect 6780 2830 7052 2864
rect 6340 2824 7052 2830
rect 7380 2864 8092 2908
rect 7380 2830 7402 2864
rect 7436 2830 7594 2864
rect 7628 2830 7786 2864
rect 7820 2830 8092 2864
rect 7380 2824 8092 2830
rect 8420 2864 9132 2908
rect 8420 2830 8442 2864
rect 8476 2830 8634 2864
rect 8668 2830 8826 2864
rect 8860 2830 9132 2864
rect 8420 2824 9132 2830
rect 9460 2864 10172 2908
rect 9460 2830 9482 2864
rect 9516 2830 9674 2864
rect 9708 2830 9866 2864
rect 9900 2830 10172 2864
rect 9460 2824 10172 2830
rect 10500 2864 11212 2908
rect 10500 2830 10522 2864
rect 10556 2830 10714 2864
rect 10748 2830 10906 2864
rect 10940 2830 11212 2864
rect 10500 2824 11212 2830
rect 11880 2864 12592 2908
rect 11880 2830 11902 2864
rect 11936 2830 12094 2864
rect 12128 2830 12286 2864
rect 12320 2830 12592 2864
rect 11880 2824 12592 2830
rect 12920 2864 13632 2908
rect 12920 2830 12942 2864
rect 12976 2830 13134 2864
rect 13168 2830 13326 2864
rect 13360 2830 13632 2864
rect 12920 2824 13632 2830
rect 13960 2864 14672 2908
rect 13960 2830 13982 2864
rect 14016 2830 14174 2864
rect 14208 2830 14366 2864
rect 14400 2830 14672 2864
rect 13960 2824 14672 2830
rect 15000 2864 15712 2908
rect 15000 2830 15022 2864
rect 15056 2830 15214 2864
rect 15248 2830 15406 2864
rect 15440 2830 15712 2864
rect 15000 2824 15712 2830
rect 16040 2864 16752 2908
rect 16040 2830 16062 2864
rect 16096 2830 16254 2864
rect 16288 2830 16446 2864
rect 16480 2830 16752 2864
rect 16040 2824 16752 2830
rect 17080 2864 17792 2908
rect 17080 2830 17102 2864
rect 17136 2830 17294 2864
rect 17328 2830 17486 2864
rect 17520 2830 17792 2864
rect 17080 2824 17792 2830
rect 18120 2864 18832 2908
rect 18120 2830 18142 2864
rect 18176 2830 18334 2864
rect 18368 2830 18526 2864
rect 18560 2830 18832 2864
rect 18120 2824 18832 2830
rect -1544 2704 -832 2748
rect -1544 2670 -1522 2704
rect -1488 2670 -1330 2704
rect -1296 2670 -1138 2704
rect -1104 2670 -832 2704
rect -1544 2664 -832 2670
rect -504 2704 208 2748
rect -504 2670 -482 2704
rect -448 2670 -290 2704
rect -256 2670 -98 2704
rect -64 2670 208 2704
rect -504 2664 208 2670
rect 536 2704 1248 2748
rect 536 2670 558 2704
rect 592 2670 750 2704
rect 784 2670 942 2704
rect 976 2670 1248 2704
rect 536 2664 1248 2670
rect 1576 2704 2288 2748
rect 1576 2670 1598 2704
rect 1632 2670 1790 2704
rect 1824 2670 1982 2704
rect 2016 2670 2288 2704
rect 1576 2664 2288 2670
rect 2616 2704 3328 2748
rect 2616 2670 2638 2704
rect 2672 2670 2830 2704
rect 2864 2670 3022 2704
rect 3056 2670 3328 2704
rect 2616 2664 3328 2670
rect -1590 2452 -1580 2632
rect -1528 2452 -1518 2632
rect -1480 2620 -1434 2632
rect -1576 2244 -1570 2452
rect -1536 2244 -1530 2452
rect -1480 2412 -1474 2620
rect -1440 2412 -1434 2620
rect -1398 2452 -1388 2632
rect -1336 2452 -1326 2632
rect -1288 2620 -1242 2632
rect -1576 2232 -1530 2244
rect -1494 2232 -1484 2412
rect -1432 2232 -1422 2412
rect -1384 2244 -1378 2452
rect -1344 2244 -1338 2452
rect -1288 2412 -1282 2620
rect -1248 2412 -1242 2620
rect -1206 2452 -1196 2632
rect -1144 2452 -1134 2632
rect -1096 2620 -1050 2632
rect -1384 2232 -1338 2244
rect -1302 2232 -1292 2412
rect -1240 2232 -1230 2412
rect -1192 2244 -1186 2452
rect -1152 2244 -1146 2452
rect -1096 2412 -1090 2620
rect -1056 2412 -1050 2620
rect -1014 2452 -1004 2632
rect -952 2452 -942 2632
rect -1192 2232 -1146 2244
rect -1110 2232 -1100 2412
rect -1048 2232 -1038 2412
rect -1000 2244 -994 2452
rect -960 2244 -954 2452
rect -1000 2232 -954 2244
rect -912 2200 -832 2664
rect -550 2452 -540 2632
rect -488 2452 -478 2632
rect -440 2620 -394 2632
rect -536 2244 -530 2452
rect -496 2244 -490 2452
rect -440 2412 -434 2620
rect -400 2412 -394 2620
rect -358 2452 -348 2632
rect -296 2452 -286 2632
rect -248 2620 -202 2632
rect -536 2232 -490 2244
rect -454 2232 -444 2412
rect -392 2232 -382 2412
rect -344 2244 -338 2452
rect -304 2244 -298 2452
rect -248 2412 -242 2620
rect -208 2412 -202 2620
rect -166 2452 -156 2632
rect -104 2452 -94 2632
rect -56 2620 -10 2632
rect -344 2232 -298 2244
rect -262 2232 -252 2412
rect -200 2232 -190 2412
rect -152 2244 -146 2452
rect -112 2244 -106 2452
rect -56 2412 -50 2620
rect -16 2412 -10 2620
rect 26 2452 36 2632
rect 88 2452 98 2632
rect -152 2232 -106 2244
rect -70 2232 -60 2412
rect -8 2232 2 2412
rect 40 2244 46 2452
rect 80 2244 86 2452
rect 40 2232 86 2244
rect 128 2200 208 2664
rect 490 2452 500 2632
rect 552 2452 562 2632
rect 600 2620 646 2632
rect 504 2244 510 2452
rect 544 2244 550 2452
rect 600 2412 606 2620
rect 640 2412 646 2620
rect 682 2452 692 2632
rect 744 2452 754 2632
rect 792 2620 838 2632
rect 504 2232 550 2244
rect 586 2232 596 2412
rect 648 2232 658 2412
rect 696 2244 702 2452
rect 736 2244 742 2452
rect 792 2412 798 2620
rect 832 2412 838 2620
rect 874 2452 884 2632
rect 936 2452 946 2632
rect 984 2620 1030 2632
rect 696 2232 742 2244
rect 778 2232 788 2412
rect 840 2232 850 2412
rect 888 2244 894 2452
rect 928 2244 934 2452
rect 984 2412 990 2620
rect 1024 2412 1030 2620
rect 1066 2452 1076 2632
rect 1128 2452 1138 2632
rect 888 2232 934 2244
rect 970 2232 980 2412
rect 1032 2232 1042 2412
rect 1080 2244 1086 2452
rect 1120 2244 1126 2452
rect 1080 2232 1126 2244
rect 1168 2200 1248 2664
rect 1530 2452 1540 2632
rect 1592 2452 1602 2632
rect 1640 2620 1686 2632
rect 1544 2244 1550 2452
rect 1584 2244 1590 2452
rect 1640 2412 1646 2620
rect 1680 2412 1686 2620
rect 1722 2452 1732 2632
rect 1784 2452 1794 2632
rect 1832 2620 1878 2632
rect 1544 2232 1590 2244
rect 1626 2232 1636 2412
rect 1688 2232 1698 2412
rect 1736 2244 1742 2452
rect 1776 2244 1782 2452
rect 1832 2412 1838 2620
rect 1872 2412 1878 2620
rect 1914 2452 1924 2632
rect 1976 2452 1986 2632
rect 2024 2620 2070 2632
rect 1736 2232 1782 2244
rect 1818 2232 1828 2412
rect 1880 2232 1890 2412
rect 1928 2244 1934 2452
rect 1968 2244 1974 2452
rect 2024 2412 2030 2620
rect 2064 2412 2070 2620
rect 2106 2452 2116 2632
rect 2168 2452 2178 2632
rect 1928 2232 1974 2244
rect 2010 2232 2020 2412
rect 2072 2232 2082 2412
rect 2120 2244 2126 2452
rect 2160 2244 2166 2452
rect 2120 2232 2166 2244
rect 2208 2200 2288 2664
rect 2570 2452 2580 2632
rect 2632 2452 2642 2632
rect 2680 2620 2726 2632
rect 2584 2244 2590 2452
rect 2624 2244 2630 2452
rect 2680 2412 2686 2620
rect 2720 2412 2726 2620
rect 2762 2452 2772 2632
rect 2824 2452 2834 2632
rect 2872 2620 2918 2632
rect 2584 2232 2630 2244
rect 2666 2232 2676 2412
rect 2728 2232 2738 2412
rect 2776 2244 2782 2452
rect 2816 2244 2822 2452
rect 2872 2412 2878 2620
rect 2912 2412 2918 2620
rect 2954 2452 2964 2632
rect 3016 2452 3026 2632
rect 3064 2620 3110 2632
rect 2776 2232 2822 2244
rect 2858 2232 2868 2412
rect 2920 2232 2930 2412
rect 2968 2244 2974 2452
rect 3008 2244 3014 2452
rect 3064 2412 3070 2620
rect 3104 2412 3110 2620
rect 3146 2452 3156 2632
rect 3208 2452 3218 2632
rect 2968 2232 3014 2244
rect 3050 2232 3060 2412
rect 3112 2232 3122 2412
rect 3160 2244 3166 2452
rect 3200 2244 3206 2452
rect 3160 2232 3206 2244
rect 3248 2200 3328 2664
rect 4214 2612 4224 2792
rect 4276 2612 4286 2792
rect 4324 2780 4370 2792
rect 4228 2404 4234 2612
rect 4268 2404 4274 2612
rect 4324 2572 4330 2780
rect 4364 2572 4370 2780
rect 4406 2612 4416 2792
rect 4468 2612 4478 2792
rect 4516 2780 4562 2792
rect 4228 2392 4274 2404
rect 4310 2392 4320 2572
rect 4372 2392 4382 2572
rect 4420 2404 4426 2612
rect 4460 2404 4466 2612
rect 4516 2572 4522 2780
rect 4556 2572 4562 2780
rect 4598 2612 4608 2792
rect 4660 2612 4670 2792
rect 4708 2780 4754 2792
rect 4420 2392 4466 2404
rect 4502 2392 4512 2572
rect 4564 2392 4574 2572
rect 4612 2404 4618 2612
rect 4652 2404 4658 2612
rect 4708 2572 4714 2780
rect 4748 2572 4754 2780
rect 4790 2612 4800 2792
rect 4852 2612 4862 2792
rect 4612 2392 4658 2404
rect 4694 2392 4704 2572
rect 4756 2392 4766 2572
rect 4804 2404 4810 2612
rect 4844 2404 4850 2612
rect 4804 2392 4850 2404
rect 4892 2360 4972 2824
rect 5254 2612 5264 2792
rect 5316 2612 5326 2792
rect 5364 2780 5410 2792
rect 5268 2404 5274 2612
rect 5308 2404 5314 2612
rect 5364 2572 5370 2780
rect 5404 2572 5410 2780
rect 5446 2612 5456 2792
rect 5508 2612 5518 2792
rect 5556 2780 5602 2792
rect 5268 2392 5314 2404
rect 5350 2392 5360 2572
rect 5412 2392 5422 2572
rect 5460 2404 5466 2612
rect 5500 2404 5506 2612
rect 5556 2572 5562 2780
rect 5596 2572 5602 2780
rect 5638 2612 5648 2792
rect 5700 2612 5710 2792
rect 5748 2780 5794 2792
rect 5460 2392 5506 2404
rect 5542 2392 5552 2572
rect 5604 2392 5614 2572
rect 5652 2404 5658 2612
rect 5692 2404 5698 2612
rect 5748 2572 5754 2780
rect 5788 2572 5794 2780
rect 5830 2612 5840 2792
rect 5892 2612 5902 2792
rect 5652 2392 5698 2404
rect 5734 2392 5744 2572
rect 5796 2392 5806 2572
rect 5844 2404 5850 2612
rect 5884 2404 5890 2612
rect 5844 2392 5890 2404
rect 5932 2360 6012 2824
rect 6294 2612 6304 2792
rect 6356 2612 6366 2792
rect 6404 2780 6450 2792
rect 6308 2404 6314 2612
rect 6348 2404 6354 2612
rect 6404 2572 6410 2780
rect 6444 2572 6450 2780
rect 6486 2612 6496 2792
rect 6548 2612 6558 2792
rect 6596 2780 6642 2792
rect 6308 2392 6354 2404
rect 6390 2392 6400 2572
rect 6452 2392 6462 2572
rect 6500 2404 6506 2612
rect 6540 2404 6546 2612
rect 6596 2572 6602 2780
rect 6636 2572 6642 2780
rect 6678 2612 6688 2792
rect 6740 2612 6750 2792
rect 6788 2780 6834 2792
rect 6500 2392 6546 2404
rect 6582 2392 6592 2572
rect 6644 2392 6654 2572
rect 6692 2404 6698 2612
rect 6732 2404 6738 2612
rect 6788 2572 6794 2780
rect 6828 2572 6834 2780
rect 6870 2612 6880 2792
rect 6932 2612 6942 2792
rect 6692 2392 6738 2404
rect 6774 2392 6784 2572
rect 6836 2392 6846 2572
rect 6884 2404 6890 2612
rect 6924 2404 6930 2612
rect 6884 2392 6930 2404
rect 6972 2360 7052 2824
rect 7334 2612 7344 2792
rect 7396 2612 7406 2792
rect 7444 2780 7490 2792
rect 7348 2404 7354 2612
rect 7388 2404 7394 2612
rect 7444 2572 7450 2780
rect 7484 2572 7490 2780
rect 7526 2612 7536 2792
rect 7588 2612 7598 2792
rect 7636 2780 7682 2792
rect 7348 2392 7394 2404
rect 7430 2392 7440 2572
rect 7492 2392 7502 2572
rect 7540 2404 7546 2612
rect 7580 2404 7586 2612
rect 7636 2572 7642 2780
rect 7676 2572 7682 2780
rect 7718 2612 7728 2792
rect 7780 2612 7790 2792
rect 7828 2780 7874 2792
rect 7540 2392 7586 2404
rect 7622 2392 7632 2572
rect 7684 2392 7694 2572
rect 7732 2404 7738 2612
rect 7772 2404 7778 2612
rect 7828 2572 7834 2780
rect 7868 2572 7874 2780
rect 7910 2612 7920 2792
rect 7972 2612 7982 2792
rect 7732 2392 7778 2404
rect 7814 2392 7824 2572
rect 7876 2392 7886 2572
rect 7924 2404 7930 2612
rect 7964 2404 7970 2612
rect 7924 2392 7970 2404
rect 8012 2360 8092 2824
rect 8374 2612 8384 2792
rect 8436 2612 8446 2792
rect 8484 2780 8530 2792
rect 8388 2404 8394 2612
rect 8428 2404 8434 2612
rect 8484 2572 8490 2780
rect 8524 2572 8530 2780
rect 8566 2612 8576 2792
rect 8628 2612 8638 2792
rect 8676 2780 8722 2792
rect 8388 2392 8434 2404
rect 8470 2392 8480 2572
rect 8532 2392 8542 2572
rect 8580 2404 8586 2612
rect 8620 2404 8626 2612
rect 8676 2572 8682 2780
rect 8716 2572 8722 2780
rect 8758 2612 8768 2792
rect 8820 2612 8830 2792
rect 8868 2780 8914 2792
rect 8580 2392 8626 2404
rect 8662 2392 8672 2572
rect 8724 2392 8734 2572
rect 8772 2404 8778 2612
rect 8812 2404 8818 2612
rect 8868 2572 8874 2780
rect 8908 2572 8914 2780
rect 8950 2612 8960 2792
rect 9012 2612 9022 2792
rect 8772 2392 8818 2404
rect 8854 2392 8864 2572
rect 8916 2392 8926 2572
rect 8964 2404 8970 2612
rect 9004 2404 9010 2612
rect 8964 2392 9010 2404
rect 9052 2360 9132 2824
rect 9414 2612 9424 2792
rect 9476 2612 9486 2792
rect 9524 2780 9570 2792
rect 9428 2404 9434 2612
rect 9468 2404 9474 2612
rect 9524 2572 9530 2780
rect 9564 2572 9570 2780
rect 9606 2612 9616 2792
rect 9668 2612 9678 2792
rect 9716 2780 9762 2792
rect 9428 2392 9474 2404
rect 9510 2392 9520 2572
rect 9572 2392 9582 2572
rect 9620 2404 9626 2612
rect 9660 2404 9666 2612
rect 9716 2572 9722 2780
rect 9756 2572 9762 2780
rect 9798 2612 9808 2792
rect 9860 2612 9870 2792
rect 9908 2780 9954 2792
rect 9620 2392 9666 2404
rect 9702 2392 9712 2572
rect 9764 2392 9774 2572
rect 9812 2404 9818 2612
rect 9852 2404 9858 2612
rect 9908 2572 9914 2780
rect 9948 2572 9954 2780
rect 9990 2612 10000 2792
rect 10052 2612 10062 2792
rect 9812 2392 9858 2404
rect 9894 2392 9904 2572
rect 9956 2392 9966 2572
rect 10004 2404 10010 2612
rect 10044 2404 10050 2612
rect 10004 2392 10050 2404
rect 10092 2360 10172 2824
rect 10454 2612 10464 2792
rect 10516 2612 10526 2792
rect 10564 2780 10610 2792
rect 10468 2404 10474 2612
rect 10508 2404 10514 2612
rect 10564 2572 10570 2780
rect 10604 2572 10610 2780
rect 10646 2612 10656 2792
rect 10708 2612 10718 2792
rect 10756 2780 10802 2792
rect 10468 2392 10514 2404
rect 10550 2392 10560 2572
rect 10612 2392 10622 2572
rect 10660 2404 10666 2612
rect 10700 2404 10706 2612
rect 10756 2572 10762 2780
rect 10796 2572 10802 2780
rect 10838 2612 10848 2792
rect 10900 2612 10910 2792
rect 10948 2780 10994 2792
rect 10660 2392 10706 2404
rect 10742 2392 10752 2572
rect 10804 2392 10814 2572
rect 10852 2404 10858 2612
rect 10892 2404 10898 2612
rect 10948 2572 10954 2780
rect 10988 2572 10994 2780
rect 11030 2612 11040 2792
rect 11092 2612 11102 2792
rect 10852 2392 10898 2404
rect 10934 2392 10944 2572
rect 10996 2392 11006 2572
rect 11044 2404 11050 2612
rect 11084 2404 11090 2612
rect 11044 2392 11090 2404
rect 11132 2360 11212 2824
rect 11834 2612 11844 2792
rect 11896 2612 11906 2792
rect 11944 2780 11990 2792
rect 11848 2404 11854 2612
rect 11888 2404 11894 2612
rect 11944 2572 11950 2780
rect 11984 2572 11990 2780
rect 12026 2612 12036 2792
rect 12088 2612 12098 2792
rect 12136 2780 12182 2792
rect 11848 2392 11894 2404
rect 11930 2392 11940 2572
rect 11992 2392 12002 2572
rect 12040 2404 12046 2612
rect 12080 2404 12086 2612
rect 12136 2572 12142 2780
rect 12176 2572 12182 2780
rect 12218 2612 12228 2792
rect 12280 2612 12290 2792
rect 12328 2780 12374 2792
rect 12040 2392 12086 2404
rect 12122 2392 12132 2572
rect 12184 2392 12194 2572
rect 12232 2404 12238 2612
rect 12272 2404 12278 2612
rect 12328 2572 12334 2780
rect 12368 2572 12374 2780
rect 12410 2612 12420 2792
rect 12472 2612 12482 2792
rect 12232 2392 12278 2404
rect 12314 2392 12324 2572
rect 12376 2392 12386 2572
rect 12424 2404 12430 2612
rect 12464 2404 12470 2612
rect 12424 2392 12470 2404
rect 12512 2360 12592 2824
rect 12874 2612 12884 2792
rect 12936 2612 12946 2792
rect 12984 2780 13030 2792
rect 12888 2404 12894 2612
rect 12928 2404 12934 2612
rect 12984 2572 12990 2780
rect 13024 2572 13030 2780
rect 13066 2612 13076 2792
rect 13128 2612 13138 2792
rect 13176 2780 13222 2792
rect 12888 2392 12934 2404
rect 12970 2392 12980 2572
rect 13032 2392 13042 2572
rect 13080 2404 13086 2612
rect 13120 2404 13126 2612
rect 13176 2572 13182 2780
rect 13216 2572 13222 2780
rect 13258 2612 13268 2792
rect 13320 2612 13330 2792
rect 13368 2780 13414 2792
rect 13080 2392 13126 2404
rect 13162 2392 13172 2572
rect 13224 2392 13234 2572
rect 13272 2404 13278 2612
rect 13312 2404 13318 2612
rect 13368 2572 13374 2780
rect 13408 2572 13414 2780
rect 13450 2612 13460 2792
rect 13512 2612 13522 2792
rect 13272 2392 13318 2404
rect 13354 2392 13364 2572
rect 13416 2392 13426 2572
rect 13464 2404 13470 2612
rect 13504 2404 13510 2612
rect 13464 2392 13510 2404
rect 13552 2360 13632 2824
rect 13914 2612 13924 2792
rect 13976 2612 13986 2792
rect 14024 2780 14070 2792
rect 13928 2404 13934 2612
rect 13968 2404 13974 2612
rect 14024 2572 14030 2780
rect 14064 2572 14070 2780
rect 14106 2612 14116 2792
rect 14168 2612 14178 2792
rect 14216 2780 14262 2792
rect 13928 2392 13974 2404
rect 14010 2392 14020 2572
rect 14072 2392 14082 2572
rect 14120 2404 14126 2612
rect 14160 2404 14166 2612
rect 14216 2572 14222 2780
rect 14256 2572 14262 2780
rect 14298 2612 14308 2792
rect 14360 2612 14370 2792
rect 14408 2780 14454 2792
rect 14120 2392 14166 2404
rect 14202 2392 14212 2572
rect 14264 2392 14274 2572
rect 14312 2404 14318 2612
rect 14352 2404 14358 2612
rect 14408 2572 14414 2780
rect 14448 2572 14454 2780
rect 14490 2612 14500 2792
rect 14552 2612 14562 2792
rect 14312 2392 14358 2404
rect 14394 2392 14404 2572
rect 14456 2392 14466 2572
rect 14504 2404 14510 2612
rect 14544 2404 14550 2612
rect 14504 2392 14550 2404
rect 14592 2360 14672 2824
rect 14954 2612 14964 2792
rect 15016 2612 15026 2792
rect 15064 2780 15110 2792
rect 14968 2404 14974 2612
rect 15008 2404 15014 2612
rect 15064 2572 15070 2780
rect 15104 2572 15110 2780
rect 15146 2612 15156 2792
rect 15208 2612 15218 2792
rect 15256 2780 15302 2792
rect 14968 2392 15014 2404
rect 15050 2392 15060 2572
rect 15112 2392 15122 2572
rect 15160 2404 15166 2612
rect 15200 2404 15206 2612
rect 15256 2572 15262 2780
rect 15296 2572 15302 2780
rect 15338 2612 15348 2792
rect 15400 2612 15410 2792
rect 15448 2780 15494 2792
rect 15160 2392 15206 2404
rect 15242 2392 15252 2572
rect 15304 2392 15314 2572
rect 15352 2404 15358 2612
rect 15392 2404 15398 2612
rect 15448 2572 15454 2780
rect 15488 2572 15494 2780
rect 15530 2612 15540 2792
rect 15592 2612 15602 2792
rect 15352 2392 15398 2404
rect 15434 2392 15444 2572
rect 15496 2392 15506 2572
rect 15544 2404 15550 2612
rect 15584 2404 15590 2612
rect 15544 2392 15590 2404
rect 15632 2360 15712 2824
rect 15994 2612 16004 2792
rect 16056 2612 16066 2792
rect 16104 2780 16150 2792
rect 16008 2404 16014 2612
rect 16048 2404 16054 2612
rect 16104 2572 16110 2780
rect 16144 2572 16150 2780
rect 16186 2612 16196 2792
rect 16248 2612 16258 2792
rect 16296 2780 16342 2792
rect 16008 2392 16054 2404
rect 16090 2392 16100 2572
rect 16152 2392 16162 2572
rect 16200 2404 16206 2612
rect 16240 2404 16246 2612
rect 16296 2572 16302 2780
rect 16336 2572 16342 2780
rect 16378 2612 16388 2792
rect 16440 2612 16450 2792
rect 16488 2780 16534 2792
rect 16200 2392 16246 2404
rect 16282 2392 16292 2572
rect 16344 2392 16354 2572
rect 16392 2404 16398 2612
rect 16432 2404 16438 2612
rect 16488 2572 16494 2780
rect 16528 2572 16534 2780
rect 16570 2612 16580 2792
rect 16632 2612 16642 2792
rect 16392 2392 16438 2404
rect 16474 2392 16484 2572
rect 16536 2392 16546 2572
rect 16584 2404 16590 2612
rect 16624 2404 16630 2612
rect 16584 2392 16630 2404
rect 16672 2360 16752 2824
rect 17034 2612 17044 2792
rect 17096 2612 17106 2792
rect 17144 2780 17190 2792
rect 17048 2404 17054 2612
rect 17088 2404 17094 2612
rect 17144 2572 17150 2780
rect 17184 2572 17190 2780
rect 17226 2612 17236 2792
rect 17288 2612 17298 2792
rect 17336 2780 17382 2792
rect 17048 2392 17094 2404
rect 17130 2392 17140 2572
rect 17192 2392 17202 2572
rect 17240 2404 17246 2612
rect 17280 2404 17286 2612
rect 17336 2572 17342 2780
rect 17376 2572 17382 2780
rect 17418 2612 17428 2792
rect 17480 2612 17490 2792
rect 17528 2780 17574 2792
rect 17240 2392 17286 2404
rect 17322 2392 17332 2572
rect 17384 2392 17394 2572
rect 17432 2404 17438 2612
rect 17472 2404 17478 2612
rect 17528 2572 17534 2780
rect 17568 2572 17574 2780
rect 17610 2612 17620 2792
rect 17672 2612 17682 2792
rect 17432 2392 17478 2404
rect 17514 2392 17524 2572
rect 17576 2392 17586 2572
rect 17624 2404 17630 2612
rect 17664 2404 17670 2612
rect 17624 2392 17670 2404
rect 17712 2360 17792 2824
rect 18074 2612 18084 2792
rect 18136 2612 18146 2792
rect 18184 2780 18230 2792
rect 18088 2404 18094 2612
rect 18128 2404 18134 2612
rect 18184 2572 18190 2780
rect 18224 2572 18230 2780
rect 18266 2612 18276 2792
rect 18328 2612 18338 2792
rect 18376 2780 18422 2792
rect 18088 2392 18134 2404
rect 18170 2392 18180 2572
rect 18232 2392 18242 2572
rect 18280 2404 18286 2612
rect 18320 2404 18326 2612
rect 18376 2572 18382 2780
rect 18416 2572 18422 2780
rect 18458 2612 18468 2792
rect 18520 2612 18530 2792
rect 18568 2780 18614 2792
rect 18280 2392 18326 2404
rect 18362 2392 18372 2572
rect 18424 2392 18434 2572
rect 18472 2404 18478 2612
rect 18512 2404 18518 2612
rect 18568 2572 18574 2780
rect 18608 2572 18614 2780
rect 18650 2612 18660 2792
rect 18712 2612 18722 2792
rect 18472 2392 18518 2404
rect 18554 2392 18564 2572
rect 18616 2392 18626 2572
rect 18664 2404 18670 2612
rect 18704 2404 18710 2612
rect 18664 2392 18710 2404
rect 18752 2360 18832 2824
rect 4320 2354 4972 2360
rect 4320 2340 4378 2354
rect -1484 2194 -832 2200
rect -1484 2160 -1426 2194
rect -1392 2160 -1234 2194
rect -1200 2160 -1042 2194
rect -1008 2160 -832 2194
rect -1484 2086 -832 2160
rect -1484 2052 -1426 2086
rect -1392 2052 -1234 2086
rect -1200 2052 -1042 2086
rect -1008 2052 -832 2086
rect -1484 2044 -832 2052
rect -444 2194 208 2200
rect -444 2160 -386 2194
rect -352 2160 -194 2194
rect -160 2160 -2 2194
rect 32 2160 208 2194
rect -444 2086 208 2160
rect -444 2052 -386 2086
rect -352 2052 -194 2086
rect -160 2052 -2 2086
rect 32 2052 208 2086
rect -444 2044 208 2052
rect 596 2194 1248 2200
rect 596 2160 654 2194
rect 688 2160 846 2194
rect 880 2160 1038 2194
rect 1072 2160 1248 2194
rect 596 2086 1248 2160
rect 596 2052 654 2086
rect 688 2052 846 2086
rect 880 2052 1038 2086
rect 1072 2052 1248 2086
rect 596 2044 1248 2052
rect 1636 2194 2288 2200
rect 1636 2160 1694 2194
rect 1728 2160 1886 2194
rect 1920 2160 2078 2194
rect 2112 2160 2288 2194
rect 1636 2086 2288 2160
rect 1636 2052 1694 2086
rect 1728 2052 1886 2086
rect 1920 2052 2078 2086
rect 2112 2052 2288 2086
rect 1636 2044 2288 2052
rect 2676 2194 3328 2200
rect 2676 2160 2734 2194
rect 2768 2160 2926 2194
rect 2960 2160 3118 2194
rect 3152 2160 3328 2194
rect 2676 2086 3328 2160
rect 2676 2052 2734 2086
rect 2768 2052 2926 2086
rect 2960 2052 3118 2086
rect 3152 2052 3328 2086
rect 2676 2044 3328 2052
rect -1576 2002 -1530 2014
rect -1576 1796 -1570 2002
rect -1536 1796 -1530 2002
rect -1494 1836 -1484 2016
rect -1432 1836 -1422 2016
rect -1384 2002 -1338 2014
rect -1590 1616 -1580 1796
rect -1528 1616 -1518 1796
rect -1480 1626 -1474 1836
rect -1440 1626 -1434 1836
rect -1384 1796 -1378 2002
rect -1344 1796 -1338 2002
rect -1302 1836 -1292 2016
rect -1240 1836 -1230 2016
rect -1192 2002 -1146 2014
rect -1576 1614 -1530 1616
rect -1480 1614 -1434 1626
rect -1398 1616 -1388 1796
rect -1336 1616 -1326 1796
rect -1288 1626 -1282 1836
rect -1248 1626 -1242 1836
rect -1192 1796 -1186 2002
rect -1152 1796 -1146 2002
rect -1110 1836 -1100 2016
rect -1048 1836 -1038 2016
rect -1000 2002 -954 2014
rect -1384 1614 -1338 1616
rect -1288 1614 -1242 1626
rect -1206 1616 -1196 1796
rect -1144 1616 -1134 1796
rect -1096 1626 -1090 1836
rect -1056 1626 -1050 1836
rect -1000 1796 -994 2002
rect -960 1796 -954 2002
rect -1192 1614 -1146 1616
rect -1096 1614 -1050 1626
rect -1014 1616 -1004 1796
rect -952 1616 -942 1796
rect -1000 1614 -954 1616
rect -1534 1580 -1476 1582
rect -1342 1580 -1284 1582
rect -1150 1580 -1092 1582
rect -912 1580 -832 2044
rect -536 2002 -490 2014
rect -536 1796 -530 2002
rect -496 1796 -490 2002
rect -454 1836 -444 2016
rect -392 1836 -382 2016
rect -344 2002 -298 2014
rect -550 1616 -540 1796
rect -488 1616 -478 1796
rect -440 1626 -434 1836
rect -400 1626 -394 1836
rect -344 1796 -338 2002
rect -304 1796 -298 2002
rect -262 1836 -252 2016
rect -200 1836 -190 2016
rect -152 2002 -106 2014
rect -536 1614 -490 1616
rect -440 1614 -394 1626
rect -358 1616 -348 1796
rect -296 1616 -286 1796
rect -248 1626 -242 1836
rect -208 1626 -202 1836
rect -152 1796 -146 2002
rect -112 1796 -106 2002
rect -70 1836 -60 2016
rect -8 1836 2 2016
rect 40 2002 86 2014
rect -344 1614 -298 1616
rect -248 1614 -202 1626
rect -166 1616 -156 1796
rect -104 1616 -94 1796
rect -56 1626 -50 1836
rect -16 1626 -10 1836
rect 40 1796 46 2002
rect 80 1796 86 2002
rect -152 1614 -106 1616
rect -56 1614 -10 1626
rect 26 1616 36 1796
rect 88 1616 98 1796
rect 40 1614 86 1616
rect -494 1580 -436 1582
rect -302 1580 -244 1582
rect -110 1580 -52 1582
rect 128 1580 208 2044
rect 504 2002 550 2014
rect 504 1796 510 2002
rect 544 1796 550 2002
rect 586 1836 596 2016
rect 648 1836 658 2016
rect 696 2002 742 2014
rect 490 1616 500 1796
rect 552 1616 562 1796
rect 600 1626 606 1836
rect 640 1626 646 1836
rect 696 1796 702 2002
rect 736 1796 742 2002
rect 778 1836 788 2016
rect 840 1836 850 2016
rect 888 2002 934 2014
rect 504 1614 550 1616
rect 600 1614 646 1626
rect 682 1616 692 1796
rect 744 1616 754 1796
rect 792 1626 798 1836
rect 832 1626 838 1836
rect 888 1796 894 2002
rect 928 1796 934 2002
rect 970 1836 980 2016
rect 1032 1836 1042 2016
rect 1080 2002 1126 2014
rect 696 1614 742 1616
rect 792 1614 838 1626
rect 874 1616 884 1796
rect 936 1616 946 1796
rect 984 1626 990 1836
rect 1024 1626 1030 1836
rect 1080 1796 1086 2002
rect 1120 1796 1126 2002
rect 888 1614 934 1616
rect 984 1614 1030 1626
rect 1066 1616 1076 1796
rect 1128 1616 1138 1796
rect 1080 1614 1126 1616
rect 546 1580 604 1582
rect 738 1580 796 1582
rect 930 1580 988 1582
rect 1168 1580 1248 2044
rect 1544 2002 1590 2014
rect 1544 1796 1550 2002
rect 1584 1796 1590 2002
rect 1626 1836 1636 2016
rect 1688 1836 1698 2016
rect 1736 2002 1782 2014
rect 1530 1616 1540 1796
rect 1592 1616 1602 1796
rect 1640 1626 1646 1836
rect 1680 1626 1686 1836
rect 1736 1796 1742 2002
rect 1776 1796 1782 2002
rect 1818 1836 1828 2016
rect 1880 1836 1890 2016
rect 1928 2002 1974 2014
rect 1544 1614 1590 1616
rect 1640 1614 1686 1626
rect 1722 1616 1732 1796
rect 1784 1616 1794 1796
rect 1832 1626 1838 1836
rect 1872 1626 1878 1836
rect 1928 1796 1934 2002
rect 1968 1796 1974 2002
rect 2010 1836 2020 2016
rect 2072 1836 2082 2016
rect 2120 2002 2166 2014
rect 1736 1614 1782 1616
rect 1832 1614 1878 1626
rect 1914 1616 1924 1796
rect 1976 1616 1986 1796
rect 2024 1626 2030 1836
rect 2064 1626 2070 1836
rect 2120 1796 2126 2002
rect 2160 1796 2166 2002
rect 1928 1614 1974 1616
rect 2024 1614 2070 1626
rect 2106 1616 2116 1796
rect 2168 1616 2178 1796
rect 2120 1614 2166 1616
rect 1586 1580 1644 1582
rect 1778 1580 1836 1582
rect 1970 1580 2028 1582
rect 2208 1580 2288 2044
rect 2584 2002 2630 2014
rect 2584 1796 2590 2002
rect 2624 1796 2630 2002
rect 2666 1836 2676 2016
rect 2728 1836 2738 2016
rect 2776 2002 2822 2014
rect 2570 1616 2580 1796
rect 2632 1616 2642 1796
rect 2680 1626 2686 1836
rect 2720 1626 2726 1836
rect 2776 1796 2782 2002
rect 2816 1796 2822 2002
rect 2858 1836 2868 2016
rect 2920 1836 2930 2016
rect 2968 2002 3014 2014
rect 2584 1614 2630 1616
rect 2680 1614 2726 1626
rect 2762 1616 2772 1796
rect 2824 1616 2834 1796
rect 2872 1626 2878 1836
rect 2912 1626 2918 1836
rect 2968 1796 2974 2002
rect 3008 1796 3014 2002
rect 3050 1836 3060 2016
rect 3112 1836 3122 2016
rect 3160 2002 3206 2014
rect 2776 1614 2822 1616
rect 2872 1614 2918 1626
rect 2954 1616 2964 1796
rect 3016 1616 3026 1796
rect 3064 1626 3070 1836
rect 3104 1626 3110 1836
rect 3160 1796 3166 2002
rect 3200 1796 3206 2002
rect 2968 1614 3014 1616
rect 3064 1614 3110 1626
rect 3146 1616 3156 1796
rect 3208 1616 3218 1796
rect 3160 1614 3206 1616
rect 2626 1580 2684 1582
rect 2818 1580 2876 1582
rect 3010 1580 3068 1582
rect 3248 1580 3328 2044
rect -1540 1576 -832 1580
rect -1540 1542 -1522 1576
rect -1488 1542 -1330 1576
rect -1296 1542 -1138 1576
rect -1104 1542 -832 1576
rect -1540 1484 -832 1542
rect -500 1576 208 1580
rect -500 1542 -482 1576
rect -448 1542 -290 1576
rect -256 1542 -98 1576
rect -64 1542 208 1576
rect -500 1484 208 1542
rect 540 1576 1248 1580
rect 540 1542 558 1576
rect 592 1542 750 1576
rect 784 1542 942 1576
rect 976 1542 1248 1576
rect 540 1484 1248 1542
rect 1580 1576 2288 1580
rect 1580 1542 1598 1576
rect 1632 1542 1790 1576
rect 1824 1542 1982 1576
rect 2016 1542 2288 1576
rect 1580 1484 2288 1542
rect 2620 1576 3328 1580
rect 2620 1542 2638 1576
rect 2672 1542 2830 1576
rect 2864 1542 3022 1576
rect 3056 1542 3328 1576
rect 2620 1484 3328 1542
rect 4000 2320 4378 2340
rect 4412 2320 4570 2354
rect 4604 2320 4762 2354
rect 4796 2340 4972 2354
rect 5360 2354 6012 2360
rect 5360 2340 5418 2354
rect 4796 2320 5418 2340
rect 5452 2320 5610 2354
rect 5644 2320 5802 2354
rect 5836 2340 6012 2354
rect 6400 2354 7052 2360
rect 6400 2340 6458 2354
rect 5836 2320 6458 2340
rect 6492 2320 6650 2354
rect 6684 2320 6842 2354
rect 6876 2340 7052 2354
rect 7440 2354 8092 2360
rect 7440 2340 7498 2354
rect 6876 2320 7498 2340
rect 7532 2320 7690 2354
rect 7724 2320 7882 2354
rect 7916 2340 8092 2354
rect 8480 2354 9132 2360
rect 8480 2340 8538 2354
rect 7916 2320 8538 2340
rect 8572 2320 8730 2354
rect 8764 2320 8922 2354
rect 8956 2340 9132 2354
rect 9520 2354 10172 2360
rect 9520 2340 9578 2354
rect 8956 2320 9578 2340
rect 9612 2320 9770 2354
rect 9804 2320 9962 2354
rect 9996 2340 10172 2354
rect 10560 2354 11212 2360
rect 10560 2340 10618 2354
rect 9996 2320 10618 2340
rect 10652 2320 10810 2354
rect 10844 2320 11002 2354
rect 11036 2340 11212 2354
rect 11940 2354 12592 2360
rect 11940 2340 11998 2354
rect 11036 2320 11998 2340
rect 12032 2320 12190 2354
rect 12224 2320 12382 2354
rect 12416 2340 12592 2354
rect 12980 2354 13632 2360
rect 12980 2340 13038 2354
rect 12416 2320 13038 2340
rect 13072 2320 13230 2354
rect 13264 2320 13422 2354
rect 13456 2340 13632 2354
rect 14020 2354 14672 2360
rect 14020 2340 14078 2354
rect 13456 2320 14078 2340
rect 14112 2320 14270 2354
rect 14304 2320 14462 2354
rect 14496 2340 14672 2354
rect 15060 2354 15712 2360
rect 15060 2340 15118 2354
rect 14496 2320 15118 2340
rect 15152 2320 15310 2354
rect 15344 2320 15502 2354
rect 15536 2340 15712 2354
rect 16100 2354 16752 2360
rect 16100 2340 16158 2354
rect 15536 2320 16158 2340
rect 16192 2320 16350 2354
rect 16384 2320 16542 2354
rect 16576 2340 16752 2354
rect 17140 2354 17792 2360
rect 17140 2340 17198 2354
rect 16576 2320 17198 2340
rect 17232 2320 17390 2354
rect 17424 2320 17582 2354
rect 17616 2340 17792 2354
rect 18180 2354 18832 2360
rect 18180 2340 18238 2354
rect 17616 2320 18238 2340
rect 18272 2320 18430 2354
rect 18464 2320 18622 2354
rect 18656 2320 18832 2354
rect 4000 2246 18832 2320
rect 4000 2224 4378 2246
rect -968 1308 -884 1484
rect 72 1308 156 1484
rect 1112 1308 1196 1484
rect 2152 1308 2236 1484
rect 3192 1308 3276 1484
rect -1532 1282 -716 1308
rect -1532 1248 -1511 1282
rect -1477 1248 -1393 1282
rect -1359 1248 -1275 1282
rect -1241 1248 -1157 1282
rect -1123 1248 -1039 1282
rect -1005 1248 -921 1282
rect -887 1248 -716 1282
rect -1532 1240 -716 1248
rect -492 1282 324 1308
rect -492 1248 -471 1282
rect -437 1248 -353 1282
rect -319 1248 -235 1282
rect -201 1248 -117 1282
rect -83 1248 1 1282
rect 35 1248 119 1282
rect 153 1248 324 1282
rect -492 1240 324 1248
rect 548 1282 1364 1308
rect 548 1248 569 1282
rect 603 1248 687 1282
rect 721 1248 805 1282
rect 839 1248 923 1282
rect 957 1248 1041 1282
rect 1075 1248 1159 1282
rect 1193 1248 1364 1282
rect 548 1240 1364 1248
rect 1588 1282 2404 1308
rect 1588 1248 1609 1282
rect 1643 1248 1727 1282
rect 1761 1248 1845 1282
rect 1879 1248 1963 1282
rect 1997 1248 2081 1282
rect 2115 1248 2199 1282
rect 2233 1248 2404 1282
rect 1588 1240 2404 1248
rect 2628 1282 3444 1308
rect 2628 1248 2649 1282
rect 2683 1248 2767 1282
rect 2801 1248 2885 1282
rect 2919 1248 3003 1282
rect 3037 1248 3121 1282
rect 3155 1248 3239 1282
rect 3273 1248 3444 1282
rect 2628 1240 3444 1248
rect -1576 1198 -1530 1210
rect -1576 988 -1570 1198
rect -1536 988 -1530 1198
rect -1470 1032 -1460 1212
rect -1408 1032 -1398 1212
rect -1340 1198 -1294 1210
rect -1590 808 -1580 988
rect -1528 808 -1518 988
rect -1458 822 -1452 1032
rect -1418 822 -1412 1032
rect -1340 988 -1334 1198
rect -1300 988 -1294 1198
rect -1234 1032 -1224 1212
rect -1172 1032 -1162 1212
rect -1104 1198 -1058 1210
rect -1458 810 -1412 822
rect -1354 808 -1344 988
rect -1292 808 -1282 988
rect -1222 822 -1216 1032
rect -1182 822 -1176 1032
rect -1104 988 -1098 1198
rect -1064 988 -1058 1198
rect -998 1032 -988 1212
rect -936 1032 -926 1212
rect -868 1198 -822 1210
rect -1222 810 -1176 822
rect -1118 808 -1108 988
rect -1056 808 -1046 988
rect -986 822 -980 1032
rect -946 822 -940 1032
rect -868 988 -862 1198
rect -828 988 -822 1198
rect -986 810 -940 822
rect -882 808 -872 988
rect -820 808 -810 988
rect -780 780 -716 1240
rect -536 1198 -490 1210
rect -536 988 -530 1198
rect -496 988 -490 1198
rect -430 1032 -420 1212
rect -368 1032 -358 1212
rect -300 1198 -254 1210
rect -550 808 -540 988
rect -488 808 -478 988
rect -418 822 -412 1032
rect -378 822 -372 1032
rect -300 988 -294 1198
rect -260 988 -254 1198
rect -194 1032 -184 1212
rect -132 1032 -122 1212
rect -64 1198 -18 1210
rect -418 810 -372 822
rect -314 808 -304 988
rect -252 808 -242 988
rect -182 822 -176 1032
rect -142 822 -136 1032
rect -64 988 -58 1198
rect -24 988 -18 1198
rect 42 1032 52 1212
rect 104 1032 114 1212
rect 172 1198 218 1210
rect -182 810 -136 822
rect -78 808 -68 988
rect -16 808 -6 988
rect 54 822 60 1032
rect 94 822 100 1032
rect 172 988 178 1198
rect 212 988 218 1198
rect 54 810 100 822
rect 158 808 168 988
rect 220 808 230 988
rect 260 780 324 1240
rect 504 1198 550 1210
rect 504 988 510 1198
rect 544 988 550 1198
rect 610 1032 620 1212
rect 672 1032 682 1212
rect 740 1198 786 1210
rect 490 808 500 988
rect 552 808 562 988
rect 622 822 628 1032
rect 662 822 668 1032
rect 740 988 746 1198
rect 780 988 786 1198
rect 846 1032 856 1212
rect 908 1032 918 1212
rect 976 1198 1022 1210
rect 622 810 668 822
rect 726 808 736 988
rect 788 808 798 988
rect 858 822 864 1032
rect 898 822 904 1032
rect 976 988 982 1198
rect 1016 988 1022 1198
rect 1082 1032 1092 1212
rect 1144 1032 1154 1212
rect 1212 1198 1258 1210
rect 858 810 904 822
rect 962 808 972 988
rect 1024 808 1034 988
rect 1094 822 1100 1032
rect 1134 822 1140 1032
rect 1212 988 1218 1198
rect 1252 988 1258 1198
rect 1094 810 1140 822
rect 1198 808 1208 988
rect 1260 808 1270 988
rect 1300 780 1364 1240
rect 1544 1198 1590 1210
rect 1544 988 1550 1198
rect 1584 988 1590 1198
rect 1650 1032 1660 1212
rect 1712 1032 1722 1212
rect 1780 1198 1826 1210
rect 1530 808 1540 988
rect 1592 808 1602 988
rect 1662 822 1668 1032
rect 1702 822 1708 1032
rect 1780 988 1786 1198
rect 1820 988 1826 1198
rect 1886 1032 1896 1212
rect 1948 1032 1958 1212
rect 2016 1198 2062 1210
rect 1662 810 1708 822
rect 1766 808 1776 988
rect 1828 808 1838 988
rect 1898 822 1904 1032
rect 1938 822 1944 1032
rect 2016 988 2022 1198
rect 2056 988 2062 1198
rect 2122 1032 2132 1212
rect 2184 1032 2194 1212
rect 2252 1198 2298 1210
rect 1898 810 1944 822
rect 2002 808 2012 988
rect 2064 808 2074 988
rect 2134 822 2140 1032
rect 2174 822 2180 1032
rect 2252 988 2258 1198
rect 2292 988 2298 1198
rect 2134 810 2180 822
rect 2238 808 2248 988
rect 2300 808 2310 988
rect 2340 780 2404 1240
rect 2584 1198 2630 1210
rect 2584 988 2590 1198
rect 2624 988 2630 1198
rect 2690 1032 2700 1212
rect 2752 1032 2762 1212
rect 2820 1198 2866 1210
rect 2570 808 2580 988
rect 2632 808 2642 988
rect 2702 822 2708 1032
rect 2742 822 2748 1032
rect 2820 988 2826 1198
rect 2860 988 2866 1198
rect 2926 1032 2936 1212
rect 2988 1032 2998 1212
rect 3056 1198 3102 1210
rect 2702 810 2748 822
rect 2806 808 2816 988
rect 2868 808 2878 988
rect 2938 822 2944 1032
rect 2978 822 2984 1032
rect 3056 988 3062 1198
rect 3096 988 3102 1198
rect 3162 1032 3172 1212
rect 3224 1032 3234 1212
rect 3292 1198 3338 1210
rect 2938 810 2984 822
rect 3042 808 3052 988
rect 3104 808 3114 988
rect 3174 822 3180 1032
rect 3214 822 3220 1032
rect 3292 988 3298 1198
rect 3332 988 3338 1198
rect 3174 810 3220 822
rect 3278 808 3288 988
rect 3340 808 3350 988
rect 3380 780 3444 1240
rect 4000 780 4156 2224
rect 4320 2212 4378 2224
rect 4412 2212 4570 2246
rect 4604 2212 4762 2246
rect 4796 2224 5418 2246
rect 4796 2212 4972 2224
rect 4320 2204 4972 2212
rect 5360 2212 5418 2224
rect 5452 2212 5610 2246
rect 5644 2212 5802 2246
rect 5836 2224 6458 2246
rect 5836 2212 6012 2224
rect 5360 2204 6012 2212
rect 6400 2212 6458 2224
rect 6492 2212 6650 2246
rect 6684 2212 6842 2246
rect 6876 2224 7498 2246
rect 6876 2212 7052 2224
rect 6400 2204 7052 2212
rect 7440 2212 7498 2224
rect 7532 2212 7690 2246
rect 7724 2212 7882 2246
rect 7916 2224 8538 2246
rect 7916 2212 8092 2224
rect 7440 2204 8092 2212
rect 8480 2212 8538 2224
rect 8572 2212 8730 2246
rect 8764 2212 8922 2246
rect 8956 2224 9578 2246
rect 8956 2212 9132 2224
rect 8480 2204 9132 2212
rect 9520 2212 9578 2224
rect 9612 2212 9770 2246
rect 9804 2212 9962 2246
rect 9996 2224 10618 2246
rect 9996 2212 10172 2224
rect 9520 2204 10172 2212
rect 10560 2212 10618 2224
rect 10652 2212 10810 2246
rect 10844 2212 11002 2246
rect 11036 2224 11998 2246
rect 11036 2212 11212 2224
rect 10560 2204 11212 2212
rect 4228 2162 4274 2174
rect 4228 1956 4234 2162
rect 4268 1956 4274 2162
rect 4310 1996 4320 2176
rect 4372 1996 4382 2176
rect 4420 2162 4466 2174
rect 4214 1776 4224 1956
rect 4276 1776 4286 1956
rect 4324 1786 4330 1996
rect 4364 1786 4370 1996
rect 4420 1956 4426 2162
rect 4460 1956 4466 2162
rect 4502 1996 4512 2176
rect 4564 1996 4574 2176
rect 4612 2162 4658 2174
rect 4228 1774 4274 1776
rect 4324 1774 4370 1786
rect 4406 1776 4416 1956
rect 4468 1776 4478 1956
rect 4516 1786 4522 1996
rect 4556 1786 4562 1996
rect 4612 1956 4618 2162
rect 4652 1956 4658 2162
rect 4694 1996 4704 2176
rect 4756 1996 4766 2176
rect 4804 2162 4850 2174
rect 4420 1774 4466 1776
rect 4516 1774 4562 1786
rect 4598 1776 4608 1956
rect 4660 1776 4670 1956
rect 4708 1786 4714 1996
rect 4748 1786 4754 1996
rect 4804 1956 4810 2162
rect 4844 1956 4850 2162
rect 4612 1774 4658 1776
rect 4708 1774 4754 1786
rect 4790 1776 4800 1956
rect 4852 1776 4862 1956
rect 4804 1774 4850 1776
rect 4270 1740 4328 1742
rect 4462 1740 4520 1742
rect 4654 1740 4712 1742
rect 4892 1740 4972 2204
rect 5268 2162 5314 2174
rect 5268 1956 5274 2162
rect 5308 1956 5314 2162
rect 5350 1996 5360 2176
rect 5412 1996 5422 2176
rect 5460 2162 5506 2174
rect 5254 1776 5264 1956
rect 5316 1776 5326 1956
rect 5364 1786 5370 1996
rect 5404 1786 5410 1996
rect 5460 1956 5466 2162
rect 5500 1956 5506 2162
rect 5542 1996 5552 2176
rect 5604 1996 5614 2176
rect 5652 2162 5698 2174
rect 5268 1774 5314 1776
rect 5364 1774 5410 1786
rect 5446 1776 5456 1956
rect 5508 1776 5518 1956
rect 5556 1786 5562 1996
rect 5596 1786 5602 1996
rect 5652 1956 5658 2162
rect 5692 1956 5698 2162
rect 5734 1996 5744 2176
rect 5796 1996 5806 2176
rect 5844 2162 5890 2174
rect 5460 1774 5506 1776
rect 5556 1774 5602 1786
rect 5638 1776 5648 1956
rect 5700 1776 5710 1956
rect 5748 1786 5754 1996
rect 5788 1786 5794 1996
rect 5844 1956 5850 2162
rect 5884 1956 5890 2162
rect 5652 1774 5698 1776
rect 5748 1774 5794 1786
rect 5830 1776 5840 1956
rect 5892 1776 5902 1956
rect 5844 1774 5890 1776
rect 5310 1740 5368 1742
rect 5502 1740 5560 1742
rect 5694 1740 5752 1742
rect 5932 1740 6012 2204
rect 6308 2162 6354 2174
rect 6308 1956 6314 2162
rect 6348 1956 6354 2162
rect 6390 1996 6400 2176
rect 6452 1996 6462 2176
rect 6500 2162 6546 2174
rect 6294 1776 6304 1956
rect 6356 1776 6366 1956
rect 6404 1786 6410 1996
rect 6444 1786 6450 1996
rect 6500 1956 6506 2162
rect 6540 1956 6546 2162
rect 6582 1996 6592 2176
rect 6644 1996 6654 2176
rect 6692 2162 6738 2174
rect 6308 1774 6354 1776
rect 6404 1774 6450 1786
rect 6486 1776 6496 1956
rect 6548 1776 6558 1956
rect 6596 1786 6602 1996
rect 6636 1786 6642 1996
rect 6692 1956 6698 2162
rect 6732 1956 6738 2162
rect 6774 1996 6784 2176
rect 6836 1996 6846 2176
rect 6884 2162 6930 2174
rect 6500 1774 6546 1776
rect 6596 1774 6642 1786
rect 6678 1776 6688 1956
rect 6740 1776 6750 1956
rect 6788 1786 6794 1996
rect 6828 1786 6834 1996
rect 6884 1956 6890 2162
rect 6924 1956 6930 2162
rect 6692 1774 6738 1776
rect 6788 1774 6834 1786
rect 6870 1776 6880 1956
rect 6932 1776 6942 1956
rect 6884 1774 6930 1776
rect 6350 1740 6408 1742
rect 6542 1740 6600 1742
rect 6734 1740 6792 1742
rect 6972 1740 7052 2204
rect 7348 2162 7394 2174
rect 7348 1956 7354 2162
rect 7388 1956 7394 2162
rect 7430 1996 7440 2176
rect 7492 1996 7502 2176
rect 7540 2162 7586 2174
rect 7334 1776 7344 1956
rect 7396 1776 7406 1956
rect 7444 1786 7450 1996
rect 7484 1786 7490 1996
rect 7540 1956 7546 2162
rect 7580 1956 7586 2162
rect 7622 1996 7632 2176
rect 7684 1996 7694 2176
rect 7732 2162 7778 2174
rect 7348 1774 7394 1776
rect 7444 1774 7490 1786
rect 7526 1776 7536 1956
rect 7588 1776 7598 1956
rect 7636 1786 7642 1996
rect 7676 1786 7682 1996
rect 7732 1956 7738 2162
rect 7772 1956 7778 2162
rect 7814 1996 7824 2176
rect 7876 1996 7886 2176
rect 7924 2162 7970 2174
rect 7540 1774 7586 1776
rect 7636 1774 7682 1786
rect 7718 1776 7728 1956
rect 7780 1776 7790 1956
rect 7828 1786 7834 1996
rect 7868 1786 7874 1996
rect 7924 1956 7930 2162
rect 7964 1956 7970 2162
rect 7732 1774 7778 1776
rect 7828 1774 7874 1786
rect 7910 1776 7920 1956
rect 7972 1776 7982 1956
rect 7924 1774 7970 1776
rect 7390 1740 7448 1742
rect 7582 1740 7640 1742
rect 7774 1740 7832 1742
rect 8012 1740 8092 2204
rect 8388 2162 8434 2174
rect 8388 1956 8394 2162
rect 8428 1956 8434 2162
rect 8470 1996 8480 2176
rect 8532 1996 8542 2176
rect 8580 2162 8626 2174
rect 8374 1776 8384 1956
rect 8436 1776 8446 1956
rect 8484 1786 8490 1996
rect 8524 1786 8530 1996
rect 8580 1956 8586 2162
rect 8620 1956 8626 2162
rect 8662 1996 8672 2176
rect 8724 1996 8734 2176
rect 8772 2162 8818 2174
rect 8388 1774 8434 1776
rect 8484 1774 8530 1786
rect 8566 1776 8576 1956
rect 8628 1776 8638 1956
rect 8676 1786 8682 1996
rect 8716 1786 8722 1996
rect 8772 1956 8778 2162
rect 8812 1956 8818 2162
rect 8854 1996 8864 2176
rect 8916 1996 8926 2176
rect 8964 2162 9010 2174
rect 8580 1774 8626 1776
rect 8676 1774 8722 1786
rect 8758 1776 8768 1956
rect 8820 1776 8830 1956
rect 8868 1786 8874 1996
rect 8908 1786 8914 1996
rect 8964 1956 8970 2162
rect 9004 1956 9010 2162
rect 8772 1774 8818 1776
rect 8868 1774 8914 1786
rect 8950 1776 8960 1956
rect 9012 1776 9022 1956
rect 8964 1774 9010 1776
rect 8430 1740 8488 1742
rect 8622 1740 8680 1742
rect 8814 1740 8872 1742
rect 9052 1740 9132 2204
rect 9428 2162 9474 2174
rect 9428 1956 9434 2162
rect 9468 1956 9474 2162
rect 9510 1996 9520 2176
rect 9572 1996 9582 2176
rect 9620 2162 9666 2174
rect 9414 1776 9424 1956
rect 9476 1776 9486 1956
rect 9524 1786 9530 1996
rect 9564 1786 9570 1996
rect 9620 1956 9626 2162
rect 9660 1956 9666 2162
rect 9702 1996 9712 2176
rect 9764 1996 9774 2176
rect 9812 2162 9858 2174
rect 9428 1774 9474 1776
rect 9524 1774 9570 1786
rect 9606 1776 9616 1956
rect 9668 1776 9678 1956
rect 9716 1786 9722 1996
rect 9756 1786 9762 1996
rect 9812 1956 9818 2162
rect 9852 1956 9858 2162
rect 9894 1996 9904 2176
rect 9956 1996 9966 2176
rect 10004 2162 10050 2174
rect 9620 1774 9666 1776
rect 9716 1774 9762 1786
rect 9798 1776 9808 1956
rect 9860 1776 9870 1956
rect 9908 1786 9914 1996
rect 9948 1786 9954 1996
rect 10004 1956 10010 2162
rect 10044 1956 10050 2162
rect 9812 1774 9858 1776
rect 9908 1774 9954 1786
rect 9990 1776 10000 1956
rect 10052 1776 10062 1956
rect 10004 1774 10050 1776
rect 9470 1740 9528 1742
rect 9662 1740 9720 1742
rect 9854 1740 9912 1742
rect 10092 1740 10172 2204
rect 10468 2162 10514 2174
rect 10468 1956 10474 2162
rect 10508 1956 10514 2162
rect 10550 1996 10560 2176
rect 10612 1996 10622 2176
rect 10660 2162 10706 2174
rect 10454 1776 10464 1956
rect 10516 1776 10526 1956
rect 10564 1786 10570 1996
rect 10604 1786 10610 1996
rect 10660 1956 10666 2162
rect 10700 1956 10706 2162
rect 10742 1996 10752 2176
rect 10804 1996 10814 2176
rect 10852 2162 10898 2174
rect 10468 1774 10514 1776
rect 10564 1774 10610 1786
rect 10646 1776 10656 1956
rect 10708 1776 10718 1956
rect 10756 1786 10762 1996
rect 10796 1786 10802 1996
rect 10852 1956 10858 2162
rect 10892 1956 10898 2162
rect 10934 1996 10944 2176
rect 10996 1996 11006 2176
rect 11044 2162 11090 2174
rect 10660 1774 10706 1776
rect 10756 1774 10802 1786
rect 10838 1776 10848 1956
rect 10900 1776 10910 1956
rect 10948 1786 10954 1996
rect 10988 1786 10994 1996
rect 11044 1956 11050 2162
rect 11084 1956 11090 2162
rect 10852 1774 10898 1776
rect 10948 1774 10994 1786
rect 11030 1776 11040 1956
rect 11092 1776 11102 1956
rect 11044 1774 11090 1776
rect 10510 1740 10568 1742
rect 10702 1740 10760 1742
rect 10894 1740 10952 1742
rect 11132 1740 11212 2204
rect 4264 1736 4972 1740
rect 4264 1702 4282 1736
rect 4316 1702 4474 1736
rect 4508 1702 4666 1736
rect 4700 1702 4972 1736
rect 4264 1644 4972 1702
rect 5304 1736 6012 1740
rect 5304 1702 5322 1736
rect 5356 1702 5514 1736
rect 5548 1702 5706 1736
rect 5740 1702 6012 1736
rect 5304 1644 6012 1702
rect 6344 1736 7052 1740
rect 6344 1702 6362 1736
rect 6396 1702 6554 1736
rect 6588 1702 6746 1736
rect 6780 1702 7052 1736
rect 6344 1644 7052 1702
rect 7384 1736 8092 1740
rect 7384 1702 7402 1736
rect 7436 1702 7594 1736
rect 7628 1702 7786 1736
rect 7820 1702 8092 1736
rect 7384 1644 8092 1702
rect 8424 1736 9132 1740
rect 8424 1702 8442 1736
rect 8476 1702 8634 1736
rect 8668 1702 8826 1736
rect 8860 1702 9132 1736
rect 8424 1644 9132 1702
rect 9464 1736 10172 1740
rect 9464 1702 9482 1736
rect 9516 1702 9674 1736
rect 9708 1702 9866 1736
rect 9900 1702 10172 1736
rect 9464 1644 10172 1702
rect 10504 1736 11212 1740
rect 10504 1702 10522 1736
rect 10556 1702 10714 1736
rect 10748 1702 10906 1736
rect 10940 1702 11212 1736
rect 10504 1644 11212 1702
rect 4836 1468 4920 1644
rect 5876 1468 5960 1644
rect 6916 1468 7000 1644
rect 7956 1468 8040 1644
rect 8996 1468 9080 1644
rect 10036 1468 10120 1644
rect 11076 1468 11160 1644
rect 4272 1442 5088 1468
rect 4272 1408 4293 1442
rect 4327 1408 4411 1442
rect 4445 1408 4529 1442
rect 4563 1408 4647 1442
rect 4681 1408 4765 1442
rect 4799 1408 4883 1442
rect 4917 1408 5088 1442
rect 4272 1400 5088 1408
rect 5312 1442 6128 1468
rect 5312 1408 5333 1442
rect 5367 1408 5451 1442
rect 5485 1408 5569 1442
rect 5603 1408 5687 1442
rect 5721 1408 5805 1442
rect 5839 1408 5923 1442
rect 5957 1408 6128 1442
rect 5312 1400 6128 1408
rect 6352 1442 7168 1468
rect 6352 1408 6373 1442
rect 6407 1408 6491 1442
rect 6525 1408 6609 1442
rect 6643 1408 6727 1442
rect 6761 1408 6845 1442
rect 6879 1408 6963 1442
rect 6997 1408 7168 1442
rect 6352 1400 7168 1408
rect 7392 1442 8208 1468
rect 7392 1408 7413 1442
rect 7447 1408 7531 1442
rect 7565 1408 7649 1442
rect 7683 1408 7767 1442
rect 7801 1408 7885 1442
rect 7919 1408 8003 1442
rect 8037 1408 8208 1442
rect 7392 1400 8208 1408
rect 8432 1442 9248 1468
rect 8432 1408 8453 1442
rect 8487 1408 8571 1442
rect 8605 1408 8689 1442
rect 8723 1408 8807 1442
rect 8841 1408 8925 1442
rect 8959 1408 9043 1442
rect 9077 1408 9248 1442
rect 8432 1400 9248 1408
rect 9472 1442 10288 1468
rect 9472 1408 9493 1442
rect 9527 1408 9611 1442
rect 9645 1408 9729 1442
rect 9763 1408 9847 1442
rect 9881 1408 9965 1442
rect 9999 1408 10083 1442
rect 10117 1408 10288 1442
rect 9472 1400 10288 1408
rect 10512 1442 11328 1468
rect 10512 1408 10533 1442
rect 10567 1408 10651 1442
rect 10685 1408 10769 1442
rect 10803 1408 10887 1442
rect 10921 1408 11005 1442
rect 11039 1408 11123 1442
rect 11157 1408 11328 1442
rect 10512 1400 11328 1408
rect 4228 1358 4274 1370
rect 4228 1148 4234 1358
rect 4268 1148 4274 1358
rect 4334 1192 4344 1372
rect 4396 1192 4406 1372
rect 4464 1358 4510 1370
rect 4214 968 4224 1148
rect 4276 968 4286 1148
rect 4346 982 4352 1192
rect 4386 982 4392 1192
rect 4464 1148 4470 1358
rect 4504 1148 4510 1358
rect 4570 1192 4580 1372
rect 4632 1192 4642 1372
rect 4700 1358 4746 1370
rect 4346 970 4392 982
rect 4450 968 4460 1148
rect 4512 968 4522 1148
rect 4582 982 4588 1192
rect 4622 982 4628 1192
rect 4700 1148 4706 1358
rect 4740 1148 4746 1358
rect 4806 1192 4816 1372
rect 4868 1192 4878 1372
rect 4936 1358 4982 1370
rect 4582 970 4628 982
rect 4686 968 4696 1148
rect 4748 968 4758 1148
rect 4818 982 4824 1192
rect 4858 982 4864 1192
rect 4936 1148 4942 1358
rect 4976 1148 4982 1358
rect 4818 970 4864 982
rect 4922 968 4932 1148
rect 4984 968 4994 1148
rect 5024 940 5088 1400
rect 5268 1358 5314 1370
rect 5268 1148 5274 1358
rect 5308 1148 5314 1358
rect 5374 1192 5384 1372
rect 5436 1192 5446 1372
rect 5504 1358 5550 1370
rect 5254 968 5264 1148
rect 5316 968 5326 1148
rect 5386 982 5392 1192
rect 5426 982 5432 1192
rect 5504 1148 5510 1358
rect 5544 1148 5550 1358
rect 5610 1192 5620 1372
rect 5672 1192 5682 1372
rect 5740 1358 5786 1370
rect 5386 970 5432 982
rect 5490 968 5500 1148
rect 5552 968 5562 1148
rect 5622 982 5628 1192
rect 5662 982 5668 1192
rect 5740 1148 5746 1358
rect 5780 1148 5786 1358
rect 5846 1192 5856 1372
rect 5908 1192 5918 1372
rect 5976 1358 6022 1370
rect 5622 970 5668 982
rect 5726 968 5736 1148
rect 5788 968 5798 1148
rect 5858 982 5864 1192
rect 5898 982 5904 1192
rect 5976 1148 5982 1358
rect 6016 1148 6022 1358
rect 5858 970 5904 982
rect 5962 968 5972 1148
rect 6024 968 6034 1148
rect 6064 940 6128 1400
rect 6308 1358 6354 1370
rect 6308 1148 6314 1358
rect 6348 1148 6354 1358
rect 6414 1192 6424 1372
rect 6476 1192 6486 1372
rect 6544 1358 6590 1370
rect 6294 968 6304 1148
rect 6356 968 6366 1148
rect 6426 982 6432 1192
rect 6466 982 6472 1192
rect 6544 1148 6550 1358
rect 6584 1148 6590 1358
rect 6650 1192 6660 1372
rect 6712 1192 6722 1372
rect 6780 1358 6826 1370
rect 6426 970 6472 982
rect 6530 968 6540 1148
rect 6592 968 6602 1148
rect 6662 982 6668 1192
rect 6702 982 6708 1192
rect 6780 1148 6786 1358
rect 6820 1148 6826 1358
rect 6886 1192 6896 1372
rect 6948 1192 6958 1372
rect 7016 1358 7062 1370
rect 6662 970 6708 982
rect 6766 968 6776 1148
rect 6828 968 6838 1148
rect 6898 982 6904 1192
rect 6938 982 6944 1192
rect 7016 1148 7022 1358
rect 7056 1148 7062 1358
rect 6898 970 6944 982
rect 7002 968 7012 1148
rect 7064 968 7074 1148
rect 7104 940 7168 1400
rect 7348 1358 7394 1370
rect 7348 1148 7354 1358
rect 7388 1148 7394 1358
rect 7454 1192 7464 1372
rect 7516 1192 7526 1372
rect 7584 1358 7630 1370
rect 7334 968 7344 1148
rect 7396 968 7406 1148
rect 7466 982 7472 1192
rect 7506 982 7512 1192
rect 7584 1148 7590 1358
rect 7624 1148 7630 1358
rect 7690 1192 7700 1372
rect 7752 1192 7762 1372
rect 7820 1358 7866 1370
rect 7466 970 7512 982
rect 7570 968 7580 1148
rect 7632 968 7642 1148
rect 7702 982 7708 1192
rect 7742 982 7748 1192
rect 7820 1148 7826 1358
rect 7860 1148 7866 1358
rect 7926 1192 7936 1372
rect 7988 1192 7998 1372
rect 8056 1358 8102 1370
rect 7702 970 7748 982
rect 7806 968 7816 1148
rect 7868 968 7878 1148
rect 7938 982 7944 1192
rect 7978 982 7984 1192
rect 8056 1148 8062 1358
rect 8096 1148 8102 1358
rect 7938 970 7984 982
rect 8042 968 8052 1148
rect 8104 968 8114 1148
rect 8144 940 8208 1400
rect 8388 1358 8434 1370
rect 8388 1148 8394 1358
rect 8428 1148 8434 1358
rect 8494 1192 8504 1372
rect 8556 1192 8566 1372
rect 8624 1358 8670 1370
rect 8374 968 8384 1148
rect 8436 968 8446 1148
rect 8506 982 8512 1192
rect 8546 982 8552 1192
rect 8624 1148 8630 1358
rect 8664 1148 8670 1358
rect 8730 1192 8740 1372
rect 8792 1192 8802 1372
rect 8860 1358 8906 1370
rect 8506 970 8552 982
rect 8610 968 8620 1148
rect 8672 968 8682 1148
rect 8742 982 8748 1192
rect 8782 982 8788 1192
rect 8860 1148 8866 1358
rect 8900 1148 8906 1358
rect 8966 1192 8976 1372
rect 9028 1192 9038 1372
rect 9096 1358 9142 1370
rect 8742 970 8788 982
rect 8846 968 8856 1148
rect 8908 968 8918 1148
rect 8978 982 8984 1192
rect 9018 982 9024 1192
rect 9096 1148 9102 1358
rect 9136 1148 9142 1358
rect 8978 970 9024 982
rect 9082 968 9092 1148
rect 9144 968 9154 1148
rect 9184 940 9248 1400
rect 9428 1358 9474 1370
rect 9428 1148 9434 1358
rect 9468 1148 9474 1358
rect 9534 1192 9544 1372
rect 9596 1192 9606 1372
rect 9664 1358 9710 1370
rect 9414 968 9424 1148
rect 9476 968 9486 1148
rect 9546 982 9552 1192
rect 9586 982 9592 1192
rect 9664 1148 9670 1358
rect 9704 1148 9710 1358
rect 9770 1192 9780 1372
rect 9832 1192 9842 1372
rect 9900 1358 9946 1370
rect 9546 970 9592 982
rect 9650 968 9660 1148
rect 9712 968 9722 1148
rect 9782 982 9788 1192
rect 9822 982 9828 1192
rect 9900 1148 9906 1358
rect 9940 1148 9946 1358
rect 10006 1192 10016 1372
rect 10068 1192 10078 1372
rect 10136 1358 10182 1370
rect 9782 970 9828 982
rect 9886 968 9896 1148
rect 9948 968 9958 1148
rect 10018 982 10024 1192
rect 10058 982 10064 1192
rect 10136 1148 10142 1358
rect 10176 1148 10182 1358
rect 10018 970 10064 982
rect 10122 968 10132 1148
rect 10184 968 10194 1148
rect 10224 940 10288 1400
rect 10468 1358 10514 1370
rect 10468 1148 10474 1358
rect 10508 1148 10514 1358
rect 10574 1192 10584 1372
rect 10636 1192 10646 1372
rect 10704 1358 10750 1370
rect 10454 968 10464 1148
rect 10516 968 10526 1148
rect 10586 982 10592 1192
rect 10626 982 10632 1192
rect 10704 1148 10710 1358
rect 10744 1148 10750 1358
rect 10810 1192 10820 1372
rect 10872 1192 10882 1372
rect 10940 1358 10986 1370
rect 10586 970 10632 982
rect 10690 968 10700 1148
rect 10752 968 10762 1148
rect 10822 982 10828 1192
rect 10862 982 10868 1192
rect 10940 1148 10946 1358
rect 10980 1148 10986 1358
rect 11046 1192 11056 1372
rect 11108 1192 11118 1372
rect 11176 1358 11222 1370
rect 10822 970 10868 982
rect 10926 968 10936 1148
rect 10988 968 10998 1148
rect 11058 982 11064 1192
rect 11098 982 11104 1192
rect 11176 1148 11182 1358
rect 11216 1148 11222 1358
rect 11058 970 11104 982
rect 11162 968 11172 1148
rect 11224 968 11234 1148
rect 11264 940 11328 1400
rect 4276 932 5088 940
rect 4276 898 4293 932
rect 4327 898 4411 932
rect 4445 898 4529 932
rect 4563 898 4647 932
rect 4681 898 4765 932
rect 4799 898 4883 932
rect 4917 898 5088 932
rect 4276 872 5088 898
rect 5316 932 6128 940
rect 5316 898 5333 932
rect 5367 898 5451 932
rect 5485 898 5569 932
rect 5603 898 5687 932
rect 5721 898 5805 932
rect 5839 898 5923 932
rect 5957 898 6128 932
rect 5316 872 6128 898
rect 6356 932 7168 940
rect 6356 898 6373 932
rect 6407 898 6491 932
rect 6525 898 6609 932
rect 6643 898 6727 932
rect 6761 898 6845 932
rect 6879 898 6963 932
rect 6997 898 7168 932
rect 6356 872 7168 898
rect 7396 932 8208 940
rect 7396 898 7413 932
rect 7447 898 7531 932
rect 7565 898 7649 932
rect 7683 898 7767 932
rect 7801 898 7885 932
rect 7919 898 8003 932
rect 8037 898 8208 932
rect 7396 872 8208 898
rect 8436 932 9248 940
rect 8436 898 8453 932
rect 8487 898 8571 932
rect 8605 898 8689 932
rect 8723 898 8807 932
rect 8841 898 8925 932
rect 8959 898 9043 932
rect 9077 898 9248 932
rect 8436 872 9248 898
rect 9476 932 10288 940
rect 9476 898 9493 932
rect 9527 898 9611 932
rect 9645 898 9729 932
rect 9763 898 9847 932
rect 9881 898 9965 932
rect 9999 898 10083 932
rect 10117 898 10288 932
rect 9476 872 10288 898
rect 10516 932 11328 940
rect 10516 898 10533 932
rect 10567 898 10651 932
rect 10685 898 10769 932
rect 10803 898 10887 932
rect 10921 898 11005 932
rect 11039 898 11123 932
rect 11157 898 11328 932
rect 10516 872 11328 898
rect -1640 772 4156 780
rect -1640 738 -1511 772
rect -1477 738 -1393 772
rect -1359 738 -1275 772
rect -1241 738 -1157 772
rect -1123 738 -1039 772
rect -1005 738 -921 772
rect -887 738 -471 772
rect -437 738 -353 772
rect -319 738 -235 772
rect -201 738 -117 772
rect -83 738 1 772
rect 35 738 119 772
rect 153 738 569 772
rect 603 738 687 772
rect 721 738 805 772
rect 839 738 923 772
rect 957 738 1041 772
rect 1075 738 1159 772
rect 1193 738 1609 772
rect 1643 738 1727 772
rect 1761 738 1845 772
rect 1879 738 1963 772
rect 1997 738 2081 772
rect 2115 738 2199 772
rect 2233 738 2649 772
rect 2683 738 2767 772
rect 2801 738 2885 772
rect 2919 738 3003 772
rect 3037 738 3121 772
rect 3155 738 3239 772
rect 3273 738 4156 772
rect -1640 660 4156 738
rect -5900 580 -4808 660
rect -4648 580 4156 660
rect 4260 624 4972 668
rect 4260 590 4282 624
rect 4316 590 4474 624
rect 4508 590 4666 624
rect 4700 590 4972 624
rect 4260 584 4972 590
rect 5300 624 6012 668
rect 5300 590 5322 624
rect 5356 590 5514 624
rect 5548 590 5706 624
rect 5740 590 6012 624
rect 5300 584 6012 590
rect 6340 624 7052 668
rect 6340 590 6362 624
rect 6396 590 6554 624
rect 6588 590 6746 624
rect 6780 590 7052 624
rect 6340 584 7052 590
rect 7380 624 8092 668
rect 7380 590 7402 624
rect 7436 590 7594 624
rect 7628 590 7786 624
rect 7820 590 8092 624
rect 7380 584 8092 590
rect 8420 624 9132 668
rect 8420 590 8442 624
rect 8476 590 8634 624
rect 8668 590 8826 624
rect 8860 590 9132 624
rect 8420 584 9132 590
rect 9460 624 10172 668
rect 9460 590 9482 624
rect 9516 590 9674 624
rect 9708 590 9866 624
rect 9900 590 10172 624
rect 9460 584 10172 590
rect 10500 624 11212 668
rect 10500 590 10522 624
rect 10556 590 10714 624
rect 10748 590 10906 624
rect 10940 590 11212 624
rect 10500 584 11212 590
rect -5900 406 -5840 580
rect 2788 492 3080 498
rect -1320 476 -1116 482
rect -1320 412 -1308 476
rect -1128 412 -1116 476
rect -1320 406 -1116 412
rect 2788 408 2800 492
rect 3068 408 3080 492
rect -6008 154 -5998 406
rect -5802 154 -5792 406
rect 2788 402 3080 408
rect 3640 156 3860 580
rect -7370 18 -6286 86
rect -7370 -16 -7352 18
rect -7318 -16 -7160 18
rect -7126 -16 -6968 18
rect -6934 -16 -6776 18
rect -6742 -16 -6584 18
rect -6550 -16 -6286 18
rect -5998 -2 -5802 154
rect 3640 76 3924 156
rect -7370 -22 -6286 -16
rect -7310 -54 -7262 -22
rect -7118 -54 -7070 -22
rect -6926 -54 -6878 -22
rect -6734 -54 -6694 -22
rect -6542 -54 -6502 -22
rect -7406 -66 -7360 -54
rect -7406 -274 -7400 -66
rect -7366 -274 -7360 -66
rect -7324 -234 -7314 -54
rect -7262 -234 -7252 -54
rect -7214 -66 -7168 -54
rect -7420 -454 -7410 -274
rect -7358 -454 -7348 -274
rect -7310 -442 -7304 -234
rect -7270 -442 -7264 -234
rect -7214 -274 -7208 -66
rect -7174 -274 -7168 -66
rect -7132 -234 -7122 -54
rect -7070 -234 -7060 -54
rect -7022 -66 -6976 -54
rect -7310 -454 -7264 -442
rect -7228 -454 -7218 -274
rect -7166 -454 -7156 -274
rect -7118 -442 -7112 -234
rect -7078 -442 -7072 -234
rect -7022 -274 -7016 -66
rect -6982 -274 -6976 -66
rect -6940 -234 -6930 -54
rect -6878 -234 -6868 -54
rect -6830 -66 -6784 -54
rect -7118 -454 -7072 -442
rect -7036 -454 -7026 -274
rect -6974 -454 -6964 -274
rect -6926 -442 -6920 -234
rect -6886 -442 -6880 -234
rect -6830 -274 -6824 -66
rect -6790 -274 -6784 -66
rect -6748 -234 -6738 -54
rect -6686 -234 -6676 -54
rect -6638 -66 -6592 -54
rect -6926 -454 -6880 -442
rect -6844 -454 -6834 -274
rect -6782 -454 -6772 -274
rect -6734 -442 -6728 -234
rect -6694 -442 -6688 -234
rect -6638 -274 -6632 -66
rect -6598 -274 -6592 -66
rect -6556 -234 -6546 -54
rect -6494 -234 -6484 -54
rect -6446 -66 -6400 -54
rect -6734 -454 -6688 -442
rect -6652 -454 -6642 -274
rect -6590 -454 -6580 -274
rect -6542 -442 -6536 -234
rect -6502 -442 -6496 -234
rect -6446 -274 -6440 -66
rect -6406 -274 -6400 -66
rect -6542 -454 -6496 -442
rect -6460 -454 -6450 -274
rect -6398 -454 -6388 -274
rect -6358 -486 -6286 -22
rect -6000 -8 -5800 -2
rect -6000 -42 -5988 -8
rect -5812 -42 -5800 -8
rect -6000 -48 -5800 -42
rect -6078 -70 -6032 -58
rect -6078 -486 -6072 -70
rect -7274 -492 -6072 -486
rect -7274 -526 -7256 -492
rect -7222 -526 -7064 -492
rect -7030 -526 -6872 -492
rect -6838 -526 -6680 -492
rect -6646 -526 -6488 -492
rect -6454 -526 -6072 -492
rect -7274 -600 -6072 -526
rect -7274 -634 -7256 -600
rect -7222 -634 -7064 -600
rect -7030 -634 -6872 -600
rect -6838 -634 -6680 -600
rect -6646 -634 -6488 -600
rect -6454 -634 -6072 -600
rect -7274 -642 -6072 -634
rect -7406 -684 -7360 -672
rect -7406 -894 -7400 -684
rect -7366 -894 -7360 -684
rect -7324 -850 -7314 -670
rect -7262 -850 -7252 -670
rect -7214 -684 -7168 -672
rect -7420 -1074 -7410 -894
rect -7358 -1074 -7348 -894
rect -7310 -1060 -7304 -850
rect -7270 -1060 -7264 -850
rect -7214 -894 -7208 -684
rect -7174 -894 -7168 -684
rect -7132 -850 -7122 -670
rect -7070 -850 -7060 -670
rect -7022 -684 -6976 -672
rect -7310 -1072 -7264 -1060
rect -7228 -1074 -7218 -894
rect -7166 -1074 -7156 -894
rect -7118 -1060 -7112 -850
rect -7078 -1060 -7072 -850
rect -7022 -894 -7016 -684
rect -6982 -894 -6976 -684
rect -6940 -850 -6930 -670
rect -6878 -850 -6868 -670
rect -6830 -684 -6784 -672
rect -7118 -1072 -7072 -1060
rect -7036 -1074 -7026 -894
rect -6974 -1074 -6964 -894
rect -6926 -1060 -6920 -850
rect -6886 -1060 -6880 -850
rect -6830 -894 -6824 -684
rect -6790 -894 -6784 -684
rect -6748 -850 -6738 -670
rect -6686 -850 -6676 -670
rect -6638 -684 -6592 -672
rect -6926 -1072 -6880 -1060
rect -6844 -1074 -6834 -894
rect -6782 -1074 -6772 -894
rect -6734 -1060 -6728 -850
rect -6694 -1060 -6688 -850
rect -6638 -894 -6632 -684
rect -6598 -894 -6592 -684
rect -6556 -850 -6546 -670
rect -6494 -850 -6484 -670
rect -6446 -684 -6400 -672
rect -6734 -1072 -6688 -1060
rect -6652 -1074 -6642 -894
rect -6590 -1074 -6580 -894
rect -6542 -1060 -6536 -850
rect -6502 -1060 -6496 -850
rect -6446 -894 -6440 -684
rect -6406 -894 -6400 -684
rect -6542 -1072 -6496 -1060
rect -6460 -1074 -6450 -894
rect -6398 -1074 -6388 -894
rect -6354 -1102 -6286 -642
rect -7374 -1110 -6286 -1102
rect -7374 -1144 -7352 -1110
rect -7318 -1144 -7160 -1110
rect -7126 -1144 -6968 -1110
rect -6934 -1144 -6776 -1110
rect -6742 -1144 -6584 -1110
rect -6550 -1144 -6286 -1110
rect -7374 -1210 -6286 -1144
rect -6078 -1638 -6072 -642
rect -6038 -486 -6032 -70
rect -5768 -70 -5722 -58
rect -5768 -486 -5762 -70
rect -6038 -642 -5762 -486
rect -6038 -1638 -6032 -642
rect -6078 -1650 -6032 -1638
rect -5768 -1638 -5762 -642
rect -5728 -1638 -5722 -70
rect 3640 -140 3712 76
rect 3912 -140 3924 76
rect 4000 100 4156 580
rect 4214 372 4224 552
rect 4276 372 4286 552
rect 4324 540 4370 552
rect 4228 164 4234 372
rect 4268 164 4274 372
rect 4324 332 4330 540
rect 4364 332 4370 540
rect 4406 372 4416 552
rect 4468 372 4478 552
rect 4516 540 4562 552
rect 4228 152 4274 164
rect 4310 152 4320 332
rect 4372 152 4382 332
rect 4420 164 4426 372
rect 4460 164 4466 372
rect 4516 332 4522 540
rect 4556 332 4562 540
rect 4598 372 4608 552
rect 4660 372 4670 552
rect 4708 540 4754 552
rect 4420 152 4466 164
rect 4502 152 4512 332
rect 4564 152 4574 332
rect 4612 164 4618 372
rect 4652 164 4658 372
rect 4708 332 4714 540
rect 4748 332 4754 540
rect 4790 372 4800 552
rect 4852 372 4862 552
rect 4612 152 4658 164
rect 4694 152 4704 332
rect 4756 152 4766 332
rect 4804 164 4810 372
rect 4844 164 4850 372
rect 4804 152 4850 164
rect 4892 120 4972 584
rect 5254 372 5264 552
rect 5316 372 5326 552
rect 5364 540 5410 552
rect 5268 164 5274 372
rect 5308 164 5314 372
rect 5364 332 5370 540
rect 5404 332 5410 540
rect 5446 372 5456 552
rect 5508 372 5518 552
rect 5556 540 5602 552
rect 5268 152 5314 164
rect 5350 152 5360 332
rect 5412 152 5422 332
rect 5460 164 5466 372
rect 5500 164 5506 372
rect 5556 332 5562 540
rect 5596 332 5602 540
rect 5638 372 5648 552
rect 5700 372 5710 552
rect 5748 540 5794 552
rect 5460 152 5506 164
rect 5542 152 5552 332
rect 5604 152 5614 332
rect 5652 164 5658 372
rect 5692 164 5698 372
rect 5748 332 5754 540
rect 5788 332 5794 540
rect 5830 372 5840 552
rect 5892 372 5902 552
rect 5652 152 5698 164
rect 5734 152 5744 332
rect 5796 152 5806 332
rect 5844 164 5850 372
rect 5884 164 5890 372
rect 5844 152 5890 164
rect 5932 120 6012 584
rect 6294 372 6304 552
rect 6356 372 6366 552
rect 6404 540 6450 552
rect 6308 164 6314 372
rect 6348 164 6354 372
rect 6404 332 6410 540
rect 6444 332 6450 540
rect 6486 372 6496 552
rect 6548 372 6558 552
rect 6596 540 6642 552
rect 6308 152 6354 164
rect 6390 152 6400 332
rect 6452 152 6462 332
rect 6500 164 6506 372
rect 6540 164 6546 372
rect 6596 332 6602 540
rect 6636 332 6642 540
rect 6678 372 6688 552
rect 6740 372 6750 552
rect 6788 540 6834 552
rect 6500 152 6546 164
rect 6582 152 6592 332
rect 6644 152 6654 332
rect 6692 164 6698 372
rect 6732 164 6738 372
rect 6788 332 6794 540
rect 6828 332 6834 540
rect 6870 372 6880 552
rect 6932 372 6942 552
rect 6692 152 6738 164
rect 6774 152 6784 332
rect 6836 152 6846 332
rect 6884 164 6890 372
rect 6924 164 6930 372
rect 6884 152 6930 164
rect 6972 120 7052 584
rect 7334 372 7344 552
rect 7396 372 7406 552
rect 7444 540 7490 552
rect 7348 164 7354 372
rect 7388 164 7394 372
rect 7444 332 7450 540
rect 7484 332 7490 540
rect 7526 372 7536 552
rect 7588 372 7598 552
rect 7636 540 7682 552
rect 7348 152 7394 164
rect 7430 152 7440 332
rect 7492 152 7502 332
rect 7540 164 7546 372
rect 7580 164 7586 372
rect 7636 332 7642 540
rect 7676 332 7682 540
rect 7718 372 7728 552
rect 7780 372 7790 552
rect 7828 540 7874 552
rect 7540 152 7586 164
rect 7622 152 7632 332
rect 7684 152 7694 332
rect 7732 164 7738 372
rect 7772 164 7778 372
rect 7828 332 7834 540
rect 7868 332 7874 540
rect 7910 372 7920 552
rect 7972 372 7982 552
rect 7732 152 7778 164
rect 7814 152 7824 332
rect 7876 152 7886 332
rect 7924 164 7930 372
rect 7964 164 7970 372
rect 7924 152 7970 164
rect 8012 120 8092 584
rect 8374 372 8384 552
rect 8436 372 8446 552
rect 8484 540 8530 552
rect 8388 164 8394 372
rect 8428 164 8434 372
rect 8484 332 8490 540
rect 8524 332 8530 540
rect 8566 372 8576 552
rect 8628 372 8638 552
rect 8676 540 8722 552
rect 8388 152 8434 164
rect 8470 152 8480 332
rect 8532 152 8542 332
rect 8580 164 8586 372
rect 8620 164 8626 372
rect 8676 332 8682 540
rect 8716 332 8722 540
rect 8758 372 8768 552
rect 8820 372 8830 552
rect 8868 540 8914 552
rect 8580 152 8626 164
rect 8662 152 8672 332
rect 8724 152 8734 332
rect 8772 164 8778 372
rect 8812 164 8818 372
rect 8868 332 8874 540
rect 8908 332 8914 540
rect 8950 372 8960 552
rect 9012 372 9022 552
rect 8772 152 8818 164
rect 8854 152 8864 332
rect 8916 152 8926 332
rect 8964 164 8970 372
rect 9004 164 9010 372
rect 8964 152 9010 164
rect 9052 120 9132 584
rect 9414 372 9424 552
rect 9476 372 9486 552
rect 9524 540 9570 552
rect 9428 164 9434 372
rect 9468 164 9474 372
rect 9524 332 9530 540
rect 9564 332 9570 540
rect 9606 372 9616 552
rect 9668 372 9678 552
rect 9716 540 9762 552
rect 9428 152 9474 164
rect 9510 152 9520 332
rect 9572 152 9582 332
rect 9620 164 9626 372
rect 9660 164 9666 372
rect 9716 332 9722 540
rect 9756 332 9762 540
rect 9798 372 9808 552
rect 9860 372 9870 552
rect 9908 540 9954 552
rect 9620 152 9666 164
rect 9702 152 9712 332
rect 9764 152 9774 332
rect 9812 164 9818 372
rect 9852 164 9858 372
rect 9908 332 9914 540
rect 9948 332 9954 540
rect 9990 372 10000 552
rect 10052 372 10062 552
rect 9812 152 9858 164
rect 9894 152 9904 332
rect 9956 152 9966 332
rect 10004 164 10010 372
rect 10044 164 10050 372
rect 10004 152 10050 164
rect 10092 120 10172 584
rect 10454 372 10464 552
rect 10516 372 10526 552
rect 10564 540 10610 552
rect 10468 164 10474 372
rect 10508 164 10514 372
rect 10564 332 10570 540
rect 10604 332 10610 540
rect 10646 372 10656 552
rect 10708 372 10718 552
rect 10756 540 10802 552
rect 10468 152 10514 164
rect 10550 152 10560 332
rect 10612 152 10622 332
rect 10660 164 10666 372
rect 10700 164 10706 372
rect 10756 332 10762 540
rect 10796 332 10802 540
rect 10838 372 10848 552
rect 10900 372 10910 552
rect 10948 540 10994 552
rect 10660 152 10706 164
rect 10742 152 10752 332
rect 10804 152 10814 332
rect 10852 164 10858 372
rect 10892 164 10898 372
rect 10948 332 10954 540
rect 10988 332 10994 540
rect 11030 372 11040 552
rect 11092 372 11102 552
rect 10852 152 10898 164
rect 10934 152 10944 332
rect 10996 152 11006 332
rect 11044 164 11050 372
rect 11084 164 11090 372
rect 11044 152 11090 164
rect 11132 120 11212 584
rect 4320 114 4972 120
rect 4320 100 4378 114
rect 4000 80 4378 100
rect 4412 80 4570 114
rect 4604 80 4762 114
rect 4796 100 4972 114
rect 5360 114 6012 120
rect 5360 100 5418 114
rect 4796 80 5418 100
rect 5452 80 5610 114
rect 5644 80 5802 114
rect 5836 100 6012 114
rect 6400 114 7052 120
rect 6400 100 6458 114
rect 5836 80 6458 100
rect 6492 80 6650 114
rect 6684 80 6842 114
rect 6876 100 7052 114
rect 7440 114 8092 120
rect 7440 100 7498 114
rect 6876 80 7498 100
rect 7532 80 7690 114
rect 7724 80 7882 114
rect 7916 100 8092 114
rect 8480 114 9132 120
rect 8480 100 8538 114
rect 7916 80 8538 100
rect 8572 80 8730 114
rect 8764 80 8922 114
rect 8956 100 9132 114
rect 9520 114 10172 120
rect 9520 100 9578 114
rect 8956 80 9578 100
rect 9612 80 9770 114
rect 9804 80 9962 114
rect 9996 100 10172 114
rect 10560 114 11212 120
rect 10560 100 10618 114
rect 9996 80 10618 100
rect 10652 80 10810 114
rect 10844 80 11002 114
rect 11036 80 11212 114
rect 4000 6 11212 80
rect 4000 -16 4378 6
rect -5768 -1650 -5722 -1638
rect -6000 -1666 -5800 -1660
rect -6000 -1700 -5988 -1666
rect -5812 -1700 -5800 -1666
rect -6000 -1706 -5800 -1700
rect -5998 -1748 -5802 -1706
rect -6198 -1754 -5778 -1748
rect -6198 -1774 -6186 -1754
rect -7406 -1818 -6186 -1774
rect -7406 -1852 -7352 -1818
rect -7318 -1852 -7160 -1818
rect -7126 -1852 -6968 -1818
rect -6934 -1834 -6186 -1818
rect -5790 -1834 -5778 -1754
rect -6934 -1840 -5778 -1834
rect -6934 -1852 -5790 -1840
rect -7406 -1858 -5790 -1852
rect -7406 -1890 -7358 -1858
rect -7214 -1890 -7166 -1858
rect -7022 -1890 -6974 -1858
rect -6830 -1890 -6782 -1858
rect -7420 -2070 -7410 -1890
rect -7358 -2070 -7348 -1890
rect -7310 -1902 -7264 -1890
rect -7406 -2278 -7400 -2070
rect -7366 -2278 -7360 -2070
rect -7310 -2110 -7304 -1902
rect -7270 -2110 -7264 -1902
rect -7228 -2070 -7218 -1890
rect -7166 -2070 -7156 -1890
rect -7118 -1902 -7072 -1890
rect -7406 -2290 -7360 -2278
rect -7324 -2290 -7314 -2110
rect -7262 -2290 -7252 -2110
rect -7214 -2278 -7208 -2070
rect -7174 -2278 -7168 -2070
rect -7118 -2110 -7112 -1902
rect -7078 -2110 -7072 -1902
rect -7036 -2070 -7026 -1890
rect -6974 -2070 -6964 -1890
rect -6926 -1902 -6880 -1890
rect -7214 -2290 -7168 -2278
rect -7132 -2290 -7122 -2110
rect -7070 -2290 -7060 -2110
rect -7022 -2278 -7016 -2070
rect -6982 -2278 -6976 -2070
rect -6926 -2110 -6920 -1902
rect -6886 -2110 -6880 -1902
rect -6844 -2070 -6834 -1890
rect -6782 -2070 -6772 -1890
rect -7022 -2290 -6976 -2278
rect -6940 -2290 -6930 -2110
rect -6878 -2290 -6868 -2110
rect -6830 -2278 -6824 -2070
rect -6790 -2278 -6784 -2070
rect -6830 -2290 -6784 -2278
rect -6742 -2322 -6662 -1858
rect 4000 -2140 4156 -16
rect 4320 -28 4378 -16
rect 4412 -28 4570 6
rect 4604 -28 4762 6
rect 4796 -16 5418 6
rect 4796 -28 4972 -16
rect 4320 -36 4972 -28
rect 5360 -28 5418 -16
rect 5452 -28 5610 6
rect 5644 -28 5802 6
rect 5836 -16 6458 6
rect 5836 -28 6012 -16
rect 5360 -36 6012 -28
rect 6400 -28 6458 -16
rect 6492 -28 6650 6
rect 6684 -28 6842 6
rect 6876 -16 7498 6
rect 6876 -28 7052 -16
rect 6400 -36 7052 -28
rect 7440 -28 7498 -16
rect 7532 -28 7690 6
rect 7724 -28 7882 6
rect 7916 -16 8538 6
rect 7916 -28 8092 -16
rect 7440 -36 8092 -28
rect 8480 -28 8538 -16
rect 8572 -28 8730 6
rect 8764 -28 8922 6
rect 8956 -16 9578 6
rect 8956 -28 9132 -16
rect 8480 -36 9132 -28
rect 9520 -28 9578 -16
rect 9612 -28 9770 6
rect 9804 -28 9962 6
rect 9996 -16 10618 6
rect 9996 -28 10172 -16
rect 9520 -36 10172 -28
rect 10560 -28 10618 -16
rect 10652 -28 10810 6
rect 10844 -28 11002 6
rect 11036 -28 11212 6
rect 10560 -36 11212 -28
rect 4228 -78 4274 -66
rect 4228 -284 4234 -78
rect 4268 -284 4274 -78
rect 4310 -244 4320 -64
rect 4372 -244 4382 -64
rect 4420 -78 4466 -66
rect 4214 -464 4224 -284
rect 4276 -464 4286 -284
rect 4324 -454 4330 -244
rect 4364 -454 4370 -244
rect 4420 -284 4426 -78
rect 4460 -284 4466 -78
rect 4502 -244 4512 -64
rect 4564 -244 4574 -64
rect 4612 -78 4658 -66
rect 4228 -466 4274 -464
rect 4324 -466 4370 -454
rect 4406 -464 4416 -284
rect 4468 -464 4478 -284
rect 4516 -454 4522 -244
rect 4556 -454 4562 -244
rect 4612 -284 4618 -78
rect 4652 -284 4658 -78
rect 4694 -244 4704 -64
rect 4756 -244 4766 -64
rect 4804 -78 4850 -66
rect 4420 -466 4466 -464
rect 4516 -466 4562 -454
rect 4598 -464 4608 -284
rect 4660 -464 4670 -284
rect 4708 -454 4714 -244
rect 4748 -454 4754 -244
rect 4804 -284 4810 -78
rect 4844 -284 4850 -78
rect 4612 -466 4658 -464
rect 4708 -466 4754 -454
rect 4790 -464 4800 -284
rect 4852 -464 4862 -284
rect 4804 -466 4850 -464
rect 4270 -500 4328 -498
rect 4462 -500 4520 -498
rect 4654 -500 4712 -498
rect 4892 -500 4972 -36
rect 5268 -78 5314 -66
rect 5268 -284 5274 -78
rect 5308 -284 5314 -78
rect 5350 -244 5360 -64
rect 5412 -244 5422 -64
rect 5460 -78 5506 -66
rect 5254 -464 5264 -284
rect 5316 -464 5326 -284
rect 5364 -454 5370 -244
rect 5404 -454 5410 -244
rect 5460 -284 5466 -78
rect 5500 -284 5506 -78
rect 5542 -244 5552 -64
rect 5604 -244 5614 -64
rect 5652 -78 5698 -66
rect 5268 -466 5314 -464
rect 5364 -466 5410 -454
rect 5446 -464 5456 -284
rect 5508 -464 5518 -284
rect 5556 -454 5562 -244
rect 5596 -454 5602 -244
rect 5652 -284 5658 -78
rect 5692 -284 5698 -78
rect 5734 -244 5744 -64
rect 5796 -244 5806 -64
rect 5844 -78 5890 -66
rect 5460 -466 5506 -464
rect 5556 -466 5602 -454
rect 5638 -464 5648 -284
rect 5700 -464 5710 -284
rect 5748 -454 5754 -244
rect 5788 -454 5794 -244
rect 5844 -284 5850 -78
rect 5884 -284 5890 -78
rect 5652 -466 5698 -464
rect 5748 -466 5794 -454
rect 5830 -464 5840 -284
rect 5892 -464 5902 -284
rect 5844 -466 5890 -464
rect 5310 -500 5368 -498
rect 5502 -500 5560 -498
rect 5694 -500 5752 -498
rect 5932 -500 6012 -36
rect 6308 -78 6354 -66
rect 6308 -284 6314 -78
rect 6348 -284 6354 -78
rect 6390 -244 6400 -64
rect 6452 -244 6462 -64
rect 6500 -78 6546 -66
rect 6294 -464 6304 -284
rect 6356 -464 6366 -284
rect 6404 -454 6410 -244
rect 6444 -454 6450 -244
rect 6500 -284 6506 -78
rect 6540 -284 6546 -78
rect 6582 -244 6592 -64
rect 6644 -244 6654 -64
rect 6692 -78 6738 -66
rect 6308 -466 6354 -464
rect 6404 -466 6450 -454
rect 6486 -464 6496 -284
rect 6548 -464 6558 -284
rect 6596 -454 6602 -244
rect 6636 -454 6642 -244
rect 6692 -284 6698 -78
rect 6732 -284 6738 -78
rect 6774 -244 6784 -64
rect 6836 -244 6846 -64
rect 6884 -78 6930 -66
rect 6500 -466 6546 -464
rect 6596 -466 6642 -454
rect 6678 -464 6688 -284
rect 6740 -464 6750 -284
rect 6788 -454 6794 -244
rect 6828 -454 6834 -244
rect 6884 -284 6890 -78
rect 6924 -284 6930 -78
rect 6692 -466 6738 -464
rect 6788 -466 6834 -454
rect 6870 -464 6880 -284
rect 6932 -464 6942 -284
rect 6884 -466 6930 -464
rect 6350 -500 6408 -498
rect 6542 -500 6600 -498
rect 6734 -500 6792 -498
rect 6972 -500 7052 -36
rect 7348 -78 7394 -66
rect 7348 -284 7354 -78
rect 7388 -284 7394 -78
rect 7430 -244 7440 -64
rect 7492 -244 7502 -64
rect 7540 -78 7586 -66
rect 7334 -464 7344 -284
rect 7396 -464 7406 -284
rect 7444 -454 7450 -244
rect 7484 -454 7490 -244
rect 7540 -284 7546 -78
rect 7580 -284 7586 -78
rect 7622 -244 7632 -64
rect 7684 -244 7694 -64
rect 7732 -78 7778 -66
rect 7348 -466 7394 -464
rect 7444 -466 7490 -454
rect 7526 -464 7536 -284
rect 7588 -464 7598 -284
rect 7636 -454 7642 -244
rect 7676 -454 7682 -244
rect 7732 -284 7738 -78
rect 7772 -284 7778 -78
rect 7814 -244 7824 -64
rect 7876 -244 7886 -64
rect 7924 -78 7970 -66
rect 7540 -466 7586 -464
rect 7636 -466 7682 -454
rect 7718 -464 7728 -284
rect 7780 -464 7790 -284
rect 7828 -454 7834 -244
rect 7868 -454 7874 -244
rect 7924 -284 7930 -78
rect 7964 -284 7970 -78
rect 7732 -466 7778 -464
rect 7828 -466 7874 -454
rect 7910 -464 7920 -284
rect 7972 -464 7982 -284
rect 7924 -466 7970 -464
rect 7390 -500 7448 -498
rect 7582 -500 7640 -498
rect 7774 -500 7832 -498
rect 8012 -500 8092 -36
rect 8388 -78 8434 -66
rect 8388 -284 8394 -78
rect 8428 -284 8434 -78
rect 8470 -244 8480 -64
rect 8532 -244 8542 -64
rect 8580 -78 8626 -66
rect 8374 -464 8384 -284
rect 8436 -464 8446 -284
rect 8484 -454 8490 -244
rect 8524 -454 8530 -244
rect 8580 -284 8586 -78
rect 8620 -284 8626 -78
rect 8662 -244 8672 -64
rect 8724 -244 8734 -64
rect 8772 -78 8818 -66
rect 8388 -466 8434 -464
rect 8484 -466 8530 -454
rect 8566 -464 8576 -284
rect 8628 -464 8638 -284
rect 8676 -454 8682 -244
rect 8716 -454 8722 -244
rect 8772 -284 8778 -78
rect 8812 -284 8818 -78
rect 8854 -244 8864 -64
rect 8916 -244 8926 -64
rect 8964 -78 9010 -66
rect 8580 -466 8626 -464
rect 8676 -466 8722 -454
rect 8758 -464 8768 -284
rect 8820 -464 8830 -284
rect 8868 -454 8874 -244
rect 8908 -454 8914 -244
rect 8964 -284 8970 -78
rect 9004 -284 9010 -78
rect 8772 -466 8818 -464
rect 8868 -466 8914 -454
rect 8950 -464 8960 -284
rect 9012 -464 9022 -284
rect 8964 -466 9010 -464
rect 8430 -500 8488 -498
rect 8622 -500 8680 -498
rect 8814 -500 8872 -498
rect 9052 -500 9132 -36
rect 9428 -78 9474 -66
rect 9428 -284 9434 -78
rect 9468 -284 9474 -78
rect 9510 -244 9520 -64
rect 9572 -244 9582 -64
rect 9620 -78 9666 -66
rect 9414 -464 9424 -284
rect 9476 -464 9486 -284
rect 9524 -454 9530 -244
rect 9564 -454 9570 -244
rect 9620 -284 9626 -78
rect 9660 -284 9666 -78
rect 9702 -244 9712 -64
rect 9764 -244 9774 -64
rect 9812 -78 9858 -66
rect 9428 -466 9474 -464
rect 9524 -466 9570 -454
rect 9606 -464 9616 -284
rect 9668 -464 9678 -284
rect 9716 -454 9722 -244
rect 9756 -454 9762 -244
rect 9812 -284 9818 -78
rect 9852 -284 9858 -78
rect 9894 -244 9904 -64
rect 9956 -244 9966 -64
rect 10004 -78 10050 -66
rect 9620 -466 9666 -464
rect 9716 -466 9762 -454
rect 9798 -464 9808 -284
rect 9860 -464 9870 -284
rect 9908 -454 9914 -244
rect 9948 -454 9954 -244
rect 10004 -284 10010 -78
rect 10044 -284 10050 -78
rect 9812 -466 9858 -464
rect 9908 -466 9954 -454
rect 9990 -464 10000 -284
rect 10052 -464 10062 -284
rect 10004 -466 10050 -464
rect 9470 -500 9528 -498
rect 9662 -500 9720 -498
rect 9854 -500 9912 -498
rect 10092 -500 10172 -36
rect 10468 -78 10514 -66
rect 10468 -284 10474 -78
rect 10508 -284 10514 -78
rect 10550 -244 10560 -64
rect 10612 -244 10622 -64
rect 10660 -78 10706 -66
rect 10454 -464 10464 -284
rect 10516 -464 10526 -284
rect 10564 -454 10570 -244
rect 10604 -454 10610 -244
rect 10660 -284 10666 -78
rect 10700 -284 10706 -78
rect 10742 -244 10752 -64
rect 10804 -244 10814 -64
rect 10852 -78 10898 -66
rect 10468 -466 10514 -464
rect 10564 -466 10610 -454
rect 10646 -464 10656 -284
rect 10708 -464 10718 -284
rect 10756 -454 10762 -244
rect 10796 -454 10802 -244
rect 10852 -284 10858 -78
rect 10892 -284 10898 -78
rect 10934 -244 10944 -64
rect 10996 -244 11006 -64
rect 11044 -78 11090 -66
rect 10660 -466 10706 -464
rect 10756 -466 10802 -454
rect 10838 -464 10848 -284
rect 10900 -464 10910 -284
rect 10948 -454 10954 -244
rect 10988 -454 10994 -244
rect 11044 -284 11050 -78
rect 11084 -284 11090 -78
rect 10852 -466 10898 -464
rect 10948 -466 10994 -454
rect 11030 -464 11040 -284
rect 11092 -464 11102 -284
rect 11044 -466 11090 -464
rect 10510 -500 10568 -498
rect 10702 -500 10760 -498
rect 10894 -500 10952 -498
rect 11132 -500 11212 -36
rect 4264 -504 4972 -500
rect 4264 -538 4282 -504
rect 4316 -538 4474 -504
rect 4508 -538 4666 -504
rect 4700 -538 4972 -504
rect 4264 -596 4972 -538
rect 5304 -504 6012 -500
rect 5304 -538 5322 -504
rect 5356 -538 5514 -504
rect 5548 -538 5706 -504
rect 5740 -538 6012 -504
rect 5304 -596 6012 -538
rect 6344 -504 7052 -500
rect 6344 -538 6362 -504
rect 6396 -538 6554 -504
rect 6588 -538 6746 -504
rect 6780 -538 7052 -504
rect 6344 -596 7052 -538
rect 7384 -504 8092 -500
rect 7384 -538 7402 -504
rect 7436 -538 7594 -504
rect 7628 -538 7786 -504
rect 7820 -538 8092 -504
rect 7384 -596 8092 -538
rect 8424 -504 9132 -500
rect 8424 -538 8442 -504
rect 8476 -538 8634 -504
rect 8668 -538 8826 -504
rect 8860 -538 9132 -504
rect 8424 -596 9132 -538
rect 9464 -504 10172 -500
rect 9464 -538 9482 -504
rect 9516 -538 9674 -504
rect 9708 -538 9866 -504
rect 9900 -538 10172 -504
rect 9464 -596 10172 -538
rect 10504 -504 11212 -500
rect 10504 -538 10522 -504
rect 10556 -538 10714 -504
rect 10748 -538 10906 -504
rect 10940 -538 11212 -504
rect 10504 -596 11212 -538
rect 11620 100 11776 2224
rect 11940 2212 11998 2224
rect 12032 2212 12190 2246
rect 12224 2212 12382 2246
rect 12416 2224 13038 2246
rect 12416 2212 12592 2224
rect 11940 2204 12592 2212
rect 12980 2212 13038 2224
rect 13072 2212 13230 2246
rect 13264 2212 13422 2246
rect 13456 2224 14078 2246
rect 13456 2212 13632 2224
rect 12980 2204 13632 2212
rect 14020 2212 14078 2224
rect 14112 2212 14270 2246
rect 14304 2212 14462 2246
rect 14496 2224 15118 2246
rect 14496 2212 14672 2224
rect 14020 2204 14672 2212
rect 15060 2212 15118 2224
rect 15152 2212 15310 2246
rect 15344 2212 15502 2246
rect 15536 2224 16158 2246
rect 15536 2212 15712 2224
rect 15060 2204 15712 2212
rect 16100 2212 16158 2224
rect 16192 2212 16350 2246
rect 16384 2212 16542 2246
rect 16576 2224 17198 2246
rect 16576 2212 16752 2224
rect 16100 2204 16752 2212
rect 17140 2212 17198 2224
rect 17232 2212 17390 2246
rect 17424 2212 17582 2246
rect 17616 2224 18238 2246
rect 17616 2212 17792 2224
rect 17140 2204 17792 2212
rect 18180 2212 18238 2224
rect 18272 2212 18430 2246
rect 18464 2212 18622 2246
rect 18656 2212 18832 2246
rect 18180 2204 18832 2212
rect 11848 2162 11894 2174
rect 11848 1956 11854 2162
rect 11888 1956 11894 2162
rect 11930 1996 11940 2176
rect 11992 1996 12002 2176
rect 12040 2162 12086 2174
rect 11834 1776 11844 1956
rect 11896 1776 11906 1956
rect 11944 1786 11950 1996
rect 11984 1786 11990 1996
rect 12040 1956 12046 2162
rect 12080 1956 12086 2162
rect 12122 1996 12132 2176
rect 12184 1996 12194 2176
rect 12232 2162 12278 2174
rect 11848 1774 11894 1776
rect 11944 1774 11990 1786
rect 12026 1776 12036 1956
rect 12088 1776 12098 1956
rect 12136 1786 12142 1996
rect 12176 1786 12182 1996
rect 12232 1956 12238 2162
rect 12272 1956 12278 2162
rect 12314 1996 12324 2176
rect 12376 1996 12386 2176
rect 12424 2162 12470 2174
rect 12040 1774 12086 1776
rect 12136 1774 12182 1786
rect 12218 1776 12228 1956
rect 12280 1776 12290 1956
rect 12328 1786 12334 1996
rect 12368 1786 12374 1996
rect 12424 1956 12430 2162
rect 12464 1956 12470 2162
rect 12232 1774 12278 1776
rect 12328 1774 12374 1786
rect 12410 1776 12420 1956
rect 12472 1776 12482 1956
rect 12424 1774 12470 1776
rect 11890 1740 11948 1742
rect 12082 1740 12140 1742
rect 12274 1740 12332 1742
rect 12512 1740 12592 2204
rect 12888 2162 12934 2174
rect 12888 1956 12894 2162
rect 12928 1956 12934 2162
rect 12970 1996 12980 2176
rect 13032 1996 13042 2176
rect 13080 2162 13126 2174
rect 12874 1776 12884 1956
rect 12936 1776 12946 1956
rect 12984 1786 12990 1996
rect 13024 1786 13030 1996
rect 13080 1956 13086 2162
rect 13120 1956 13126 2162
rect 13162 1996 13172 2176
rect 13224 1996 13234 2176
rect 13272 2162 13318 2174
rect 12888 1774 12934 1776
rect 12984 1774 13030 1786
rect 13066 1776 13076 1956
rect 13128 1776 13138 1956
rect 13176 1786 13182 1996
rect 13216 1786 13222 1996
rect 13272 1956 13278 2162
rect 13312 1956 13318 2162
rect 13354 1996 13364 2176
rect 13416 1996 13426 2176
rect 13464 2162 13510 2174
rect 13080 1774 13126 1776
rect 13176 1774 13222 1786
rect 13258 1776 13268 1956
rect 13320 1776 13330 1956
rect 13368 1786 13374 1996
rect 13408 1786 13414 1996
rect 13464 1956 13470 2162
rect 13504 1956 13510 2162
rect 13272 1774 13318 1776
rect 13368 1774 13414 1786
rect 13450 1776 13460 1956
rect 13512 1776 13522 1956
rect 13464 1774 13510 1776
rect 12930 1740 12988 1742
rect 13122 1740 13180 1742
rect 13314 1740 13372 1742
rect 13552 1740 13632 2204
rect 13928 2162 13974 2174
rect 13928 1956 13934 2162
rect 13968 1956 13974 2162
rect 14010 1996 14020 2176
rect 14072 1996 14082 2176
rect 14120 2162 14166 2174
rect 13914 1776 13924 1956
rect 13976 1776 13986 1956
rect 14024 1786 14030 1996
rect 14064 1786 14070 1996
rect 14120 1956 14126 2162
rect 14160 1956 14166 2162
rect 14202 1996 14212 2176
rect 14264 1996 14274 2176
rect 14312 2162 14358 2174
rect 13928 1774 13974 1776
rect 14024 1774 14070 1786
rect 14106 1776 14116 1956
rect 14168 1776 14178 1956
rect 14216 1786 14222 1996
rect 14256 1786 14262 1996
rect 14312 1956 14318 2162
rect 14352 1956 14358 2162
rect 14394 1996 14404 2176
rect 14456 1996 14466 2176
rect 14504 2162 14550 2174
rect 14120 1774 14166 1776
rect 14216 1774 14262 1786
rect 14298 1776 14308 1956
rect 14360 1776 14370 1956
rect 14408 1786 14414 1996
rect 14448 1786 14454 1996
rect 14504 1956 14510 2162
rect 14544 1956 14550 2162
rect 14312 1774 14358 1776
rect 14408 1774 14454 1786
rect 14490 1776 14500 1956
rect 14552 1776 14562 1956
rect 14504 1774 14550 1776
rect 13970 1740 14028 1742
rect 14162 1740 14220 1742
rect 14354 1740 14412 1742
rect 14592 1740 14672 2204
rect 14968 2162 15014 2174
rect 14968 1956 14974 2162
rect 15008 1956 15014 2162
rect 15050 1996 15060 2176
rect 15112 1996 15122 2176
rect 15160 2162 15206 2174
rect 14954 1776 14964 1956
rect 15016 1776 15026 1956
rect 15064 1786 15070 1996
rect 15104 1786 15110 1996
rect 15160 1956 15166 2162
rect 15200 1956 15206 2162
rect 15242 1996 15252 2176
rect 15304 1996 15314 2176
rect 15352 2162 15398 2174
rect 14968 1774 15014 1776
rect 15064 1774 15110 1786
rect 15146 1776 15156 1956
rect 15208 1776 15218 1956
rect 15256 1786 15262 1996
rect 15296 1786 15302 1996
rect 15352 1956 15358 2162
rect 15392 1956 15398 2162
rect 15434 1996 15444 2176
rect 15496 1996 15506 2176
rect 15544 2162 15590 2174
rect 15160 1774 15206 1776
rect 15256 1774 15302 1786
rect 15338 1776 15348 1956
rect 15400 1776 15410 1956
rect 15448 1786 15454 1996
rect 15488 1786 15494 1996
rect 15544 1956 15550 2162
rect 15584 1956 15590 2162
rect 15352 1774 15398 1776
rect 15448 1774 15494 1786
rect 15530 1776 15540 1956
rect 15592 1776 15602 1956
rect 15544 1774 15590 1776
rect 15010 1740 15068 1742
rect 15202 1740 15260 1742
rect 15394 1740 15452 1742
rect 15632 1740 15712 2204
rect 16008 2162 16054 2174
rect 16008 1956 16014 2162
rect 16048 1956 16054 2162
rect 16090 1996 16100 2176
rect 16152 1996 16162 2176
rect 16200 2162 16246 2174
rect 15994 1776 16004 1956
rect 16056 1776 16066 1956
rect 16104 1786 16110 1996
rect 16144 1786 16150 1996
rect 16200 1956 16206 2162
rect 16240 1956 16246 2162
rect 16282 1996 16292 2176
rect 16344 1996 16354 2176
rect 16392 2162 16438 2174
rect 16008 1774 16054 1776
rect 16104 1774 16150 1786
rect 16186 1776 16196 1956
rect 16248 1776 16258 1956
rect 16296 1786 16302 1996
rect 16336 1786 16342 1996
rect 16392 1956 16398 2162
rect 16432 1956 16438 2162
rect 16474 1996 16484 2176
rect 16536 1996 16546 2176
rect 16584 2162 16630 2174
rect 16200 1774 16246 1776
rect 16296 1774 16342 1786
rect 16378 1776 16388 1956
rect 16440 1776 16450 1956
rect 16488 1786 16494 1996
rect 16528 1786 16534 1996
rect 16584 1956 16590 2162
rect 16624 1956 16630 2162
rect 16392 1774 16438 1776
rect 16488 1774 16534 1786
rect 16570 1776 16580 1956
rect 16632 1776 16642 1956
rect 16584 1774 16630 1776
rect 16050 1740 16108 1742
rect 16242 1740 16300 1742
rect 16434 1740 16492 1742
rect 16672 1740 16752 2204
rect 17048 2162 17094 2174
rect 17048 1956 17054 2162
rect 17088 1956 17094 2162
rect 17130 1996 17140 2176
rect 17192 1996 17202 2176
rect 17240 2162 17286 2174
rect 17034 1776 17044 1956
rect 17096 1776 17106 1956
rect 17144 1786 17150 1996
rect 17184 1786 17190 1996
rect 17240 1956 17246 2162
rect 17280 1956 17286 2162
rect 17322 1996 17332 2176
rect 17384 1996 17394 2176
rect 17432 2162 17478 2174
rect 17048 1774 17094 1776
rect 17144 1774 17190 1786
rect 17226 1776 17236 1956
rect 17288 1776 17298 1956
rect 17336 1786 17342 1996
rect 17376 1786 17382 1996
rect 17432 1956 17438 2162
rect 17472 1956 17478 2162
rect 17514 1996 17524 2176
rect 17576 1996 17586 2176
rect 17624 2162 17670 2174
rect 17240 1774 17286 1776
rect 17336 1774 17382 1786
rect 17418 1776 17428 1956
rect 17480 1776 17490 1956
rect 17528 1786 17534 1996
rect 17568 1786 17574 1996
rect 17624 1956 17630 2162
rect 17664 1956 17670 2162
rect 17432 1774 17478 1776
rect 17528 1774 17574 1786
rect 17610 1776 17620 1956
rect 17672 1776 17682 1956
rect 17624 1774 17670 1776
rect 17090 1740 17148 1742
rect 17282 1740 17340 1742
rect 17474 1740 17532 1742
rect 17712 1740 17792 2204
rect 18088 2162 18134 2174
rect 18088 1956 18094 2162
rect 18128 1956 18134 2162
rect 18170 1996 18180 2176
rect 18232 1996 18242 2176
rect 18280 2162 18326 2174
rect 18074 1776 18084 1956
rect 18136 1776 18146 1956
rect 18184 1786 18190 1996
rect 18224 1786 18230 1996
rect 18280 1956 18286 2162
rect 18320 1956 18326 2162
rect 18362 1996 18372 2176
rect 18424 1996 18434 2176
rect 18472 2162 18518 2174
rect 18088 1774 18134 1776
rect 18184 1774 18230 1786
rect 18266 1776 18276 1956
rect 18328 1776 18338 1956
rect 18376 1786 18382 1996
rect 18416 1786 18422 1996
rect 18472 1956 18478 2162
rect 18512 1956 18518 2162
rect 18554 1996 18564 2176
rect 18616 1996 18626 2176
rect 18664 2162 18710 2174
rect 18280 1774 18326 1776
rect 18376 1774 18422 1786
rect 18458 1776 18468 1956
rect 18520 1776 18530 1956
rect 18568 1786 18574 1996
rect 18608 1786 18614 1996
rect 18664 1956 18670 2162
rect 18704 1956 18710 2162
rect 18472 1774 18518 1776
rect 18568 1774 18614 1786
rect 18650 1776 18660 1956
rect 18712 1776 18722 1956
rect 18664 1774 18710 1776
rect 18130 1740 18188 1742
rect 18322 1740 18380 1742
rect 18514 1740 18572 1742
rect 18752 1740 18832 2204
rect 11884 1736 12592 1740
rect 11884 1702 11902 1736
rect 11936 1702 12094 1736
rect 12128 1702 12286 1736
rect 12320 1702 12592 1736
rect 11884 1644 12592 1702
rect 12924 1736 13632 1740
rect 12924 1702 12942 1736
rect 12976 1702 13134 1736
rect 13168 1702 13326 1736
rect 13360 1702 13632 1736
rect 12924 1644 13632 1702
rect 13964 1736 14672 1740
rect 13964 1702 13982 1736
rect 14016 1702 14174 1736
rect 14208 1702 14366 1736
rect 14400 1702 14672 1736
rect 13964 1644 14672 1702
rect 15004 1736 15712 1740
rect 15004 1702 15022 1736
rect 15056 1702 15214 1736
rect 15248 1702 15406 1736
rect 15440 1702 15712 1736
rect 15004 1644 15712 1702
rect 16044 1736 16752 1740
rect 16044 1702 16062 1736
rect 16096 1702 16254 1736
rect 16288 1702 16446 1736
rect 16480 1702 16752 1736
rect 16044 1644 16752 1702
rect 17084 1736 17792 1740
rect 17084 1702 17102 1736
rect 17136 1702 17294 1736
rect 17328 1702 17486 1736
rect 17520 1702 17792 1736
rect 17084 1644 17792 1702
rect 18124 1736 18832 1740
rect 18124 1702 18142 1736
rect 18176 1702 18334 1736
rect 18368 1702 18526 1736
rect 18560 1702 18832 1736
rect 18124 1644 18832 1702
rect 12456 1468 12540 1644
rect 13496 1468 13580 1644
rect 14536 1468 14620 1644
rect 15576 1468 15660 1644
rect 16616 1468 16700 1644
rect 17656 1468 17740 1644
rect 18696 1468 18780 1644
rect 11892 1442 12708 1468
rect 11892 1408 11913 1442
rect 11947 1408 12031 1442
rect 12065 1408 12149 1442
rect 12183 1408 12267 1442
rect 12301 1408 12385 1442
rect 12419 1408 12503 1442
rect 12537 1408 12708 1442
rect 11892 1400 12708 1408
rect 12932 1442 13748 1468
rect 12932 1408 12953 1442
rect 12987 1408 13071 1442
rect 13105 1408 13189 1442
rect 13223 1408 13307 1442
rect 13341 1408 13425 1442
rect 13459 1408 13543 1442
rect 13577 1408 13748 1442
rect 12932 1400 13748 1408
rect 13972 1442 14788 1468
rect 13972 1408 13993 1442
rect 14027 1408 14111 1442
rect 14145 1408 14229 1442
rect 14263 1408 14347 1442
rect 14381 1408 14465 1442
rect 14499 1408 14583 1442
rect 14617 1408 14788 1442
rect 13972 1400 14788 1408
rect 15012 1442 15828 1468
rect 15012 1408 15033 1442
rect 15067 1408 15151 1442
rect 15185 1408 15269 1442
rect 15303 1408 15387 1442
rect 15421 1408 15505 1442
rect 15539 1408 15623 1442
rect 15657 1408 15828 1442
rect 15012 1400 15828 1408
rect 16052 1442 16868 1468
rect 16052 1408 16073 1442
rect 16107 1408 16191 1442
rect 16225 1408 16309 1442
rect 16343 1408 16427 1442
rect 16461 1408 16545 1442
rect 16579 1408 16663 1442
rect 16697 1408 16868 1442
rect 16052 1400 16868 1408
rect 17092 1442 17908 1468
rect 17092 1408 17113 1442
rect 17147 1408 17231 1442
rect 17265 1408 17349 1442
rect 17383 1408 17467 1442
rect 17501 1408 17585 1442
rect 17619 1408 17703 1442
rect 17737 1408 17908 1442
rect 17092 1400 17908 1408
rect 18132 1442 18948 1468
rect 18132 1408 18153 1442
rect 18187 1408 18271 1442
rect 18305 1408 18389 1442
rect 18423 1408 18507 1442
rect 18541 1408 18625 1442
rect 18659 1408 18743 1442
rect 18777 1408 18948 1442
rect 18132 1400 18948 1408
rect 11848 1358 11894 1370
rect 11848 1148 11854 1358
rect 11888 1148 11894 1358
rect 11954 1192 11964 1372
rect 12016 1192 12026 1372
rect 12084 1358 12130 1370
rect 11834 968 11844 1148
rect 11896 968 11906 1148
rect 11966 982 11972 1192
rect 12006 982 12012 1192
rect 12084 1148 12090 1358
rect 12124 1148 12130 1358
rect 12190 1192 12200 1372
rect 12252 1192 12262 1372
rect 12320 1358 12366 1370
rect 11966 970 12012 982
rect 12070 968 12080 1148
rect 12132 968 12142 1148
rect 12202 982 12208 1192
rect 12242 982 12248 1192
rect 12320 1148 12326 1358
rect 12360 1148 12366 1358
rect 12426 1192 12436 1372
rect 12488 1192 12498 1372
rect 12556 1358 12602 1370
rect 12202 970 12248 982
rect 12306 968 12316 1148
rect 12368 968 12378 1148
rect 12438 982 12444 1192
rect 12478 982 12484 1192
rect 12556 1148 12562 1358
rect 12596 1148 12602 1358
rect 12438 970 12484 982
rect 12542 968 12552 1148
rect 12604 968 12614 1148
rect 12644 940 12708 1400
rect 12888 1358 12934 1370
rect 12888 1148 12894 1358
rect 12928 1148 12934 1358
rect 12994 1192 13004 1372
rect 13056 1192 13066 1372
rect 13124 1358 13170 1370
rect 12874 968 12884 1148
rect 12936 968 12946 1148
rect 13006 982 13012 1192
rect 13046 982 13052 1192
rect 13124 1148 13130 1358
rect 13164 1148 13170 1358
rect 13230 1192 13240 1372
rect 13292 1192 13302 1372
rect 13360 1358 13406 1370
rect 13006 970 13052 982
rect 13110 968 13120 1148
rect 13172 968 13182 1148
rect 13242 982 13248 1192
rect 13282 982 13288 1192
rect 13360 1148 13366 1358
rect 13400 1148 13406 1358
rect 13466 1192 13476 1372
rect 13528 1192 13538 1372
rect 13596 1358 13642 1370
rect 13242 970 13288 982
rect 13346 968 13356 1148
rect 13408 968 13418 1148
rect 13478 982 13484 1192
rect 13518 982 13524 1192
rect 13596 1148 13602 1358
rect 13636 1148 13642 1358
rect 13478 970 13524 982
rect 13582 968 13592 1148
rect 13644 968 13654 1148
rect 13684 940 13748 1400
rect 13928 1358 13974 1370
rect 13928 1148 13934 1358
rect 13968 1148 13974 1358
rect 14034 1192 14044 1372
rect 14096 1192 14106 1372
rect 14164 1358 14210 1370
rect 13914 968 13924 1148
rect 13976 968 13986 1148
rect 14046 982 14052 1192
rect 14086 982 14092 1192
rect 14164 1148 14170 1358
rect 14204 1148 14210 1358
rect 14270 1192 14280 1372
rect 14332 1192 14342 1372
rect 14400 1358 14446 1370
rect 14046 970 14092 982
rect 14150 968 14160 1148
rect 14212 968 14222 1148
rect 14282 982 14288 1192
rect 14322 982 14328 1192
rect 14400 1148 14406 1358
rect 14440 1148 14446 1358
rect 14506 1192 14516 1372
rect 14568 1192 14578 1372
rect 14636 1358 14682 1370
rect 14282 970 14328 982
rect 14386 968 14396 1148
rect 14448 968 14458 1148
rect 14518 982 14524 1192
rect 14558 982 14564 1192
rect 14636 1148 14642 1358
rect 14676 1148 14682 1358
rect 14518 970 14564 982
rect 14622 968 14632 1148
rect 14684 968 14694 1148
rect 14724 940 14788 1400
rect 14968 1358 15014 1370
rect 14968 1148 14974 1358
rect 15008 1148 15014 1358
rect 15074 1192 15084 1372
rect 15136 1192 15146 1372
rect 15204 1358 15250 1370
rect 14954 968 14964 1148
rect 15016 968 15026 1148
rect 15086 982 15092 1192
rect 15126 982 15132 1192
rect 15204 1148 15210 1358
rect 15244 1148 15250 1358
rect 15310 1192 15320 1372
rect 15372 1192 15382 1372
rect 15440 1358 15486 1370
rect 15086 970 15132 982
rect 15190 968 15200 1148
rect 15252 968 15262 1148
rect 15322 982 15328 1192
rect 15362 982 15368 1192
rect 15440 1148 15446 1358
rect 15480 1148 15486 1358
rect 15546 1192 15556 1372
rect 15608 1192 15618 1372
rect 15676 1358 15722 1370
rect 15322 970 15368 982
rect 15426 968 15436 1148
rect 15488 968 15498 1148
rect 15558 982 15564 1192
rect 15598 982 15604 1192
rect 15676 1148 15682 1358
rect 15716 1148 15722 1358
rect 15558 970 15604 982
rect 15662 968 15672 1148
rect 15724 968 15734 1148
rect 15764 940 15828 1400
rect 16008 1358 16054 1370
rect 16008 1148 16014 1358
rect 16048 1148 16054 1358
rect 16114 1192 16124 1372
rect 16176 1192 16186 1372
rect 16244 1358 16290 1370
rect 15994 968 16004 1148
rect 16056 968 16066 1148
rect 16126 982 16132 1192
rect 16166 982 16172 1192
rect 16244 1148 16250 1358
rect 16284 1148 16290 1358
rect 16350 1192 16360 1372
rect 16412 1192 16422 1372
rect 16480 1358 16526 1370
rect 16126 970 16172 982
rect 16230 968 16240 1148
rect 16292 968 16302 1148
rect 16362 982 16368 1192
rect 16402 982 16408 1192
rect 16480 1148 16486 1358
rect 16520 1148 16526 1358
rect 16586 1192 16596 1372
rect 16648 1192 16658 1372
rect 16716 1358 16762 1370
rect 16362 970 16408 982
rect 16466 968 16476 1148
rect 16528 968 16538 1148
rect 16598 982 16604 1192
rect 16638 982 16644 1192
rect 16716 1148 16722 1358
rect 16756 1148 16762 1358
rect 16598 970 16644 982
rect 16702 968 16712 1148
rect 16764 968 16774 1148
rect 16804 940 16868 1400
rect 17048 1358 17094 1370
rect 17048 1148 17054 1358
rect 17088 1148 17094 1358
rect 17154 1192 17164 1372
rect 17216 1192 17226 1372
rect 17284 1358 17330 1370
rect 17034 968 17044 1148
rect 17096 968 17106 1148
rect 17166 982 17172 1192
rect 17206 982 17212 1192
rect 17284 1148 17290 1358
rect 17324 1148 17330 1358
rect 17390 1192 17400 1372
rect 17452 1192 17462 1372
rect 17520 1358 17566 1370
rect 17166 970 17212 982
rect 17270 968 17280 1148
rect 17332 968 17342 1148
rect 17402 982 17408 1192
rect 17442 982 17448 1192
rect 17520 1148 17526 1358
rect 17560 1148 17566 1358
rect 17626 1192 17636 1372
rect 17688 1192 17698 1372
rect 17756 1358 17802 1370
rect 17402 970 17448 982
rect 17506 968 17516 1148
rect 17568 968 17578 1148
rect 17638 982 17644 1192
rect 17678 982 17684 1192
rect 17756 1148 17762 1358
rect 17796 1148 17802 1358
rect 17638 970 17684 982
rect 17742 968 17752 1148
rect 17804 968 17814 1148
rect 17844 940 17908 1400
rect 18088 1358 18134 1370
rect 18088 1148 18094 1358
rect 18128 1148 18134 1358
rect 18194 1192 18204 1372
rect 18256 1192 18266 1372
rect 18324 1358 18370 1370
rect 18074 968 18084 1148
rect 18136 968 18146 1148
rect 18206 982 18212 1192
rect 18246 982 18252 1192
rect 18324 1148 18330 1358
rect 18364 1148 18370 1358
rect 18430 1192 18440 1372
rect 18492 1192 18502 1372
rect 18560 1358 18606 1370
rect 18206 970 18252 982
rect 18310 968 18320 1148
rect 18372 968 18382 1148
rect 18442 982 18448 1192
rect 18482 982 18488 1192
rect 18560 1148 18566 1358
rect 18600 1148 18606 1358
rect 18666 1192 18676 1372
rect 18728 1192 18738 1372
rect 18796 1358 18842 1370
rect 18442 970 18488 982
rect 18546 968 18556 1148
rect 18608 968 18618 1148
rect 18678 982 18684 1192
rect 18718 982 18724 1192
rect 18796 1148 18802 1358
rect 18836 1148 18842 1358
rect 18678 970 18724 982
rect 18782 968 18792 1148
rect 18844 968 18854 1148
rect 18884 940 18948 1400
rect 11896 932 12708 940
rect 11896 898 11913 932
rect 11947 898 12031 932
rect 12065 898 12149 932
rect 12183 898 12267 932
rect 12301 898 12385 932
rect 12419 898 12503 932
rect 12537 898 12708 932
rect 11896 872 12708 898
rect 12936 932 13748 940
rect 12936 898 12953 932
rect 12987 898 13071 932
rect 13105 898 13189 932
rect 13223 898 13307 932
rect 13341 898 13425 932
rect 13459 898 13543 932
rect 13577 898 13748 932
rect 12936 872 13748 898
rect 13976 932 14788 940
rect 13976 898 13993 932
rect 14027 898 14111 932
rect 14145 898 14229 932
rect 14263 898 14347 932
rect 14381 898 14465 932
rect 14499 898 14583 932
rect 14617 898 14788 932
rect 13976 872 14788 898
rect 15016 932 15828 940
rect 15016 898 15033 932
rect 15067 898 15151 932
rect 15185 898 15269 932
rect 15303 898 15387 932
rect 15421 898 15505 932
rect 15539 898 15623 932
rect 15657 898 15828 932
rect 15016 872 15828 898
rect 16056 932 16868 940
rect 16056 898 16073 932
rect 16107 898 16191 932
rect 16225 898 16309 932
rect 16343 898 16427 932
rect 16461 898 16545 932
rect 16579 898 16663 932
rect 16697 898 16868 932
rect 16056 872 16868 898
rect 17096 932 17908 940
rect 17096 898 17113 932
rect 17147 898 17231 932
rect 17265 898 17349 932
rect 17383 898 17467 932
rect 17501 898 17585 932
rect 17619 898 17703 932
rect 17737 898 17908 932
rect 17096 872 17908 898
rect 18136 932 18948 940
rect 18136 898 18153 932
rect 18187 898 18271 932
rect 18305 898 18389 932
rect 18423 898 18507 932
rect 18541 898 18625 932
rect 18659 898 18743 932
rect 18777 898 18948 932
rect 18136 872 18948 898
rect 11880 624 12592 668
rect 11880 590 11902 624
rect 11936 590 12094 624
rect 12128 590 12286 624
rect 12320 590 12592 624
rect 11880 584 12592 590
rect 12920 624 13632 668
rect 12920 590 12942 624
rect 12976 590 13134 624
rect 13168 590 13326 624
rect 13360 590 13632 624
rect 12920 584 13632 590
rect 13960 624 14672 668
rect 13960 590 13982 624
rect 14016 590 14174 624
rect 14208 590 14366 624
rect 14400 590 14672 624
rect 13960 584 14672 590
rect 15000 624 15712 668
rect 15000 590 15022 624
rect 15056 590 15214 624
rect 15248 590 15406 624
rect 15440 590 15712 624
rect 15000 584 15712 590
rect 16040 624 16752 668
rect 16040 590 16062 624
rect 16096 590 16254 624
rect 16288 590 16446 624
rect 16480 590 16752 624
rect 16040 584 16752 590
rect 17080 624 17792 668
rect 17080 590 17102 624
rect 17136 590 17294 624
rect 17328 590 17486 624
rect 17520 590 17792 624
rect 17080 584 17792 590
rect 18120 624 18832 668
rect 18120 590 18142 624
rect 18176 590 18334 624
rect 18368 590 18526 624
rect 18560 590 18832 624
rect 18120 584 18832 590
rect 11834 372 11844 552
rect 11896 372 11906 552
rect 11944 540 11990 552
rect 11848 164 11854 372
rect 11888 164 11894 372
rect 11944 332 11950 540
rect 11984 332 11990 540
rect 12026 372 12036 552
rect 12088 372 12098 552
rect 12136 540 12182 552
rect 11848 152 11894 164
rect 11930 152 11940 332
rect 11992 152 12002 332
rect 12040 164 12046 372
rect 12080 164 12086 372
rect 12136 332 12142 540
rect 12176 332 12182 540
rect 12218 372 12228 552
rect 12280 372 12290 552
rect 12328 540 12374 552
rect 12040 152 12086 164
rect 12122 152 12132 332
rect 12184 152 12194 332
rect 12232 164 12238 372
rect 12272 164 12278 372
rect 12328 332 12334 540
rect 12368 332 12374 540
rect 12410 372 12420 552
rect 12472 372 12482 552
rect 12232 152 12278 164
rect 12314 152 12324 332
rect 12376 152 12386 332
rect 12424 164 12430 372
rect 12464 164 12470 372
rect 12424 152 12470 164
rect 12512 120 12592 584
rect 12874 372 12884 552
rect 12936 372 12946 552
rect 12984 540 13030 552
rect 12888 164 12894 372
rect 12928 164 12934 372
rect 12984 332 12990 540
rect 13024 332 13030 540
rect 13066 372 13076 552
rect 13128 372 13138 552
rect 13176 540 13222 552
rect 12888 152 12934 164
rect 12970 152 12980 332
rect 13032 152 13042 332
rect 13080 164 13086 372
rect 13120 164 13126 372
rect 13176 332 13182 540
rect 13216 332 13222 540
rect 13258 372 13268 552
rect 13320 372 13330 552
rect 13368 540 13414 552
rect 13080 152 13126 164
rect 13162 152 13172 332
rect 13224 152 13234 332
rect 13272 164 13278 372
rect 13312 164 13318 372
rect 13368 332 13374 540
rect 13408 332 13414 540
rect 13450 372 13460 552
rect 13512 372 13522 552
rect 13272 152 13318 164
rect 13354 152 13364 332
rect 13416 152 13426 332
rect 13464 164 13470 372
rect 13504 164 13510 372
rect 13464 152 13510 164
rect 13552 120 13632 584
rect 13914 372 13924 552
rect 13976 372 13986 552
rect 14024 540 14070 552
rect 13928 164 13934 372
rect 13968 164 13974 372
rect 14024 332 14030 540
rect 14064 332 14070 540
rect 14106 372 14116 552
rect 14168 372 14178 552
rect 14216 540 14262 552
rect 13928 152 13974 164
rect 14010 152 14020 332
rect 14072 152 14082 332
rect 14120 164 14126 372
rect 14160 164 14166 372
rect 14216 332 14222 540
rect 14256 332 14262 540
rect 14298 372 14308 552
rect 14360 372 14370 552
rect 14408 540 14454 552
rect 14120 152 14166 164
rect 14202 152 14212 332
rect 14264 152 14274 332
rect 14312 164 14318 372
rect 14352 164 14358 372
rect 14408 332 14414 540
rect 14448 332 14454 540
rect 14490 372 14500 552
rect 14552 372 14562 552
rect 14312 152 14358 164
rect 14394 152 14404 332
rect 14456 152 14466 332
rect 14504 164 14510 372
rect 14544 164 14550 372
rect 14504 152 14550 164
rect 14592 120 14672 584
rect 14954 372 14964 552
rect 15016 372 15026 552
rect 15064 540 15110 552
rect 14968 164 14974 372
rect 15008 164 15014 372
rect 15064 332 15070 540
rect 15104 332 15110 540
rect 15146 372 15156 552
rect 15208 372 15218 552
rect 15256 540 15302 552
rect 14968 152 15014 164
rect 15050 152 15060 332
rect 15112 152 15122 332
rect 15160 164 15166 372
rect 15200 164 15206 372
rect 15256 332 15262 540
rect 15296 332 15302 540
rect 15338 372 15348 552
rect 15400 372 15410 552
rect 15448 540 15494 552
rect 15160 152 15206 164
rect 15242 152 15252 332
rect 15304 152 15314 332
rect 15352 164 15358 372
rect 15392 164 15398 372
rect 15448 332 15454 540
rect 15488 332 15494 540
rect 15530 372 15540 552
rect 15592 372 15602 552
rect 15352 152 15398 164
rect 15434 152 15444 332
rect 15496 152 15506 332
rect 15544 164 15550 372
rect 15584 164 15590 372
rect 15544 152 15590 164
rect 15632 120 15712 584
rect 15994 372 16004 552
rect 16056 372 16066 552
rect 16104 540 16150 552
rect 16008 164 16014 372
rect 16048 164 16054 372
rect 16104 332 16110 540
rect 16144 332 16150 540
rect 16186 372 16196 552
rect 16248 372 16258 552
rect 16296 540 16342 552
rect 16008 152 16054 164
rect 16090 152 16100 332
rect 16152 152 16162 332
rect 16200 164 16206 372
rect 16240 164 16246 372
rect 16296 332 16302 540
rect 16336 332 16342 540
rect 16378 372 16388 552
rect 16440 372 16450 552
rect 16488 540 16534 552
rect 16200 152 16246 164
rect 16282 152 16292 332
rect 16344 152 16354 332
rect 16392 164 16398 372
rect 16432 164 16438 372
rect 16488 332 16494 540
rect 16528 332 16534 540
rect 16570 372 16580 552
rect 16632 372 16642 552
rect 16392 152 16438 164
rect 16474 152 16484 332
rect 16536 152 16546 332
rect 16584 164 16590 372
rect 16624 164 16630 372
rect 16584 152 16630 164
rect 16672 120 16752 584
rect 17034 372 17044 552
rect 17096 372 17106 552
rect 17144 540 17190 552
rect 17048 164 17054 372
rect 17088 164 17094 372
rect 17144 332 17150 540
rect 17184 332 17190 540
rect 17226 372 17236 552
rect 17288 372 17298 552
rect 17336 540 17382 552
rect 17048 152 17094 164
rect 17130 152 17140 332
rect 17192 152 17202 332
rect 17240 164 17246 372
rect 17280 164 17286 372
rect 17336 332 17342 540
rect 17376 332 17382 540
rect 17418 372 17428 552
rect 17480 372 17490 552
rect 17528 540 17574 552
rect 17240 152 17286 164
rect 17322 152 17332 332
rect 17384 152 17394 332
rect 17432 164 17438 372
rect 17472 164 17478 372
rect 17528 332 17534 540
rect 17568 332 17574 540
rect 17610 372 17620 552
rect 17672 372 17682 552
rect 17432 152 17478 164
rect 17514 152 17524 332
rect 17576 152 17586 332
rect 17624 164 17630 372
rect 17664 164 17670 372
rect 17624 152 17670 164
rect 17712 120 17792 584
rect 18074 372 18084 552
rect 18136 372 18146 552
rect 18184 540 18230 552
rect 18088 164 18094 372
rect 18128 164 18134 372
rect 18184 332 18190 540
rect 18224 332 18230 540
rect 18266 372 18276 552
rect 18328 372 18338 552
rect 18376 540 18422 552
rect 18088 152 18134 164
rect 18170 152 18180 332
rect 18232 152 18242 332
rect 18280 164 18286 372
rect 18320 164 18326 372
rect 18376 332 18382 540
rect 18416 332 18422 540
rect 18458 372 18468 552
rect 18520 372 18530 552
rect 18568 540 18614 552
rect 18280 152 18326 164
rect 18362 152 18372 332
rect 18424 152 18434 332
rect 18472 164 18478 372
rect 18512 164 18518 372
rect 18568 332 18574 540
rect 18608 332 18614 540
rect 18650 372 18660 552
rect 18712 372 18722 552
rect 18472 152 18518 164
rect 18554 152 18564 332
rect 18616 152 18626 332
rect 18664 164 18670 372
rect 18704 164 18710 372
rect 18664 152 18710 164
rect 18752 120 18832 584
rect 11940 114 12592 120
rect 11940 100 11998 114
rect 11620 80 11998 100
rect 12032 80 12190 114
rect 12224 80 12382 114
rect 12416 100 12592 114
rect 12980 114 13632 120
rect 12980 100 13038 114
rect 12416 80 13038 100
rect 13072 80 13230 114
rect 13264 80 13422 114
rect 13456 100 13632 114
rect 14020 114 14672 120
rect 14020 100 14078 114
rect 13456 80 14078 100
rect 14112 80 14270 114
rect 14304 80 14462 114
rect 14496 100 14672 114
rect 15060 114 15712 120
rect 15060 100 15118 114
rect 14496 80 15118 100
rect 15152 80 15310 114
rect 15344 80 15502 114
rect 15536 100 15712 114
rect 16100 114 16752 120
rect 16100 100 16158 114
rect 15536 80 16158 100
rect 16192 80 16350 114
rect 16384 80 16542 114
rect 16576 100 16752 114
rect 17140 114 17792 120
rect 17140 100 17198 114
rect 16576 80 17198 100
rect 17232 80 17390 114
rect 17424 80 17582 114
rect 17616 100 17792 114
rect 18180 114 18832 120
rect 18180 100 18238 114
rect 17616 80 18238 100
rect 18272 80 18430 114
rect 18464 80 18622 114
rect 18656 80 18832 114
rect 11620 6 18832 80
rect 11620 -16 11998 6
rect 4836 -772 4920 -596
rect 5876 -772 5960 -596
rect 6916 -772 7000 -596
rect 7956 -772 8040 -596
rect 8996 -772 9080 -596
rect 10036 -772 10120 -596
rect 11076 -772 11160 -596
rect 4272 -798 5088 -772
rect 4272 -832 4293 -798
rect 4327 -832 4411 -798
rect 4445 -832 4529 -798
rect 4563 -832 4647 -798
rect 4681 -832 4765 -798
rect 4799 -832 4883 -798
rect 4917 -832 5088 -798
rect 4272 -840 5088 -832
rect 5312 -798 6128 -772
rect 5312 -832 5333 -798
rect 5367 -832 5451 -798
rect 5485 -832 5569 -798
rect 5603 -832 5687 -798
rect 5721 -832 5805 -798
rect 5839 -832 5923 -798
rect 5957 -832 6128 -798
rect 5312 -840 6128 -832
rect 6352 -798 7168 -772
rect 6352 -832 6373 -798
rect 6407 -832 6491 -798
rect 6525 -832 6609 -798
rect 6643 -832 6727 -798
rect 6761 -832 6845 -798
rect 6879 -832 6963 -798
rect 6997 -832 7168 -798
rect 6352 -840 7168 -832
rect 7392 -798 8208 -772
rect 7392 -832 7413 -798
rect 7447 -832 7531 -798
rect 7565 -832 7649 -798
rect 7683 -832 7767 -798
rect 7801 -832 7885 -798
rect 7919 -832 8003 -798
rect 8037 -832 8208 -798
rect 7392 -840 8208 -832
rect 8432 -798 9248 -772
rect 8432 -832 8453 -798
rect 8487 -832 8571 -798
rect 8605 -832 8689 -798
rect 8723 -832 8807 -798
rect 8841 -832 8925 -798
rect 8959 -832 9043 -798
rect 9077 -832 9248 -798
rect 8432 -840 9248 -832
rect 9472 -798 10288 -772
rect 9472 -832 9493 -798
rect 9527 -832 9611 -798
rect 9645 -832 9729 -798
rect 9763 -832 9847 -798
rect 9881 -832 9965 -798
rect 9999 -832 10083 -798
rect 10117 -832 10288 -798
rect 9472 -840 10288 -832
rect 10512 -798 11328 -772
rect 10512 -832 10533 -798
rect 10567 -832 10651 -798
rect 10685 -832 10769 -798
rect 10803 -832 10887 -798
rect 10921 -832 11005 -798
rect 11039 -832 11123 -798
rect 11157 -832 11328 -798
rect 10512 -840 11328 -832
rect 4228 -882 4274 -870
rect 4228 -1092 4234 -882
rect 4268 -1092 4274 -882
rect 4334 -1048 4344 -868
rect 4396 -1048 4406 -868
rect 4464 -882 4510 -870
rect 4214 -1272 4224 -1092
rect 4276 -1272 4286 -1092
rect 4346 -1258 4352 -1048
rect 4386 -1258 4392 -1048
rect 4464 -1092 4470 -882
rect 4504 -1092 4510 -882
rect 4570 -1048 4580 -868
rect 4632 -1048 4642 -868
rect 4700 -882 4746 -870
rect 4346 -1270 4392 -1258
rect 4450 -1272 4460 -1092
rect 4512 -1272 4522 -1092
rect 4582 -1258 4588 -1048
rect 4622 -1258 4628 -1048
rect 4700 -1092 4706 -882
rect 4740 -1092 4746 -882
rect 4806 -1048 4816 -868
rect 4868 -1048 4878 -868
rect 4936 -882 4982 -870
rect 4582 -1270 4628 -1258
rect 4686 -1272 4696 -1092
rect 4748 -1272 4758 -1092
rect 4818 -1258 4824 -1048
rect 4858 -1258 4864 -1048
rect 4936 -1092 4942 -882
rect 4976 -1092 4982 -882
rect 4818 -1270 4864 -1258
rect 4922 -1272 4932 -1092
rect 4984 -1272 4994 -1092
rect 5024 -1300 5088 -840
rect 5268 -882 5314 -870
rect 5268 -1092 5274 -882
rect 5308 -1092 5314 -882
rect 5374 -1048 5384 -868
rect 5436 -1048 5446 -868
rect 5504 -882 5550 -870
rect 5254 -1272 5264 -1092
rect 5316 -1272 5326 -1092
rect 5386 -1258 5392 -1048
rect 5426 -1258 5432 -1048
rect 5504 -1092 5510 -882
rect 5544 -1092 5550 -882
rect 5610 -1048 5620 -868
rect 5672 -1048 5682 -868
rect 5740 -882 5786 -870
rect 5386 -1270 5432 -1258
rect 5490 -1272 5500 -1092
rect 5552 -1272 5562 -1092
rect 5622 -1258 5628 -1048
rect 5662 -1258 5668 -1048
rect 5740 -1092 5746 -882
rect 5780 -1092 5786 -882
rect 5846 -1048 5856 -868
rect 5908 -1048 5918 -868
rect 5976 -882 6022 -870
rect 5622 -1270 5668 -1258
rect 5726 -1272 5736 -1092
rect 5788 -1272 5798 -1092
rect 5858 -1258 5864 -1048
rect 5898 -1258 5904 -1048
rect 5976 -1092 5982 -882
rect 6016 -1092 6022 -882
rect 5858 -1270 5904 -1258
rect 5962 -1272 5972 -1092
rect 6024 -1272 6034 -1092
rect 6064 -1300 6128 -840
rect 6308 -882 6354 -870
rect 6308 -1092 6314 -882
rect 6348 -1092 6354 -882
rect 6414 -1048 6424 -868
rect 6476 -1048 6486 -868
rect 6544 -882 6590 -870
rect 6294 -1272 6304 -1092
rect 6356 -1272 6366 -1092
rect 6426 -1258 6432 -1048
rect 6466 -1258 6472 -1048
rect 6544 -1092 6550 -882
rect 6584 -1092 6590 -882
rect 6650 -1048 6660 -868
rect 6712 -1048 6722 -868
rect 6780 -882 6826 -870
rect 6426 -1270 6472 -1258
rect 6530 -1272 6540 -1092
rect 6592 -1272 6602 -1092
rect 6662 -1258 6668 -1048
rect 6702 -1258 6708 -1048
rect 6780 -1092 6786 -882
rect 6820 -1092 6826 -882
rect 6886 -1048 6896 -868
rect 6948 -1048 6958 -868
rect 7016 -882 7062 -870
rect 6662 -1270 6708 -1258
rect 6766 -1272 6776 -1092
rect 6828 -1272 6838 -1092
rect 6898 -1258 6904 -1048
rect 6938 -1258 6944 -1048
rect 7016 -1092 7022 -882
rect 7056 -1092 7062 -882
rect 6898 -1270 6944 -1258
rect 7002 -1272 7012 -1092
rect 7064 -1272 7074 -1092
rect 7104 -1300 7168 -840
rect 7348 -882 7394 -870
rect 7348 -1092 7354 -882
rect 7388 -1092 7394 -882
rect 7454 -1048 7464 -868
rect 7516 -1048 7526 -868
rect 7584 -882 7630 -870
rect 7334 -1272 7344 -1092
rect 7396 -1272 7406 -1092
rect 7466 -1258 7472 -1048
rect 7506 -1258 7512 -1048
rect 7584 -1092 7590 -882
rect 7624 -1092 7630 -882
rect 7690 -1048 7700 -868
rect 7752 -1048 7762 -868
rect 7820 -882 7866 -870
rect 7466 -1270 7512 -1258
rect 7570 -1272 7580 -1092
rect 7632 -1272 7642 -1092
rect 7702 -1258 7708 -1048
rect 7742 -1258 7748 -1048
rect 7820 -1092 7826 -882
rect 7860 -1092 7866 -882
rect 7926 -1048 7936 -868
rect 7988 -1048 7998 -868
rect 8056 -882 8102 -870
rect 7702 -1270 7748 -1258
rect 7806 -1272 7816 -1092
rect 7868 -1272 7878 -1092
rect 7938 -1258 7944 -1048
rect 7978 -1258 7984 -1048
rect 8056 -1092 8062 -882
rect 8096 -1092 8102 -882
rect 7938 -1270 7984 -1258
rect 8042 -1272 8052 -1092
rect 8104 -1272 8114 -1092
rect 8144 -1300 8208 -840
rect 8388 -882 8434 -870
rect 8388 -1092 8394 -882
rect 8428 -1092 8434 -882
rect 8494 -1048 8504 -868
rect 8556 -1048 8566 -868
rect 8624 -882 8670 -870
rect 8374 -1272 8384 -1092
rect 8436 -1272 8446 -1092
rect 8506 -1258 8512 -1048
rect 8546 -1258 8552 -1048
rect 8624 -1092 8630 -882
rect 8664 -1092 8670 -882
rect 8730 -1048 8740 -868
rect 8792 -1048 8802 -868
rect 8860 -882 8906 -870
rect 8506 -1270 8552 -1258
rect 8610 -1272 8620 -1092
rect 8672 -1272 8682 -1092
rect 8742 -1258 8748 -1048
rect 8782 -1258 8788 -1048
rect 8860 -1092 8866 -882
rect 8900 -1092 8906 -882
rect 8966 -1048 8976 -868
rect 9028 -1048 9038 -868
rect 9096 -882 9142 -870
rect 8742 -1270 8788 -1258
rect 8846 -1272 8856 -1092
rect 8908 -1272 8918 -1092
rect 8978 -1258 8984 -1048
rect 9018 -1258 9024 -1048
rect 9096 -1092 9102 -882
rect 9136 -1092 9142 -882
rect 8978 -1270 9024 -1258
rect 9082 -1272 9092 -1092
rect 9144 -1272 9154 -1092
rect 9184 -1300 9248 -840
rect 9428 -882 9474 -870
rect 9428 -1092 9434 -882
rect 9468 -1092 9474 -882
rect 9534 -1048 9544 -868
rect 9596 -1048 9606 -868
rect 9664 -882 9710 -870
rect 9414 -1272 9424 -1092
rect 9476 -1272 9486 -1092
rect 9546 -1258 9552 -1048
rect 9586 -1258 9592 -1048
rect 9664 -1092 9670 -882
rect 9704 -1092 9710 -882
rect 9770 -1048 9780 -868
rect 9832 -1048 9842 -868
rect 9900 -882 9946 -870
rect 9546 -1270 9592 -1258
rect 9650 -1272 9660 -1092
rect 9712 -1272 9722 -1092
rect 9782 -1258 9788 -1048
rect 9822 -1258 9828 -1048
rect 9900 -1092 9906 -882
rect 9940 -1092 9946 -882
rect 10006 -1048 10016 -868
rect 10068 -1048 10078 -868
rect 10136 -882 10182 -870
rect 9782 -1270 9828 -1258
rect 9886 -1272 9896 -1092
rect 9948 -1272 9958 -1092
rect 10018 -1258 10024 -1048
rect 10058 -1258 10064 -1048
rect 10136 -1092 10142 -882
rect 10176 -1092 10182 -882
rect 10018 -1270 10064 -1258
rect 10122 -1272 10132 -1092
rect 10184 -1272 10194 -1092
rect 10224 -1300 10288 -840
rect 10468 -882 10514 -870
rect 10468 -1092 10474 -882
rect 10508 -1092 10514 -882
rect 10574 -1048 10584 -868
rect 10636 -1048 10646 -868
rect 10704 -882 10750 -870
rect 10454 -1272 10464 -1092
rect 10516 -1272 10526 -1092
rect 10586 -1258 10592 -1048
rect 10626 -1258 10632 -1048
rect 10704 -1092 10710 -882
rect 10744 -1092 10750 -882
rect 10810 -1048 10820 -868
rect 10872 -1048 10882 -868
rect 10940 -882 10986 -870
rect 10586 -1270 10632 -1258
rect 10690 -1272 10700 -1092
rect 10752 -1272 10762 -1092
rect 10822 -1258 10828 -1048
rect 10862 -1258 10868 -1048
rect 10940 -1092 10946 -882
rect 10980 -1092 10986 -882
rect 11046 -1048 11056 -868
rect 11108 -1048 11118 -868
rect 11176 -882 11222 -870
rect 10822 -1270 10868 -1258
rect 10926 -1272 10936 -1092
rect 10988 -1272 10998 -1092
rect 11058 -1258 11064 -1048
rect 11098 -1258 11104 -1048
rect 11176 -1092 11182 -882
rect 11216 -1092 11222 -882
rect 11058 -1270 11104 -1258
rect 11162 -1272 11172 -1092
rect 11224 -1272 11234 -1092
rect 11264 -1300 11328 -840
rect 4276 -1308 5088 -1300
rect 4276 -1342 4293 -1308
rect 4327 -1342 4411 -1308
rect 4445 -1342 4529 -1308
rect 4563 -1342 4647 -1308
rect 4681 -1342 4765 -1308
rect 4799 -1342 4883 -1308
rect 4917 -1342 5088 -1308
rect 4276 -1368 5088 -1342
rect 5316 -1308 6128 -1300
rect 5316 -1342 5333 -1308
rect 5367 -1342 5451 -1308
rect 5485 -1342 5569 -1308
rect 5603 -1342 5687 -1308
rect 5721 -1342 5805 -1308
rect 5839 -1342 5923 -1308
rect 5957 -1342 6128 -1308
rect 5316 -1368 6128 -1342
rect 6356 -1308 7168 -1300
rect 6356 -1342 6373 -1308
rect 6407 -1342 6491 -1308
rect 6525 -1342 6609 -1308
rect 6643 -1342 6727 -1308
rect 6761 -1342 6845 -1308
rect 6879 -1342 6963 -1308
rect 6997 -1342 7168 -1308
rect 6356 -1368 7168 -1342
rect 7396 -1308 8208 -1300
rect 7396 -1342 7413 -1308
rect 7447 -1342 7531 -1308
rect 7565 -1342 7649 -1308
rect 7683 -1342 7767 -1308
rect 7801 -1342 7885 -1308
rect 7919 -1342 8003 -1308
rect 8037 -1342 8208 -1308
rect 7396 -1368 8208 -1342
rect 8436 -1308 9248 -1300
rect 8436 -1342 8453 -1308
rect 8487 -1342 8571 -1308
rect 8605 -1342 8689 -1308
rect 8723 -1342 8807 -1308
rect 8841 -1342 8925 -1308
rect 8959 -1342 9043 -1308
rect 9077 -1342 9248 -1308
rect 8436 -1368 9248 -1342
rect 9476 -1308 10288 -1300
rect 9476 -1342 9493 -1308
rect 9527 -1342 9611 -1308
rect 9645 -1342 9729 -1308
rect 9763 -1342 9847 -1308
rect 9881 -1342 9965 -1308
rect 9999 -1342 10083 -1308
rect 10117 -1342 10288 -1308
rect 9476 -1368 10288 -1342
rect 10516 -1308 11328 -1300
rect 10516 -1342 10533 -1308
rect 10567 -1342 10651 -1308
rect 10685 -1342 10769 -1308
rect 10803 -1342 10887 -1308
rect 10921 -1342 11005 -1308
rect 11039 -1342 11123 -1308
rect 11157 -1342 11328 -1308
rect 10516 -1368 11328 -1342
rect 4260 -1616 4972 -1572
rect 4260 -1650 4282 -1616
rect 4316 -1650 4474 -1616
rect 4508 -1650 4666 -1616
rect 4700 -1650 4972 -1616
rect 4260 -1656 4972 -1650
rect 5300 -1616 6012 -1572
rect 5300 -1650 5322 -1616
rect 5356 -1650 5514 -1616
rect 5548 -1650 5706 -1616
rect 5740 -1650 6012 -1616
rect 5300 -1656 6012 -1650
rect 6340 -1616 7052 -1572
rect 6340 -1650 6362 -1616
rect 6396 -1650 6554 -1616
rect 6588 -1650 6746 -1616
rect 6780 -1650 7052 -1616
rect 6340 -1656 7052 -1650
rect 7380 -1616 8092 -1572
rect 7380 -1650 7402 -1616
rect 7436 -1650 7594 -1616
rect 7628 -1650 7786 -1616
rect 7820 -1650 8092 -1616
rect 7380 -1656 8092 -1650
rect 8420 -1616 9132 -1572
rect 8420 -1650 8442 -1616
rect 8476 -1650 8634 -1616
rect 8668 -1650 8826 -1616
rect 8860 -1650 9132 -1616
rect 8420 -1656 9132 -1650
rect 4214 -1868 4224 -1688
rect 4276 -1868 4286 -1688
rect 4324 -1700 4370 -1688
rect 4228 -2076 4234 -1868
rect 4268 -2076 4274 -1868
rect 4324 -1908 4330 -1700
rect 4364 -1908 4370 -1700
rect 4406 -1868 4416 -1688
rect 4468 -1868 4478 -1688
rect 4516 -1700 4562 -1688
rect 4228 -2088 4274 -2076
rect 4310 -2088 4320 -1908
rect 4372 -2088 4382 -1908
rect 4420 -2076 4426 -1868
rect 4460 -2076 4466 -1868
rect 4516 -1908 4522 -1700
rect 4556 -1908 4562 -1700
rect 4598 -1868 4608 -1688
rect 4660 -1868 4670 -1688
rect 4708 -1700 4754 -1688
rect 4420 -2088 4466 -2076
rect 4502 -2088 4512 -1908
rect 4564 -2088 4574 -1908
rect 4612 -2076 4618 -1868
rect 4652 -2076 4658 -1868
rect 4708 -1908 4714 -1700
rect 4748 -1908 4754 -1700
rect 4790 -1868 4800 -1688
rect 4852 -1868 4862 -1688
rect 4612 -2088 4658 -2076
rect 4694 -2088 4704 -1908
rect 4756 -2088 4766 -1908
rect 4804 -2076 4810 -1868
rect 4844 -2076 4850 -1868
rect 4804 -2088 4850 -2076
rect 4892 -2120 4972 -1656
rect 5254 -1868 5264 -1688
rect 5316 -1868 5326 -1688
rect 5364 -1700 5410 -1688
rect 5268 -2076 5274 -1868
rect 5308 -2076 5314 -1868
rect 5364 -1908 5370 -1700
rect 5404 -1908 5410 -1700
rect 5446 -1868 5456 -1688
rect 5508 -1868 5518 -1688
rect 5556 -1700 5602 -1688
rect 5268 -2088 5314 -2076
rect 5350 -2088 5360 -1908
rect 5412 -2088 5422 -1908
rect 5460 -2076 5466 -1868
rect 5500 -2076 5506 -1868
rect 5556 -1908 5562 -1700
rect 5596 -1908 5602 -1700
rect 5638 -1868 5648 -1688
rect 5700 -1868 5710 -1688
rect 5748 -1700 5794 -1688
rect 5460 -2088 5506 -2076
rect 5542 -2088 5552 -1908
rect 5604 -2088 5614 -1908
rect 5652 -2076 5658 -1868
rect 5692 -2076 5698 -1868
rect 5748 -1908 5754 -1700
rect 5788 -1908 5794 -1700
rect 5830 -1868 5840 -1688
rect 5892 -1868 5902 -1688
rect 5652 -2088 5698 -2076
rect 5734 -2088 5744 -1908
rect 5796 -2088 5806 -1908
rect 5844 -2076 5850 -1868
rect 5884 -2076 5890 -1868
rect 5844 -2088 5890 -2076
rect 5932 -2120 6012 -1656
rect 6294 -1868 6304 -1688
rect 6356 -1868 6366 -1688
rect 6404 -1700 6450 -1688
rect 6308 -2076 6314 -1868
rect 6348 -2076 6354 -1868
rect 6404 -1908 6410 -1700
rect 6444 -1908 6450 -1700
rect 6486 -1868 6496 -1688
rect 6548 -1868 6558 -1688
rect 6596 -1700 6642 -1688
rect 6308 -2088 6354 -2076
rect 6390 -2088 6400 -1908
rect 6452 -2088 6462 -1908
rect 6500 -2076 6506 -1868
rect 6540 -2076 6546 -1868
rect 6596 -1908 6602 -1700
rect 6636 -1908 6642 -1700
rect 6678 -1868 6688 -1688
rect 6740 -1868 6750 -1688
rect 6788 -1700 6834 -1688
rect 6500 -2088 6546 -2076
rect 6582 -2088 6592 -1908
rect 6644 -2088 6654 -1908
rect 6692 -2076 6698 -1868
rect 6732 -2076 6738 -1868
rect 6788 -1908 6794 -1700
rect 6828 -1908 6834 -1700
rect 6870 -1868 6880 -1688
rect 6932 -1868 6942 -1688
rect 6692 -2088 6738 -2076
rect 6774 -2088 6784 -1908
rect 6836 -2088 6846 -1908
rect 6884 -2076 6890 -1868
rect 6924 -2076 6930 -1868
rect 6884 -2088 6930 -2076
rect 6972 -2120 7052 -1656
rect 7334 -1868 7344 -1688
rect 7396 -1868 7406 -1688
rect 7444 -1700 7490 -1688
rect 7348 -2076 7354 -1868
rect 7388 -2076 7394 -1868
rect 7444 -1908 7450 -1700
rect 7484 -1908 7490 -1700
rect 7526 -1868 7536 -1688
rect 7588 -1868 7598 -1688
rect 7636 -1700 7682 -1688
rect 7348 -2088 7394 -2076
rect 7430 -2088 7440 -1908
rect 7492 -2088 7502 -1908
rect 7540 -2076 7546 -1868
rect 7580 -2076 7586 -1868
rect 7636 -1908 7642 -1700
rect 7676 -1908 7682 -1700
rect 7718 -1868 7728 -1688
rect 7780 -1868 7790 -1688
rect 7828 -1700 7874 -1688
rect 7540 -2088 7586 -2076
rect 7622 -2088 7632 -1908
rect 7684 -2088 7694 -1908
rect 7732 -2076 7738 -1868
rect 7772 -2076 7778 -1868
rect 7828 -1908 7834 -1700
rect 7868 -1908 7874 -1700
rect 7910 -1868 7920 -1688
rect 7972 -1868 7982 -1688
rect 7732 -2088 7778 -2076
rect 7814 -2088 7824 -1908
rect 7876 -2088 7886 -1908
rect 7924 -2076 7930 -1868
rect 7964 -2076 7970 -1868
rect 7924 -2088 7970 -2076
rect 8012 -2120 8092 -1656
rect 8374 -1868 8384 -1688
rect 8436 -1868 8446 -1688
rect 8484 -1700 8530 -1688
rect 8388 -2076 8394 -1868
rect 8428 -2076 8434 -1868
rect 8484 -1908 8490 -1700
rect 8524 -1908 8530 -1700
rect 8566 -1868 8576 -1688
rect 8628 -1868 8638 -1688
rect 8676 -1700 8722 -1688
rect 8388 -2088 8434 -2076
rect 8470 -2088 8480 -1908
rect 8532 -2088 8542 -1908
rect 8580 -2076 8586 -1868
rect 8620 -2076 8626 -1868
rect 8676 -1908 8682 -1700
rect 8716 -1908 8722 -1700
rect 8758 -1868 8768 -1688
rect 8820 -1868 8830 -1688
rect 8868 -1700 8914 -1688
rect 8580 -2088 8626 -2076
rect 8662 -2088 8672 -1908
rect 8724 -2088 8734 -1908
rect 8772 -2076 8778 -1868
rect 8812 -2076 8818 -1868
rect 8868 -1908 8874 -1700
rect 8908 -1908 8914 -1700
rect 8950 -1868 8960 -1688
rect 9012 -1868 9022 -1688
rect 8772 -2088 8818 -2076
rect 8854 -2088 8864 -1908
rect 8916 -2088 8926 -1908
rect 8964 -2076 8970 -1868
rect 9004 -2076 9010 -1868
rect 8964 -2088 9010 -2076
rect 9052 -2120 9132 -1656
rect 4320 -2126 4972 -2120
rect 4320 -2140 4378 -2126
rect 4000 -2160 4378 -2140
rect 4412 -2160 4570 -2126
rect 4604 -2160 4762 -2126
rect 4796 -2140 4972 -2126
rect 5360 -2126 6012 -2120
rect 5360 -2140 5418 -2126
rect 4796 -2160 5418 -2140
rect 5452 -2160 5610 -2126
rect 5644 -2160 5802 -2126
rect 5836 -2140 6012 -2126
rect 6400 -2126 7052 -2120
rect 6400 -2140 6458 -2126
rect 5836 -2160 6458 -2140
rect 6492 -2160 6650 -2126
rect 6684 -2160 6842 -2126
rect 6876 -2140 7052 -2126
rect 7440 -2126 8092 -2120
rect 7440 -2140 7498 -2126
rect 6876 -2160 7498 -2140
rect 7532 -2160 7690 -2126
rect 7724 -2160 7882 -2126
rect 7916 -2140 8092 -2126
rect 8480 -2126 9132 -2120
rect 8480 -2140 8538 -2126
rect 7916 -2160 8538 -2140
rect 8572 -2160 8730 -2126
rect 8764 -2160 8922 -2126
rect 8956 -2160 9132 -2126
rect 4000 -2234 9132 -2160
rect 4000 -2256 4378 -2234
rect 4320 -2268 4378 -2256
rect 4412 -2268 4570 -2234
rect 4604 -2268 4762 -2234
rect 4796 -2256 5418 -2234
rect 4796 -2268 4972 -2256
rect 4320 -2276 4972 -2268
rect 5360 -2268 5418 -2256
rect 5452 -2268 5610 -2234
rect 5644 -2268 5802 -2234
rect 5836 -2256 6458 -2234
rect 5836 -2268 6012 -2256
rect 5360 -2276 6012 -2268
rect 6400 -2268 6458 -2256
rect 6492 -2268 6650 -2234
rect 6684 -2268 6842 -2234
rect 6876 -2256 7498 -2234
rect 6876 -2268 7052 -2256
rect 6400 -2276 7052 -2268
rect 7440 -2268 7498 -2256
rect 7532 -2268 7690 -2234
rect 7724 -2268 7882 -2234
rect 7916 -2256 8538 -2234
rect 7916 -2268 8092 -2256
rect 7440 -2276 8092 -2268
rect 8480 -2268 8538 -2256
rect 8572 -2268 8730 -2234
rect 8764 -2268 8922 -2234
rect 8956 -2268 9132 -2234
rect 11620 -2140 11776 -16
rect 11940 -28 11998 -16
rect 12032 -28 12190 6
rect 12224 -28 12382 6
rect 12416 -16 13038 6
rect 12416 -28 12592 -16
rect 11940 -36 12592 -28
rect 12980 -28 13038 -16
rect 13072 -28 13230 6
rect 13264 -28 13422 6
rect 13456 -16 14078 6
rect 13456 -28 13632 -16
rect 12980 -36 13632 -28
rect 14020 -28 14078 -16
rect 14112 -28 14270 6
rect 14304 -28 14462 6
rect 14496 -16 15118 6
rect 14496 -28 14672 -16
rect 14020 -36 14672 -28
rect 15060 -28 15118 -16
rect 15152 -28 15310 6
rect 15344 -28 15502 6
rect 15536 -16 16158 6
rect 15536 -28 15712 -16
rect 15060 -36 15712 -28
rect 16100 -28 16158 -16
rect 16192 -28 16350 6
rect 16384 -28 16542 6
rect 16576 -16 17198 6
rect 16576 -28 16752 -16
rect 16100 -36 16752 -28
rect 17140 -28 17198 -16
rect 17232 -28 17390 6
rect 17424 -28 17582 6
rect 17616 -16 18238 6
rect 17616 -28 17792 -16
rect 17140 -36 17792 -28
rect 18180 -28 18238 -16
rect 18272 -28 18430 6
rect 18464 -28 18622 6
rect 18656 -28 18832 6
rect 18180 -36 18832 -28
rect 11848 -78 11894 -66
rect 11848 -284 11854 -78
rect 11888 -284 11894 -78
rect 11930 -244 11940 -64
rect 11992 -244 12002 -64
rect 12040 -78 12086 -66
rect 11834 -464 11844 -284
rect 11896 -464 11906 -284
rect 11944 -454 11950 -244
rect 11984 -454 11990 -244
rect 12040 -284 12046 -78
rect 12080 -284 12086 -78
rect 12122 -244 12132 -64
rect 12184 -244 12194 -64
rect 12232 -78 12278 -66
rect 11848 -466 11894 -464
rect 11944 -466 11990 -454
rect 12026 -464 12036 -284
rect 12088 -464 12098 -284
rect 12136 -454 12142 -244
rect 12176 -454 12182 -244
rect 12232 -284 12238 -78
rect 12272 -284 12278 -78
rect 12314 -244 12324 -64
rect 12376 -244 12386 -64
rect 12424 -78 12470 -66
rect 12040 -466 12086 -464
rect 12136 -466 12182 -454
rect 12218 -464 12228 -284
rect 12280 -464 12290 -284
rect 12328 -454 12334 -244
rect 12368 -454 12374 -244
rect 12424 -284 12430 -78
rect 12464 -284 12470 -78
rect 12232 -466 12278 -464
rect 12328 -466 12374 -454
rect 12410 -464 12420 -284
rect 12472 -464 12482 -284
rect 12424 -466 12470 -464
rect 11890 -500 11948 -498
rect 12082 -500 12140 -498
rect 12274 -500 12332 -498
rect 12512 -500 12592 -36
rect 12888 -78 12934 -66
rect 12888 -284 12894 -78
rect 12928 -284 12934 -78
rect 12970 -244 12980 -64
rect 13032 -244 13042 -64
rect 13080 -78 13126 -66
rect 12874 -464 12884 -284
rect 12936 -464 12946 -284
rect 12984 -454 12990 -244
rect 13024 -454 13030 -244
rect 13080 -284 13086 -78
rect 13120 -284 13126 -78
rect 13162 -244 13172 -64
rect 13224 -244 13234 -64
rect 13272 -78 13318 -66
rect 12888 -466 12934 -464
rect 12984 -466 13030 -454
rect 13066 -464 13076 -284
rect 13128 -464 13138 -284
rect 13176 -454 13182 -244
rect 13216 -454 13222 -244
rect 13272 -284 13278 -78
rect 13312 -284 13318 -78
rect 13354 -244 13364 -64
rect 13416 -244 13426 -64
rect 13464 -78 13510 -66
rect 13080 -466 13126 -464
rect 13176 -466 13222 -454
rect 13258 -464 13268 -284
rect 13320 -464 13330 -284
rect 13368 -454 13374 -244
rect 13408 -454 13414 -244
rect 13464 -284 13470 -78
rect 13504 -284 13510 -78
rect 13272 -466 13318 -464
rect 13368 -466 13414 -454
rect 13450 -464 13460 -284
rect 13512 -464 13522 -284
rect 13464 -466 13510 -464
rect 12930 -500 12988 -498
rect 13122 -500 13180 -498
rect 13314 -500 13372 -498
rect 13552 -500 13632 -36
rect 13928 -78 13974 -66
rect 13928 -284 13934 -78
rect 13968 -284 13974 -78
rect 14010 -244 14020 -64
rect 14072 -244 14082 -64
rect 14120 -78 14166 -66
rect 13914 -464 13924 -284
rect 13976 -464 13986 -284
rect 14024 -454 14030 -244
rect 14064 -454 14070 -244
rect 14120 -284 14126 -78
rect 14160 -284 14166 -78
rect 14202 -244 14212 -64
rect 14264 -244 14274 -64
rect 14312 -78 14358 -66
rect 13928 -466 13974 -464
rect 14024 -466 14070 -454
rect 14106 -464 14116 -284
rect 14168 -464 14178 -284
rect 14216 -454 14222 -244
rect 14256 -454 14262 -244
rect 14312 -284 14318 -78
rect 14352 -284 14358 -78
rect 14394 -244 14404 -64
rect 14456 -244 14466 -64
rect 14504 -78 14550 -66
rect 14120 -466 14166 -464
rect 14216 -466 14262 -454
rect 14298 -464 14308 -284
rect 14360 -464 14370 -284
rect 14408 -454 14414 -244
rect 14448 -454 14454 -244
rect 14504 -284 14510 -78
rect 14544 -284 14550 -78
rect 14312 -466 14358 -464
rect 14408 -466 14454 -454
rect 14490 -464 14500 -284
rect 14552 -464 14562 -284
rect 14504 -466 14550 -464
rect 13970 -500 14028 -498
rect 14162 -500 14220 -498
rect 14354 -500 14412 -498
rect 14592 -500 14672 -36
rect 14968 -78 15014 -66
rect 14968 -284 14974 -78
rect 15008 -284 15014 -78
rect 15050 -244 15060 -64
rect 15112 -244 15122 -64
rect 15160 -78 15206 -66
rect 14954 -464 14964 -284
rect 15016 -464 15026 -284
rect 15064 -454 15070 -244
rect 15104 -454 15110 -244
rect 15160 -284 15166 -78
rect 15200 -284 15206 -78
rect 15242 -244 15252 -64
rect 15304 -244 15314 -64
rect 15352 -78 15398 -66
rect 14968 -466 15014 -464
rect 15064 -466 15110 -454
rect 15146 -464 15156 -284
rect 15208 -464 15218 -284
rect 15256 -454 15262 -244
rect 15296 -454 15302 -244
rect 15352 -284 15358 -78
rect 15392 -284 15398 -78
rect 15434 -244 15444 -64
rect 15496 -244 15506 -64
rect 15544 -78 15590 -66
rect 15160 -466 15206 -464
rect 15256 -466 15302 -454
rect 15338 -464 15348 -284
rect 15400 -464 15410 -284
rect 15448 -454 15454 -244
rect 15488 -454 15494 -244
rect 15544 -284 15550 -78
rect 15584 -284 15590 -78
rect 15352 -466 15398 -464
rect 15448 -466 15494 -454
rect 15530 -464 15540 -284
rect 15592 -464 15602 -284
rect 15544 -466 15590 -464
rect 15010 -500 15068 -498
rect 15202 -500 15260 -498
rect 15394 -500 15452 -498
rect 15632 -500 15712 -36
rect 16008 -78 16054 -66
rect 16008 -284 16014 -78
rect 16048 -284 16054 -78
rect 16090 -244 16100 -64
rect 16152 -244 16162 -64
rect 16200 -78 16246 -66
rect 15994 -464 16004 -284
rect 16056 -464 16066 -284
rect 16104 -454 16110 -244
rect 16144 -454 16150 -244
rect 16200 -284 16206 -78
rect 16240 -284 16246 -78
rect 16282 -244 16292 -64
rect 16344 -244 16354 -64
rect 16392 -78 16438 -66
rect 16008 -466 16054 -464
rect 16104 -466 16150 -454
rect 16186 -464 16196 -284
rect 16248 -464 16258 -284
rect 16296 -454 16302 -244
rect 16336 -454 16342 -244
rect 16392 -284 16398 -78
rect 16432 -284 16438 -78
rect 16474 -244 16484 -64
rect 16536 -244 16546 -64
rect 16584 -78 16630 -66
rect 16200 -466 16246 -464
rect 16296 -466 16342 -454
rect 16378 -464 16388 -284
rect 16440 -464 16450 -284
rect 16488 -454 16494 -244
rect 16528 -454 16534 -244
rect 16584 -284 16590 -78
rect 16624 -284 16630 -78
rect 16392 -466 16438 -464
rect 16488 -466 16534 -454
rect 16570 -464 16580 -284
rect 16632 -464 16642 -284
rect 16584 -466 16630 -464
rect 16050 -500 16108 -498
rect 16242 -500 16300 -498
rect 16434 -500 16492 -498
rect 16672 -500 16752 -36
rect 17048 -78 17094 -66
rect 17048 -284 17054 -78
rect 17088 -284 17094 -78
rect 17130 -244 17140 -64
rect 17192 -244 17202 -64
rect 17240 -78 17286 -66
rect 17034 -464 17044 -284
rect 17096 -464 17106 -284
rect 17144 -454 17150 -244
rect 17184 -454 17190 -244
rect 17240 -284 17246 -78
rect 17280 -284 17286 -78
rect 17322 -244 17332 -64
rect 17384 -244 17394 -64
rect 17432 -78 17478 -66
rect 17048 -466 17094 -464
rect 17144 -466 17190 -454
rect 17226 -464 17236 -284
rect 17288 -464 17298 -284
rect 17336 -454 17342 -244
rect 17376 -454 17382 -244
rect 17432 -284 17438 -78
rect 17472 -284 17478 -78
rect 17514 -244 17524 -64
rect 17576 -244 17586 -64
rect 17624 -78 17670 -66
rect 17240 -466 17286 -464
rect 17336 -466 17382 -454
rect 17418 -464 17428 -284
rect 17480 -464 17490 -284
rect 17528 -454 17534 -244
rect 17568 -454 17574 -244
rect 17624 -284 17630 -78
rect 17664 -284 17670 -78
rect 17432 -466 17478 -464
rect 17528 -466 17574 -454
rect 17610 -464 17620 -284
rect 17672 -464 17682 -284
rect 17624 -466 17670 -464
rect 17090 -500 17148 -498
rect 17282 -500 17340 -498
rect 17474 -500 17532 -498
rect 17712 -500 17792 -36
rect 18088 -78 18134 -66
rect 18088 -284 18094 -78
rect 18128 -284 18134 -78
rect 18170 -244 18180 -64
rect 18232 -244 18242 -64
rect 18280 -78 18326 -66
rect 18074 -464 18084 -284
rect 18136 -464 18146 -284
rect 18184 -454 18190 -244
rect 18224 -454 18230 -244
rect 18280 -284 18286 -78
rect 18320 -284 18326 -78
rect 18362 -244 18372 -64
rect 18424 -244 18434 -64
rect 18472 -78 18518 -66
rect 18088 -466 18134 -464
rect 18184 -466 18230 -454
rect 18266 -464 18276 -284
rect 18328 -464 18338 -284
rect 18376 -454 18382 -244
rect 18416 -454 18422 -244
rect 18472 -284 18478 -78
rect 18512 -284 18518 -78
rect 18554 -244 18564 -64
rect 18616 -244 18626 -64
rect 18664 -78 18710 -66
rect 18280 -466 18326 -464
rect 18376 -466 18422 -454
rect 18458 -464 18468 -284
rect 18520 -464 18530 -284
rect 18568 -454 18574 -244
rect 18608 -454 18614 -244
rect 18664 -284 18670 -78
rect 18704 -284 18710 -78
rect 18472 -466 18518 -464
rect 18568 -466 18614 -454
rect 18650 -464 18660 -284
rect 18712 -464 18722 -284
rect 18664 -466 18710 -464
rect 18130 -500 18188 -498
rect 18322 -500 18380 -498
rect 18514 -500 18572 -498
rect 18752 -500 18832 -36
rect 11884 -504 12592 -500
rect 11884 -538 11902 -504
rect 11936 -538 12094 -504
rect 12128 -538 12286 -504
rect 12320 -538 12592 -504
rect 11884 -596 12592 -538
rect 12924 -504 13632 -500
rect 12924 -538 12942 -504
rect 12976 -538 13134 -504
rect 13168 -538 13326 -504
rect 13360 -538 13632 -504
rect 12924 -596 13632 -538
rect 13964 -504 14672 -500
rect 13964 -538 13982 -504
rect 14016 -538 14174 -504
rect 14208 -538 14366 -504
rect 14400 -538 14672 -504
rect 13964 -596 14672 -538
rect 15004 -504 15712 -500
rect 15004 -538 15022 -504
rect 15056 -538 15214 -504
rect 15248 -538 15406 -504
rect 15440 -538 15712 -504
rect 15004 -596 15712 -538
rect 16044 -504 16752 -500
rect 16044 -538 16062 -504
rect 16096 -538 16254 -504
rect 16288 -538 16446 -504
rect 16480 -538 16752 -504
rect 16044 -596 16752 -538
rect 17084 -504 17792 -500
rect 17084 -538 17102 -504
rect 17136 -538 17294 -504
rect 17328 -538 17486 -504
rect 17520 -538 17792 -504
rect 17084 -596 17792 -538
rect 18124 -504 18832 -500
rect 18124 -538 18142 -504
rect 18176 -538 18334 -504
rect 18368 -538 18526 -504
rect 18560 -538 18832 -504
rect 18124 -596 18832 -538
rect 12456 -772 12540 -596
rect 13496 -772 13580 -596
rect 14536 -772 14620 -596
rect 15576 -772 15660 -596
rect 16616 -772 16700 -596
rect 17656 -772 17740 -596
rect 18696 -772 18780 -596
rect 11892 -798 12708 -772
rect 11892 -832 11913 -798
rect 11947 -832 12031 -798
rect 12065 -832 12149 -798
rect 12183 -832 12267 -798
rect 12301 -832 12385 -798
rect 12419 -832 12503 -798
rect 12537 -832 12708 -798
rect 11892 -840 12708 -832
rect 12932 -798 13748 -772
rect 12932 -832 12953 -798
rect 12987 -832 13071 -798
rect 13105 -832 13189 -798
rect 13223 -832 13307 -798
rect 13341 -832 13425 -798
rect 13459 -832 13543 -798
rect 13577 -832 13748 -798
rect 12932 -840 13748 -832
rect 13972 -798 14788 -772
rect 13972 -832 13993 -798
rect 14027 -832 14111 -798
rect 14145 -832 14229 -798
rect 14263 -832 14347 -798
rect 14381 -832 14465 -798
rect 14499 -832 14583 -798
rect 14617 -832 14788 -798
rect 13972 -840 14788 -832
rect 15012 -798 15828 -772
rect 15012 -832 15033 -798
rect 15067 -832 15151 -798
rect 15185 -832 15269 -798
rect 15303 -832 15387 -798
rect 15421 -832 15505 -798
rect 15539 -832 15623 -798
rect 15657 -832 15828 -798
rect 15012 -840 15828 -832
rect 16052 -798 16868 -772
rect 16052 -832 16073 -798
rect 16107 -832 16191 -798
rect 16225 -832 16309 -798
rect 16343 -832 16427 -798
rect 16461 -832 16545 -798
rect 16579 -832 16663 -798
rect 16697 -832 16868 -798
rect 16052 -840 16868 -832
rect 17092 -798 17908 -772
rect 17092 -832 17113 -798
rect 17147 -832 17231 -798
rect 17265 -832 17349 -798
rect 17383 -832 17467 -798
rect 17501 -832 17585 -798
rect 17619 -832 17703 -798
rect 17737 -832 17908 -798
rect 17092 -840 17908 -832
rect 18132 -798 18948 -772
rect 18132 -832 18153 -798
rect 18187 -832 18271 -798
rect 18305 -832 18389 -798
rect 18423 -832 18507 -798
rect 18541 -832 18625 -798
rect 18659 -832 18743 -798
rect 18777 -832 18948 -798
rect 18132 -840 18948 -832
rect 11848 -882 11894 -870
rect 11848 -1092 11854 -882
rect 11888 -1092 11894 -882
rect 11954 -1048 11964 -868
rect 12016 -1048 12026 -868
rect 12084 -882 12130 -870
rect 11834 -1272 11844 -1092
rect 11896 -1272 11906 -1092
rect 11966 -1258 11972 -1048
rect 12006 -1258 12012 -1048
rect 12084 -1092 12090 -882
rect 12124 -1092 12130 -882
rect 12190 -1048 12200 -868
rect 12252 -1048 12262 -868
rect 12320 -882 12366 -870
rect 11966 -1270 12012 -1258
rect 12070 -1272 12080 -1092
rect 12132 -1272 12142 -1092
rect 12202 -1258 12208 -1048
rect 12242 -1258 12248 -1048
rect 12320 -1092 12326 -882
rect 12360 -1092 12366 -882
rect 12426 -1048 12436 -868
rect 12488 -1048 12498 -868
rect 12556 -882 12602 -870
rect 12202 -1270 12248 -1258
rect 12306 -1272 12316 -1092
rect 12368 -1272 12378 -1092
rect 12438 -1258 12444 -1048
rect 12478 -1258 12484 -1048
rect 12556 -1092 12562 -882
rect 12596 -1092 12602 -882
rect 12438 -1270 12484 -1258
rect 12542 -1272 12552 -1092
rect 12604 -1272 12614 -1092
rect 12644 -1300 12708 -840
rect 12888 -882 12934 -870
rect 12888 -1092 12894 -882
rect 12928 -1092 12934 -882
rect 12994 -1048 13004 -868
rect 13056 -1048 13066 -868
rect 13124 -882 13170 -870
rect 12874 -1272 12884 -1092
rect 12936 -1272 12946 -1092
rect 13006 -1258 13012 -1048
rect 13046 -1258 13052 -1048
rect 13124 -1092 13130 -882
rect 13164 -1092 13170 -882
rect 13230 -1048 13240 -868
rect 13292 -1048 13302 -868
rect 13360 -882 13406 -870
rect 13006 -1270 13052 -1258
rect 13110 -1272 13120 -1092
rect 13172 -1272 13182 -1092
rect 13242 -1258 13248 -1048
rect 13282 -1258 13288 -1048
rect 13360 -1092 13366 -882
rect 13400 -1092 13406 -882
rect 13466 -1048 13476 -868
rect 13528 -1048 13538 -868
rect 13596 -882 13642 -870
rect 13242 -1270 13288 -1258
rect 13346 -1272 13356 -1092
rect 13408 -1272 13418 -1092
rect 13478 -1258 13484 -1048
rect 13518 -1258 13524 -1048
rect 13596 -1092 13602 -882
rect 13636 -1092 13642 -882
rect 13478 -1270 13524 -1258
rect 13582 -1272 13592 -1092
rect 13644 -1272 13654 -1092
rect 13684 -1300 13748 -840
rect 13928 -882 13974 -870
rect 13928 -1092 13934 -882
rect 13968 -1092 13974 -882
rect 14034 -1048 14044 -868
rect 14096 -1048 14106 -868
rect 14164 -882 14210 -870
rect 13914 -1272 13924 -1092
rect 13976 -1272 13986 -1092
rect 14046 -1258 14052 -1048
rect 14086 -1258 14092 -1048
rect 14164 -1092 14170 -882
rect 14204 -1092 14210 -882
rect 14270 -1048 14280 -868
rect 14332 -1048 14342 -868
rect 14400 -882 14446 -870
rect 14046 -1270 14092 -1258
rect 14150 -1272 14160 -1092
rect 14212 -1272 14222 -1092
rect 14282 -1258 14288 -1048
rect 14322 -1258 14328 -1048
rect 14400 -1092 14406 -882
rect 14440 -1092 14446 -882
rect 14506 -1048 14516 -868
rect 14568 -1048 14578 -868
rect 14636 -882 14682 -870
rect 14282 -1270 14328 -1258
rect 14386 -1272 14396 -1092
rect 14448 -1272 14458 -1092
rect 14518 -1258 14524 -1048
rect 14558 -1258 14564 -1048
rect 14636 -1092 14642 -882
rect 14676 -1092 14682 -882
rect 14518 -1270 14564 -1258
rect 14622 -1272 14632 -1092
rect 14684 -1272 14694 -1092
rect 14724 -1300 14788 -840
rect 14968 -882 15014 -870
rect 14968 -1092 14974 -882
rect 15008 -1092 15014 -882
rect 15074 -1048 15084 -868
rect 15136 -1048 15146 -868
rect 15204 -882 15250 -870
rect 14954 -1272 14964 -1092
rect 15016 -1272 15026 -1092
rect 15086 -1258 15092 -1048
rect 15126 -1258 15132 -1048
rect 15204 -1092 15210 -882
rect 15244 -1092 15250 -882
rect 15310 -1048 15320 -868
rect 15372 -1048 15382 -868
rect 15440 -882 15486 -870
rect 15086 -1270 15132 -1258
rect 15190 -1272 15200 -1092
rect 15252 -1272 15262 -1092
rect 15322 -1258 15328 -1048
rect 15362 -1258 15368 -1048
rect 15440 -1092 15446 -882
rect 15480 -1092 15486 -882
rect 15546 -1048 15556 -868
rect 15608 -1048 15618 -868
rect 15676 -882 15722 -870
rect 15322 -1270 15368 -1258
rect 15426 -1272 15436 -1092
rect 15488 -1272 15498 -1092
rect 15558 -1258 15564 -1048
rect 15598 -1258 15604 -1048
rect 15676 -1092 15682 -882
rect 15716 -1092 15722 -882
rect 15558 -1270 15604 -1258
rect 15662 -1272 15672 -1092
rect 15724 -1272 15734 -1092
rect 15764 -1300 15828 -840
rect 16008 -882 16054 -870
rect 16008 -1092 16014 -882
rect 16048 -1092 16054 -882
rect 16114 -1048 16124 -868
rect 16176 -1048 16186 -868
rect 16244 -882 16290 -870
rect 15994 -1272 16004 -1092
rect 16056 -1272 16066 -1092
rect 16126 -1258 16132 -1048
rect 16166 -1258 16172 -1048
rect 16244 -1092 16250 -882
rect 16284 -1092 16290 -882
rect 16350 -1048 16360 -868
rect 16412 -1048 16422 -868
rect 16480 -882 16526 -870
rect 16126 -1270 16172 -1258
rect 16230 -1272 16240 -1092
rect 16292 -1272 16302 -1092
rect 16362 -1258 16368 -1048
rect 16402 -1258 16408 -1048
rect 16480 -1092 16486 -882
rect 16520 -1092 16526 -882
rect 16586 -1048 16596 -868
rect 16648 -1048 16658 -868
rect 16716 -882 16762 -870
rect 16362 -1270 16408 -1258
rect 16466 -1272 16476 -1092
rect 16528 -1272 16538 -1092
rect 16598 -1258 16604 -1048
rect 16638 -1258 16644 -1048
rect 16716 -1092 16722 -882
rect 16756 -1092 16762 -882
rect 16598 -1270 16644 -1258
rect 16702 -1272 16712 -1092
rect 16764 -1272 16774 -1092
rect 16804 -1300 16868 -840
rect 17048 -882 17094 -870
rect 17048 -1092 17054 -882
rect 17088 -1092 17094 -882
rect 17154 -1048 17164 -868
rect 17216 -1048 17226 -868
rect 17284 -882 17330 -870
rect 17034 -1272 17044 -1092
rect 17096 -1272 17106 -1092
rect 17166 -1258 17172 -1048
rect 17206 -1258 17212 -1048
rect 17284 -1092 17290 -882
rect 17324 -1092 17330 -882
rect 17390 -1048 17400 -868
rect 17452 -1048 17462 -868
rect 17520 -882 17566 -870
rect 17166 -1270 17212 -1258
rect 17270 -1272 17280 -1092
rect 17332 -1272 17342 -1092
rect 17402 -1258 17408 -1048
rect 17442 -1258 17448 -1048
rect 17520 -1092 17526 -882
rect 17560 -1092 17566 -882
rect 17626 -1048 17636 -868
rect 17688 -1048 17698 -868
rect 17756 -882 17802 -870
rect 17402 -1270 17448 -1258
rect 17506 -1272 17516 -1092
rect 17568 -1272 17578 -1092
rect 17638 -1258 17644 -1048
rect 17678 -1258 17684 -1048
rect 17756 -1092 17762 -882
rect 17796 -1092 17802 -882
rect 17638 -1270 17684 -1258
rect 17742 -1272 17752 -1092
rect 17804 -1272 17814 -1092
rect 17844 -1300 17908 -840
rect 18088 -882 18134 -870
rect 18088 -1092 18094 -882
rect 18128 -1092 18134 -882
rect 18194 -1048 18204 -868
rect 18256 -1048 18266 -868
rect 18324 -882 18370 -870
rect 18074 -1272 18084 -1092
rect 18136 -1272 18146 -1092
rect 18206 -1258 18212 -1048
rect 18246 -1258 18252 -1048
rect 18324 -1092 18330 -882
rect 18364 -1092 18370 -882
rect 18430 -1048 18440 -868
rect 18492 -1048 18502 -868
rect 18560 -882 18606 -870
rect 18206 -1270 18252 -1258
rect 18310 -1272 18320 -1092
rect 18372 -1272 18382 -1092
rect 18442 -1258 18448 -1048
rect 18482 -1258 18488 -1048
rect 18560 -1092 18566 -882
rect 18600 -1092 18606 -882
rect 18666 -1048 18676 -868
rect 18728 -1048 18738 -868
rect 18796 -882 18842 -870
rect 18442 -1270 18488 -1258
rect 18546 -1272 18556 -1092
rect 18608 -1272 18618 -1092
rect 18678 -1258 18684 -1048
rect 18718 -1258 18724 -1048
rect 18796 -1092 18802 -882
rect 18836 -1092 18842 -882
rect 18678 -1270 18724 -1258
rect 18782 -1272 18792 -1092
rect 18844 -1272 18854 -1092
rect 18884 -1300 18948 -840
rect 11896 -1308 12708 -1300
rect 11896 -1342 11913 -1308
rect 11947 -1342 12031 -1308
rect 12065 -1342 12149 -1308
rect 12183 -1342 12267 -1308
rect 12301 -1342 12385 -1308
rect 12419 -1342 12503 -1308
rect 12537 -1342 12708 -1308
rect 11896 -1368 12708 -1342
rect 12936 -1308 13748 -1300
rect 12936 -1342 12953 -1308
rect 12987 -1342 13071 -1308
rect 13105 -1342 13189 -1308
rect 13223 -1342 13307 -1308
rect 13341 -1342 13425 -1308
rect 13459 -1342 13543 -1308
rect 13577 -1342 13748 -1308
rect 12936 -1368 13748 -1342
rect 13976 -1308 14788 -1300
rect 13976 -1342 13993 -1308
rect 14027 -1342 14111 -1308
rect 14145 -1342 14229 -1308
rect 14263 -1342 14347 -1308
rect 14381 -1342 14465 -1308
rect 14499 -1342 14583 -1308
rect 14617 -1342 14788 -1308
rect 13976 -1368 14788 -1342
rect 15016 -1308 15828 -1300
rect 15016 -1342 15033 -1308
rect 15067 -1342 15151 -1308
rect 15185 -1342 15269 -1308
rect 15303 -1342 15387 -1308
rect 15421 -1342 15505 -1308
rect 15539 -1342 15623 -1308
rect 15657 -1342 15828 -1308
rect 15016 -1368 15828 -1342
rect 16056 -1308 16868 -1300
rect 16056 -1342 16073 -1308
rect 16107 -1342 16191 -1308
rect 16225 -1342 16309 -1308
rect 16343 -1342 16427 -1308
rect 16461 -1342 16545 -1308
rect 16579 -1342 16663 -1308
rect 16697 -1342 16868 -1308
rect 16056 -1368 16868 -1342
rect 17096 -1308 17908 -1300
rect 17096 -1342 17113 -1308
rect 17147 -1342 17231 -1308
rect 17265 -1342 17349 -1308
rect 17383 -1342 17467 -1308
rect 17501 -1342 17585 -1308
rect 17619 -1342 17703 -1308
rect 17737 -1342 17908 -1308
rect 17096 -1368 17908 -1342
rect 18136 -1308 18948 -1300
rect 18136 -1342 18153 -1308
rect 18187 -1342 18271 -1308
rect 18305 -1342 18389 -1308
rect 18423 -1342 18507 -1308
rect 18541 -1342 18625 -1308
rect 18659 -1342 18743 -1308
rect 18777 -1342 18948 -1308
rect 18136 -1368 18948 -1342
rect 11880 -1616 12592 -1572
rect 11880 -1650 11902 -1616
rect 11936 -1650 12094 -1616
rect 12128 -1650 12286 -1616
rect 12320 -1650 12592 -1616
rect 11880 -1656 12592 -1650
rect 12920 -1616 13632 -1572
rect 12920 -1650 12942 -1616
rect 12976 -1650 13134 -1616
rect 13168 -1650 13326 -1616
rect 13360 -1650 13632 -1616
rect 12920 -1656 13632 -1650
rect 13960 -1616 14672 -1572
rect 13960 -1650 13982 -1616
rect 14016 -1650 14174 -1616
rect 14208 -1650 14366 -1616
rect 14400 -1650 14672 -1616
rect 13960 -1656 14672 -1650
rect 15000 -1616 15712 -1572
rect 15000 -1650 15022 -1616
rect 15056 -1650 15214 -1616
rect 15248 -1650 15406 -1616
rect 15440 -1650 15712 -1616
rect 15000 -1656 15712 -1650
rect 16040 -1616 16752 -1572
rect 16040 -1650 16062 -1616
rect 16096 -1650 16254 -1616
rect 16288 -1650 16446 -1616
rect 16480 -1650 16752 -1616
rect 16040 -1656 16752 -1650
rect 11834 -1868 11844 -1688
rect 11896 -1868 11906 -1688
rect 11944 -1700 11990 -1688
rect 11848 -2076 11854 -1868
rect 11888 -2076 11894 -1868
rect 11944 -1908 11950 -1700
rect 11984 -1908 11990 -1700
rect 12026 -1868 12036 -1688
rect 12088 -1868 12098 -1688
rect 12136 -1700 12182 -1688
rect 11848 -2088 11894 -2076
rect 11930 -2088 11940 -1908
rect 11992 -2088 12002 -1908
rect 12040 -2076 12046 -1868
rect 12080 -2076 12086 -1868
rect 12136 -1908 12142 -1700
rect 12176 -1908 12182 -1700
rect 12218 -1868 12228 -1688
rect 12280 -1868 12290 -1688
rect 12328 -1700 12374 -1688
rect 12040 -2088 12086 -2076
rect 12122 -2088 12132 -1908
rect 12184 -2088 12194 -1908
rect 12232 -2076 12238 -1868
rect 12272 -2076 12278 -1868
rect 12328 -1908 12334 -1700
rect 12368 -1908 12374 -1700
rect 12410 -1868 12420 -1688
rect 12472 -1868 12482 -1688
rect 12232 -2088 12278 -2076
rect 12314 -2088 12324 -1908
rect 12376 -2088 12386 -1908
rect 12424 -2076 12430 -1868
rect 12464 -2076 12470 -1868
rect 12424 -2088 12470 -2076
rect 12512 -2120 12592 -1656
rect 12874 -1868 12884 -1688
rect 12936 -1868 12946 -1688
rect 12984 -1700 13030 -1688
rect 12888 -2076 12894 -1868
rect 12928 -2076 12934 -1868
rect 12984 -1908 12990 -1700
rect 13024 -1908 13030 -1700
rect 13066 -1868 13076 -1688
rect 13128 -1868 13138 -1688
rect 13176 -1700 13222 -1688
rect 12888 -2088 12934 -2076
rect 12970 -2088 12980 -1908
rect 13032 -2088 13042 -1908
rect 13080 -2076 13086 -1868
rect 13120 -2076 13126 -1868
rect 13176 -1908 13182 -1700
rect 13216 -1908 13222 -1700
rect 13258 -1868 13268 -1688
rect 13320 -1868 13330 -1688
rect 13368 -1700 13414 -1688
rect 13080 -2088 13126 -2076
rect 13162 -2088 13172 -1908
rect 13224 -2088 13234 -1908
rect 13272 -2076 13278 -1868
rect 13312 -2076 13318 -1868
rect 13368 -1908 13374 -1700
rect 13408 -1908 13414 -1700
rect 13450 -1868 13460 -1688
rect 13512 -1868 13522 -1688
rect 13272 -2088 13318 -2076
rect 13354 -2088 13364 -1908
rect 13416 -2088 13426 -1908
rect 13464 -2076 13470 -1868
rect 13504 -2076 13510 -1868
rect 13464 -2088 13510 -2076
rect 13552 -2120 13632 -1656
rect 13914 -1868 13924 -1688
rect 13976 -1868 13986 -1688
rect 14024 -1700 14070 -1688
rect 13928 -2076 13934 -1868
rect 13968 -2076 13974 -1868
rect 14024 -1908 14030 -1700
rect 14064 -1908 14070 -1700
rect 14106 -1868 14116 -1688
rect 14168 -1868 14178 -1688
rect 14216 -1700 14262 -1688
rect 13928 -2088 13974 -2076
rect 14010 -2088 14020 -1908
rect 14072 -2088 14082 -1908
rect 14120 -2076 14126 -1868
rect 14160 -2076 14166 -1868
rect 14216 -1908 14222 -1700
rect 14256 -1908 14262 -1700
rect 14298 -1868 14308 -1688
rect 14360 -1868 14370 -1688
rect 14408 -1700 14454 -1688
rect 14120 -2088 14166 -2076
rect 14202 -2088 14212 -1908
rect 14264 -2088 14274 -1908
rect 14312 -2076 14318 -1868
rect 14352 -2076 14358 -1868
rect 14408 -1908 14414 -1700
rect 14448 -1908 14454 -1700
rect 14490 -1868 14500 -1688
rect 14552 -1868 14562 -1688
rect 14312 -2088 14358 -2076
rect 14394 -2088 14404 -1908
rect 14456 -2088 14466 -1908
rect 14504 -2076 14510 -1868
rect 14544 -2076 14550 -1868
rect 14504 -2088 14550 -2076
rect 14592 -2120 14672 -1656
rect 14954 -1868 14964 -1688
rect 15016 -1868 15026 -1688
rect 15064 -1700 15110 -1688
rect 14968 -2076 14974 -1868
rect 15008 -2076 15014 -1868
rect 15064 -1908 15070 -1700
rect 15104 -1908 15110 -1700
rect 15146 -1868 15156 -1688
rect 15208 -1868 15218 -1688
rect 15256 -1700 15302 -1688
rect 14968 -2088 15014 -2076
rect 15050 -2088 15060 -1908
rect 15112 -2088 15122 -1908
rect 15160 -2076 15166 -1868
rect 15200 -2076 15206 -1868
rect 15256 -1908 15262 -1700
rect 15296 -1908 15302 -1700
rect 15338 -1868 15348 -1688
rect 15400 -1868 15410 -1688
rect 15448 -1700 15494 -1688
rect 15160 -2088 15206 -2076
rect 15242 -2088 15252 -1908
rect 15304 -2088 15314 -1908
rect 15352 -2076 15358 -1868
rect 15392 -2076 15398 -1868
rect 15448 -1908 15454 -1700
rect 15488 -1908 15494 -1700
rect 15530 -1868 15540 -1688
rect 15592 -1868 15602 -1688
rect 15352 -2088 15398 -2076
rect 15434 -2088 15444 -1908
rect 15496 -2088 15506 -1908
rect 15544 -2076 15550 -1868
rect 15584 -2076 15590 -1868
rect 15544 -2088 15590 -2076
rect 15632 -2120 15712 -1656
rect 15994 -1868 16004 -1688
rect 16056 -1868 16066 -1688
rect 16104 -1700 16150 -1688
rect 16008 -2076 16014 -1868
rect 16048 -2076 16054 -1868
rect 16104 -1908 16110 -1700
rect 16144 -1908 16150 -1700
rect 16186 -1868 16196 -1688
rect 16248 -1868 16258 -1688
rect 16296 -1700 16342 -1688
rect 16008 -2088 16054 -2076
rect 16090 -2088 16100 -1908
rect 16152 -2088 16162 -1908
rect 16200 -2076 16206 -1868
rect 16240 -2076 16246 -1868
rect 16296 -1908 16302 -1700
rect 16336 -1908 16342 -1700
rect 16378 -1868 16388 -1688
rect 16440 -1868 16450 -1688
rect 16488 -1700 16534 -1688
rect 16200 -2088 16246 -2076
rect 16282 -2088 16292 -1908
rect 16344 -2088 16354 -1908
rect 16392 -2076 16398 -1868
rect 16432 -2076 16438 -1868
rect 16488 -1908 16494 -1700
rect 16528 -1908 16534 -1700
rect 16570 -1868 16580 -1688
rect 16632 -1868 16642 -1688
rect 16392 -2088 16438 -2076
rect 16474 -2088 16484 -1908
rect 16536 -2088 16546 -1908
rect 16584 -2076 16590 -1868
rect 16624 -2076 16630 -1868
rect 16584 -2088 16630 -2076
rect 16672 -2120 16752 -1656
rect 11940 -2126 12592 -2120
rect 11940 -2140 11998 -2126
rect 11620 -2160 11998 -2140
rect 12032 -2160 12190 -2126
rect 12224 -2160 12382 -2126
rect 12416 -2140 12592 -2126
rect 12980 -2126 13632 -2120
rect 12980 -2140 13038 -2126
rect 12416 -2160 13038 -2140
rect 13072 -2160 13230 -2126
rect 13264 -2160 13422 -2126
rect 13456 -2140 13632 -2126
rect 14020 -2126 14672 -2120
rect 14020 -2140 14078 -2126
rect 13456 -2160 14078 -2140
rect 14112 -2160 14270 -2126
rect 14304 -2160 14462 -2126
rect 14496 -2140 14672 -2126
rect 15060 -2126 15712 -2120
rect 15060 -2140 15118 -2126
rect 14496 -2160 15118 -2140
rect 15152 -2160 15310 -2126
rect 15344 -2160 15502 -2126
rect 15536 -2140 15712 -2126
rect 16100 -2126 16752 -2120
rect 16100 -2140 16158 -2126
rect 15536 -2160 16158 -2140
rect 16192 -2160 16350 -2126
rect 16384 -2160 16542 -2126
rect 16576 -2160 16752 -2126
rect 11620 -2234 16752 -2160
rect 11620 -2256 11998 -2234
rect 8480 -2276 9132 -2268
rect 11940 -2268 11998 -2256
rect 12032 -2268 12190 -2234
rect 12224 -2268 12382 -2234
rect 12416 -2256 13038 -2234
rect 12416 -2268 12592 -2256
rect 11940 -2276 12592 -2268
rect 12980 -2268 13038 -2256
rect 13072 -2268 13230 -2234
rect 13264 -2268 13422 -2234
rect 13456 -2256 14078 -2234
rect 13456 -2268 13632 -2256
rect 12980 -2276 13632 -2268
rect 14020 -2268 14078 -2256
rect 14112 -2268 14270 -2234
rect 14304 -2268 14462 -2234
rect 14496 -2256 15118 -2234
rect 14496 -2268 14672 -2256
rect 14020 -2276 14672 -2268
rect 15060 -2268 15118 -2256
rect 15152 -2268 15310 -2234
rect 15344 -2268 15502 -2234
rect 15536 -2256 16158 -2234
rect 15536 -2268 15712 -2256
rect 15060 -2276 15712 -2268
rect 16100 -2268 16158 -2256
rect 16192 -2268 16350 -2234
rect 16384 -2268 16542 -2234
rect 16576 -2268 16752 -2234
rect 16100 -2276 16752 -2268
rect -7314 -2328 -6662 -2322
rect -7314 -2362 -7256 -2328
rect -7222 -2362 -7064 -2328
rect -7030 -2362 -6872 -2328
rect -6838 -2362 -6662 -2328
rect -7314 -2436 -6662 -2362
rect -7314 -2470 -7256 -2436
rect -7222 -2470 -7064 -2436
rect -7030 -2470 -6872 -2436
rect -6838 -2470 -6662 -2436
rect -7314 -2478 -6662 -2470
rect -7406 -2520 -7360 -2508
rect -7406 -2726 -7400 -2520
rect -7366 -2726 -7360 -2520
rect -7324 -2686 -7314 -2506
rect -7262 -2686 -7252 -2506
rect -7214 -2520 -7168 -2508
rect -7420 -2906 -7410 -2726
rect -7358 -2906 -7348 -2726
rect -7310 -2896 -7304 -2686
rect -7270 -2896 -7264 -2686
rect -7214 -2726 -7208 -2520
rect -7174 -2726 -7168 -2520
rect -7132 -2686 -7122 -2506
rect -7070 -2686 -7060 -2506
rect -7022 -2520 -6976 -2508
rect -7406 -2908 -7360 -2906
rect -7310 -2908 -7264 -2896
rect -7228 -2906 -7218 -2726
rect -7166 -2906 -7156 -2726
rect -7118 -2896 -7112 -2686
rect -7078 -2896 -7072 -2686
rect -7022 -2726 -7016 -2520
rect -6982 -2726 -6976 -2520
rect -6940 -2686 -6930 -2506
rect -6878 -2686 -6868 -2506
rect -6830 -2520 -6784 -2508
rect -7214 -2908 -7168 -2906
rect -7118 -2908 -7072 -2896
rect -7036 -2906 -7026 -2726
rect -6974 -2906 -6964 -2726
rect -6926 -2896 -6920 -2686
rect -6886 -2896 -6880 -2686
rect -6830 -2726 -6824 -2520
rect -6790 -2726 -6784 -2520
rect -7022 -2908 -6976 -2906
rect -6926 -2908 -6880 -2896
rect -6844 -2906 -6834 -2726
rect -6782 -2906 -6772 -2726
rect -6830 -2908 -6784 -2906
rect -7364 -2942 -7306 -2940
rect -7172 -2942 -7114 -2940
rect -6980 -2942 -6922 -2940
rect -6742 -2942 -6662 -2478
rect 4228 -2318 4274 -2306
rect 4228 -2524 4234 -2318
rect 4268 -2524 4274 -2318
rect 4310 -2484 4320 -2304
rect 4372 -2484 4382 -2304
rect 4420 -2318 4466 -2306
rect 4214 -2704 4224 -2524
rect 4276 -2704 4286 -2524
rect 4324 -2694 4330 -2484
rect 4364 -2694 4370 -2484
rect 4420 -2524 4426 -2318
rect 4460 -2524 4466 -2318
rect 4502 -2484 4512 -2304
rect 4564 -2484 4574 -2304
rect 4612 -2318 4658 -2306
rect 4228 -2706 4274 -2704
rect 4324 -2706 4370 -2694
rect 4406 -2704 4416 -2524
rect 4468 -2704 4478 -2524
rect 4516 -2694 4522 -2484
rect 4556 -2694 4562 -2484
rect 4612 -2524 4618 -2318
rect 4652 -2524 4658 -2318
rect 4694 -2484 4704 -2304
rect 4756 -2484 4766 -2304
rect 4804 -2318 4850 -2306
rect 4420 -2706 4466 -2704
rect 4516 -2706 4562 -2694
rect 4598 -2704 4608 -2524
rect 4660 -2704 4670 -2524
rect 4708 -2694 4714 -2484
rect 4748 -2694 4754 -2484
rect 4804 -2524 4810 -2318
rect 4844 -2524 4850 -2318
rect 4612 -2706 4658 -2704
rect 4708 -2706 4754 -2694
rect 4790 -2704 4800 -2524
rect 4852 -2704 4862 -2524
rect 4804 -2706 4850 -2704
rect 4270 -2740 4328 -2738
rect 4462 -2740 4520 -2738
rect 4654 -2740 4712 -2738
rect 4892 -2740 4972 -2276
rect 5268 -2318 5314 -2306
rect 5268 -2524 5274 -2318
rect 5308 -2524 5314 -2318
rect 5350 -2484 5360 -2304
rect 5412 -2484 5422 -2304
rect 5460 -2318 5506 -2306
rect 5254 -2704 5264 -2524
rect 5316 -2704 5326 -2524
rect 5364 -2694 5370 -2484
rect 5404 -2694 5410 -2484
rect 5460 -2524 5466 -2318
rect 5500 -2524 5506 -2318
rect 5542 -2484 5552 -2304
rect 5604 -2484 5614 -2304
rect 5652 -2318 5698 -2306
rect 5268 -2706 5314 -2704
rect 5364 -2706 5410 -2694
rect 5446 -2704 5456 -2524
rect 5508 -2704 5518 -2524
rect 5556 -2694 5562 -2484
rect 5596 -2694 5602 -2484
rect 5652 -2524 5658 -2318
rect 5692 -2524 5698 -2318
rect 5734 -2484 5744 -2304
rect 5796 -2484 5806 -2304
rect 5844 -2318 5890 -2306
rect 5460 -2706 5506 -2704
rect 5556 -2706 5602 -2694
rect 5638 -2704 5648 -2524
rect 5700 -2704 5710 -2524
rect 5748 -2694 5754 -2484
rect 5788 -2694 5794 -2484
rect 5844 -2524 5850 -2318
rect 5884 -2524 5890 -2318
rect 5652 -2706 5698 -2704
rect 5748 -2706 5794 -2694
rect 5830 -2704 5840 -2524
rect 5892 -2704 5902 -2524
rect 5844 -2706 5890 -2704
rect 5310 -2740 5368 -2738
rect 5502 -2740 5560 -2738
rect 5694 -2740 5752 -2738
rect 5932 -2740 6012 -2276
rect 6308 -2318 6354 -2306
rect 6308 -2524 6314 -2318
rect 6348 -2524 6354 -2318
rect 6390 -2484 6400 -2304
rect 6452 -2484 6462 -2304
rect 6500 -2318 6546 -2306
rect 6294 -2704 6304 -2524
rect 6356 -2704 6366 -2524
rect 6404 -2694 6410 -2484
rect 6444 -2694 6450 -2484
rect 6500 -2524 6506 -2318
rect 6540 -2524 6546 -2318
rect 6582 -2484 6592 -2304
rect 6644 -2484 6654 -2304
rect 6692 -2318 6738 -2306
rect 6308 -2706 6354 -2704
rect 6404 -2706 6450 -2694
rect 6486 -2704 6496 -2524
rect 6548 -2704 6558 -2524
rect 6596 -2694 6602 -2484
rect 6636 -2694 6642 -2484
rect 6692 -2524 6698 -2318
rect 6732 -2524 6738 -2318
rect 6774 -2484 6784 -2304
rect 6836 -2484 6846 -2304
rect 6884 -2318 6930 -2306
rect 6500 -2706 6546 -2704
rect 6596 -2706 6642 -2694
rect 6678 -2704 6688 -2524
rect 6740 -2704 6750 -2524
rect 6788 -2694 6794 -2484
rect 6828 -2694 6834 -2484
rect 6884 -2524 6890 -2318
rect 6924 -2524 6930 -2318
rect 6692 -2706 6738 -2704
rect 6788 -2706 6834 -2694
rect 6870 -2704 6880 -2524
rect 6932 -2704 6942 -2524
rect 6884 -2706 6930 -2704
rect 6350 -2740 6408 -2738
rect 6542 -2740 6600 -2738
rect 6734 -2740 6792 -2738
rect 6972 -2740 7052 -2276
rect 7348 -2318 7394 -2306
rect 7348 -2524 7354 -2318
rect 7388 -2524 7394 -2318
rect 7430 -2484 7440 -2304
rect 7492 -2484 7502 -2304
rect 7540 -2318 7586 -2306
rect 7334 -2704 7344 -2524
rect 7396 -2704 7406 -2524
rect 7444 -2694 7450 -2484
rect 7484 -2694 7490 -2484
rect 7540 -2524 7546 -2318
rect 7580 -2524 7586 -2318
rect 7622 -2484 7632 -2304
rect 7684 -2484 7694 -2304
rect 7732 -2318 7778 -2306
rect 7348 -2706 7394 -2704
rect 7444 -2706 7490 -2694
rect 7526 -2704 7536 -2524
rect 7588 -2704 7598 -2524
rect 7636 -2694 7642 -2484
rect 7676 -2694 7682 -2484
rect 7732 -2524 7738 -2318
rect 7772 -2524 7778 -2318
rect 7814 -2484 7824 -2304
rect 7876 -2484 7886 -2304
rect 7924 -2318 7970 -2306
rect 7540 -2706 7586 -2704
rect 7636 -2706 7682 -2694
rect 7718 -2704 7728 -2524
rect 7780 -2704 7790 -2524
rect 7828 -2694 7834 -2484
rect 7868 -2694 7874 -2484
rect 7924 -2524 7930 -2318
rect 7964 -2524 7970 -2318
rect 7732 -2706 7778 -2704
rect 7828 -2706 7874 -2694
rect 7910 -2704 7920 -2524
rect 7972 -2704 7982 -2524
rect 7924 -2706 7970 -2704
rect 7390 -2740 7448 -2738
rect 7582 -2740 7640 -2738
rect 7774 -2740 7832 -2738
rect 8012 -2740 8092 -2276
rect 8388 -2318 8434 -2306
rect 8388 -2524 8394 -2318
rect 8428 -2524 8434 -2318
rect 8470 -2484 8480 -2304
rect 8532 -2484 8542 -2304
rect 8580 -2318 8626 -2306
rect 8374 -2704 8384 -2524
rect 8436 -2704 8446 -2524
rect 8484 -2694 8490 -2484
rect 8524 -2694 8530 -2484
rect 8580 -2524 8586 -2318
rect 8620 -2524 8626 -2318
rect 8662 -2484 8672 -2304
rect 8724 -2484 8734 -2304
rect 8772 -2318 8818 -2306
rect 8388 -2706 8434 -2704
rect 8484 -2706 8530 -2694
rect 8566 -2704 8576 -2524
rect 8628 -2704 8638 -2524
rect 8676 -2694 8682 -2484
rect 8716 -2694 8722 -2484
rect 8772 -2524 8778 -2318
rect 8812 -2524 8818 -2318
rect 8854 -2484 8864 -2304
rect 8916 -2484 8926 -2304
rect 8964 -2318 9010 -2306
rect 8580 -2706 8626 -2704
rect 8676 -2706 8722 -2694
rect 8758 -2704 8768 -2524
rect 8820 -2704 8830 -2524
rect 8868 -2694 8874 -2484
rect 8908 -2694 8914 -2484
rect 8964 -2524 8970 -2318
rect 9004 -2524 9010 -2318
rect 8772 -2706 8818 -2704
rect 8868 -2706 8914 -2694
rect 8950 -2704 8960 -2524
rect 9012 -2704 9022 -2524
rect 8964 -2706 9010 -2704
rect 8430 -2740 8488 -2738
rect 8622 -2740 8680 -2738
rect 8814 -2740 8872 -2738
rect 9052 -2740 9132 -2276
rect 11848 -2318 11894 -2306
rect 11848 -2524 11854 -2318
rect 11888 -2524 11894 -2318
rect 11930 -2484 11940 -2304
rect 11992 -2484 12002 -2304
rect 12040 -2318 12086 -2306
rect 11834 -2704 11844 -2524
rect 11896 -2704 11906 -2524
rect 11944 -2694 11950 -2484
rect 11984 -2694 11990 -2484
rect 12040 -2524 12046 -2318
rect 12080 -2524 12086 -2318
rect 12122 -2484 12132 -2304
rect 12184 -2484 12194 -2304
rect 12232 -2318 12278 -2306
rect 11848 -2706 11894 -2704
rect 11944 -2706 11990 -2694
rect 12026 -2704 12036 -2524
rect 12088 -2704 12098 -2524
rect 12136 -2694 12142 -2484
rect 12176 -2694 12182 -2484
rect 12232 -2524 12238 -2318
rect 12272 -2524 12278 -2318
rect 12314 -2484 12324 -2304
rect 12376 -2484 12386 -2304
rect 12424 -2318 12470 -2306
rect 12040 -2706 12086 -2704
rect 12136 -2706 12182 -2694
rect 12218 -2704 12228 -2524
rect 12280 -2704 12290 -2524
rect 12328 -2694 12334 -2484
rect 12368 -2694 12374 -2484
rect 12424 -2524 12430 -2318
rect 12464 -2524 12470 -2318
rect 12232 -2706 12278 -2704
rect 12328 -2706 12374 -2694
rect 12410 -2704 12420 -2524
rect 12472 -2704 12482 -2524
rect 12424 -2706 12470 -2704
rect 11890 -2740 11948 -2738
rect 12082 -2740 12140 -2738
rect 12274 -2740 12332 -2738
rect 12512 -2740 12592 -2276
rect 12888 -2318 12934 -2306
rect 12888 -2524 12894 -2318
rect 12928 -2524 12934 -2318
rect 12970 -2484 12980 -2304
rect 13032 -2484 13042 -2304
rect 13080 -2318 13126 -2306
rect 12874 -2704 12884 -2524
rect 12936 -2704 12946 -2524
rect 12984 -2694 12990 -2484
rect 13024 -2694 13030 -2484
rect 13080 -2524 13086 -2318
rect 13120 -2524 13126 -2318
rect 13162 -2484 13172 -2304
rect 13224 -2484 13234 -2304
rect 13272 -2318 13318 -2306
rect 12888 -2706 12934 -2704
rect 12984 -2706 13030 -2694
rect 13066 -2704 13076 -2524
rect 13128 -2704 13138 -2524
rect 13176 -2694 13182 -2484
rect 13216 -2694 13222 -2484
rect 13272 -2524 13278 -2318
rect 13312 -2524 13318 -2318
rect 13354 -2484 13364 -2304
rect 13416 -2484 13426 -2304
rect 13464 -2318 13510 -2306
rect 13080 -2706 13126 -2704
rect 13176 -2706 13222 -2694
rect 13258 -2704 13268 -2524
rect 13320 -2704 13330 -2524
rect 13368 -2694 13374 -2484
rect 13408 -2694 13414 -2484
rect 13464 -2524 13470 -2318
rect 13504 -2524 13510 -2318
rect 13272 -2706 13318 -2704
rect 13368 -2706 13414 -2694
rect 13450 -2704 13460 -2524
rect 13512 -2704 13522 -2524
rect 13464 -2706 13510 -2704
rect 12930 -2740 12988 -2738
rect 13122 -2740 13180 -2738
rect 13314 -2740 13372 -2738
rect 13552 -2740 13632 -2276
rect 13928 -2318 13974 -2306
rect 13928 -2524 13934 -2318
rect 13968 -2524 13974 -2318
rect 14010 -2484 14020 -2304
rect 14072 -2484 14082 -2304
rect 14120 -2318 14166 -2306
rect 13914 -2704 13924 -2524
rect 13976 -2704 13986 -2524
rect 14024 -2694 14030 -2484
rect 14064 -2694 14070 -2484
rect 14120 -2524 14126 -2318
rect 14160 -2524 14166 -2318
rect 14202 -2484 14212 -2304
rect 14264 -2484 14274 -2304
rect 14312 -2318 14358 -2306
rect 13928 -2706 13974 -2704
rect 14024 -2706 14070 -2694
rect 14106 -2704 14116 -2524
rect 14168 -2704 14178 -2524
rect 14216 -2694 14222 -2484
rect 14256 -2694 14262 -2484
rect 14312 -2524 14318 -2318
rect 14352 -2524 14358 -2318
rect 14394 -2484 14404 -2304
rect 14456 -2484 14466 -2304
rect 14504 -2318 14550 -2306
rect 14120 -2706 14166 -2704
rect 14216 -2706 14262 -2694
rect 14298 -2704 14308 -2524
rect 14360 -2704 14370 -2524
rect 14408 -2694 14414 -2484
rect 14448 -2694 14454 -2484
rect 14504 -2524 14510 -2318
rect 14544 -2524 14550 -2318
rect 14312 -2706 14358 -2704
rect 14408 -2706 14454 -2694
rect 14490 -2704 14500 -2524
rect 14552 -2704 14562 -2524
rect 14504 -2706 14550 -2704
rect 13970 -2740 14028 -2738
rect 14162 -2740 14220 -2738
rect 14354 -2740 14412 -2738
rect 14592 -2740 14672 -2276
rect 14968 -2318 15014 -2306
rect 14968 -2524 14974 -2318
rect 15008 -2524 15014 -2318
rect 15050 -2484 15060 -2304
rect 15112 -2484 15122 -2304
rect 15160 -2318 15206 -2306
rect 14954 -2704 14964 -2524
rect 15016 -2704 15026 -2524
rect 15064 -2694 15070 -2484
rect 15104 -2694 15110 -2484
rect 15160 -2524 15166 -2318
rect 15200 -2524 15206 -2318
rect 15242 -2484 15252 -2304
rect 15304 -2484 15314 -2304
rect 15352 -2318 15398 -2306
rect 14968 -2706 15014 -2704
rect 15064 -2706 15110 -2694
rect 15146 -2704 15156 -2524
rect 15208 -2704 15218 -2524
rect 15256 -2694 15262 -2484
rect 15296 -2694 15302 -2484
rect 15352 -2524 15358 -2318
rect 15392 -2524 15398 -2318
rect 15434 -2484 15444 -2304
rect 15496 -2484 15506 -2304
rect 15544 -2318 15590 -2306
rect 15160 -2706 15206 -2704
rect 15256 -2706 15302 -2694
rect 15338 -2704 15348 -2524
rect 15400 -2704 15410 -2524
rect 15448 -2694 15454 -2484
rect 15488 -2694 15494 -2484
rect 15544 -2524 15550 -2318
rect 15584 -2524 15590 -2318
rect 15352 -2706 15398 -2704
rect 15448 -2706 15494 -2694
rect 15530 -2704 15540 -2524
rect 15592 -2704 15602 -2524
rect 15544 -2706 15590 -2704
rect 15010 -2740 15068 -2738
rect 15202 -2740 15260 -2738
rect 15394 -2740 15452 -2738
rect 15632 -2740 15712 -2276
rect 16008 -2318 16054 -2306
rect 16008 -2524 16014 -2318
rect 16048 -2524 16054 -2318
rect 16090 -2484 16100 -2304
rect 16152 -2484 16162 -2304
rect 16200 -2318 16246 -2306
rect 15994 -2704 16004 -2524
rect 16056 -2704 16066 -2524
rect 16104 -2694 16110 -2484
rect 16144 -2694 16150 -2484
rect 16200 -2524 16206 -2318
rect 16240 -2524 16246 -2318
rect 16282 -2484 16292 -2304
rect 16344 -2484 16354 -2304
rect 16392 -2318 16438 -2306
rect 16008 -2706 16054 -2704
rect 16104 -2706 16150 -2694
rect 16186 -2704 16196 -2524
rect 16248 -2704 16258 -2524
rect 16296 -2694 16302 -2484
rect 16336 -2694 16342 -2484
rect 16392 -2524 16398 -2318
rect 16432 -2524 16438 -2318
rect 16474 -2484 16484 -2304
rect 16536 -2484 16546 -2304
rect 16584 -2318 16630 -2306
rect 16200 -2706 16246 -2704
rect 16296 -2706 16342 -2694
rect 16378 -2704 16388 -2524
rect 16440 -2704 16450 -2524
rect 16488 -2694 16494 -2484
rect 16528 -2694 16534 -2484
rect 16584 -2524 16590 -2318
rect 16624 -2524 16630 -2318
rect 16392 -2706 16438 -2704
rect 16488 -2706 16534 -2694
rect 16570 -2704 16580 -2524
rect 16632 -2704 16642 -2524
rect 16584 -2706 16630 -2704
rect 16050 -2740 16108 -2738
rect 16242 -2740 16300 -2738
rect 16434 -2740 16492 -2738
rect 16672 -2740 16752 -2276
rect 4264 -2744 4972 -2740
rect 4264 -2778 4282 -2744
rect 4316 -2778 4474 -2744
rect 4508 -2778 4666 -2744
rect 4700 -2778 4972 -2744
rect 4264 -2836 4972 -2778
rect 5304 -2744 6012 -2740
rect 5304 -2778 5322 -2744
rect 5356 -2778 5514 -2744
rect 5548 -2778 5706 -2744
rect 5740 -2778 6012 -2744
rect 5304 -2836 6012 -2778
rect 6344 -2744 7052 -2740
rect 6344 -2778 6362 -2744
rect 6396 -2778 6554 -2744
rect 6588 -2778 6746 -2744
rect 6780 -2778 7052 -2744
rect 6344 -2836 7052 -2778
rect 7384 -2744 8092 -2740
rect 7384 -2778 7402 -2744
rect 7436 -2778 7594 -2744
rect 7628 -2778 7786 -2744
rect 7820 -2778 8092 -2744
rect 7384 -2836 8092 -2778
rect 8424 -2744 9132 -2740
rect 8424 -2778 8442 -2744
rect 8476 -2778 8634 -2744
rect 8668 -2778 8826 -2744
rect 8860 -2778 9132 -2744
rect 8424 -2836 9132 -2778
rect 11884 -2744 12592 -2740
rect 11884 -2778 11902 -2744
rect 11936 -2778 12094 -2744
rect 12128 -2778 12286 -2744
rect 12320 -2778 12592 -2744
rect 11884 -2836 12592 -2778
rect 12924 -2744 13632 -2740
rect 12924 -2778 12942 -2744
rect 12976 -2778 13134 -2744
rect 13168 -2778 13326 -2744
rect 13360 -2778 13632 -2744
rect 12924 -2836 13632 -2778
rect 13964 -2744 14672 -2740
rect 13964 -2778 13982 -2744
rect 14016 -2778 14174 -2744
rect 14208 -2778 14366 -2744
rect 14400 -2778 14672 -2744
rect 13964 -2836 14672 -2778
rect 15004 -2744 15712 -2740
rect 15004 -2778 15022 -2744
rect 15056 -2778 15214 -2744
rect 15248 -2778 15406 -2744
rect 15440 -2778 15712 -2744
rect 15004 -2836 15712 -2778
rect 16044 -2744 16752 -2740
rect 16044 -2778 16062 -2744
rect 16096 -2778 16254 -2744
rect 16288 -2778 16446 -2744
rect 16480 -2778 16752 -2744
rect 16044 -2836 16752 -2778
rect -7370 -2946 -6662 -2942
rect -7370 -2980 -7352 -2946
rect -7318 -2980 -7160 -2946
rect -7126 -2980 -6968 -2946
rect -6934 -2980 -6662 -2946
rect -7370 -3038 -6662 -2980
rect 4836 -3012 4920 -2836
rect 5876 -3012 5960 -2836
rect 6916 -3012 7000 -2836
rect 7956 -3012 8040 -2836
rect 8996 -3012 9080 -2836
rect 12456 -3012 12540 -2836
rect 13496 -3012 13580 -2836
rect 14536 -3012 14620 -2836
rect 15576 -3012 15660 -2836
rect 16616 -3012 16700 -2836
rect 4272 -3038 5088 -3012
rect -6798 -3214 -6714 -3038
rect 4272 -3072 4293 -3038
rect 4327 -3072 4411 -3038
rect 4445 -3072 4529 -3038
rect 4563 -3072 4647 -3038
rect 4681 -3072 4765 -3038
rect 4799 -3072 4883 -3038
rect 4917 -3072 5088 -3038
rect 4272 -3080 5088 -3072
rect 5312 -3038 6128 -3012
rect 5312 -3072 5333 -3038
rect 5367 -3072 5451 -3038
rect 5485 -3072 5569 -3038
rect 5603 -3072 5687 -3038
rect 5721 -3072 5805 -3038
rect 5839 -3072 5923 -3038
rect 5957 -3072 6128 -3038
rect 5312 -3080 6128 -3072
rect 6352 -3038 7168 -3012
rect 6352 -3072 6373 -3038
rect 6407 -3072 6491 -3038
rect 6525 -3072 6609 -3038
rect 6643 -3072 6727 -3038
rect 6761 -3072 6845 -3038
rect 6879 -3072 6963 -3038
rect 6997 -3072 7168 -3038
rect 6352 -3080 7168 -3072
rect 7392 -3038 8208 -3012
rect 7392 -3072 7413 -3038
rect 7447 -3072 7531 -3038
rect 7565 -3072 7649 -3038
rect 7683 -3072 7767 -3038
rect 7801 -3072 7885 -3038
rect 7919 -3072 8003 -3038
rect 8037 -3072 8208 -3038
rect 7392 -3080 8208 -3072
rect 8432 -3038 9248 -3012
rect 8432 -3072 8453 -3038
rect 8487 -3072 8571 -3038
rect 8605 -3072 8689 -3038
rect 8723 -3072 8807 -3038
rect 8841 -3072 8925 -3038
rect 8959 -3072 9043 -3038
rect 9077 -3072 9248 -3038
rect 8432 -3080 9248 -3072
rect 11892 -3038 12708 -3012
rect 11892 -3072 11913 -3038
rect 11947 -3072 12031 -3038
rect 12065 -3072 12149 -3038
rect 12183 -3072 12267 -3038
rect 12301 -3072 12385 -3038
rect 12419 -3072 12503 -3038
rect 12537 -3072 12708 -3038
rect 11892 -3080 12708 -3072
rect 12932 -3038 13748 -3012
rect 12932 -3072 12953 -3038
rect 12987 -3072 13071 -3038
rect 13105 -3072 13189 -3038
rect 13223 -3072 13307 -3038
rect 13341 -3072 13425 -3038
rect 13459 -3072 13543 -3038
rect 13577 -3072 13748 -3038
rect 12932 -3080 13748 -3072
rect 13972 -3038 14788 -3012
rect 13972 -3072 13993 -3038
rect 14027 -3072 14111 -3038
rect 14145 -3072 14229 -3038
rect 14263 -3072 14347 -3038
rect 14381 -3072 14465 -3038
rect 14499 -3072 14583 -3038
rect 14617 -3072 14788 -3038
rect 13972 -3080 14788 -3072
rect 15012 -3038 15828 -3012
rect 15012 -3072 15033 -3038
rect 15067 -3072 15151 -3038
rect 15185 -3072 15269 -3038
rect 15303 -3072 15387 -3038
rect 15421 -3072 15505 -3038
rect 15539 -3072 15623 -3038
rect 15657 -3072 15828 -3038
rect 15012 -3080 15828 -3072
rect 16052 -3038 16868 -3012
rect 16052 -3072 16073 -3038
rect 16107 -3072 16191 -3038
rect 16225 -3072 16309 -3038
rect 16343 -3072 16427 -3038
rect 16461 -3072 16545 -3038
rect 16579 -3072 16663 -3038
rect 16697 -3072 16868 -3038
rect 16052 -3080 16868 -3072
rect 4228 -3122 4274 -3110
rect -7362 -3240 -6546 -3214
rect -7362 -3274 -7341 -3240
rect -7307 -3274 -7223 -3240
rect -7189 -3274 -7105 -3240
rect -7071 -3274 -6987 -3240
rect -6953 -3274 -6869 -3240
rect -6835 -3274 -6751 -3240
rect -6717 -3274 -6546 -3240
rect -7362 -3282 -6546 -3274
rect -7406 -3324 -7360 -3312
rect -7406 -3534 -7400 -3324
rect -7366 -3534 -7360 -3324
rect -7300 -3490 -7290 -3310
rect -7238 -3490 -7228 -3310
rect -7170 -3324 -7124 -3312
rect -7420 -3714 -7410 -3534
rect -7358 -3714 -7348 -3534
rect -7288 -3700 -7282 -3490
rect -7248 -3700 -7242 -3490
rect -7170 -3534 -7164 -3324
rect -7130 -3534 -7124 -3324
rect -7064 -3490 -7054 -3310
rect -7002 -3490 -6992 -3310
rect -6934 -3324 -6888 -3312
rect -7288 -3712 -7242 -3700
rect -7184 -3714 -7174 -3534
rect -7122 -3714 -7112 -3534
rect -7052 -3700 -7046 -3490
rect -7012 -3700 -7006 -3490
rect -6934 -3534 -6928 -3324
rect -6894 -3534 -6888 -3324
rect -6828 -3490 -6818 -3310
rect -6766 -3490 -6756 -3310
rect -6698 -3324 -6652 -3312
rect -7052 -3712 -7006 -3700
rect -6948 -3714 -6938 -3534
rect -6886 -3714 -6876 -3534
rect -6816 -3700 -6810 -3490
rect -6776 -3700 -6770 -3490
rect -6698 -3534 -6692 -3324
rect -6658 -3534 -6652 -3324
rect -6816 -3712 -6770 -3700
rect -6712 -3714 -6702 -3534
rect -6650 -3714 -6640 -3534
rect -6610 -3742 -6546 -3282
rect 4228 -3332 4234 -3122
rect 4268 -3332 4274 -3122
rect 4334 -3288 4344 -3108
rect 4396 -3288 4406 -3108
rect 4464 -3122 4510 -3110
rect 4214 -3512 4224 -3332
rect 4276 -3512 4286 -3332
rect 4346 -3498 4352 -3288
rect 4386 -3498 4392 -3288
rect 4464 -3332 4470 -3122
rect 4504 -3332 4510 -3122
rect 4570 -3288 4580 -3108
rect 4632 -3288 4642 -3108
rect 4700 -3122 4746 -3110
rect 4346 -3510 4392 -3498
rect 4450 -3512 4460 -3332
rect 4512 -3512 4522 -3332
rect 4582 -3498 4588 -3288
rect 4622 -3498 4628 -3288
rect 4700 -3332 4706 -3122
rect 4740 -3332 4746 -3122
rect 4806 -3288 4816 -3108
rect 4868 -3288 4878 -3108
rect 4936 -3122 4982 -3110
rect 4582 -3510 4628 -3498
rect 4686 -3512 4696 -3332
rect 4748 -3512 4758 -3332
rect 4818 -3498 4824 -3288
rect 4858 -3498 4864 -3288
rect 4936 -3332 4942 -3122
rect 4976 -3332 4982 -3122
rect 4818 -3510 4864 -3498
rect 4922 -3512 4932 -3332
rect 4984 -3512 4994 -3332
rect 5024 -3540 5088 -3080
rect 5268 -3122 5314 -3110
rect 5268 -3332 5274 -3122
rect 5308 -3332 5314 -3122
rect 5374 -3288 5384 -3108
rect 5436 -3288 5446 -3108
rect 5504 -3122 5550 -3110
rect 5254 -3512 5264 -3332
rect 5316 -3512 5326 -3332
rect 5386 -3498 5392 -3288
rect 5426 -3498 5432 -3288
rect 5504 -3332 5510 -3122
rect 5544 -3332 5550 -3122
rect 5610 -3288 5620 -3108
rect 5672 -3288 5682 -3108
rect 5740 -3122 5786 -3110
rect 5386 -3510 5432 -3498
rect 5490 -3512 5500 -3332
rect 5552 -3512 5562 -3332
rect 5622 -3498 5628 -3288
rect 5662 -3498 5668 -3288
rect 5740 -3332 5746 -3122
rect 5780 -3332 5786 -3122
rect 5846 -3288 5856 -3108
rect 5908 -3288 5918 -3108
rect 5976 -3122 6022 -3110
rect 5622 -3510 5668 -3498
rect 5726 -3512 5736 -3332
rect 5788 -3512 5798 -3332
rect 5858 -3498 5864 -3288
rect 5898 -3498 5904 -3288
rect 5976 -3332 5982 -3122
rect 6016 -3332 6022 -3122
rect 5858 -3510 5904 -3498
rect 5962 -3512 5972 -3332
rect 6024 -3512 6034 -3332
rect 6064 -3540 6128 -3080
rect 6308 -3122 6354 -3110
rect 6308 -3332 6314 -3122
rect 6348 -3332 6354 -3122
rect 6414 -3288 6424 -3108
rect 6476 -3288 6486 -3108
rect 6544 -3122 6590 -3110
rect 6294 -3512 6304 -3332
rect 6356 -3512 6366 -3332
rect 6426 -3498 6432 -3288
rect 6466 -3498 6472 -3288
rect 6544 -3332 6550 -3122
rect 6584 -3332 6590 -3122
rect 6650 -3288 6660 -3108
rect 6712 -3288 6722 -3108
rect 6780 -3122 6826 -3110
rect 6426 -3510 6472 -3498
rect 6530 -3512 6540 -3332
rect 6592 -3512 6602 -3332
rect 6662 -3498 6668 -3288
rect 6702 -3498 6708 -3288
rect 6780 -3332 6786 -3122
rect 6820 -3332 6826 -3122
rect 6886 -3288 6896 -3108
rect 6948 -3288 6958 -3108
rect 7016 -3122 7062 -3110
rect 6662 -3510 6708 -3498
rect 6766 -3512 6776 -3332
rect 6828 -3512 6838 -3332
rect 6898 -3498 6904 -3288
rect 6938 -3498 6944 -3288
rect 7016 -3332 7022 -3122
rect 7056 -3332 7062 -3122
rect 6898 -3510 6944 -3498
rect 7002 -3512 7012 -3332
rect 7064 -3512 7074 -3332
rect 7104 -3540 7168 -3080
rect 7348 -3122 7394 -3110
rect 7348 -3332 7354 -3122
rect 7388 -3332 7394 -3122
rect 7454 -3288 7464 -3108
rect 7516 -3288 7526 -3108
rect 7584 -3122 7630 -3110
rect 7334 -3512 7344 -3332
rect 7396 -3512 7406 -3332
rect 7466 -3498 7472 -3288
rect 7506 -3498 7512 -3288
rect 7584 -3332 7590 -3122
rect 7624 -3332 7630 -3122
rect 7690 -3288 7700 -3108
rect 7752 -3288 7762 -3108
rect 7820 -3122 7866 -3110
rect 7466 -3510 7512 -3498
rect 7570 -3512 7580 -3332
rect 7632 -3512 7642 -3332
rect 7702 -3498 7708 -3288
rect 7742 -3498 7748 -3288
rect 7820 -3332 7826 -3122
rect 7860 -3332 7866 -3122
rect 7926 -3288 7936 -3108
rect 7988 -3288 7998 -3108
rect 8056 -3122 8102 -3110
rect 7702 -3510 7748 -3498
rect 7806 -3512 7816 -3332
rect 7868 -3512 7878 -3332
rect 7938 -3498 7944 -3288
rect 7978 -3498 7984 -3288
rect 8056 -3332 8062 -3122
rect 8096 -3332 8102 -3122
rect 7938 -3510 7984 -3498
rect 8042 -3512 8052 -3332
rect 8104 -3512 8114 -3332
rect 8144 -3540 8208 -3080
rect 8388 -3122 8434 -3110
rect 8388 -3332 8394 -3122
rect 8428 -3332 8434 -3122
rect 8494 -3288 8504 -3108
rect 8556 -3288 8566 -3108
rect 8624 -3122 8670 -3110
rect 8374 -3512 8384 -3332
rect 8436 -3512 8446 -3332
rect 8506 -3498 8512 -3288
rect 8546 -3498 8552 -3288
rect 8624 -3332 8630 -3122
rect 8664 -3332 8670 -3122
rect 8730 -3288 8740 -3108
rect 8792 -3288 8802 -3108
rect 8860 -3122 8906 -3110
rect 8506 -3510 8552 -3498
rect 8610 -3512 8620 -3332
rect 8672 -3512 8682 -3332
rect 8742 -3498 8748 -3288
rect 8782 -3498 8788 -3288
rect 8860 -3332 8866 -3122
rect 8900 -3332 8906 -3122
rect 8966 -3288 8976 -3108
rect 9028 -3288 9038 -3108
rect 9096 -3122 9142 -3110
rect 8742 -3510 8788 -3498
rect 8846 -3512 8856 -3332
rect 8908 -3512 8918 -3332
rect 8978 -3498 8984 -3288
rect 9018 -3498 9024 -3288
rect 9096 -3332 9102 -3122
rect 9136 -3332 9142 -3122
rect 8978 -3510 9024 -3498
rect 9082 -3512 9092 -3332
rect 9144 -3512 9154 -3332
rect 9184 -3540 9248 -3080
rect 11848 -3122 11894 -3110
rect 11848 -3332 11854 -3122
rect 11888 -3332 11894 -3122
rect 11954 -3288 11964 -3108
rect 12016 -3288 12026 -3108
rect 12084 -3122 12130 -3110
rect 11834 -3512 11844 -3332
rect 11896 -3512 11906 -3332
rect 11966 -3498 11972 -3288
rect 12006 -3498 12012 -3288
rect 12084 -3332 12090 -3122
rect 12124 -3332 12130 -3122
rect 12190 -3288 12200 -3108
rect 12252 -3288 12262 -3108
rect 12320 -3122 12366 -3110
rect 11966 -3510 12012 -3498
rect 12070 -3512 12080 -3332
rect 12132 -3512 12142 -3332
rect 12202 -3498 12208 -3288
rect 12242 -3498 12248 -3288
rect 12320 -3332 12326 -3122
rect 12360 -3332 12366 -3122
rect 12426 -3288 12436 -3108
rect 12488 -3288 12498 -3108
rect 12556 -3122 12602 -3110
rect 12202 -3510 12248 -3498
rect 12306 -3512 12316 -3332
rect 12368 -3512 12378 -3332
rect 12438 -3498 12444 -3288
rect 12478 -3498 12484 -3288
rect 12556 -3332 12562 -3122
rect 12596 -3332 12602 -3122
rect 12438 -3510 12484 -3498
rect 12542 -3512 12552 -3332
rect 12604 -3512 12614 -3332
rect 12644 -3540 12708 -3080
rect 12888 -3122 12934 -3110
rect 12888 -3332 12894 -3122
rect 12928 -3332 12934 -3122
rect 12994 -3288 13004 -3108
rect 13056 -3288 13066 -3108
rect 13124 -3122 13170 -3110
rect 12874 -3512 12884 -3332
rect 12936 -3512 12946 -3332
rect 13006 -3498 13012 -3288
rect 13046 -3498 13052 -3288
rect 13124 -3332 13130 -3122
rect 13164 -3332 13170 -3122
rect 13230 -3288 13240 -3108
rect 13292 -3288 13302 -3108
rect 13360 -3122 13406 -3110
rect 13006 -3510 13052 -3498
rect 13110 -3512 13120 -3332
rect 13172 -3512 13182 -3332
rect 13242 -3498 13248 -3288
rect 13282 -3498 13288 -3288
rect 13360 -3332 13366 -3122
rect 13400 -3332 13406 -3122
rect 13466 -3288 13476 -3108
rect 13528 -3288 13538 -3108
rect 13596 -3122 13642 -3110
rect 13242 -3510 13288 -3498
rect 13346 -3512 13356 -3332
rect 13408 -3512 13418 -3332
rect 13478 -3498 13484 -3288
rect 13518 -3498 13524 -3288
rect 13596 -3332 13602 -3122
rect 13636 -3332 13642 -3122
rect 13478 -3510 13524 -3498
rect 13582 -3512 13592 -3332
rect 13644 -3512 13654 -3332
rect 13684 -3540 13748 -3080
rect 13928 -3122 13974 -3110
rect 13928 -3332 13934 -3122
rect 13968 -3332 13974 -3122
rect 14034 -3288 14044 -3108
rect 14096 -3288 14106 -3108
rect 14164 -3122 14210 -3110
rect 13914 -3512 13924 -3332
rect 13976 -3512 13986 -3332
rect 14046 -3498 14052 -3288
rect 14086 -3498 14092 -3288
rect 14164 -3332 14170 -3122
rect 14204 -3332 14210 -3122
rect 14270 -3288 14280 -3108
rect 14332 -3288 14342 -3108
rect 14400 -3122 14446 -3110
rect 14046 -3510 14092 -3498
rect 14150 -3512 14160 -3332
rect 14212 -3512 14222 -3332
rect 14282 -3498 14288 -3288
rect 14322 -3498 14328 -3288
rect 14400 -3332 14406 -3122
rect 14440 -3332 14446 -3122
rect 14506 -3288 14516 -3108
rect 14568 -3288 14578 -3108
rect 14636 -3122 14682 -3110
rect 14282 -3510 14328 -3498
rect 14386 -3512 14396 -3332
rect 14448 -3512 14458 -3332
rect 14518 -3498 14524 -3288
rect 14558 -3498 14564 -3288
rect 14636 -3332 14642 -3122
rect 14676 -3332 14682 -3122
rect 14518 -3510 14564 -3498
rect 14622 -3512 14632 -3332
rect 14684 -3512 14694 -3332
rect 14724 -3540 14788 -3080
rect 14968 -3122 15014 -3110
rect 14968 -3332 14974 -3122
rect 15008 -3332 15014 -3122
rect 15074 -3288 15084 -3108
rect 15136 -3288 15146 -3108
rect 15204 -3122 15250 -3110
rect 14954 -3512 14964 -3332
rect 15016 -3512 15026 -3332
rect 15086 -3498 15092 -3288
rect 15126 -3498 15132 -3288
rect 15204 -3332 15210 -3122
rect 15244 -3332 15250 -3122
rect 15310 -3288 15320 -3108
rect 15372 -3288 15382 -3108
rect 15440 -3122 15486 -3110
rect 15086 -3510 15132 -3498
rect 15190 -3512 15200 -3332
rect 15252 -3512 15262 -3332
rect 15322 -3498 15328 -3288
rect 15362 -3498 15368 -3288
rect 15440 -3332 15446 -3122
rect 15480 -3332 15486 -3122
rect 15546 -3288 15556 -3108
rect 15608 -3288 15618 -3108
rect 15676 -3122 15722 -3110
rect 15322 -3510 15368 -3498
rect 15426 -3512 15436 -3332
rect 15488 -3512 15498 -3332
rect 15558 -3498 15564 -3288
rect 15598 -3498 15604 -3288
rect 15676 -3332 15682 -3122
rect 15716 -3332 15722 -3122
rect 15558 -3510 15604 -3498
rect 15662 -3512 15672 -3332
rect 15724 -3512 15734 -3332
rect 15764 -3540 15828 -3080
rect 16008 -3122 16054 -3110
rect 16008 -3332 16014 -3122
rect 16048 -3332 16054 -3122
rect 16114 -3288 16124 -3108
rect 16176 -3288 16186 -3108
rect 16244 -3122 16290 -3110
rect 15994 -3512 16004 -3332
rect 16056 -3512 16066 -3332
rect 16126 -3498 16132 -3288
rect 16166 -3498 16172 -3288
rect 16244 -3332 16250 -3122
rect 16284 -3332 16290 -3122
rect 16350 -3288 16360 -3108
rect 16412 -3288 16422 -3108
rect 16480 -3122 16526 -3110
rect 16126 -3510 16172 -3498
rect 16230 -3512 16240 -3332
rect 16292 -3512 16302 -3332
rect 16362 -3498 16368 -3288
rect 16402 -3498 16408 -3288
rect 16480 -3332 16486 -3122
rect 16520 -3332 16526 -3122
rect 16586 -3288 16596 -3108
rect 16648 -3288 16658 -3108
rect 16716 -3122 16762 -3110
rect 16362 -3510 16408 -3498
rect 16466 -3512 16476 -3332
rect 16528 -3512 16538 -3332
rect 16598 -3498 16604 -3288
rect 16638 -3498 16644 -3288
rect 16716 -3332 16722 -3122
rect 16756 -3332 16762 -3122
rect 16598 -3510 16644 -3498
rect 16702 -3512 16712 -3332
rect 16764 -3512 16774 -3332
rect 16804 -3540 16868 -3080
rect 4276 -3548 5088 -3540
rect 4276 -3582 4293 -3548
rect 4327 -3582 4411 -3548
rect 4445 -3582 4529 -3548
rect 4563 -3582 4647 -3548
rect 4681 -3582 4765 -3548
rect 4799 -3582 4883 -3548
rect 4917 -3582 5088 -3548
rect 4276 -3608 5088 -3582
rect 5316 -3548 6128 -3540
rect 5316 -3582 5333 -3548
rect 5367 -3582 5451 -3548
rect 5485 -3582 5569 -3548
rect 5603 -3582 5687 -3548
rect 5721 -3582 5805 -3548
rect 5839 -3582 5923 -3548
rect 5957 -3582 6128 -3548
rect 5316 -3608 6128 -3582
rect 6356 -3548 7168 -3540
rect 6356 -3582 6373 -3548
rect 6407 -3582 6491 -3548
rect 6525 -3582 6609 -3548
rect 6643 -3582 6727 -3548
rect 6761 -3582 6845 -3548
rect 6879 -3582 6963 -3548
rect 6997 -3582 7168 -3548
rect 6356 -3608 7168 -3582
rect 7396 -3548 8208 -3540
rect 7396 -3582 7413 -3548
rect 7447 -3582 7531 -3548
rect 7565 -3582 7649 -3548
rect 7683 -3582 7767 -3548
rect 7801 -3582 7885 -3548
rect 7919 -3582 8003 -3548
rect 8037 -3582 8208 -3548
rect 7396 -3608 8208 -3582
rect 8436 -3548 9248 -3540
rect 8436 -3582 8453 -3548
rect 8487 -3582 8571 -3548
rect 8605 -3582 8689 -3548
rect 8723 -3582 8807 -3548
rect 8841 -3582 8925 -3548
rect 8959 -3582 9043 -3548
rect 9077 -3582 9248 -3548
rect 8436 -3608 9248 -3582
rect 11896 -3548 12708 -3540
rect 11896 -3582 11913 -3548
rect 11947 -3582 12031 -3548
rect 12065 -3582 12149 -3548
rect 12183 -3582 12267 -3548
rect 12301 -3582 12385 -3548
rect 12419 -3582 12503 -3548
rect 12537 -3582 12708 -3548
rect 11896 -3608 12708 -3582
rect 12936 -3548 13748 -3540
rect 12936 -3582 12953 -3548
rect 12987 -3582 13071 -3548
rect 13105 -3582 13189 -3548
rect 13223 -3582 13307 -3548
rect 13341 -3582 13425 -3548
rect 13459 -3582 13543 -3548
rect 13577 -3582 13748 -3548
rect 12936 -3608 13748 -3582
rect 13976 -3548 14788 -3540
rect 13976 -3582 13993 -3548
rect 14027 -3582 14111 -3548
rect 14145 -3582 14229 -3548
rect 14263 -3582 14347 -3548
rect 14381 -3582 14465 -3548
rect 14499 -3582 14583 -3548
rect 14617 -3582 14788 -3548
rect 13976 -3608 14788 -3582
rect 15016 -3548 15828 -3540
rect 15016 -3582 15033 -3548
rect 15067 -3582 15151 -3548
rect 15185 -3582 15269 -3548
rect 15303 -3582 15387 -3548
rect 15421 -3582 15505 -3548
rect 15539 -3582 15623 -3548
rect 15657 -3582 15828 -3548
rect 15016 -3608 15828 -3582
rect 16056 -3548 16868 -3540
rect 16056 -3582 16073 -3548
rect 16107 -3582 16191 -3548
rect 16225 -3582 16309 -3548
rect 16343 -3582 16427 -3548
rect 16461 -3582 16545 -3548
rect 16579 -3582 16663 -3548
rect 16697 -3582 16868 -3548
rect 16056 -3608 16868 -3582
rect -7358 -3750 -6546 -3742
rect -7358 -3784 -7341 -3750
rect -7307 -3784 -7223 -3750
rect -7189 -3784 -7105 -3750
rect -7071 -3784 -6987 -3750
rect -6953 -3784 -6869 -3750
rect -6835 -3784 -6751 -3750
rect -6717 -3784 -6546 -3750
rect -7358 -3810 -6546 -3784
rect 4912 -3720 5236 -3714
rect 4912 -3840 4924 -3720
rect 5224 -3840 5236 -3720
rect 4912 -3846 5236 -3840
rect 8552 -3720 8876 -3714
rect 8552 -3840 8564 -3720
rect 8864 -3840 8876 -3720
rect 8552 -3846 8876 -3840
rect 12532 -3720 12856 -3714
rect 12532 -3840 12544 -3720
rect 12844 -3840 12856 -3720
rect 12532 -3846 12856 -3840
rect 16172 -3720 16496 -3714
rect 16172 -3840 16184 -3720
rect 16484 -3840 16496 -3720
rect 16172 -3846 16496 -3840
rect -7242 -3862 -6938 -3856
rect -7242 -3982 -7230 -3862
rect -6950 -3982 -6938 -3862
rect -7242 -3988 -6938 -3982
<< via1 >>
rect -28 6584 384 6588
rect -1456 6187 -1418 6580
rect -1418 6187 -1168 6580
rect -1168 6187 -1044 6580
rect -28 6192 94 6584
rect 94 6192 344 6584
rect 344 6192 384 6584
rect 2772 6584 3184 6588
rect -1456 6184 -1044 6187
rect 1344 6187 1382 6580
rect 1382 6187 1632 6580
rect 1632 6187 1756 6580
rect 2772 6192 2894 6584
rect 2894 6192 3144 6584
rect 3144 6192 3184 6584
rect 1344 6184 1756 6187
rect -916 5368 -790 5744
rect -790 5368 -662 5744
rect -662 5368 -412 5744
rect -412 5368 -284 5744
rect -284 5368 -144 5744
rect 1884 5368 2010 5744
rect 2010 5368 2138 5744
rect 2138 5368 2388 5744
rect 2388 5368 2516 5744
rect 2516 5368 2656 5744
rect -28 5216 384 5220
rect -1456 4819 -1418 5212
rect -1418 4819 -1168 5212
rect -1168 4819 -1044 5212
rect -28 4824 94 5216
rect 94 4824 344 5216
rect 344 4824 384 5216
rect 2772 5216 3184 5220
rect -1456 4816 -1044 4819
rect 1344 4819 1382 5212
rect 1382 4819 1632 5212
rect 1632 4819 1756 5212
rect 2772 4824 2894 5216
rect 2894 4824 3144 5216
rect 3144 4824 3184 5216
rect 4520 5452 4572 5468
rect 4520 5284 4530 5452
rect 4530 5284 4564 5452
rect 4564 5284 4572 5452
rect 4424 5076 4434 5248
rect 4434 5076 4468 5248
rect 4468 5076 4476 5248
rect 4424 5064 4476 5076
rect 4712 5452 4764 5468
rect 4712 5284 4722 5452
rect 4722 5284 4756 5452
rect 4756 5284 4764 5452
rect 4616 5076 4626 5248
rect 4626 5076 4660 5248
rect 4660 5076 4668 5248
rect 4616 5064 4668 5076
rect 4904 5452 4956 5468
rect 4904 5284 4914 5452
rect 4914 5284 4948 5452
rect 4948 5284 4956 5452
rect 4808 5076 4818 5248
rect 4818 5076 4852 5248
rect 4852 5076 4860 5248
rect 4808 5064 4860 5076
rect 5096 5452 5148 5468
rect 5096 5284 5106 5452
rect 5106 5284 5140 5452
rect 5140 5284 5148 5452
rect 5000 5076 5010 5248
rect 5010 5076 5044 5248
rect 5044 5076 5052 5248
rect 5000 5064 5052 5076
rect 5288 5452 5340 5468
rect 5288 5284 5298 5452
rect 5298 5284 5332 5452
rect 5332 5284 5340 5452
rect 5192 5076 5202 5248
rect 5202 5076 5236 5248
rect 5236 5076 5244 5248
rect 5192 5064 5244 5076
rect 5480 5452 5532 5468
rect 5480 5284 5490 5452
rect 5490 5284 5524 5452
rect 5524 5284 5532 5452
rect 5384 5076 5394 5248
rect 5394 5076 5428 5248
rect 5428 5076 5436 5248
rect 5384 5064 5436 5076
rect 5672 5452 5724 5468
rect 5672 5284 5682 5452
rect 5682 5284 5716 5452
rect 5716 5284 5724 5452
rect 5576 5076 5586 5248
rect 5586 5076 5620 5248
rect 5620 5076 5628 5248
rect 5576 5064 5628 5076
rect 5864 5452 5916 5468
rect 5864 5284 5874 5452
rect 5874 5284 5908 5452
rect 5908 5284 5916 5452
rect 5768 5076 5778 5248
rect 5778 5076 5812 5248
rect 5812 5076 5820 5248
rect 5768 5064 5820 5076
rect 6056 5452 6108 5468
rect 6056 5284 6066 5452
rect 6066 5284 6100 5452
rect 6100 5284 6108 5452
rect 5960 5076 5970 5248
rect 5970 5076 6004 5248
rect 6004 5076 6012 5248
rect 5960 5064 6012 5076
rect 6248 5452 6300 5468
rect 6248 5284 6258 5452
rect 6258 5284 6292 5452
rect 6292 5284 6300 5452
rect 6152 5076 6162 5248
rect 6162 5076 6196 5248
rect 6196 5076 6204 5248
rect 6152 5064 6204 5076
rect 6440 5452 6492 5468
rect 6440 5284 6450 5452
rect 6450 5284 6484 5452
rect 6484 5284 6492 5452
rect 6344 5076 6354 5248
rect 6354 5076 6388 5248
rect 6388 5076 6396 5248
rect 6344 5064 6396 5076
rect 6632 5452 6684 5468
rect 6632 5284 6642 5452
rect 6642 5284 6676 5452
rect 6676 5284 6684 5452
rect 6536 5076 6546 5248
rect 6546 5076 6580 5248
rect 6580 5076 6588 5248
rect 6536 5064 6588 5076
rect 6824 5452 6876 5468
rect 6824 5284 6834 5452
rect 6834 5284 6868 5452
rect 6868 5284 6876 5452
rect 6728 5076 6738 5248
rect 6738 5076 6772 5248
rect 6772 5076 6780 5248
rect 6728 5064 6780 5076
rect 7016 5452 7068 5468
rect 7016 5284 7026 5452
rect 7026 5284 7060 5452
rect 7060 5284 7068 5452
rect 6920 5076 6930 5248
rect 6930 5076 6964 5248
rect 6964 5076 6972 5248
rect 6920 5064 6972 5076
rect 7208 5452 7260 5468
rect 7208 5284 7218 5452
rect 7218 5284 7252 5452
rect 7252 5284 7260 5452
rect 7112 5076 7122 5248
rect 7122 5076 7156 5248
rect 7156 5076 7164 5248
rect 7112 5064 7164 5076
rect 7304 5076 7314 5248
rect 7314 5076 7348 5248
rect 7348 5076 7356 5248
rect 7304 5064 7356 5076
rect 8160 5452 8212 5468
rect 8160 5284 8170 5452
rect 8170 5284 8204 5452
rect 8204 5284 8212 5452
rect 8064 5076 8074 5248
rect 8074 5076 8108 5248
rect 8108 5076 8116 5248
rect 8064 5064 8116 5076
rect 8352 5452 8404 5468
rect 8352 5284 8362 5452
rect 8362 5284 8396 5452
rect 8396 5284 8404 5452
rect 8256 5076 8266 5248
rect 8266 5076 8300 5248
rect 8300 5076 8308 5248
rect 8256 5064 8308 5076
rect 8544 5452 8596 5468
rect 8544 5284 8554 5452
rect 8554 5284 8588 5452
rect 8588 5284 8596 5452
rect 8448 5076 8458 5248
rect 8458 5076 8492 5248
rect 8492 5076 8500 5248
rect 8448 5064 8500 5076
rect 8736 5452 8788 5468
rect 8736 5284 8746 5452
rect 8746 5284 8780 5452
rect 8780 5284 8788 5452
rect 8640 5076 8650 5248
rect 8650 5076 8684 5248
rect 8684 5076 8692 5248
rect 8640 5064 8692 5076
rect 8928 5452 8980 5468
rect 8928 5284 8938 5452
rect 8938 5284 8972 5452
rect 8972 5284 8980 5452
rect 8832 5076 8842 5248
rect 8842 5076 8876 5248
rect 8876 5076 8884 5248
rect 8832 5064 8884 5076
rect 9120 5452 9172 5468
rect 9120 5284 9130 5452
rect 9130 5284 9164 5452
rect 9164 5284 9172 5452
rect 9024 5076 9034 5248
rect 9034 5076 9068 5248
rect 9068 5076 9076 5248
rect 9024 5064 9076 5076
rect 9312 5452 9364 5468
rect 9312 5284 9322 5452
rect 9322 5284 9356 5452
rect 9356 5284 9364 5452
rect 9216 5076 9226 5248
rect 9226 5076 9260 5248
rect 9260 5076 9268 5248
rect 9216 5064 9268 5076
rect 9504 5452 9556 5468
rect 9504 5284 9514 5452
rect 9514 5284 9548 5452
rect 9548 5284 9556 5452
rect 9408 5076 9418 5248
rect 9418 5076 9452 5248
rect 9452 5076 9460 5248
rect 9408 5064 9460 5076
rect 9696 5452 9748 5468
rect 9696 5284 9706 5452
rect 9706 5284 9740 5452
rect 9740 5284 9748 5452
rect 9600 5076 9610 5248
rect 9610 5076 9644 5248
rect 9644 5076 9652 5248
rect 9600 5064 9652 5076
rect 9888 5452 9940 5468
rect 9888 5284 9898 5452
rect 9898 5284 9932 5452
rect 9932 5284 9940 5452
rect 9792 5076 9802 5248
rect 9802 5076 9836 5248
rect 9836 5076 9844 5248
rect 9792 5064 9844 5076
rect 10080 5452 10132 5468
rect 10080 5284 10090 5452
rect 10090 5284 10124 5452
rect 10124 5284 10132 5452
rect 9984 5076 9994 5248
rect 9994 5076 10028 5248
rect 10028 5076 10036 5248
rect 9984 5064 10036 5076
rect 10272 5452 10324 5468
rect 10272 5284 10282 5452
rect 10282 5284 10316 5452
rect 10316 5284 10324 5452
rect 10176 5076 10186 5248
rect 10186 5076 10220 5248
rect 10220 5076 10228 5248
rect 10176 5064 10228 5076
rect 10464 5452 10516 5468
rect 10464 5284 10474 5452
rect 10474 5284 10508 5452
rect 10508 5284 10516 5452
rect 10368 5076 10378 5248
rect 10378 5076 10412 5248
rect 10412 5076 10420 5248
rect 10368 5064 10420 5076
rect 10656 5452 10708 5468
rect 10656 5284 10666 5452
rect 10666 5284 10700 5452
rect 10700 5284 10708 5452
rect 10560 5076 10570 5248
rect 10570 5076 10604 5248
rect 10604 5076 10612 5248
rect 10560 5064 10612 5076
rect 10848 5452 10900 5468
rect 10848 5284 10858 5452
rect 10858 5284 10892 5452
rect 10892 5284 10900 5452
rect 10752 5076 10762 5248
rect 10762 5076 10796 5248
rect 10796 5076 10804 5248
rect 10752 5064 10804 5076
rect 12140 5452 12192 5468
rect 12140 5284 12150 5452
rect 12150 5284 12184 5452
rect 12184 5284 12192 5452
rect 10944 5076 10954 5248
rect 10954 5076 10988 5248
rect 10988 5076 10996 5248
rect 10944 5064 10996 5076
rect 12044 5076 12054 5248
rect 12054 5076 12088 5248
rect 12088 5076 12096 5248
rect 12044 5064 12096 5076
rect 12332 5452 12384 5468
rect 12332 5284 12342 5452
rect 12342 5284 12376 5452
rect 12376 5284 12384 5452
rect 12236 5076 12246 5248
rect 12246 5076 12280 5248
rect 12280 5076 12288 5248
rect 12236 5064 12288 5076
rect 12524 5452 12576 5468
rect 12524 5284 12534 5452
rect 12534 5284 12568 5452
rect 12568 5284 12576 5452
rect 12428 5076 12438 5248
rect 12438 5076 12472 5248
rect 12472 5076 12480 5248
rect 12428 5064 12480 5076
rect 12716 5452 12768 5468
rect 12716 5284 12726 5452
rect 12726 5284 12760 5452
rect 12760 5284 12768 5452
rect 12620 5076 12630 5248
rect 12630 5076 12664 5248
rect 12664 5076 12672 5248
rect 12620 5064 12672 5076
rect 12908 5452 12960 5468
rect 12908 5284 12918 5452
rect 12918 5284 12952 5452
rect 12952 5284 12960 5452
rect 12812 5076 12822 5248
rect 12822 5076 12856 5248
rect 12856 5076 12864 5248
rect 12812 5064 12864 5076
rect 13100 5452 13152 5468
rect 13100 5284 13110 5452
rect 13110 5284 13144 5452
rect 13144 5284 13152 5452
rect 13004 5076 13014 5248
rect 13014 5076 13048 5248
rect 13048 5076 13056 5248
rect 13004 5064 13056 5076
rect 13292 5452 13344 5468
rect 13292 5284 13302 5452
rect 13302 5284 13336 5452
rect 13336 5284 13344 5452
rect 13196 5076 13206 5248
rect 13206 5076 13240 5248
rect 13240 5076 13248 5248
rect 13196 5064 13248 5076
rect 13484 5452 13536 5468
rect 13484 5284 13494 5452
rect 13494 5284 13528 5452
rect 13528 5284 13536 5452
rect 13388 5076 13398 5248
rect 13398 5076 13432 5248
rect 13432 5076 13440 5248
rect 13388 5064 13440 5076
rect 13676 5452 13728 5468
rect 13676 5284 13686 5452
rect 13686 5284 13720 5452
rect 13720 5284 13728 5452
rect 13580 5076 13590 5248
rect 13590 5076 13624 5248
rect 13624 5076 13632 5248
rect 13580 5064 13632 5076
rect 13868 5452 13920 5468
rect 13868 5284 13878 5452
rect 13878 5284 13912 5452
rect 13912 5284 13920 5452
rect 13772 5076 13782 5248
rect 13782 5076 13816 5248
rect 13816 5076 13824 5248
rect 13772 5064 13824 5076
rect 14060 5452 14112 5468
rect 14060 5284 14070 5452
rect 14070 5284 14104 5452
rect 14104 5284 14112 5452
rect 13964 5076 13974 5248
rect 13974 5076 14008 5248
rect 14008 5076 14016 5248
rect 13964 5064 14016 5076
rect 14252 5452 14304 5468
rect 14252 5284 14262 5452
rect 14262 5284 14296 5452
rect 14296 5284 14304 5452
rect 14156 5076 14166 5248
rect 14166 5076 14200 5248
rect 14200 5076 14208 5248
rect 14156 5064 14208 5076
rect 14444 5452 14496 5468
rect 14444 5284 14454 5452
rect 14454 5284 14488 5452
rect 14488 5284 14496 5452
rect 14348 5076 14358 5248
rect 14358 5076 14392 5248
rect 14392 5076 14400 5248
rect 14348 5064 14400 5076
rect 14636 5452 14688 5468
rect 14636 5284 14646 5452
rect 14646 5284 14680 5452
rect 14680 5284 14688 5452
rect 14540 5076 14550 5248
rect 14550 5076 14584 5248
rect 14584 5076 14592 5248
rect 14540 5064 14592 5076
rect 14828 5452 14880 5468
rect 14828 5284 14838 5452
rect 14838 5284 14872 5452
rect 14872 5284 14880 5452
rect 14732 5076 14742 5248
rect 14742 5076 14776 5248
rect 14776 5076 14784 5248
rect 14732 5064 14784 5076
rect 15080 5420 15540 5780
rect 14924 5076 14934 5248
rect 14934 5076 14968 5248
rect 14968 5076 14976 5248
rect 14924 5064 14976 5076
rect 15780 5452 15832 5468
rect 15780 5284 15790 5452
rect 15790 5284 15824 5452
rect 15824 5284 15832 5452
rect 15684 5076 15694 5248
rect 15694 5076 15728 5248
rect 15728 5076 15736 5248
rect 15684 5064 15736 5076
rect 15972 5452 16024 5468
rect 15972 5284 15982 5452
rect 15982 5284 16016 5452
rect 16016 5284 16024 5452
rect 15876 5076 15886 5248
rect 15886 5076 15920 5248
rect 15920 5076 15928 5248
rect 15876 5064 15928 5076
rect 16164 5452 16216 5468
rect 16164 5284 16174 5452
rect 16174 5284 16208 5452
rect 16208 5284 16216 5452
rect 16068 5076 16078 5248
rect 16078 5076 16112 5248
rect 16112 5076 16120 5248
rect 16068 5064 16120 5076
rect 16356 5452 16408 5468
rect 16356 5284 16366 5452
rect 16366 5284 16400 5452
rect 16400 5284 16408 5452
rect 16260 5076 16270 5248
rect 16270 5076 16304 5248
rect 16304 5076 16312 5248
rect 16260 5064 16312 5076
rect 16548 5452 16600 5468
rect 16548 5284 16558 5452
rect 16558 5284 16592 5452
rect 16592 5284 16600 5452
rect 16452 5076 16462 5248
rect 16462 5076 16496 5248
rect 16496 5076 16504 5248
rect 16452 5064 16504 5076
rect 16740 5452 16792 5468
rect 16740 5284 16750 5452
rect 16750 5284 16784 5452
rect 16784 5284 16792 5452
rect 16644 5076 16654 5248
rect 16654 5076 16688 5248
rect 16688 5076 16696 5248
rect 16644 5064 16696 5076
rect 16932 5452 16984 5468
rect 16932 5284 16942 5452
rect 16942 5284 16976 5452
rect 16976 5284 16984 5452
rect 16836 5076 16846 5248
rect 16846 5076 16880 5248
rect 16880 5076 16888 5248
rect 16836 5064 16888 5076
rect 17124 5452 17176 5468
rect 17124 5284 17134 5452
rect 17134 5284 17168 5452
rect 17168 5284 17176 5452
rect 17028 5076 17038 5248
rect 17038 5076 17072 5248
rect 17072 5076 17080 5248
rect 17028 5064 17080 5076
rect 17316 5452 17368 5468
rect 17316 5284 17326 5452
rect 17326 5284 17360 5452
rect 17360 5284 17368 5452
rect 17220 5076 17230 5248
rect 17230 5076 17264 5248
rect 17264 5076 17272 5248
rect 17220 5064 17272 5076
rect 17508 5452 17560 5468
rect 17508 5284 17518 5452
rect 17518 5284 17552 5452
rect 17552 5284 17560 5452
rect 17412 5076 17422 5248
rect 17422 5076 17456 5248
rect 17456 5076 17464 5248
rect 17412 5064 17464 5076
rect 17700 5452 17752 5468
rect 17700 5284 17710 5452
rect 17710 5284 17744 5452
rect 17744 5284 17752 5452
rect 17604 5076 17614 5248
rect 17614 5076 17648 5248
rect 17648 5076 17656 5248
rect 17604 5064 17656 5076
rect 17892 5452 17944 5468
rect 17892 5284 17902 5452
rect 17902 5284 17936 5452
rect 17936 5284 17944 5452
rect 17796 5076 17806 5248
rect 17806 5076 17840 5248
rect 17840 5076 17848 5248
rect 17796 5064 17848 5076
rect 18084 5452 18136 5468
rect 18084 5284 18094 5452
rect 18094 5284 18128 5452
rect 18128 5284 18136 5452
rect 17988 5076 17998 5248
rect 17998 5076 18032 5248
rect 18032 5076 18040 5248
rect 17988 5064 18040 5076
rect 18276 5452 18328 5468
rect 18276 5284 18286 5452
rect 18286 5284 18320 5452
rect 18320 5284 18328 5452
rect 18180 5076 18190 5248
rect 18190 5076 18224 5248
rect 18224 5076 18232 5248
rect 18180 5064 18232 5076
rect 18468 5452 18520 5468
rect 18468 5284 18478 5452
rect 18478 5284 18512 5452
rect 18512 5284 18520 5452
rect 18372 5076 18382 5248
rect 18382 5076 18416 5248
rect 18416 5076 18424 5248
rect 18372 5064 18424 5076
rect 18564 5076 18574 5248
rect 18574 5076 18608 5248
rect 18608 5076 18616 5248
rect 18564 5064 18616 5076
rect 1344 4816 1756 4819
rect 4520 4834 4572 4848
rect 4520 4664 4530 4834
rect 4530 4664 4564 4834
rect 4564 4664 4572 4834
rect 4424 4458 4434 4628
rect 4434 4458 4468 4628
rect 4468 4458 4476 4628
rect 4424 4444 4476 4458
rect 4712 4834 4764 4848
rect 4712 4664 4722 4834
rect 4722 4664 4756 4834
rect 4756 4664 4764 4834
rect 4616 4458 4626 4628
rect 4626 4458 4660 4628
rect 4660 4458 4668 4628
rect 4616 4444 4668 4458
rect 4904 4834 4956 4848
rect 4904 4664 4914 4834
rect 4914 4664 4948 4834
rect 4948 4664 4956 4834
rect 4808 4458 4818 4628
rect 4818 4458 4852 4628
rect 4852 4458 4860 4628
rect 4808 4444 4860 4458
rect 5096 4834 5148 4848
rect 5096 4664 5106 4834
rect 5106 4664 5140 4834
rect 5140 4664 5148 4834
rect 5000 4458 5010 4628
rect 5010 4458 5044 4628
rect 5044 4458 5052 4628
rect 5000 4444 5052 4458
rect 5288 4834 5340 4848
rect 5288 4664 5298 4834
rect 5298 4664 5332 4834
rect 5332 4664 5340 4834
rect 5192 4458 5202 4628
rect 5202 4458 5236 4628
rect 5236 4458 5244 4628
rect 5192 4444 5244 4458
rect 5480 4834 5532 4848
rect 5480 4664 5490 4834
rect 5490 4664 5524 4834
rect 5524 4664 5532 4834
rect 5384 4458 5394 4628
rect 5394 4458 5428 4628
rect 5428 4458 5436 4628
rect 5384 4444 5436 4458
rect 5672 4834 5724 4848
rect 5672 4664 5682 4834
rect 5682 4664 5716 4834
rect 5716 4664 5724 4834
rect 5576 4458 5586 4628
rect 5586 4458 5620 4628
rect 5620 4458 5628 4628
rect 5576 4444 5628 4458
rect 5864 4834 5916 4848
rect 5864 4664 5874 4834
rect 5874 4664 5908 4834
rect 5908 4664 5916 4834
rect 5768 4458 5778 4628
rect 5778 4458 5812 4628
rect 5812 4458 5820 4628
rect 5768 4444 5820 4458
rect 6056 4834 6108 4848
rect 6056 4664 6066 4834
rect 6066 4664 6100 4834
rect 6100 4664 6108 4834
rect 5960 4458 5970 4628
rect 5970 4458 6004 4628
rect 6004 4458 6012 4628
rect 5960 4444 6012 4458
rect 6248 4834 6300 4848
rect 6248 4664 6258 4834
rect 6258 4664 6292 4834
rect 6292 4664 6300 4834
rect 6152 4458 6162 4628
rect 6162 4458 6196 4628
rect 6196 4458 6204 4628
rect 6152 4444 6204 4458
rect 6440 4834 6492 4848
rect 6440 4664 6450 4834
rect 6450 4664 6484 4834
rect 6484 4664 6492 4834
rect 6344 4458 6354 4628
rect 6354 4458 6388 4628
rect 6388 4458 6396 4628
rect 6344 4444 6396 4458
rect 6632 4834 6684 4848
rect 6632 4664 6642 4834
rect 6642 4664 6676 4834
rect 6676 4664 6684 4834
rect 6536 4458 6546 4628
rect 6546 4458 6580 4628
rect 6580 4458 6588 4628
rect 6536 4444 6588 4458
rect 6824 4834 6876 4848
rect 6824 4664 6834 4834
rect 6834 4664 6868 4834
rect 6868 4664 6876 4834
rect 6728 4458 6738 4628
rect 6738 4458 6772 4628
rect 6772 4458 6780 4628
rect 6728 4444 6780 4458
rect 7016 4834 7068 4848
rect 7016 4664 7026 4834
rect 7026 4664 7060 4834
rect 7060 4664 7068 4834
rect 6920 4458 6930 4628
rect 6930 4458 6964 4628
rect 6964 4458 6972 4628
rect 6920 4444 6972 4458
rect 7208 4834 7260 4848
rect 7208 4664 7218 4834
rect 7218 4664 7252 4834
rect 7252 4664 7260 4834
rect 7112 4458 7122 4628
rect 7122 4458 7156 4628
rect 7156 4458 7164 4628
rect 7112 4444 7164 4458
rect 7304 4458 7314 4628
rect 7314 4458 7348 4628
rect 7348 4458 7356 4628
rect 7304 4444 7356 4458
rect 8160 4834 8212 4848
rect 8160 4664 8170 4834
rect 8170 4664 8204 4834
rect 8204 4664 8212 4834
rect 8064 4458 8074 4628
rect 8074 4458 8108 4628
rect 8108 4458 8116 4628
rect 8064 4444 8116 4458
rect 8352 4834 8404 4848
rect 8352 4664 8362 4834
rect 8362 4664 8396 4834
rect 8396 4664 8404 4834
rect 8256 4458 8266 4628
rect 8266 4458 8300 4628
rect 8300 4458 8308 4628
rect 8256 4444 8308 4458
rect 8544 4834 8596 4848
rect 8544 4664 8554 4834
rect 8554 4664 8588 4834
rect 8588 4664 8596 4834
rect 8448 4458 8458 4628
rect 8458 4458 8492 4628
rect 8492 4458 8500 4628
rect 8448 4444 8500 4458
rect 8736 4834 8788 4848
rect 8736 4664 8746 4834
rect 8746 4664 8780 4834
rect 8780 4664 8788 4834
rect 8640 4458 8650 4628
rect 8650 4458 8684 4628
rect 8684 4458 8692 4628
rect 8640 4444 8692 4458
rect 8928 4834 8980 4848
rect 8928 4664 8938 4834
rect 8938 4664 8972 4834
rect 8972 4664 8980 4834
rect 8832 4458 8842 4628
rect 8842 4458 8876 4628
rect 8876 4458 8884 4628
rect 8832 4444 8884 4458
rect 9120 4834 9172 4848
rect 9120 4664 9130 4834
rect 9130 4664 9164 4834
rect 9164 4664 9172 4834
rect 9024 4458 9034 4628
rect 9034 4458 9068 4628
rect 9068 4458 9076 4628
rect 9024 4444 9076 4458
rect 9312 4834 9364 4848
rect 9312 4664 9322 4834
rect 9322 4664 9356 4834
rect 9356 4664 9364 4834
rect 9216 4458 9226 4628
rect 9226 4458 9260 4628
rect 9260 4458 9268 4628
rect 9216 4444 9268 4458
rect 9504 4834 9556 4848
rect 9504 4664 9514 4834
rect 9514 4664 9548 4834
rect 9548 4664 9556 4834
rect 9408 4458 9418 4628
rect 9418 4458 9452 4628
rect 9452 4458 9460 4628
rect 9408 4444 9460 4458
rect 9696 4834 9748 4848
rect 9696 4664 9706 4834
rect 9706 4664 9740 4834
rect 9740 4664 9748 4834
rect 9600 4458 9610 4628
rect 9610 4458 9644 4628
rect 9644 4458 9652 4628
rect 9600 4444 9652 4458
rect 9888 4834 9940 4848
rect 9888 4664 9898 4834
rect 9898 4664 9932 4834
rect 9932 4664 9940 4834
rect 9792 4458 9802 4628
rect 9802 4458 9836 4628
rect 9836 4458 9844 4628
rect 9792 4444 9844 4458
rect 10080 4834 10132 4848
rect 10080 4664 10090 4834
rect 10090 4664 10124 4834
rect 10124 4664 10132 4834
rect 9984 4458 9994 4628
rect 9994 4458 10028 4628
rect 10028 4458 10036 4628
rect 9984 4444 10036 4458
rect 10272 4834 10324 4848
rect 10272 4664 10282 4834
rect 10282 4664 10316 4834
rect 10316 4664 10324 4834
rect 10176 4458 10186 4628
rect 10186 4458 10220 4628
rect 10220 4458 10228 4628
rect 10176 4444 10228 4458
rect 10464 4834 10516 4848
rect 10464 4664 10474 4834
rect 10474 4664 10508 4834
rect 10508 4664 10516 4834
rect 10368 4458 10378 4628
rect 10378 4458 10412 4628
rect 10412 4458 10420 4628
rect 10368 4444 10420 4458
rect 10656 4834 10708 4848
rect 10656 4664 10666 4834
rect 10666 4664 10700 4834
rect 10700 4664 10708 4834
rect 10560 4458 10570 4628
rect 10570 4458 10604 4628
rect 10604 4458 10612 4628
rect 10560 4444 10612 4458
rect 10848 4834 10900 4848
rect 10848 4664 10858 4834
rect 10858 4664 10892 4834
rect 10892 4664 10900 4834
rect 10752 4458 10762 4628
rect 10762 4458 10796 4628
rect 10796 4458 10804 4628
rect 10752 4444 10804 4458
rect 12140 4834 12192 4848
rect 12140 4664 12150 4834
rect 12150 4664 12184 4834
rect 12184 4664 12192 4834
rect 10944 4458 10954 4628
rect 10954 4458 10988 4628
rect 10988 4458 10996 4628
rect 10944 4444 10996 4458
rect 12044 4458 12054 4628
rect 12054 4458 12088 4628
rect 12088 4458 12096 4628
rect 12044 4444 12096 4458
rect 12332 4834 12384 4848
rect 12332 4664 12342 4834
rect 12342 4664 12376 4834
rect 12376 4664 12384 4834
rect 12236 4458 12246 4628
rect 12246 4458 12280 4628
rect 12280 4458 12288 4628
rect 12236 4444 12288 4458
rect 12524 4834 12576 4848
rect 12524 4664 12534 4834
rect 12534 4664 12568 4834
rect 12568 4664 12576 4834
rect 12428 4458 12438 4628
rect 12438 4458 12472 4628
rect 12472 4458 12480 4628
rect 12428 4444 12480 4458
rect 12716 4834 12768 4848
rect 12716 4664 12726 4834
rect 12726 4664 12760 4834
rect 12760 4664 12768 4834
rect 12620 4458 12630 4628
rect 12630 4458 12664 4628
rect 12664 4458 12672 4628
rect 12620 4444 12672 4458
rect 12908 4834 12960 4848
rect 12908 4664 12918 4834
rect 12918 4664 12952 4834
rect 12952 4664 12960 4834
rect 12812 4458 12822 4628
rect 12822 4458 12856 4628
rect 12856 4458 12864 4628
rect 12812 4444 12864 4458
rect 13100 4834 13152 4848
rect 13100 4664 13110 4834
rect 13110 4664 13144 4834
rect 13144 4664 13152 4834
rect 13004 4458 13014 4628
rect 13014 4458 13048 4628
rect 13048 4458 13056 4628
rect 13004 4444 13056 4458
rect 13292 4834 13344 4848
rect 13292 4664 13302 4834
rect 13302 4664 13336 4834
rect 13336 4664 13344 4834
rect 13196 4458 13206 4628
rect 13206 4458 13240 4628
rect 13240 4458 13248 4628
rect 13196 4444 13248 4458
rect 13484 4834 13536 4848
rect 13484 4664 13494 4834
rect 13494 4664 13528 4834
rect 13528 4664 13536 4834
rect 13388 4458 13398 4628
rect 13398 4458 13432 4628
rect 13432 4458 13440 4628
rect 13388 4444 13440 4458
rect 13676 4834 13728 4848
rect 13676 4664 13686 4834
rect 13686 4664 13720 4834
rect 13720 4664 13728 4834
rect 13580 4458 13590 4628
rect 13590 4458 13624 4628
rect 13624 4458 13632 4628
rect 13580 4444 13632 4458
rect 13868 4834 13920 4848
rect 13868 4664 13878 4834
rect 13878 4664 13912 4834
rect 13912 4664 13920 4834
rect 13772 4458 13782 4628
rect 13782 4458 13816 4628
rect 13816 4458 13824 4628
rect 13772 4444 13824 4458
rect 14060 4834 14112 4848
rect 14060 4664 14070 4834
rect 14070 4664 14104 4834
rect 14104 4664 14112 4834
rect 13964 4458 13974 4628
rect 13974 4458 14008 4628
rect 14008 4458 14016 4628
rect 13964 4444 14016 4458
rect 14252 4834 14304 4848
rect 14252 4664 14262 4834
rect 14262 4664 14296 4834
rect 14296 4664 14304 4834
rect 14156 4458 14166 4628
rect 14166 4458 14200 4628
rect 14200 4458 14208 4628
rect 14156 4444 14208 4458
rect 14444 4834 14496 4848
rect 14444 4664 14454 4834
rect 14454 4664 14488 4834
rect 14488 4664 14496 4834
rect 14348 4458 14358 4628
rect 14358 4458 14392 4628
rect 14392 4458 14400 4628
rect 14348 4444 14400 4458
rect 14636 4834 14688 4848
rect 14636 4664 14646 4834
rect 14646 4664 14680 4834
rect 14680 4664 14688 4834
rect 14540 4458 14550 4628
rect 14550 4458 14584 4628
rect 14584 4458 14592 4628
rect 14540 4444 14592 4458
rect 14828 4834 14880 4848
rect 14828 4664 14838 4834
rect 14838 4664 14872 4834
rect 14872 4664 14880 4834
rect 14732 4458 14742 4628
rect 14742 4458 14776 4628
rect 14776 4458 14784 4628
rect 14732 4444 14784 4458
rect 14924 4458 14934 4628
rect 14934 4458 14968 4628
rect 14968 4458 14976 4628
rect 14924 4444 14976 4458
rect 15780 4834 15832 4848
rect 15780 4664 15790 4834
rect 15790 4664 15824 4834
rect 15824 4664 15832 4834
rect 15684 4458 15694 4628
rect 15694 4458 15728 4628
rect 15728 4458 15736 4628
rect 15684 4444 15736 4458
rect 15972 4834 16024 4848
rect 15972 4664 15982 4834
rect 15982 4664 16016 4834
rect 16016 4664 16024 4834
rect 15876 4458 15886 4628
rect 15886 4458 15920 4628
rect 15920 4458 15928 4628
rect 15876 4444 15928 4458
rect 16164 4834 16216 4848
rect 16164 4664 16174 4834
rect 16174 4664 16208 4834
rect 16208 4664 16216 4834
rect 16068 4458 16078 4628
rect 16078 4458 16112 4628
rect 16112 4458 16120 4628
rect 16068 4444 16120 4458
rect 16356 4834 16408 4848
rect 16356 4664 16366 4834
rect 16366 4664 16400 4834
rect 16400 4664 16408 4834
rect 16260 4458 16270 4628
rect 16270 4458 16304 4628
rect 16304 4458 16312 4628
rect 16260 4444 16312 4458
rect 16548 4834 16600 4848
rect 16548 4664 16558 4834
rect 16558 4664 16592 4834
rect 16592 4664 16600 4834
rect 16452 4458 16462 4628
rect 16462 4458 16496 4628
rect 16496 4458 16504 4628
rect 16452 4444 16504 4458
rect 16740 4834 16792 4848
rect 16740 4664 16750 4834
rect 16750 4664 16784 4834
rect 16784 4664 16792 4834
rect 16644 4458 16654 4628
rect 16654 4458 16688 4628
rect 16688 4458 16696 4628
rect 16644 4444 16696 4458
rect 16932 4834 16984 4848
rect 16932 4664 16942 4834
rect 16942 4664 16976 4834
rect 16976 4664 16984 4834
rect 16836 4458 16846 4628
rect 16846 4458 16880 4628
rect 16880 4458 16888 4628
rect 16836 4444 16888 4458
rect 17124 4834 17176 4848
rect 17124 4664 17134 4834
rect 17134 4664 17168 4834
rect 17168 4664 17176 4834
rect 17028 4458 17038 4628
rect 17038 4458 17072 4628
rect 17072 4458 17080 4628
rect 17028 4444 17080 4458
rect 17316 4834 17368 4848
rect 17316 4664 17326 4834
rect 17326 4664 17360 4834
rect 17360 4664 17368 4834
rect 17220 4458 17230 4628
rect 17230 4458 17264 4628
rect 17264 4458 17272 4628
rect 17220 4444 17272 4458
rect 17508 4834 17560 4848
rect 17508 4664 17518 4834
rect 17518 4664 17552 4834
rect 17552 4664 17560 4834
rect 17412 4458 17422 4628
rect 17422 4458 17456 4628
rect 17456 4458 17464 4628
rect 17412 4444 17464 4458
rect 17700 4834 17752 4848
rect 17700 4664 17710 4834
rect 17710 4664 17744 4834
rect 17744 4664 17752 4834
rect 17604 4458 17614 4628
rect 17614 4458 17648 4628
rect 17648 4458 17656 4628
rect 17604 4444 17656 4458
rect 17892 4834 17944 4848
rect 17892 4664 17902 4834
rect 17902 4664 17936 4834
rect 17936 4664 17944 4834
rect 17796 4458 17806 4628
rect 17806 4458 17840 4628
rect 17840 4458 17848 4628
rect 17796 4444 17848 4458
rect 18084 4834 18136 4848
rect 18084 4664 18094 4834
rect 18094 4664 18128 4834
rect 18128 4664 18136 4834
rect 17988 4458 17998 4628
rect 17998 4458 18032 4628
rect 18032 4458 18040 4628
rect 17988 4444 18040 4458
rect 18276 4834 18328 4848
rect 18276 4664 18286 4834
rect 18286 4664 18320 4834
rect 18320 4664 18328 4834
rect 18180 4458 18190 4628
rect 18190 4458 18224 4628
rect 18224 4458 18232 4628
rect 18180 4444 18232 4458
rect 18468 4834 18520 4848
rect 18468 4664 18478 4834
rect 18478 4664 18512 4834
rect 18512 4664 18520 4834
rect 18372 4458 18382 4628
rect 18382 4458 18416 4628
rect 18416 4458 18424 4628
rect 18372 4444 18424 4458
rect 18564 4458 18574 4628
rect 18574 4458 18608 4628
rect 18608 4458 18616 4628
rect 18564 4444 18616 4458
rect -916 3996 -790 4372
rect -790 3996 -662 4372
rect -662 3996 -412 4372
rect -412 3996 -284 4372
rect -284 3996 -144 4372
rect 1884 3996 2010 4372
rect 2010 3996 2138 4372
rect 2138 3996 2388 4372
rect 2388 3996 2516 4372
rect 2516 3996 2656 4372
rect 4520 4216 4572 4232
rect 4520 4048 4530 4216
rect 4530 4048 4564 4216
rect 4564 4048 4572 4216
rect 4424 3840 4434 4012
rect 4434 3840 4468 4012
rect 4468 3840 4476 4012
rect 4424 3828 4476 3840
rect 4712 4216 4764 4232
rect 4712 4048 4722 4216
rect 4722 4048 4756 4216
rect 4756 4048 4764 4216
rect 4616 3840 4626 4012
rect 4626 3840 4660 4012
rect 4660 3840 4668 4012
rect 4616 3828 4668 3840
rect 4904 4216 4956 4232
rect 4904 4048 4914 4216
rect 4914 4048 4948 4216
rect 4948 4048 4956 4216
rect 4808 3840 4818 4012
rect 4818 3840 4852 4012
rect 4852 3840 4860 4012
rect 4808 3828 4860 3840
rect 5096 4216 5148 4232
rect 5096 4048 5106 4216
rect 5106 4048 5140 4216
rect 5140 4048 5148 4216
rect 5000 3840 5010 4012
rect 5010 3840 5044 4012
rect 5044 3840 5052 4012
rect 5000 3828 5052 3840
rect 5288 4216 5340 4232
rect 5288 4048 5298 4216
rect 5298 4048 5332 4216
rect 5332 4048 5340 4216
rect 5192 3840 5202 4012
rect 5202 3840 5236 4012
rect 5236 3840 5244 4012
rect 5192 3828 5244 3840
rect 5480 4216 5532 4232
rect 5480 4048 5490 4216
rect 5490 4048 5524 4216
rect 5524 4048 5532 4216
rect 5384 3840 5394 4012
rect 5394 3840 5428 4012
rect 5428 3840 5436 4012
rect 5384 3828 5436 3840
rect 5672 4216 5724 4232
rect 5672 4048 5682 4216
rect 5682 4048 5716 4216
rect 5716 4048 5724 4216
rect 5576 3840 5586 4012
rect 5586 3840 5620 4012
rect 5620 3840 5628 4012
rect 5576 3828 5628 3840
rect 5864 4216 5916 4232
rect 5864 4048 5874 4216
rect 5874 4048 5908 4216
rect 5908 4048 5916 4216
rect 5768 3840 5778 4012
rect 5778 3840 5812 4012
rect 5812 3840 5820 4012
rect 5768 3828 5820 3840
rect 6056 4216 6108 4232
rect 6056 4048 6066 4216
rect 6066 4048 6100 4216
rect 6100 4048 6108 4216
rect 5960 3840 5970 4012
rect 5970 3840 6004 4012
rect 6004 3840 6012 4012
rect 5960 3828 6012 3840
rect 6248 4216 6300 4232
rect 6248 4048 6258 4216
rect 6258 4048 6292 4216
rect 6292 4048 6300 4216
rect 6152 3840 6162 4012
rect 6162 3840 6196 4012
rect 6196 3840 6204 4012
rect 6152 3828 6204 3840
rect 6440 4216 6492 4232
rect 6440 4048 6450 4216
rect 6450 4048 6484 4216
rect 6484 4048 6492 4216
rect 6344 3840 6354 4012
rect 6354 3840 6388 4012
rect 6388 3840 6396 4012
rect 6344 3828 6396 3840
rect 6632 4216 6684 4232
rect 6632 4048 6642 4216
rect 6642 4048 6676 4216
rect 6676 4048 6684 4216
rect 6536 3840 6546 4012
rect 6546 3840 6580 4012
rect 6580 3840 6588 4012
rect 6536 3828 6588 3840
rect 6824 4216 6876 4232
rect 6824 4048 6834 4216
rect 6834 4048 6868 4216
rect 6868 4048 6876 4216
rect 6728 3840 6738 4012
rect 6738 3840 6772 4012
rect 6772 3840 6780 4012
rect 6728 3828 6780 3840
rect 7016 4216 7068 4232
rect 7016 4048 7026 4216
rect 7026 4048 7060 4216
rect 7060 4048 7068 4216
rect 6920 3840 6930 4012
rect 6930 3840 6964 4012
rect 6964 3840 6972 4012
rect 6920 3828 6972 3840
rect 7208 4216 7260 4232
rect 7208 4048 7218 4216
rect 7218 4048 7252 4216
rect 7252 4048 7260 4216
rect 7112 3840 7122 4012
rect 7122 3840 7156 4012
rect 7156 3840 7164 4012
rect 7112 3828 7164 3840
rect 7304 3840 7314 4012
rect 7314 3840 7348 4012
rect 7348 3840 7356 4012
rect 7304 3828 7356 3840
rect 8160 4216 8212 4232
rect 8160 4048 8170 4216
rect 8170 4048 8204 4216
rect 8204 4048 8212 4216
rect 8064 3840 8074 4012
rect 8074 3840 8108 4012
rect 8108 3840 8116 4012
rect 8064 3828 8116 3840
rect 8352 4216 8404 4232
rect 8352 4048 8362 4216
rect 8362 4048 8396 4216
rect 8396 4048 8404 4216
rect 8256 3840 8266 4012
rect 8266 3840 8300 4012
rect 8300 3840 8308 4012
rect 8256 3828 8308 3840
rect 8544 4216 8596 4232
rect 8544 4048 8554 4216
rect 8554 4048 8588 4216
rect 8588 4048 8596 4216
rect 8448 3840 8458 4012
rect 8458 3840 8492 4012
rect 8492 3840 8500 4012
rect 8448 3828 8500 3840
rect 8736 4216 8788 4232
rect 8736 4048 8746 4216
rect 8746 4048 8780 4216
rect 8780 4048 8788 4216
rect 8640 3840 8650 4012
rect 8650 3840 8684 4012
rect 8684 3840 8692 4012
rect 8640 3828 8692 3840
rect 8928 4216 8980 4232
rect 8928 4048 8938 4216
rect 8938 4048 8972 4216
rect 8972 4048 8980 4216
rect 8832 3840 8842 4012
rect 8842 3840 8876 4012
rect 8876 3840 8884 4012
rect 8832 3828 8884 3840
rect 9120 4216 9172 4232
rect 9120 4048 9130 4216
rect 9130 4048 9164 4216
rect 9164 4048 9172 4216
rect 9024 3840 9034 4012
rect 9034 3840 9068 4012
rect 9068 3840 9076 4012
rect 9024 3828 9076 3840
rect 9312 4216 9364 4232
rect 9312 4048 9322 4216
rect 9322 4048 9356 4216
rect 9356 4048 9364 4216
rect 9216 3840 9226 4012
rect 9226 3840 9260 4012
rect 9260 3840 9268 4012
rect 9216 3828 9268 3840
rect 9504 4216 9556 4232
rect 9504 4048 9514 4216
rect 9514 4048 9548 4216
rect 9548 4048 9556 4216
rect 9408 3840 9418 4012
rect 9418 3840 9452 4012
rect 9452 3840 9460 4012
rect 9408 3828 9460 3840
rect 9696 4216 9748 4232
rect 9696 4048 9706 4216
rect 9706 4048 9740 4216
rect 9740 4048 9748 4216
rect 9600 3840 9610 4012
rect 9610 3840 9644 4012
rect 9644 3840 9652 4012
rect 9600 3828 9652 3840
rect 9888 4216 9940 4232
rect 9888 4048 9898 4216
rect 9898 4048 9932 4216
rect 9932 4048 9940 4216
rect 9792 3840 9802 4012
rect 9802 3840 9836 4012
rect 9836 3840 9844 4012
rect 9792 3828 9844 3840
rect 10080 4216 10132 4232
rect 10080 4048 10090 4216
rect 10090 4048 10124 4216
rect 10124 4048 10132 4216
rect 9984 3840 9994 4012
rect 9994 3840 10028 4012
rect 10028 3840 10036 4012
rect 9984 3828 10036 3840
rect 10272 4216 10324 4232
rect 10272 4048 10282 4216
rect 10282 4048 10316 4216
rect 10316 4048 10324 4216
rect 10176 3840 10186 4012
rect 10186 3840 10220 4012
rect 10220 3840 10228 4012
rect 10176 3828 10228 3840
rect 10464 4216 10516 4232
rect 10464 4048 10474 4216
rect 10474 4048 10508 4216
rect 10508 4048 10516 4216
rect 10368 3840 10378 4012
rect 10378 3840 10412 4012
rect 10412 3840 10420 4012
rect 10368 3828 10420 3840
rect 10656 4216 10708 4232
rect 10656 4048 10666 4216
rect 10666 4048 10700 4216
rect 10700 4048 10708 4216
rect 10560 3840 10570 4012
rect 10570 3840 10604 4012
rect 10604 3840 10612 4012
rect 10560 3828 10612 3840
rect 10848 4216 10900 4232
rect 10848 4048 10858 4216
rect 10858 4048 10892 4216
rect 10892 4048 10900 4216
rect 10752 3840 10762 4012
rect 10762 3840 10796 4012
rect 10796 3840 10804 4012
rect 10752 3828 10804 3840
rect 12140 4216 12192 4232
rect 12140 4048 12150 4216
rect 12150 4048 12184 4216
rect 12184 4048 12192 4216
rect 10944 3840 10954 4012
rect 10954 3840 10988 4012
rect 10988 3840 10996 4012
rect 10944 3828 10996 3840
rect 12044 3840 12054 4012
rect 12054 3840 12088 4012
rect 12088 3840 12096 4012
rect 12044 3828 12096 3840
rect 12332 4216 12384 4232
rect 12332 4048 12342 4216
rect 12342 4048 12376 4216
rect 12376 4048 12384 4216
rect 12236 3840 12246 4012
rect 12246 3840 12280 4012
rect 12280 3840 12288 4012
rect 12236 3828 12288 3840
rect 12524 4216 12576 4232
rect 12524 4048 12534 4216
rect 12534 4048 12568 4216
rect 12568 4048 12576 4216
rect 12428 3840 12438 4012
rect 12438 3840 12472 4012
rect 12472 3840 12480 4012
rect 12428 3828 12480 3840
rect 12716 4216 12768 4232
rect 12716 4048 12726 4216
rect 12726 4048 12760 4216
rect 12760 4048 12768 4216
rect 12620 3840 12630 4012
rect 12630 3840 12664 4012
rect 12664 3840 12672 4012
rect 12620 3828 12672 3840
rect 12908 4216 12960 4232
rect 12908 4048 12918 4216
rect 12918 4048 12952 4216
rect 12952 4048 12960 4216
rect 12812 3840 12822 4012
rect 12822 3840 12856 4012
rect 12856 3840 12864 4012
rect 12812 3828 12864 3840
rect 13100 4216 13152 4232
rect 13100 4048 13110 4216
rect 13110 4048 13144 4216
rect 13144 4048 13152 4216
rect 13004 3840 13014 4012
rect 13014 3840 13048 4012
rect 13048 3840 13056 4012
rect 13004 3828 13056 3840
rect 13292 4216 13344 4232
rect 13292 4048 13302 4216
rect 13302 4048 13336 4216
rect 13336 4048 13344 4216
rect 13196 3840 13206 4012
rect 13206 3840 13240 4012
rect 13240 3840 13248 4012
rect 13196 3828 13248 3840
rect 13484 4216 13536 4232
rect 13484 4048 13494 4216
rect 13494 4048 13528 4216
rect 13528 4048 13536 4216
rect 13388 3840 13398 4012
rect 13398 3840 13432 4012
rect 13432 3840 13440 4012
rect 13388 3828 13440 3840
rect 13676 4216 13728 4232
rect 13676 4048 13686 4216
rect 13686 4048 13720 4216
rect 13720 4048 13728 4216
rect 13580 3840 13590 4012
rect 13590 3840 13624 4012
rect 13624 3840 13632 4012
rect 13580 3828 13632 3840
rect 13868 4216 13920 4232
rect 13868 4048 13878 4216
rect 13878 4048 13912 4216
rect 13912 4048 13920 4216
rect 13772 3840 13782 4012
rect 13782 3840 13816 4012
rect 13816 3840 13824 4012
rect 13772 3828 13824 3840
rect 14060 4216 14112 4232
rect 14060 4048 14070 4216
rect 14070 4048 14104 4216
rect 14104 4048 14112 4216
rect 13964 3840 13974 4012
rect 13974 3840 14008 4012
rect 14008 3840 14016 4012
rect 13964 3828 14016 3840
rect 14252 4216 14304 4232
rect 14252 4048 14262 4216
rect 14262 4048 14296 4216
rect 14296 4048 14304 4216
rect 14156 3840 14166 4012
rect 14166 3840 14200 4012
rect 14200 3840 14208 4012
rect 14156 3828 14208 3840
rect 14444 4216 14496 4232
rect 14444 4048 14454 4216
rect 14454 4048 14488 4216
rect 14488 4048 14496 4216
rect 14348 3840 14358 4012
rect 14358 3840 14392 4012
rect 14392 3840 14400 4012
rect 14348 3828 14400 3840
rect 14636 4216 14688 4232
rect 14636 4048 14646 4216
rect 14646 4048 14680 4216
rect 14680 4048 14688 4216
rect 14540 3840 14550 4012
rect 14550 3840 14584 4012
rect 14584 3840 14592 4012
rect 14540 3828 14592 3840
rect 14828 4216 14880 4232
rect 14828 4048 14838 4216
rect 14838 4048 14872 4216
rect 14872 4048 14880 4216
rect 14732 3840 14742 4012
rect 14742 3840 14776 4012
rect 14776 3840 14784 4012
rect 14732 3828 14784 3840
rect 14924 3840 14934 4012
rect 14934 3840 14968 4012
rect 14968 3840 14976 4012
rect 14924 3828 14976 3840
rect 15780 4216 15832 4232
rect 15780 4048 15790 4216
rect 15790 4048 15824 4216
rect 15824 4048 15832 4216
rect 15684 3840 15694 4012
rect 15694 3840 15728 4012
rect 15728 3840 15736 4012
rect 15684 3828 15736 3840
rect 15972 4216 16024 4232
rect 15972 4048 15982 4216
rect 15982 4048 16016 4216
rect 16016 4048 16024 4216
rect 15876 3840 15886 4012
rect 15886 3840 15920 4012
rect 15920 3840 15928 4012
rect 15876 3828 15928 3840
rect 16164 4216 16216 4232
rect 16164 4048 16174 4216
rect 16174 4048 16208 4216
rect 16208 4048 16216 4216
rect 16068 3840 16078 4012
rect 16078 3840 16112 4012
rect 16112 3840 16120 4012
rect 16068 3828 16120 3840
rect 16356 4216 16408 4232
rect 16356 4048 16366 4216
rect 16366 4048 16400 4216
rect 16400 4048 16408 4216
rect 16260 3840 16270 4012
rect 16270 3840 16304 4012
rect 16304 3840 16312 4012
rect 16260 3828 16312 3840
rect 16548 4216 16600 4232
rect 16548 4048 16558 4216
rect 16558 4048 16592 4216
rect 16592 4048 16600 4216
rect 16452 3840 16462 4012
rect 16462 3840 16496 4012
rect 16496 3840 16504 4012
rect 16452 3828 16504 3840
rect 16740 4216 16792 4232
rect 16740 4048 16750 4216
rect 16750 4048 16784 4216
rect 16784 4048 16792 4216
rect 16644 3840 16654 4012
rect 16654 3840 16688 4012
rect 16688 3840 16696 4012
rect 16644 3828 16696 3840
rect 16932 4216 16984 4232
rect 16932 4048 16942 4216
rect 16942 4048 16976 4216
rect 16976 4048 16984 4216
rect 16836 3840 16846 4012
rect 16846 3840 16880 4012
rect 16880 3840 16888 4012
rect 16836 3828 16888 3840
rect 17124 4216 17176 4232
rect 17124 4048 17134 4216
rect 17134 4048 17168 4216
rect 17168 4048 17176 4216
rect 17028 3840 17038 4012
rect 17038 3840 17072 4012
rect 17072 3840 17080 4012
rect 17028 3828 17080 3840
rect 17316 4216 17368 4232
rect 17316 4048 17326 4216
rect 17326 4048 17360 4216
rect 17360 4048 17368 4216
rect 17220 3840 17230 4012
rect 17230 3840 17264 4012
rect 17264 3840 17272 4012
rect 17220 3828 17272 3840
rect 17508 4216 17560 4232
rect 17508 4048 17518 4216
rect 17518 4048 17552 4216
rect 17552 4048 17560 4216
rect 17412 3840 17422 4012
rect 17422 3840 17456 4012
rect 17456 3840 17464 4012
rect 17412 3828 17464 3840
rect 17700 4216 17752 4232
rect 17700 4048 17710 4216
rect 17710 4048 17744 4216
rect 17744 4048 17752 4216
rect 17604 3840 17614 4012
rect 17614 3840 17648 4012
rect 17648 3840 17656 4012
rect 17604 3828 17656 3840
rect 17892 4216 17944 4232
rect 17892 4048 17902 4216
rect 17902 4048 17936 4216
rect 17936 4048 17944 4216
rect 17796 3840 17806 4012
rect 17806 3840 17840 4012
rect 17840 3840 17848 4012
rect 17796 3828 17848 3840
rect 18084 4216 18136 4232
rect 18084 4048 18094 4216
rect 18094 4048 18128 4216
rect 18128 4048 18136 4216
rect 17988 3840 17998 4012
rect 17998 3840 18032 4012
rect 18032 3840 18040 4012
rect 17988 3828 18040 3840
rect 18276 4216 18328 4232
rect 18276 4048 18286 4216
rect 18286 4048 18320 4216
rect 18320 4048 18328 4216
rect 18180 3840 18190 4012
rect 18190 3840 18224 4012
rect 18224 3840 18232 4012
rect 18180 3828 18232 3840
rect 18468 4216 18520 4232
rect 18468 4048 18478 4216
rect 18478 4048 18512 4216
rect 18512 4048 18520 4216
rect 18372 3840 18382 4012
rect 18382 3840 18416 4012
rect 18416 3840 18424 4012
rect 18372 3828 18424 3840
rect 18564 3840 18574 4012
rect 18574 3840 18608 4012
rect 18608 3840 18616 4012
rect 18564 3828 18616 3840
rect -944 3598 -892 3608
rect -944 3428 -934 3598
rect -934 3428 -900 3598
rect -900 3428 -892 3598
rect -1040 3222 -1030 3392
rect -1030 3222 -996 3392
rect -996 3222 -988 3392
rect -1040 3212 -988 3222
rect -752 3598 -700 3608
rect -752 3428 -742 3598
rect -742 3428 -708 3598
rect -708 3428 -700 3598
rect -848 3222 -838 3392
rect -838 3222 -804 3392
rect -804 3222 -796 3392
rect -848 3212 -796 3222
rect -560 3598 -508 3608
rect -560 3428 -550 3598
rect -550 3428 -516 3598
rect -516 3428 -508 3598
rect -656 3222 -646 3392
rect -646 3222 -612 3392
rect -612 3222 -604 3392
rect -656 3212 -604 3222
rect -368 3598 -316 3608
rect -368 3428 -358 3598
rect -358 3428 -324 3598
rect -324 3428 -316 3598
rect -464 3222 -454 3392
rect -454 3222 -420 3392
rect -420 3222 -412 3392
rect -464 3212 -412 3222
rect -176 3598 -124 3608
rect -176 3428 -166 3598
rect -166 3428 -132 3598
rect -132 3428 -124 3598
rect -272 3222 -262 3392
rect -262 3222 -228 3392
rect -228 3222 -220 3392
rect -272 3212 -220 3222
rect -80 3222 -70 3392
rect -70 3222 -36 3392
rect -36 3222 -28 3392
rect -80 3212 -28 3222
rect 1856 3598 1908 3608
rect 1856 3428 1866 3598
rect 1866 3428 1900 3598
rect 1900 3428 1908 3598
rect 1760 3222 1770 3392
rect 1770 3222 1804 3392
rect 1804 3222 1812 3392
rect 1760 3212 1812 3222
rect 2048 3598 2100 3608
rect 2048 3428 2058 3598
rect 2058 3428 2092 3598
rect 2092 3428 2100 3598
rect 1952 3222 1962 3392
rect 1962 3222 1996 3392
rect 1996 3222 2004 3392
rect 1952 3212 2004 3222
rect 2240 3598 2292 3608
rect 2240 3428 2250 3598
rect 2250 3428 2284 3598
rect 2284 3428 2292 3598
rect 2144 3222 2154 3392
rect 2154 3222 2188 3392
rect 2188 3222 2196 3392
rect 2144 3212 2196 3222
rect 2432 3598 2484 3608
rect 2432 3428 2442 3598
rect 2442 3428 2476 3598
rect 2476 3428 2484 3598
rect 2336 3222 2346 3392
rect 2346 3222 2380 3392
rect 2380 3222 2388 3392
rect 2336 3212 2388 3222
rect 2624 3598 2676 3608
rect 2624 3428 2634 3598
rect 2634 3428 2668 3598
rect 2668 3428 2676 3598
rect 2528 3222 2538 3392
rect 2538 3222 2572 3392
rect 2572 3222 2580 3392
rect 2528 3212 2580 3222
rect 2720 3222 2730 3392
rect 2730 3222 2764 3392
rect 2764 3222 2772 3392
rect 2720 3212 2772 3222
rect 4520 3598 4572 3612
rect 4520 3428 4530 3598
rect 4530 3428 4564 3598
rect 4564 3428 4572 3598
rect 4424 3222 4434 3392
rect 4434 3222 4468 3392
rect 4468 3222 4476 3392
rect 4424 3208 4476 3222
rect 4712 3598 4764 3612
rect 4712 3428 4722 3598
rect 4722 3428 4756 3598
rect 4756 3428 4764 3598
rect 4616 3222 4626 3392
rect 4626 3222 4660 3392
rect 4660 3222 4668 3392
rect 4616 3208 4668 3222
rect 4904 3598 4956 3612
rect 4904 3428 4914 3598
rect 4914 3428 4948 3598
rect 4948 3428 4956 3598
rect 4808 3222 4818 3392
rect 4818 3222 4852 3392
rect 4852 3222 4860 3392
rect 4808 3208 4860 3222
rect 5096 3598 5148 3612
rect 5096 3428 5106 3598
rect 5106 3428 5140 3598
rect 5140 3428 5148 3598
rect 5000 3222 5010 3392
rect 5010 3222 5044 3392
rect 5044 3222 5052 3392
rect 5000 3208 5052 3222
rect 5288 3598 5340 3612
rect 5288 3428 5298 3598
rect 5298 3428 5332 3598
rect 5332 3428 5340 3598
rect 5192 3222 5202 3392
rect 5202 3222 5236 3392
rect 5236 3222 5244 3392
rect 5192 3208 5244 3222
rect 5480 3598 5532 3612
rect 5480 3428 5490 3598
rect 5490 3428 5524 3598
rect 5524 3428 5532 3598
rect 5384 3222 5394 3392
rect 5394 3222 5428 3392
rect 5428 3222 5436 3392
rect 5384 3208 5436 3222
rect 5672 3598 5724 3612
rect 5672 3428 5682 3598
rect 5682 3428 5716 3598
rect 5716 3428 5724 3598
rect 5576 3222 5586 3392
rect 5586 3222 5620 3392
rect 5620 3222 5628 3392
rect 5576 3208 5628 3222
rect 5864 3598 5916 3612
rect 5864 3428 5874 3598
rect 5874 3428 5908 3598
rect 5908 3428 5916 3598
rect 5768 3222 5778 3392
rect 5778 3222 5812 3392
rect 5812 3222 5820 3392
rect 5768 3208 5820 3222
rect 6056 3598 6108 3612
rect 6056 3428 6066 3598
rect 6066 3428 6100 3598
rect 6100 3428 6108 3598
rect 5960 3222 5970 3392
rect 5970 3222 6004 3392
rect 6004 3222 6012 3392
rect 5960 3208 6012 3222
rect 6248 3598 6300 3612
rect 6248 3428 6258 3598
rect 6258 3428 6292 3598
rect 6292 3428 6300 3598
rect 6152 3222 6162 3392
rect 6162 3222 6196 3392
rect 6196 3222 6204 3392
rect 6152 3208 6204 3222
rect 6440 3598 6492 3612
rect 6440 3428 6450 3598
rect 6450 3428 6484 3598
rect 6484 3428 6492 3598
rect 6344 3222 6354 3392
rect 6354 3222 6388 3392
rect 6388 3222 6396 3392
rect 6344 3208 6396 3222
rect 6632 3598 6684 3612
rect 6632 3428 6642 3598
rect 6642 3428 6676 3598
rect 6676 3428 6684 3598
rect 6536 3222 6546 3392
rect 6546 3222 6580 3392
rect 6580 3222 6588 3392
rect 6536 3208 6588 3222
rect 6824 3598 6876 3612
rect 6824 3428 6834 3598
rect 6834 3428 6868 3598
rect 6868 3428 6876 3598
rect 6728 3222 6738 3392
rect 6738 3222 6772 3392
rect 6772 3222 6780 3392
rect 6728 3208 6780 3222
rect 7016 3598 7068 3612
rect 7016 3428 7026 3598
rect 7026 3428 7060 3598
rect 7060 3428 7068 3598
rect 6920 3222 6930 3392
rect 6930 3222 6964 3392
rect 6964 3222 6972 3392
rect 6920 3208 6972 3222
rect 7208 3598 7260 3612
rect 7208 3428 7218 3598
rect 7218 3428 7252 3598
rect 7252 3428 7260 3598
rect 7112 3222 7122 3392
rect 7122 3222 7156 3392
rect 7156 3222 7164 3392
rect 7112 3208 7164 3222
rect 7304 3222 7314 3392
rect 7314 3222 7348 3392
rect 7348 3222 7356 3392
rect 7304 3208 7356 3222
rect 8160 3598 8212 3612
rect 8160 3428 8170 3598
rect 8170 3428 8204 3598
rect 8204 3428 8212 3598
rect 8064 3222 8074 3392
rect 8074 3222 8108 3392
rect 8108 3222 8116 3392
rect 8064 3208 8116 3222
rect 8352 3598 8404 3612
rect 8352 3428 8362 3598
rect 8362 3428 8396 3598
rect 8396 3428 8404 3598
rect 8256 3222 8266 3392
rect 8266 3222 8300 3392
rect 8300 3222 8308 3392
rect 8256 3208 8308 3222
rect 8544 3598 8596 3612
rect 8544 3428 8554 3598
rect 8554 3428 8588 3598
rect 8588 3428 8596 3598
rect 8448 3222 8458 3392
rect 8458 3222 8492 3392
rect 8492 3222 8500 3392
rect 8448 3208 8500 3222
rect 8736 3598 8788 3612
rect 8736 3428 8746 3598
rect 8746 3428 8780 3598
rect 8780 3428 8788 3598
rect 8640 3222 8650 3392
rect 8650 3222 8684 3392
rect 8684 3222 8692 3392
rect 8640 3208 8692 3222
rect 8928 3598 8980 3612
rect 8928 3428 8938 3598
rect 8938 3428 8972 3598
rect 8972 3428 8980 3598
rect 8832 3222 8842 3392
rect 8842 3222 8876 3392
rect 8876 3222 8884 3392
rect 8832 3208 8884 3222
rect 9120 3598 9172 3612
rect 9120 3428 9130 3598
rect 9130 3428 9164 3598
rect 9164 3428 9172 3598
rect 9024 3222 9034 3392
rect 9034 3222 9068 3392
rect 9068 3222 9076 3392
rect 9024 3208 9076 3222
rect 9312 3598 9364 3612
rect 9312 3428 9322 3598
rect 9322 3428 9356 3598
rect 9356 3428 9364 3598
rect 9216 3222 9226 3392
rect 9226 3222 9260 3392
rect 9260 3222 9268 3392
rect 9216 3208 9268 3222
rect 9504 3598 9556 3612
rect 9504 3428 9514 3598
rect 9514 3428 9548 3598
rect 9548 3428 9556 3598
rect 9408 3222 9418 3392
rect 9418 3222 9452 3392
rect 9452 3222 9460 3392
rect 9408 3208 9460 3222
rect 9696 3598 9748 3612
rect 9696 3428 9706 3598
rect 9706 3428 9740 3598
rect 9740 3428 9748 3598
rect 9600 3222 9610 3392
rect 9610 3222 9644 3392
rect 9644 3222 9652 3392
rect 9600 3208 9652 3222
rect 9888 3598 9940 3612
rect 9888 3428 9898 3598
rect 9898 3428 9932 3598
rect 9932 3428 9940 3598
rect 9792 3222 9802 3392
rect 9802 3222 9836 3392
rect 9836 3222 9844 3392
rect 9792 3208 9844 3222
rect 10080 3598 10132 3612
rect 10080 3428 10090 3598
rect 10090 3428 10124 3598
rect 10124 3428 10132 3598
rect 9984 3222 9994 3392
rect 9994 3222 10028 3392
rect 10028 3222 10036 3392
rect 9984 3208 10036 3222
rect 10272 3598 10324 3612
rect 10272 3428 10282 3598
rect 10282 3428 10316 3598
rect 10316 3428 10324 3598
rect 10176 3222 10186 3392
rect 10186 3222 10220 3392
rect 10220 3222 10228 3392
rect 10176 3208 10228 3222
rect 10464 3598 10516 3612
rect 10464 3428 10474 3598
rect 10474 3428 10508 3598
rect 10508 3428 10516 3598
rect 10368 3222 10378 3392
rect 10378 3222 10412 3392
rect 10412 3222 10420 3392
rect 10368 3208 10420 3222
rect 10656 3598 10708 3612
rect 10656 3428 10666 3598
rect 10666 3428 10700 3598
rect 10700 3428 10708 3598
rect 10560 3222 10570 3392
rect 10570 3222 10604 3392
rect 10604 3222 10612 3392
rect 10560 3208 10612 3222
rect 10848 3598 10900 3612
rect 10848 3428 10858 3598
rect 10858 3428 10892 3598
rect 10892 3428 10900 3598
rect 10752 3222 10762 3392
rect 10762 3222 10796 3392
rect 10796 3222 10804 3392
rect 10752 3208 10804 3222
rect 12140 3598 12192 3612
rect 12140 3428 12150 3598
rect 12150 3428 12184 3598
rect 12184 3428 12192 3598
rect 10944 3222 10954 3392
rect 10954 3222 10988 3392
rect 10988 3222 10996 3392
rect 10944 3208 10996 3222
rect 12044 3222 12054 3392
rect 12054 3222 12088 3392
rect 12088 3222 12096 3392
rect 12044 3208 12096 3222
rect 12332 3598 12384 3612
rect 12332 3428 12342 3598
rect 12342 3428 12376 3598
rect 12376 3428 12384 3598
rect 12236 3222 12246 3392
rect 12246 3222 12280 3392
rect 12280 3222 12288 3392
rect 12236 3208 12288 3222
rect 12524 3598 12576 3612
rect 12524 3428 12534 3598
rect 12534 3428 12568 3598
rect 12568 3428 12576 3598
rect 12428 3222 12438 3392
rect 12438 3222 12472 3392
rect 12472 3222 12480 3392
rect 12428 3208 12480 3222
rect 12716 3598 12768 3612
rect 12716 3428 12726 3598
rect 12726 3428 12760 3598
rect 12760 3428 12768 3598
rect 12620 3222 12630 3392
rect 12630 3222 12664 3392
rect 12664 3222 12672 3392
rect 12620 3208 12672 3222
rect 12908 3598 12960 3612
rect 12908 3428 12918 3598
rect 12918 3428 12952 3598
rect 12952 3428 12960 3598
rect 12812 3222 12822 3392
rect 12822 3222 12856 3392
rect 12856 3222 12864 3392
rect 12812 3208 12864 3222
rect 13100 3598 13152 3612
rect 13100 3428 13110 3598
rect 13110 3428 13144 3598
rect 13144 3428 13152 3598
rect 13004 3222 13014 3392
rect 13014 3222 13048 3392
rect 13048 3222 13056 3392
rect 13004 3208 13056 3222
rect 13292 3598 13344 3612
rect 13292 3428 13302 3598
rect 13302 3428 13336 3598
rect 13336 3428 13344 3598
rect 13196 3222 13206 3392
rect 13206 3222 13240 3392
rect 13240 3222 13248 3392
rect 13196 3208 13248 3222
rect 13484 3598 13536 3612
rect 13484 3428 13494 3598
rect 13494 3428 13528 3598
rect 13528 3428 13536 3598
rect 13388 3222 13398 3392
rect 13398 3222 13432 3392
rect 13432 3222 13440 3392
rect 13388 3208 13440 3222
rect 13676 3598 13728 3612
rect 13676 3428 13686 3598
rect 13686 3428 13720 3598
rect 13720 3428 13728 3598
rect 13580 3222 13590 3392
rect 13590 3222 13624 3392
rect 13624 3222 13632 3392
rect 13580 3208 13632 3222
rect 13868 3598 13920 3612
rect 13868 3428 13878 3598
rect 13878 3428 13912 3598
rect 13912 3428 13920 3598
rect 13772 3222 13782 3392
rect 13782 3222 13816 3392
rect 13816 3222 13824 3392
rect 13772 3208 13824 3222
rect 14060 3598 14112 3612
rect 14060 3428 14070 3598
rect 14070 3428 14104 3598
rect 14104 3428 14112 3598
rect 13964 3222 13974 3392
rect 13974 3222 14008 3392
rect 14008 3222 14016 3392
rect 13964 3208 14016 3222
rect 14252 3598 14304 3612
rect 14252 3428 14262 3598
rect 14262 3428 14296 3598
rect 14296 3428 14304 3598
rect 14156 3222 14166 3392
rect 14166 3222 14200 3392
rect 14200 3222 14208 3392
rect 14156 3208 14208 3222
rect 14444 3598 14496 3612
rect 14444 3428 14454 3598
rect 14454 3428 14488 3598
rect 14488 3428 14496 3598
rect 14348 3222 14358 3392
rect 14358 3222 14392 3392
rect 14392 3222 14400 3392
rect 14348 3208 14400 3222
rect 14636 3598 14688 3612
rect 14636 3428 14646 3598
rect 14646 3428 14680 3598
rect 14680 3428 14688 3598
rect 14540 3222 14550 3392
rect 14550 3222 14584 3392
rect 14584 3222 14592 3392
rect 14540 3208 14592 3222
rect 14828 3598 14880 3612
rect 14828 3428 14838 3598
rect 14838 3428 14872 3598
rect 14872 3428 14880 3598
rect 14732 3222 14742 3392
rect 14742 3222 14776 3392
rect 14776 3222 14784 3392
rect 14732 3208 14784 3222
rect 14924 3222 14934 3392
rect 14934 3222 14968 3392
rect 14968 3222 14976 3392
rect 14924 3208 14976 3222
rect 15780 3598 15832 3612
rect 15780 3428 15790 3598
rect 15790 3428 15824 3598
rect 15824 3428 15832 3598
rect 15684 3222 15694 3392
rect 15694 3222 15728 3392
rect 15728 3222 15736 3392
rect 15684 3208 15736 3222
rect 15972 3598 16024 3612
rect 15972 3428 15982 3598
rect 15982 3428 16016 3598
rect 16016 3428 16024 3598
rect 15876 3222 15886 3392
rect 15886 3222 15920 3392
rect 15920 3222 15928 3392
rect 15876 3208 15928 3222
rect 16164 3598 16216 3612
rect 16164 3428 16174 3598
rect 16174 3428 16208 3598
rect 16208 3428 16216 3598
rect 16068 3222 16078 3392
rect 16078 3222 16112 3392
rect 16112 3222 16120 3392
rect 16068 3208 16120 3222
rect 16356 3598 16408 3612
rect 16356 3428 16366 3598
rect 16366 3428 16400 3598
rect 16400 3428 16408 3598
rect 16260 3222 16270 3392
rect 16270 3222 16304 3392
rect 16304 3222 16312 3392
rect 16260 3208 16312 3222
rect 16548 3598 16600 3612
rect 16548 3428 16558 3598
rect 16558 3428 16592 3598
rect 16592 3428 16600 3598
rect 16452 3222 16462 3392
rect 16462 3222 16496 3392
rect 16496 3222 16504 3392
rect 16452 3208 16504 3222
rect 16740 3598 16792 3612
rect 16740 3428 16750 3598
rect 16750 3428 16784 3598
rect 16784 3428 16792 3598
rect 16644 3222 16654 3392
rect 16654 3222 16688 3392
rect 16688 3222 16696 3392
rect 16644 3208 16696 3222
rect 16932 3598 16984 3612
rect 16932 3428 16942 3598
rect 16942 3428 16976 3598
rect 16976 3428 16984 3598
rect 16836 3222 16846 3392
rect 16846 3222 16880 3392
rect 16880 3222 16888 3392
rect 16836 3208 16888 3222
rect 17124 3598 17176 3612
rect 17124 3428 17134 3598
rect 17134 3428 17168 3598
rect 17168 3428 17176 3598
rect 17028 3222 17038 3392
rect 17038 3222 17072 3392
rect 17072 3222 17080 3392
rect 17028 3208 17080 3222
rect 17316 3598 17368 3612
rect 17316 3428 17326 3598
rect 17326 3428 17360 3598
rect 17360 3428 17368 3598
rect 17220 3222 17230 3392
rect 17230 3222 17264 3392
rect 17264 3222 17272 3392
rect 17220 3208 17272 3222
rect 17508 3598 17560 3612
rect 17508 3428 17518 3598
rect 17518 3428 17552 3598
rect 17552 3428 17560 3598
rect 17412 3222 17422 3392
rect 17422 3222 17456 3392
rect 17456 3222 17464 3392
rect 17412 3208 17464 3222
rect 17700 3598 17752 3612
rect 17700 3428 17710 3598
rect 17710 3428 17744 3598
rect 17744 3428 17752 3598
rect 17604 3222 17614 3392
rect 17614 3222 17648 3392
rect 17648 3222 17656 3392
rect 17604 3208 17656 3222
rect 17892 3598 17944 3612
rect 17892 3428 17902 3598
rect 17902 3428 17936 3598
rect 17936 3428 17944 3598
rect 17796 3222 17806 3392
rect 17806 3222 17840 3392
rect 17840 3222 17848 3392
rect 17796 3208 17848 3222
rect 18084 3598 18136 3612
rect 18084 3428 18094 3598
rect 18094 3428 18128 3598
rect 18128 3428 18136 3598
rect 17988 3222 17998 3392
rect 17998 3222 18032 3392
rect 18032 3222 18040 3392
rect 17988 3208 18040 3222
rect 18276 3598 18328 3612
rect 18276 3428 18286 3598
rect 18286 3428 18320 3598
rect 18320 3428 18328 3598
rect 18180 3222 18190 3392
rect 18190 3222 18224 3392
rect 18224 3222 18232 3392
rect 18180 3208 18232 3222
rect 18468 3598 18520 3612
rect 18468 3428 18478 3598
rect 18478 3428 18512 3598
rect 18512 3428 18520 3598
rect 18372 3222 18382 3392
rect 18382 3222 18416 3392
rect 18416 3222 18424 3392
rect 18372 3208 18424 3222
rect 18564 3222 18574 3392
rect 18574 3222 18608 3392
rect 18608 3222 18616 3392
rect 18564 3208 18616 3222
rect -1580 2620 -1528 2632
rect -1580 2452 -1570 2620
rect -1570 2452 -1536 2620
rect -1536 2452 -1528 2620
rect -1388 2620 -1336 2632
rect -1388 2452 -1378 2620
rect -1378 2452 -1344 2620
rect -1344 2452 -1336 2620
rect -1484 2244 -1474 2412
rect -1474 2244 -1440 2412
rect -1440 2244 -1432 2412
rect -1484 2232 -1432 2244
rect -1196 2620 -1144 2632
rect -1196 2452 -1186 2620
rect -1186 2452 -1152 2620
rect -1152 2452 -1144 2620
rect -1292 2244 -1282 2412
rect -1282 2244 -1248 2412
rect -1248 2244 -1240 2412
rect -1292 2232 -1240 2244
rect -1004 2620 -952 2632
rect -1004 2452 -994 2620
rect -994 2452 -960 2620
rect -960 2452 -952 2620
rect -1100 2244 -1090 2412
rect -1090 2244 -1056 2412
rect -1056 2244 -1048 2412
rect -1100 2232 -1048 2244
rect -540 2620 -488 2632
rect -540 2452 -530 2620
rect -530 2452 -496 2620
rect -496 2452 -488 2620
rect -348 2620 -296 2632
rect -348 2452 -338 2620
rect -338 2452 -304 2620
rect -304 2452 -296 2620
rect -444 2244 -434 2412
rect -434 2244 -400 2412
rect -400 2244 -392 2412
rect -444 2232 -392 2244
rect -156 2620 -104 2632
rect -156 2452 -146 2620
rect -146 2452 -112 2620
rect -112 2452 -104 2620
rect -252 2244 -242 2412
rect -242 2244 -208 2412
rect -208 2244 -200 2412
rect -252 2232 -200 2244
rect 36 2620 88 2632
rect 36 2452 46 2620
rect 46 2452 80 2620
rect 80 2452 88 2620
rect -60 2244 -50 2412
rect -50 2244 -16 2412
rect -16 2244 -8 2412
rect -60 2232 -8 2244
rect 500 2620 552 2632
rect 500 2452 510 2620
rect 510 2452 544 2620
rect 544 2452 552 2620
rect 692 2620 744 2632
rect 692 2452 702 2620
rect 702 2452 736 2620
rect 736 2452 744 2620
rect 596 2244 606 2412
rect 606 2244 640 2412
rect 640 2244 648 2412
rect 596 2232 648 2244
rect 884 2620 936 2632
rect 884 2452 894 2620
rect 894 2452 928 2620
rect 928 2452 936 2620
rect 788 2244 798 2412
rect 798 2244 832 2412
rect 832 2244 840 2412
rect 788 2232 840 2244
rect 1076 2620 1128 2632
rect 1076 2452 1086 2620
rect 1086 2452 1120 2620
rect 1120 2452 1128 2620
rect 980 2244 990 2412
rect 990 2244 1024 2412
rect 1024 2244 1032 2412
rect 980 2232 1032 2244
rect 1540 2620 1592 2632
rect 1540 2452 1550 2620
rect 1550 2452 1584 2620
rect 1584 2452 1592 2620
rect 1732 2620 1784 2632
rect 1732 2452 1742 2620
rect 1742 2452 1776 2620
rect 1776 2452 1784 2620
rect 1636 2244 1646 2412
rect 1646 2244 1680 2412
rect 1680 2244 1688 2412
rect 1636 2232 1688 2244
rect 1924 2620 1976 2632
rect 1924 2452 1934 2620
rect 1934 2452 1968 2620
rect 1968 2452 1976 2620
rect 1828 2244 1838 2412
rect 1838 2244 1872 2412
rect 1872 2244 1880 2412
rect 1828 2232 1880 2244
rect 2116 2620 2168 2632
rect 2116 2452 2126 2620
rect 2126 2452 2160 2620
rect 2160 2452 2168 2620
rect 2020 2244 2030 2412
rect 2030 2244 2064 2412
rect 2064 2244 2072 2412
rect 2020 2232 2072 2244
rect 2580 2620 2632 2632
rect 2580 2452 2590 2620
rect 2590 2452 2624 2620
rect 2624 2452 2632 2620
rect 2772 2620 2824 2632
rect 2772 2452 2782 2620
rect 2782 2452 2816 2620
rect 2816 2452 2824 2620
rect 2676 2244 2686 2412
rect 2686 2244 2720 2412
rect 2720 2244 2728 2412
rect 2676 2232 2728 2244
rect 2964 2620 3016 2632
rect 2964 2452 2974 2620
rect 2974 2452 3008 2620
rect 3008 2452 3016 2620
rect 2868 2244 2878 2412
rect 2878 2244 2912 2412
rect 2912 2244 2920 2412
rect 2868 2232 2920 2244
rect 3156 2620 3208 2632
rect 3156 2452 3166 2620
rect 3166 2452 3200 2620
rect 3200 2452 3208 2620
rect 3060 2244 3070 2412
rect 3070 2244 3104 2412
rect 3104 2244 3112 2412
rect 3060 2232 3112 2244
rect 4224 2780 4276 2792
rect 4224 2612 4234 2780
rect 4234 2612 4268 2780
rect 4268 2612 4276 2780
rect 4416 2780 4468 2792
rect 4416 2612 4426 2780
rect 4426 2612 4460 2780
rect 4460 2612 4468 2780
rect 4320 2404 4330 2572
rect 4330 2404 4364 2572
rect 4364 2404 4372 2572
rect 4320 2392 4372 2404
rect 4608 2780 4660 2792
rect 4608 2612 4618 2780
rect 4618 2612 4652 2780
rect 4652 2612 4660 2780
rect 4512 2404 4522 2572
rect 4522 2404 4556 2572
rect 4556 2404 4564 2572
rect 4512 2392 4564 2404
rect 4800 2780 4852 2792
rect 4800 2612 4810 2780
rect 4810 2612 4844 2780
rect 4844 2612 4852 2780
rect 4704 2404 4714 2572
rect 4714 2404 4748 2572
rect 4748 2404 4756 2572
rect 4704 2392 4756 2404
rect 5264 2780 5316 2792
rect 5264 2612 5274 2780
rect 5274 2612 5308 2780
rect 5308 2612 5316 2780
rect 5456 2780 5508 2792
rect 5456 2612 5466 2780
rect 5466 2612 5500 2780
rect 5500 2612 5508 2780
rect 5360 2404 5370 2572
rect 5370 2404 5404 2572
rect 5404 2404 5412 2572
rect 5360 2392 5412 2404
rect 5648 2780 5700 2792
rect 5648 2612 5658 2780
rect 5658 2612 5692 2780
rect 5692 2612 5700 2780
rect 5552 2404 5562 2572
rect 5562 2404 5596 2572
rect 5596 2404 5604 2572
rect 5552 2392 5604 2404
rect 5840 2780 5892 2792
rect 5840 2612 5850 2780
rect 5850 2612 5884 2780
rect 5884 2612 5892 2780
rect 5744 2404 5754 2572
rect 5754 2404 5788 2572
rect 5788 2404 5796 2572
rect 5744 2392 5796 2404
rect 6304 2780 6356 2792
rect 6304 2612 6314 2780
rect 6314 2612 6348 2780
rect 6348 2612 6356 2780
rect 6496 2780 6548 2792
rect 6496 2612 6506 2780
rect 6506 2612 6540 2780
rect 6540 2612 6548 2780
rect 6400 2404 6410 2572
rect 6410 2404 6444 2572
rect 6444 2404 6452 2572
rect 6400 2392 6452 2404
rect 6688 2780 6740 2792
rect 6688 2612 6698 2780
rect 6698 2612 6732 2780
rect 6732 2612 6740 2780
rect 6592 2404 6602 2572
rect 6602 2404 6636 2572
rect 6636 2404 6644 2572
rect 6592 2392 6644 2404
rect 6880 2780 6932 2792
rect 6880 2612 6890 2780
rect 6890 2612 6924 2780
rect 6924 2612 6932 2780
rect 6784 2404 6794 2572
rect 6794 2404 6828 2572
rect 6828 2404 6836 2572
rect 6784 2392 6836 2404
rect 7344 2780 7396 2792
rect 7344 2612 7354 2780
rect 7354 2612 7388 2780
rect 7388 2612 7396 2780
rect 7536 2780 7588 2792
rect 7536 2612 7546 2780
rect 7546 2612 7580 2780
rect 7580 2612 7588 2780
rect 7440 2404 7450 2572
rect 7450 2404 7484 2572
rect 7484 2404 7492 2572
rect 7440 2392 7492 2404
rect 7728 2780 7780 2792
rect 7728 2612 7738 2780
rect 7738 2612 7772 2780
rect 7772 2612 7780 2780
rect 7632 2404 7642 2572
rect 7642 2404 7676 2572
rect 7676 2404 7684 2572
rect 7632 2392 7684 2404
rect 7920 2780 7972 2792
rect 7920 2612 7930 2780
rect 7930 2612 7964 2780
rect 7964 2612 7972 2780
rect 7824 2404 7834 2572
rect 7834 2404 7868 2572
rect 7868 2404 7876 2572
rect 7824 2392 7876 2404
rect 8384 2780 8436 2792
rect 8384 2612 8394 2780
rect 8394 2612 8428 2780
rect 8428 2612 8436 2780
rect 8576 2780 8628 2792
rect 8576 2612 8586 2780
rect 8586 2612 8620 2780
rect 8620 2612 8628 2780
rect 8480 2404 8490 2572
rect 8490 2404 8524 2572
rect 8524 2404 8532 2572
rect 8480 2392 8532 2404
rect 8768 2780 8820 2792
rect 8768 2612 8778 2780
rect 8778 2612 8812 2780
rect 8812 2612 8820 2780
rect 8672 2404 8682 2572
rect 8682 2404 8716 2572
rect 8716 2404 8724 2572
rect 8672 2392 8724 2404
rect 8960 2780 9012 2792
rect 8960 2612 8970 2780
rect 8970 2612 9004 2780
rect 9004 2612 9012 2780
rect 8864 2404 8874 2572
rect 8874 2404 8908 2572
rect 8908 2404 8916 2572
rect 8864 2392 8916 2404
rect 9424 2780 9476 2792
rect 9424 2612 9434 2780
rect 9434 2612 9468 2780
rect 9468 2612 9476 2780
rect 9616 2780 9668 2792
rect 9616 2612 9626 2780
rect 9626 2612 9660 2780
rect 9660 2612 9668 2780
rect 9520 2404 9530 2572
rect 9530 2404 9564 2572
rect 9564 2404 9572 2572
rect 9520 2392 9572 2404
rect 9808 2780 9860 2792
rect 9808 2612 9818 2780
rect 9818 2612 9852 2780
rect 9852 2612 9860 2780
rect 9712 2404 9722 2572
rect 9722 2404 9756 2572
rect 9756 2404 9764 2572
rect 9712 2392 9764 2404
rect 10000 2780 10052 2792
rect 10000 2612 10010 2780
rect 10010 2612 10044 2780
rect 10044 2612 10052 2780
rect 9904 2404 9914 2572
rect 9914 2404 9948 2572
rect 9948 2404 9956 2572
rect 9904 2392 9956 2404
rect 10464 2780 10516 2792
rect 10464 2612 10474 2780
rect 10474 2612 10508 2780
rect 10508 2612 10516 2780
rect 10656 2780 10708 2792
rect 10656 2612 10666 2780
rect 10666 2612 10700 2780
rect 10700 2612 10708 2780
rect 10560 2404 10570 2572
rect 10570 2404 10604 2572
rect 10604 2404 10612 2572
rect 10560 2392 10612 2404
rect 10848 2780 10900 2792
rect 10848 2612 10858 2780
rect 10858 2612 10892 2780
rect 10892 2612 10900 2780
rect 10752 2404 10762 2572
rect 10762 2404 10796 2572
rect 10796 2404 10804 2572
rect 10752 2392 10804 2404
rect 11040 2780 11092 2792
rect 11040 2612 11050 2780
rect 11050 2612 11084 2780
rect 11084 2612 11092 2780
rect 10944 2404 10954 2572
rect 10954 2404 10988 2572
rect 10988 2404 10996 2572
rect 10944 2392 10996 2404
rect 11844 2780 11896 2792
rect 11844 2612 11854 2780
rect 11854 2612 11888 2780
rect 11888 2612 11896 2780
rect 12036 2780 12088 2792
rect 12036 2612 12046 2780
rect 12046 2612 12080 2780
rect 12080 2612 12088 2780
rect 11940 2404 11950 2572
rect 11950 2404 11984 2572
rect 11984 2404 11992 2572
rect 11940 2392 11992 2404
rect 12228 2780 12280 2792
rect 12228 2612 12238 2780
rect 12238 2612 12272 2780
rect 12272 2612 12280 2780
rect 12132 2404 12142 2572
rect 12142 2404 12176 2572
rect 12176 2404 12184 2572
rect 12132 2392 12184 2404
rect 12420 2780 12472 2792
rect 12420 2612 12430 2780
rect 12430 2612 12464 2780
rect 12464 2612 12472 2780
rect 12324 2404 12334 2572
rect 12334 2404 12368 2572
rect 12368 2404 12376 2572
rect 12324 2392 12376 2404
rect 12884 2780 12936 2792
rect 12884 2612 12894 2780
rect 12894 2612 12928 2780
rect 12928 2612 12936 2780
rect 13076 2780 13128 2792
rect 13076 2612 13086 2780
rect 13086 2612 13120 2780
rect 13120 2612 13128 2780
rect 12980 2404 12990 2572
rect 12990 2404 13024 2572
rect 13024 2404 13032 2572
rect 12980 2392 13032 2404
rect 13268 2780 13320 2792
rect 13268 2612 13278 2780
rect 13278 2612 13312 2780
rect 13312 2612 13320 2780
rect 13172 2404 13182 2572
rect 13182 2404 13216 2572
rect 13216 2404 13224 2572
rect 13172 2392 13224 2404
rect 13460 2780 13512 2792
rect 13460 2612 13470 2780
rect 13470 2612 13504 2780
rect 13504 2612 13512 2780
rect 13364 2404 13374 2572
rect 13374 2404 13408 2572
rect 13408 2404 13416 2572
rect 13364 2392 13416 2404
rect 13924 2780 13976 2792
rect 13924 2612 13934 2780
rect 13934 2612 13968 2780
rect 13968 2612 13976 2780
rect 14116 2780 14168 2792
rect 14116 2612 14126 2780
rect 14126 2612 14160 2780
rect 14160 2612 14168 2780
rect 14020 2404 14030 2572
rect 14030 2404 14064 2572
rect 14064 2404 14072 2572
rect 14020 2392 14072 2404
rect 14308 2780 14360 2792
rect 14308 2612 14318 2780
rect 14318 2612 14352 2780
rect 14352 2612 14360 2780
rect 14212 2404 14222 2572
rect 14222 2404 14256 2572
rect 14256 2404 14264 2572
rect 14212 2392 14264 2404
rect 14500 2780 14552 2792
rect 14500 2612 14510 2780
rect 14510 2612 14544 2780
rect 14544 2612 14552 2780
rect 14404 2404 14414 2572
rect 14414 2404 14448 2572
rect 14448 2404 14456 2572
rect 14404 2392 14456 2404
rect 14964 2780 15016 2792
rect 14964 2612 14974 2780
rect 14974 2612 15008 2780
rect 15008 2612 15016 2780
rect 15156 2780 15208 2792
rect 15156 2612 15166 2780
rect 15166 2612 15200 2780
rect 15200 2612 15208 2780
rect 15060 2404 15070 2572
rect 15070 2404 15104 2572
rect 15104 2404 15112 2572
rect 15060 2392 15112 2404
rect 15348 2780 15400 2792
rect 15348 2612 15358 2780
rect 15358 2612 15392 2780
rect 15392 2612 15400 2780
rect 15252 2404 15262 2572
rect 15262 2404 15296 2572
rect 15296 2404 15304 2572
rect 15252 2392 15304 2404
rect 15540 2780 15592 2792
rect 15540 2612 15550 2780
rect 15550 2612 15584 2780
rect 15584 2612 15592 2780
rect 15444 2404 15454 2572
rect 15454 2404 15488 2572
rect 15488 2404 15496 2572
rect 15444 2392 15496 2404
rect 16004 2780 16056 2792
rect 16004 2612 16014 2780
rect 16014 2612 16048 2780
rect 16048 2612 16056 2780
rect 16196 2780 16248 2792
rect 16196 2612 16206 2780
rect 16206 2612 16240 2780
rect 16240 2612 16248 2780
rect 16100 2404 16110 2572
rect 16110 2404 16144 2572
rect 16144 2404 16152 2572
rect 16100 2392 16152 2404
rect 16388 2780 16440 2792
rect 16388 2612 16398 2780
rect 16398 2612 16432 2780
rect 16432 2612 16440 2780
rect 16292 2404 16302 2572
rect 16302 2404 16336 2572
rect 16336 2404 16344 2572
rect 16292 2392 16344 2404
rect 16580 2780 16632 2792
rect 16580 2612 16590 2780
rect 16590 2612 16624 2780
rect 16624 2612 16632 2780
rect 16484 2404 16494 2572
rect 16494 2404 16528 2572
rect 16528 2404 16536 2572
rect 16484 2392 16536 2404
rect 17044 2780 17096 2792
rect 17044 2612 17054 2780
rect 17054 2612 17088 2780
rect 17088 2612 17096 2780
rect 17236 2780 17288 2792
rect 17236 2612 17246 2780
rect 17246 2612 17280 2780
rect 17280 2612 17288 2780
rect 17140 2404 17150 2572
rect 17150 2404 17184 2572
rect 17184 2404 17192 2572
rect 17140 2392 17192 2404
rect 17428 2780 17480 2792
rect 17428 2612 17438 2780
rect 17438 2612 17472 2780
rect 17472 2612 17480 2780
rect 17332 2404 17342 2572
rect 17342 2404 17376 2572
rect 17376 2404 17384 2572
rect 17332 2392 17384 2404
rect 17620 2780 17672 2792
rect 17620 2612 17630 2780
rect 17630 2612 17664 2780
rect 17664 2612 17672 2780
rect 17524 2404 17534 2572
rect 17534 2404 17568 2572
rect 17568 2404 17576 2572
rect 17524 2392 17576 2404
rect 18084 2780 18136 2792
rect 18084 2612 18094 2780
rect 18094 2612 18128 2780
rect 18128 2612 18136 2780
rect 18276 2780 18328 2792
rect 18276 2612 18286 2780
rect 18286 2612 18320 2780
rect 18320 2612 18328 2780
rect 18180 2404 18190 2572
rect 18190 2404 18224 2572
rect 18224 2404 18232 2572
rect 18180 2392 18232 2404
rect 18468 2780 18520 2792
rect 18468 2612 18478 2780
rect 18478 2612 18512 2780
rect 18512 2612 18520 2780
rect 18372 2404 18382 2572
rect 18382 2404 18416 2572
rect 18416 2404 18424 2572
rect 18372 2392 18424 2404
rect 18660 2780 18712 2792
rect 18660 2612 18670 2780
rect 18670 2612 18704 2780
rect 18704 2612 18712 2780
rect 18564 2404 18574 2572
rect 18574 2404 18608 2572
rect 18608 2404 18616 2572
rect 18564 2392 18616 2404
rect -1484 2002 -1432 2016
rect -1484 1836 -1474 2002
rect -1474 1836 -1440 2002
rect -1440 1836 -1432 2002
rect -1580 1626 -1570 1796
rect -1570 1626 -1536 1796
rect -1536 1626 -1528 1796
rect -1580 1616 -1528 1626
rect -1292 2002 -1240 2016
rect -1292 1836 -1282 2002
rect -1282 1836 -1248 2002
rect -1248 1836 -1240 2002
rect -1388 1626 -1378 1796
rect -1378 1626 -1344 1796
rect -1344 1626 -1336 1796
rect -1388 1616 -1336 1626
rect -1100 2002 -1048 2016
rect -1100 1836 -1090 2002
rect -1090 1836 -1056 2002
rect -1056 1836 -1048 2002
rect -1196 1626 -1186 1796
rect -1186 1626 -1152 1796
rect -1152 1626 -1144 1796
rect -1196 1616 -1144 1626
rect -1004 1626 -994 1796
rect -994 1626 -960 1796
rect -960 1626 -952 1796
rect -1004 1616 -952 1626
rect -444 2002 -392 2016
rect -444 1836 -434 2002
rect -434 1836 -400 2002
rect -400 1836 -392 2002
rect -540 1626 -530 1796
rect -530 1626 -496 1796
rect -496 1626 -488 1796
rect -540 1616 -488 1626
rect -252 2002 -200 2016
rect -252 1836 -242 2002
rect -242 1836 -208 2002
rect -208 1836 -200 2002
rect -348 1626 -338 1796
rect -338 1626 -304 1796
rect -304 1626 -296 1796
rect -348 1616 -296 1626
rect -60 2002 -8 2016
rect -60 1836 -50 2002
rect -50 1836 -16 2002
rect -16 1836 -8 2002
rect -156 1626 -146 1796
rect -146 1626 -112 1796
rect -112 1626 -104 1796
rect -156 1616 -104 1626
rect 36 1626 46 1796
rect 46 1626 80 1796
rect 80 1626 88 1796
rect 36 1616 88 1626
rect 596 2002 648 2016
rect 596 1836 606 2002
rect 606 1836 640 2002
rect 640 1836 648 2002
rect 500 1626 510 1796
rect 510 1626 544 1796
rect 544 1626 552 1796
rect 500 1616 552 1626
rect 788 2002 840 2016
rect 788 1836 798 2002
rect 798 1836 832 2002
rect 832 1836 840 2002
rect 692 1626 702 1796
rect 702 1626 736 1796
rect 736 1626 744 1796
rect 692 1616 744 1626
rect 980 2002 1032 2016
rect 980 1836 990 2002
rect 990 1836 1024 2002
rect 1024 1836 1032 2002
rect 884 1626 894 1796
rect 894 1626 928 1796
rect 928 1626 936 1796
rect 884 1616 936 1626
rect 1076 1626 1086 1796
rect 1086 1626 1120 1796
rect 1120 1626 1128 1796
rect 1076 1616 1128 1626
rect 1636 2002 1688 2016
rect 1636 1836 1646 2002
rect 1646 1836 1680 2002
rect 1680 1836 1688 2002
rect 1540 1626 1550 1796
rect 1550 1626 1584 1796
rect 1584 1626 1592 1796
rect 1540 1616 1592 1626
rect 1828 2002 1880 2016
rect 1828 1836 1838 2002
rect 1838 1836 1872 2002
rect 1872 1836 1880 2002
rect 1732 1626 1742 1796
rect 1742 1626 1776 1796
rect 1776 1626 1784 1796
rect 1732 1616 1784 1626
rect 2020 2002 2072 2016
rect 2020 1836 2030 2002
rect 2030 1836 2064 2002
rect 2064 1836 2072 2002
rect 1924 1626 1934 1796
rect 1934 1626 1968 1796
rect 1968 1626 1976 1796
rect 1924 1616 1976 1626
rect 2116 1626 2126 1796
rect 2126 1626 2160 1796
rect 2160 1626 2168 1796
rect 2116 1616 2168 1626
rect 2676 2002 2728 2016
rect 2676 1836 2686 2002
rect 2686 1836 2720 2002
rect 2720 1836 2728 2002
rect 2580 1626 2590 1796
rect 2590 1626 2624 1796
rect 2624 1626 2632 1796
rect 2580 1616 2632 1626
rect 2868 2002 2920 2016
rect 2868 1836 2878 2002
rect 2878 1836 2912 2002
rect 2912 1836 2920 2002
rect 2772 1626 2782 1796
rect 2782 1626 2816 1796
rect 2816 1626 2824 1796
rect 2772 1616 2824 1626
rect 3060 2002 3112 2016
rect 3060 1836 3070 2002
rect 3070 1836 3104 2002
rect 3104 1836 3112 2002
rect 2964 1626 2974 1796
rect 2974 1626 3008 1796
rect 3008 1626 3016 1796
rect 2964 1616 3016 1626
rect 3156 1626 3166 1796
rect 3166 1626 3200 1796
rect 3200 1626 3208 1796
rect 3156 1616 3208 1626
rect -1460 1198 -1408 1212
rect -1460 1032 -1452 1198
rect -1452 1032 -1418 1198
rect -1418 1032 -1408 1198
rect -1580 822 -1570 988
rect -1570 822 -1536 988
rect -1536 822 -1528 988
rect -1580 808 -1528 822
rect -1224 1198 -1172 1212
rect -1224 1032 -1216 1198
rect -1216 1032 -1182 1198
rect -1182 1032 -1172 1198
rect -1344 822 -1334 988
rect -1334 822 -1300 988
rect -1300 822 -1292 988
rect -1344 808 -1292 822
rect -988 1198 -936 1212
rect -988 1032 -980 1198
rect -980 1032 -946 1198
rect -946 1032 -936 1198
rect -1108 822 -1098 988
rect -1098 822 -1064 988
rect -1064 822 -1056 988
rect -1108 808 -1056 822
rect -872 822 -862 988
rect -862 822 -828 988
rect -828 822 -820 988
rect -872 808 -820 822
rect -420 1198 -368 1212
rect -420 1032 -412 1198
rect -412 1032 -378 1198
rect -378 1032 -368 1198
rect -540 822 -530 988
rect -530 822 -496 988
rect -496 822 -488 988
rect -540 808 -488 822
rect -184 1198 -132 1212
rect -184 1032 -176 1198
rect -176 1032 -142 1198
rect -142 1032 -132 1198
rect -304 822 -294 988
rect -294 822 -260 988
rect -260 822 -252 988
rect -304 808 -252 822
rect 52 1198 104 1212
rect 52 1032 60 1198
rect 60 1032 94 1198
rect 94 1032 104 1198
rect -68 822 -58 988
rect -58 822 -24 988
rect -24 822 -16 988
rect -68 808 -16 822
rect 168 822 178 988
rect 178 822 212 988
rect 212 822 220 988
rect 168 808 220 822
rect 620 1198 672 1212
rect 620 1032 628 1198
rect 628 1032 662 1198
rect 662 1032 672 1198
rect 500 822 510 988
rect 510 822 544 988
rect 544 822 552 988
rect 500 808 552 822
rect 856 1198 908 1212
rect 856 1032 864 1198
rect 864 1032 898 1198
rect 898 1032 908 1198
rect 736 822 746 988
rect 746 822 780 988
rect 780 822 788 988
rect 736 808 788 822
rect 1092 1198 1144 1212
rect 1092 1032 1100 1198
rect 1100 1032 1134 1198
rect 1134 1032 1144 1198
rect 972 822 982 988
rect 982 822 1016 988
rect 1016 822 1024 988
rect 972 808 1024 822
rect 1208 822 1218 988
rect 1218 822 1252 988
rect 1252 822 1260 988
rect 1208 808 1260 822
rect 1660 1198 1712 1212
rect 1660 1032 1668 1198
rect 1668 1032 1702 1198
rect 1702 1032 1712 1198
rect 1540 822 1550 988
rect 1550 822 1584 988
rect 1584 822 1592 988
rect 1540 808 1592 822
rect 1896 1198 1948 1212
rect 1896 1032 1904 1198
rect 1904 1032 1938 1198
rect 1938 1032 1948 1198
rect 1776 822 1786 988
rect 1786 822 1820 988
rect 1820 822 1828 988
rect 1776 808 1828 822
rect 2132 1198 2184 1212
rect 2132 1032 2140 1198
rect 2140 1032 2174 1198
rect 2174 1032 2184 1198
rect 2012 822 2022 988
rect 2022 822 2056 988
rect 2056 822 2064 988
rect 2012 808 2064 822
rect 2248 822 2258 988
rect 2258 822 2292 988
rect 2292 822 2300 988
rect 2248 808 2300 822
rect 2700 1198 2752 1212
rect 2700 1032 2708 1198
rect 2708 1032 2742 1198
rect 2742 1032 2752 1198
rect 2580 822 2590 988
rect 2590 822 2624 988
rect 2624 822 2632 988
rect 2580 808 2632 822
rect 2936 1198 2988 1212
rect 2936 1032 2944 1198
rect 2944 1032 2978 1198
rect 2978 1032 2988 1198
rect 2816 822 2826 988
rect 2826 822 2860 988
rect 2860 822 2868 988
rect 2816 808 2868 822
rect 3172 1198 3224 1212
rect 3172 1032 3180 1198
rect 3180 1032 3214 1198
rect 3214 1032 3224 1198
rect 3052 822 3062 988
rect 3062 822 3096 988
rect 3096 822 3104 988
rect 3052 808 3104 822
rect 3288 822 3298 988
rect 3298 822 3332 988
rect 3332 822 3340 988
rect 3288 808 3340 822
rect 4320 2162 4372 2176
rect 4320 1996 4330 2162
rect 4330 1996 4364 2162
rect 4364 1996 4372 2162
rect 4224 1786 4234 1956
rect 4234 1786 4268 1956
rect 4268 1786 4276 1956
rect 4224 1776 4276 1786
rect 4512 2162 4564 2176
rect 4512 1996 4522 2162
rect 4522 1996 4556 2162
rect 4556 1996 4564 2162
rect 4416 1786 4426 1956
rect 4426 1786 4460 1956
rect 4460 1786 4468 1956
rect 4416 1776 4468 1786
rect 4704 2162 4756 2176
rect 4704 1996 4714 2162
rect 4714 1996 4748 2162
rect 4748 1996 4756 2162
rect 4608 1786 4618 1956
rect 4618 1786 4652 1956
rect 4652 1786 4660 1956
rect 4608 1776 4660 1786
rect 4800 1786 4810 1956
rect 4810 1786 4844 1956
rect 4844 1786 4852 1956
rect 4800 1776 4852 1786
rect 5360 2162 5412 2176
rect 5360 1996 5370 2162
rect 5370 1996 5404 2162
rect 5404 1996 5412 2162
rect 5264 1786 5274 1956
rect 5274 1786 5308 1956
rect 5308 1786 5316 1956
rect 5264 1776 5316 1786
rect 5552 2162 5604 2176
rect 5552 1996 5562 2162
rect 5562 1996 5596 2162
rect 5596 1996 5604 2162
rect 5456 1786 5466 1956
rect 5466 1786 5500 1956
rect 5500 1786 5508 1956
rect 5456 1776 5508 1786
rect 5744 2162 5796 2176
rect 5744 1996 5754 2162
rect 5754 1996 5788 2162
rect 5788 1996 5796 2162
rect 5648 1786 5658 1956
rect 5658 1786 5692 1956
rect 5692 1786 5700 1956
rect 5648 1776 5700 1786
rect 5840 1786 5850 1956
rect 5850 1786 5884 1956
rect 5884 1786 5892 1956
rect 5840 1776 5892 1786
rect 6400 2162 6452 2176
rect 6400 1996 6410 2162
rect 6410 1996 6444 2162
rect 6444 1996 6452 2162
rect 6304 1786 6314 1956
rect 6314 1786 6348 1956
rect 6348 1786 6356 1956
rect 6304 1776 6356 1786
rect 6592 2162 6644 2176
rect 6592 1996 6602 2162
rect 6602 1996 6636 2162
rect 6636 1996 6644 2162
rect 6496 1786 6506 1956
rect 6506 1786 6540 1956
rect 6540 1786 6548 1956
rect 6496 1776 6548 1786
rect 6784 2162 6836 2176
rect 6784 1996 6794 2162
rect 6794 1996 6828 2162
rect 6828 1996 6836 2162
rect 6688 1786 6698 1956
rect 6698 1786 6732 1956
rect 6732 1786 6740 1956
rect 6688 1776 6740 1786
rect 6880 1786 6890 1956
rect 6890 1786 6924 1956
rect 6924 1786 6932 1956
rect 6880 1776 6932 1786
rect 7440 2162 7492 2176
rect 7440 1996 7450 2162
rect 7450 1996 7484 2162
rect 7484 1996 7492 2162
rect 7344 1786 7354 1956
rect 7354 1786 7388 1956
rect 7388 1786 7396 1956
rect 7344 1776 7396 1786
rect 7632 2162 7684 2176
rect 7632 1996 7642 2162
rect 7642 1996 7676 2162
rect 7676 1996 7684 2162
rect 7536 1786 7546 1956
rect 7546 1786 7580 1956
rect 7580 1786 7588 1956
rect 7536 1776 7588 1786
rect 7824 2162 7876 2176
rect 7824 1996 7834 2162
rect 7834 1996 7868 2162
rect 7868 1996 7876 2162
rect 7728 1786 7738 1956
rect 7738 1786 7772 1956
rect 7772 1786 7780 1956
rect 7728 1776 7780 1786
rect 7920 1786 7930 1956
rect 7930 1786 7964 1956
rect 7964 1786 7972 1956
rect 7920 1776 7972 1786
rect 8480 2162 8532 2176
rect 8480 1996 8490 2162
rect 8490 1996 8524 2162
rect 8524 1996 8532 2162
rect 8384 1786 8394 1956
rect 8394 1786 8428 1956
rect 8428 1786 8436 1956
rect 8384 1776 8436 1786
rect 8672 2162 8724 2176
rect 8672 1996 8682 2162
rect 8682 1996 8716 2162
rect 8716 1996 8724 2162
rect 8576 1786 8586 1956
rect 8586 1786 8620 1956
rect 8620 1786 8628 1956
rect 8576 1776 8628 1786
rect 8864 2162 8916 2176
rect 8864 1996 8874 2162
rect 8874 1996 8908 2162
rect 8908 1996 8916 2162
rect 8768 1786 8778 1956
rect 8778 1786 8812 1956
rect 8812 1786 8820 1956
rect 8768 1776 8820 1786
rect 8960 1786 8970 1956
rect 8970 1786 9004 1956
rect 9004 1786 9012 1956
rect 8960 1776 9012 1786
rect 9520 2162 9572 2176
rect 9520 1996 9530 2162
rect 9530 1996 9564 2162
rect 9564 1996 9572 2162
rect 9424 1786 9434 1956
rect 9434 1786 9468 1956
rect 9468 1786 9476 1956
rect 9424 1776 9476 1786
rect 9712 2162 9764 2176
rect 9712 1996 9722 2162
rect 9722 1996 9756 2162
rect 9756 1996 9764 2162
rect 9616 1786 9626 1956
rect 9626 1786 9660 1956
rect 9660 1786 9668 1956
rect 9616 1776 9668 1786
rect 9904 2162 9956 2176
rect 9904 1996 9914 2162
rect 9914 1996 9948 2162
rect 9948 1996 9956 2162
rect 9808 1786 9818 1956
rect 9818 1786 9852 1956
rect 9852 1786 9860 1956
rect 9808 1776 9860 1786
rect 10000 1786 10010 1956
rect 10010 1786 10044 1956
rect 10044 1786 10052 1956
rect 10000 1776 10052 1786
rect 10560 2162 10612 2176
rect 10560 1996 10570 2162
rect 10570 1996 10604 2162
rect 10604 1996 10612 2162
rect 10464 1786 10474 1956
rect 10474 1786 10508 1956
rect 10508 1786 10516 1956
rect 10464 1776 10516 1786
rect 10752 2162 10804 2176
rect 10752 1996 10762 2162
rect 10762 1996 10796 2162
rect 10796 1996 10804 2162
rect 10656 1786 10666 1956
rect 10666 1786 10700 1956
rect 10700 1786 10708 1956
rect 10656 1776 10708 1786
rect 10944 2162 10996 2176
rect 10944 1996 10954 2162
rect 10954 1996 10988 2162
rect 10988 1996 10996 2162
rect 10848 1786 10858 1956
rect 10858 1786 10892 1956
rect 10892 1786 10900 1956
rect 10848 1776 10900 1786
rect 11040 1786 11050 1956
rect 11050 1786 11084 1956
rect 11084 1786 11092 1956
rect 11040 1776 11092 1786
rect 4344 1358 4396 1372
rect 4344 1192 4352 1358
rect 4352 1192 4386 1358
rect 4386 1192 4396 1358
rect 4224 982 4234 1148
rect 4234 982 4268 1148
rect 4268 982 4276 1148
rect 4224 968 4276 982
rect 4580 1358 4632 1372
rect 4580 1192 4588 1358
rect 4588 1192 4622 1358
rect 4622 1192 4632 1358
rect 4460 982 4470 1148
rect 4470 982 4504 1148
rect 4504 982 4512 1148
rect 4460 968 4512 982
rect 4816 1358 4868 1372
rect 4816 1192 4824 1358
rect 4824 1192 4858 1358
rect 4858 1192 4868 1358
rect 4696 982 4706 1148
rect 4706 982 4740 1148
rect 4740 982 4748 1148
rect 4696 968 4748 982
rect 4932 982 4942 1148
rect 4942 982 4976 1148
rect 4976 982 4984 1148
rect 4932 968 4984 982
rect 5384 1358 5436 1372
rect 5384 1192 5392 1358
rect 5392 1192 5426 1358
rect 5426 1192 5436 1358
rect 5264 982 5274 1148
rect 5274 982 5308 1148
rect 5308 982 5316 1148
rect 5264 968 5316 982
rect 5620 1358 5672 1372
rect 5620 1192 5628 1358
rect 5628 1192 5662 1358
rect 5662 1192 5672 1358
rect 5500 982 5510 1148
rect 5510 982 5544 1148
rect 5544 982 5552 1148
rect 5500 968 5552 982
rect 5856 1358 5908 1372
rect 5856 1192 5864 1358
rect 5864 1192 5898 1358
rect 5898 1192 5908 1358
rect 5736 982 5746 1148
rect 5746 982 5780 1148
rect 5780 982 5788 1148
rect 5736 968 5788 982
rect 5972 982 5982 1148
rect 5982 982 6016 1148
rect 6016 982 6024 1148
rect 5972 968 6024 982
rect 6424 1358 6476 1372
rect 6424 1192 6432 1358
rect 6432 1192 6466 1358
rect 6466 1192 6476 1358
rect 6304 982 6314 1148
rect 6314 982 6348 1148
rect 6348 982 6356 1148
rect 6304 968 6356 982
rect 6660 1358 6712 1372
rect 6660 1192 6668 1358
rect 6668 1192 6702 1358
rect 6702 1192 6712 1358
rect 6540 982 6550 1148
rect 6550 982 6584 1148
rect 6584 982 6592 1148
rect 6540 968 6592 982
rect 6896 1358 6948 1372
rect 6896 1192 6904 1358
rect 6904 1192 6938 1358
rect 6938 1192 6948 1358
rect 6776 982 6786 1148
rect 6786 982 6820 1148
rect 6820 982 6828 1148
rect 6776 968 6828 982
rect 7012 982 7022 1148
rect 7022 982 7056 1148
rect 7056 982 7064 1148
rect 7012 968 7064 982
rect 7464 1358 7516 1372
rect 7464 1192 7472 1358
rect 7472 1192 7506 1358
rect 7506 1192 7516 1358
rect 7344 982 7354 1148
rect 7354 982 7388 1148
rect 7388 982 7396 1148
rect 7344 968 7396 982
rect 7700 1358 7752 1372
rect 7700 1192 7708 1358
rect 7708 1192 7742 1358
rect 7742 1192 7752 1358
rect 7580 982 7590 1148
rect 7590 982 7624 1148
rect 7624 982 7632 1148
rect 7580 968 7632 982
rect 7936 1358 7988 1372
rect 7936 1192 7944 1358
rect 7944 1192 7978 1358
rect 7978 1192 7988 1358
rect 7816 982 7826 1148
rect 7826 982 7860 1148
rect 7860 982 7868 1148
rect 7816 968 7868 982
rect 8052 982 8062 1148
rect 8062 982 8096 1148
rect 8096 982 8104 1148
rect 8052 968 8104 982
rect 8504 1358 8556 1372
rect 8504 1192 8512 1358
rect 8512 1192 8546 1358
rect 8546 1192 8556 1358
rect 8384 982 8394 1148
rect 8394 982 8428 1148
rect 8428 982 8436 1148
rect 8384 968 8436 982
rect 8740 1358 8792 1372
rect 8740 1192 8748 1358
rect 8748 1192 8782 1358
rect 8782 1192 8792 1358
rect 8620 982 8630 1148
rect 8630 982 8664 1148
rect 8664 982 8672 1148
rect 8620 968 8672 982
rect 8976 1358 9028 1372
rect 8976 1192 8984 1358
rect 8984 1192 9018 1358
rect 9018 1192 9028 1358
rect 8856 982 8866 1148
rect 8866 982 8900 1148
rect 8900 982 8908 1148
rect 8856 968 8908 982
rect 9092 982 9102 1148
rect 9102 982 9136 1148
rect 9136 982 9144 1148
rect 9092 968 9144 982
rect 9544 1358 9596 1372
rect 9544 1192 9552 1358
rect 9552 1192 9586 1358
rect 9586 1192 9596 1358
rect 9424 982 9434 1148
rect 9434 982 9468 1148
rect 9468 982 9476 1148
rect 9424 968 9476 982
rect 9780 1358 9832 1372
rect 9780 1192 9788 1358
rect 9788 1192 9822 1358
rect 9822 1192 9832 1358
rect 9660 982 9670 1148
rect 9670 982 9704 1148
rect 9704 982 9712 1148
rect 9660 968 9712 982
rect 10016 1358 10068 1372
rect 10016 1192 10024 1358
rect 10024 1192 10058 1358
rect 10058 1192 10068 1358
rect 9896 982 9906 1148
rect 9906 982 9940 1148
rect 9940 982 9948 1148
rect 9896 968 9948 982
rect 10132 982 10142 1148
rect 10142 982 10176 1148
rect 10176 982 10184 1148
rect 10132 968 10184 982
rect 10584 1358 10636 1372
rect 10584 1192 10592 1358
rect 10592 1192 10626 1358
rect 10626 1192 10636 1358
rect 10464 982 10474 1148
rect 10474 982 10508 1148
rect 10508 982 10516 1148
rect 10464 968 10516 982
rect 10820 1358 10872 1372
rect 10820 1192 10828 1358
rect 10828 1192 10862 1358
rect 10862 1192 10872 1358
rect 10700 982 10710 1148
rect 10710 982 10744 1148
rect 10744 982 10752 1148
rect 10700 968 10752 982
rect 11056 1358 11108 1372
rect 11056 1192 11064 1358
rect 11064 1192 11098 1358
rect 11098 1192 11108 1358
rect 10936 982 10946 1148
rect 10946 982 10980 1148
rect 10980 982 10988 1148
rect 10936 968 10988 982
rect 11172 982 11182 1148
rect 11182 982 11216 1148
rect 11216 982 11224 1148
rect 11172 968 11224 982
rect -1308 412 -1128 476
rect 2800 408 3068 492
rect -5998 154 -5802 406
rect -7314 -66 -7262 -54
rect -7314 -234 -7304 -66
rect -7304 -234 -7270 -66
rect -7270 -234 -7262 -66
rect -7410 -442 -7400 -274
rect -7400 -442 -7366 -274
rect -7366 -442 -7358 -274
rect -7410 -454 -7358 -442
rect -7122 -66 -7070 -54
rect -7122 -234 -7112 -66
rect -7112 -234 -7078 -66
rect -7078 -234 -7070 -66
rect -7218 -442 -7208 -274
rect -7208 -442 -7174 -274
rect -7174 -442 -7166 -274
rect -7218 -454 -7166 -442
rect -6930 -66 -6878 -54
rect -6930 -234 -6920 -66
rect -6920 -234 -6886 -66
rect -6886 -234 -6878 -66
rect -7026 -442 -7016 -274
rect -7016 -442 -6982 -274
rect -6982 -442 -6974 -274
rect -7026 -454 -6974 -442
rect -6738 -66 -6686 -54
rect -6738 -234 -6728 -66
rect -6728 -234 -6694 -66
rect -6694 -234 -6686 -66
rect -6834 -442 -6824 -274
rect -6824 -442 -6790 -274
rect -6790 -442 -6782 -274
rect -6834 -454 -6782 -442
rect -6546 -66 -6494 -54
rect -6546 -234 -6536 -66
rect -6536 -234 -6502 -66
rect -6502 -234 -6494 -66
rect -6642 -442 -6632 -274
rect -6632 -442 -6598 -274
rect -6598 -442 -6590 -274
rect -6642 -454 -6590 -442
rect -6450 -442 -6440 -274
rect -6440 -442 -6406 -274
rect -6406 -442 -6398 -274
rect -6450 -454 -6398 -442
rect -7314 -684 -7262 -670
rect -7314 -850 -7304 -684
rect -7304 -850 -7270 -684
rect -7270 -850 -7262 -684
rect -7410 -1060 -7400 -894
rect -7400 -1060 -7366 -894
rect -7366 -1060 -7358 -894
rect -7410 -1074 -7358 -1060
rect -7122 -684 -7070 -670
rect -7122 -850 -7112 -684
rect -7112 -850 -7078 -684
rect -7078 -850 -7070 -684
rect -7218 -1060 -7208 -894
rect -7208 -1060 -7174 -894
rect -7174 -1060 -7166 -894
rect -7218 -1074 -7166 -1060
rect -6930 -684 -6878 -670
rect -6930 -850 -6920 -684
rect -6920 -850 -6886 -684
rect -6886 -850 -6878 -684
rect -7026 -1060 -7016 -894
rect -7016 -1060 -6982 -894
rect -6982 -1060 -6974 -894
rect -7026 -1074 -6974 -1060
rect -6738 -684 -6686 -670
rect -6738 -850 -6728 -684
rect -6728 -850 -6694 -684
rect -6694 -850 -6686 -684
rect -6834 -1060 -6824 -894
rect -6824 -1060 -6790 -894
rect -6790 -1060 -6782 -894
rect -6834 -1074 -6782 -1060
rect -6546 -684 -6494 -670
rect -6546 -850 -6536 -684
rect -6536 -850 -6502 -684
rect -6502 -850 -6494 -684
rect -6642 -1060 -6632 -894
rect -6632 -1060 -6598 -894
rect -6598 -1060 -6590 -894
rect -6642 -1074 -6590 -1060
rect -6450 -1060 -6440 -894
rect -6440 -1060 -6406 -894
rect -6406 -1060 -6398 -894
rect -6450 -1074 -6398 -1060
rect 3712 -140 3912 76
rect 4224 540 4276 552
rect 4224 372 4234 540
rect 4234 372 4268 540
rect 4268 372 4276 540
rect 4416 540 4468 552
rect 4416 372 4426 540
rect 4426 372 4460 540
rect 4460 372 4468 540
rect 4320 164 4330 332
rect 4330 164 4364 332
rect 4364 164 4372 332
rect 4320 152 4372 164
rect 4608 540 4660 552
rect 4608 372 4618 540
rect 4618 372 4652 540
rect 4652 372 4660 540
rect 4512 164 4522 332
rect 4522 164 4556 332
rect 4556 164 4564 332
rect 4512 152 4564 164
rect 4800 540 4852 552
rect 4800 372 4810 540
rect 4810 372 4844 540
rect 4844 372 4852 540
rect 4704 164 4714 332
rect 4714 164 4748 332
rect 4748 164 4756 332
rect 4704 152 4756 164
rect 5264 540 5316 552
rect 5264 372 5274 540
rect 5274 372 5308 540
rect 5308 372 5316 540
rect 5456 540 5508 552
rect 5456 372 5466 540
rect 5466 372 5500 540
rect 5500 372 5508 540
rect 5360 164 5370 332
rect 5370 164 5404 332
rect 5404 164 5412 332
rect 5360 152 5412 164
rect 5648 540 5700 552
rect 5648 372 5658 540
rect 5658 372 5692 540
rect 5692 372 5700 540
rect 5552 164 5562 332
rect 5562 164 5596 332
rect 5596 164 5604 332
rect 5552 152 5604 164
rect 5840 540 5892 552
rect 5840 372 5850 540
rect 5850 372 5884 540
rect 5884 372 5892 540
rect 5744 164 5754 332
rect 5754 164 5788 332
rect 5788 164 5796 332
rect 5744 152 5796 164
rect 6304 540 6356 552
rect 6304 372 6314 540
rect 6314 372 6348 540
rect 6348 372 6356 540
rect 6496 540 6548 552
rect 6496 372 6506 540
rect 6506 372 6540 540
rect 6540 372 6548 540
rect 6400 164 6410 332
rect 6410 164 6444 332
rect 6444 164 6452 332
rect 6400 152 6452 164
rect 6688 540 6740 552
rect 6688 372 6698 540
rect 6698 372 6732 540
rect 6732 372 6740 540
rect 6592 164 6602 332
rect 6602 164 6636 332
rect 6636 164 6644 332
rect 6592 152 6644 164
rect 6880 540 6932 552
rect 6880 372 6890 540
rect 6890 372 6924 540
rect 6924 372 6932 540
rect 6784 164 6794 332
rect 6794 164 6828 332
rect 6828 164 6836 332
rect 6784 152 6836 164
rect 7344 540 7396 552
rect 7344 372 7354 540
rect 7354 372 7388 540
rect 7388 372 7396 540
rect 7536 540 7588 552
rect 7536 372 7546 540
rect 7546 372 7580 540
rect 7580 372 7588 540
rect 7440 164 7450 332
rect 7450 164 7484 332
rect 7484 164 7492 332
rect 7440 152 7492 164
rect 7728 540 7780 552
rect 7728 372 7738 540
rect 7738 372 7772 540
rect 7772 372 7780 540
rect 7632 164 7642 332
rect 7642 164 7676 332
rect 7676 164 7684 332
rect 7632 152 7684 164
rect 7920 540 7972 552
rect 7920 372 7930 540
rect 7930 372 7964 540
rect 7964 372 7972 540
rect 7824 164 7834 332
rect 7834 164 7868 332
rect 7868 164 7876 332
rect 7824 152 7876 164
rect 8384 540 8436 552
rect 8384 372 8394 540
rect 8394 372 8428 540
rect 8428 372 8436 540
rect 8576 540 8628 552
rect 8576 372 8586 540
rect 8586 372 8620 540
rect 8620 372 8628 540
rect 8480 164 8490 332
rect 8490 164 8524 332
rect 8524 164 8532 332
rect 8480 152 8532 164
rect 8768 540 8820 552
rect 8768 372 8778 540
rect 8778 372 8812 540
rect 8812 372 8820 540
rect 8672 164 8682 332
rect 8682 164 8716 332
rect 8716 164 8724 332
rect 8672 152 8724 164
rect 8960 540 9012 552
rect 8960 372 8970 540
rect 8970 372 9004 540
rect 9004 372 9012 540
rect 8864 164 8874 332
rect 8874 164 8908 332
rect 8908 164 8916 332
rect 8864 152 8916 164
rect 9424 540 9476 552
rect 9424 372 9434 540
rect 9434 372 9468 540
rect 9468 372 9476 540
rect 9616 540 9668 552
rect 9616 372 9626 540
rect 9626 372 9660 540
rect 9660 372 9668 540
rect 9520 164 9530 332
rect 9530 164 9564 332
rect 9564 164 9572 332
rect 9520 152 9572 164
rect 9808 540 9860 552
rect 9808 372 9818 540
rect 9818 372 9852 540
rect 9852 372 9860 540
rect 9712 164 9722 332
rect 9722 164 9756 332
rect 9756 164 9764 332
rect 9712 152 9764 164
rect 10000 540 10052 552
rect 10000 372 10010 540
rect 10010 372 10044 540
rect 10044 372 10052 540
rect 9904 164 9914 332
rect 9914 164 9948 332
rect 9948 164 9956 332
rect 9904 152 9956 164
rect 10464 540 10516 552
rect 10464 372 10474 540
rect 10474 372 10508 540
rect 10508 372 10516 540
rect 10656 540 10708 552
rect 10656 372 10666 540
rect 10666 372 10700 540
rect 10700 372 10708 540
rect 10560 164 10570 332
rect 10570 164 10604 332
rect 10604 164 10612 332
rect 10560 152 10612 164
rect 10848 540 10900 552
rect 10848 372 10858 540
rect 10858 372 10892 540
rect 10892 372 10900 540
rect 10752 164 10762 332
rect 10762 164 10796 332
rect 10796 164 10804 332
rect 10752 152 10804 164
rect 11040 540 11092 552
rect 11040 372 11050 540
rect 11050 372 11084 540
rect 11084 372 11092 540
rect 10944 164 10954 332
rect 10954 164 10988 332
rect 10988 164 10996 332
rect 10944 152 10996 164
rect -7410 -1902 -7358 -1890
rect -7410 -2070 -7400 -1902
rect -7400 -2070 -7366 -1902
rect -7366 -2070 -7358 -1902
rect -7218 -1902 -7166 -1890
rect -7218 -2070 -7208 -1902
rect -7208 -2070 -7174 -1902
rect -7174 -2070 -7166 -1902
rect -7314 -2278 -7304 -2110
rect -7304 -2278 -7270 -2110
rect -7270 -2278 -7262 -2110
rect -7314 -2290 -7262 -2278
rect -7026 -1902 -6974 -1890
rect -7026 -2070 -7016 -1902
rect -7016 -2070 -6982 -1902
rect -6982 -2070 -6974 -1902
rect -7122 -2278 -7112 -2110
rect -7112 -2278 -7078 -2110
rect -7078 -2278 -7070 -2110
rect -7122 -2290 -7070 -2278
rect -6834 -1902 -6782 -1890
rect -6834 -2070 -6824 -1902
rect -6824 -2070 -6790 -1902
rect -6790 -2070 -6782 -1902
rect -6930 -2278 -6920 -2110
rect -6920 -2278 -6886 -2110
rect -6886 -2278 -6878 -2110
rect -6930 -2290 -6878 -2278
rect 4320 -78 4372 -64
rect 4320 -244 4330 -78
rect 4330 -244 4364 -78
rect 4364 -244 4372 -78
rect 4224 -454 4234 -284
rect 4234 -454 4268 -284
rect 4268 -454 4276 -284
rect 4224 -464 4276 -454
rect 4512 -78 4564 -64
rect 4512 -244 4522 -78
rect 4522 -244 4556 -78
rect 4556 -244 4564 -78
rect 4416 -454 4426 -284
rect 4426 -454 4460 -284
rect 4460 -454 4468 -284
rect 4416 -464 4468 -454
rect 4704 -78 4756 -64
rect 4704 -244 4714 -78
rect 4714 -244 4748 -78
rect 4748 -244 4756 -78
rect 4608 -454 4618 -284
rect 4618 -454 4652 -284
rect 4652 -454 4660 -284
rect 4608 -464 4660 -454
rect 4800 -454 4810 -284
rect 4810 -454 4844 -284
rect 4844 -454 4852 -284
rect 4800 -464 4852 -454
rect 5360 -78 5412 -64
rect 5360 -244 5370 -78
rect 5370 -244 5404 -78
rect 5404 -244 5412 -78
rect 5264 -454 5274 -284
rect 5274 -454 5308 -284
rect 5308 -454 5316 -284
rect 5264 -464 5316 -454
rect 5552 -78 5604 -64
rect 5552 -244 5562 -78
rect 5562 -244 5596 -78
rect 5596 -244 5604 -78
rect 5456 -454 5466 -284
rect 5466 -454 5500 -284
rect 5500 -454 5508 -284
rect 5456 -464 5508 -454
rect 5744 -78 5796 -64
rect 5744 -244 5754 -78
rect 5754 -244 5788 -78
rect 5788 -244 5796 -78
rect 5648 -454 5658 -284
rect 5658 -454 5692 -284
rect 5692 -454 5700 -284
rect 5648 -464 5700 -454
rect 5840 -454 5850 -284
rect 5850 -454 5884 -284
rect 5884 -454 5892 -284
rect 5840 -464 5892 -454
rect 6400 -78 6452 -64
rect 6400 -244 6410 -78
rect 6410 -244 6444 -78
rect 6444 -244 6452 -78
rect 6304 -454 6314 -284
rect 6314 -454 6348 -284
rect 6348 -454 6356 -284
rect 6304 -464 6356 -454
rect 6592 -78 6644 -64
rect 6592 -244 6602 -78
rect 6602 -244 6636 -78
rect 6636 -244 6644 -78
rect 6496 -454 6506 -284
rect 6506 -454 6540 -284
rect 6540 -454 6548 -284
rect 6496 -464 6548 -454
rect 6784 -78 6836 -64
rect 6784 -244 6794 -78
rect 6794 -244 6828 -78
rect 6828 -244 6836 -78
rect 6688 -454 6698 -284
rect 6698 -454 6732 -284
rect 6732 -454 6740 -284
rect 6688 -464 6740 -454
rect 6880 -454 6890 -284
rect 6890 -454 6924 -284
rect 6924 -454 6932 -284
rect 6880 -464 6932 -454
rect 7440 -78 7492 -64
rect 7440 -244 7450 -78
rect 7450 -244 7484 -78
rect 7484 -244 7492 -78
rect 7344 -454 7354 -284
rect 7354 -454 7388 -284
rect 7388 -454 7396 -284
rect 7344 -464 7396 -454
rect 7632 -78 7684 -64
rect 7632 -244 7642 -78
rect 7642 -244 7676 -78
rect 7676 -244 7684 -78
rect 7536 -454 7546 -284
rect 7546 -454 7580 -284
rect 7580 -454 7588 -284
rect 7536 -464 7588 -454
rect 7824 -78 7876 -64
rect 7824 -244 7834 -78
rect 7834 -244 7868 -78
rect 7868 -244 7876 -78
rect 7728 -454 7738 -284
rect 7738 -454 7772 -284
rect 7772 -454 7780 -284
rect 7728 -464 7780 -454
rect 7920 -454 7930 -284
rect 7930 -454 7964 -284
rect 7964 -454 7972 -284
rect 7920 -464 7972 -454
rect 8480 -78 8532 -64
rect 8480 -244 8490 -78
rect 8490 -244 8524 -78
rect 8524 -244 8532 -78
rect 8384 -454 8394 -284
rect 8394 -454 8428 -284
rect 8428 -454 8436 -284
rect 8384 -464 8436 -454
rect 8672 -78 8724 -64
rect 8672 -244 8682 -78
rect 8682 -244 8716 -78
rect 8716 -244 8724 -78
rect 8576 -454 8586 -284
rect 8586 -454 8620 -284
rect 8620 -454 8628 -284
rect 8576 -464 8628 -454
rect 8864 -78 8916 -64
rect 8864 -244 8874 -78
rect 8874 -244 8908 -78
rect 8908 -244 8916 -78
rect 8768 -454 8778 -284
rect 8778 -454 8812 -284
rect 8812 -454 8820 -284
rect 8768 -464 8820 -454
rect 8960 -454 8970 -284
rect 8970 -454 9004 -284
rect 9004 -454 9012 -284
rect 8960 -464 9012 -454
rect 9520 -78 9572 -64
rect 9520 -244 9530 -78
rect 9530 -244 9564 -78
rect 9564 -244 9572 -78
rect 9424 -454 9434 -284
rect 9434 -454 9468 -284
rect 9468 -454 9476 -284
rect 9424 -464 9476 -454
rect 9712 -78 9764 -64
rect 9712 -244 9722 -78
rect 9722 -244 9756 -78
rect 9756 -244 9764 -78
rect 9616 -454 9626 -284
rect 9626 -454 9660 -284
rect 9660 -454 9668 -284
rect 9616 -464 9668 -454
rect 9904 -78 9956 -64
rect 9904 -244 9914 -78
rect 9914 -244 9948 -78
rect 9948 -244 9956 -78
rect 9808 -454 9818 -284
rect 9818 -454 9852 -284
rect 9852 -454 9860 -284
rect 9808 -464 9860 -454
rect 10000 -454 10010 -284
rect 10010 -454 10044 -284
rect 10044 -454 10052 -284
rect 10000 -464 10052 -454
rect 10560 -78 10612 -64
rect 10560 -244 10570 -78
rect 10570 -244 10604 -78
rect 10604 -244 10612 -78
rect 10464 -454 10474 -284
rect 10474 -454 10508 -284
rect 10508 -454 10516 -284
rect 10464 -464 10516 -454
rect 10752 -78 10804 -64
rect 10752 -244 10762 -78
rect 10762 -244 10796 -78
rect 10796 -244 10804 -78
rect 10656 -454 10666 -284
rect 10666 -454 10700 -284
rect 10700 -454 10708 -284
rect 10656 -464 10708 -454
rect 10944 -78 10996 -64
rect 10944 -244 10954 -78
rect 10954 -244 10988 -78
rect 10988 -244 10996 -78
rect 10848 -454 10858 -284
rect 10858 -454 10892 -284
rect 10892 -454 10900 -284
rect 10848 -464 10900 -454
rect 11040 -454 11050 -284
rect 11050 -454 11084 -284
rect 11084 -454 11092 -284
rect 11040 -464 11092 -454
rect 11940 2162 11992 2176
rect 11940 1996 11950 2162
rect 11950 1996 11984 2162
rect 11984 1996 11992 2162
rect 11844 1786 11854 1956
rect 11854 1786 11888 1956
rect 11888 1786 11896 1956
rect 11844 1776 11896 1786
rect 12132 2162 12184 2176
rect 12132 1996 12142 2162
rect 12142 1996 12176 2162
rect 12176 1996 12184 2162
rect 12036 1786 12046 1956
rect 12046 1786 12080 1956
rect 12080 1786 12088 1956
rect 12036 1776 12088 1786
rect 12324 2162 12376 2176
rect 12324 1996 12334 2162
rect 12334 1996 12368 2162
rect 12368 1996 12376 2162
rect 12228 1786 12238 1956
rect 12238 1786 12272 1956
rect 12272 1786 12280 1956
rect 12228 1776 12280 1786
rect 12420 1786 12430 1956
rect 12430 1786 12464 1956
rect 12464 1786 12472 1956
rect 12420 1776 12472 1786
rect 12980 2162 13032 2176
rect 12980 1996 12990 2162
rect 12990 1996 13024 2162
rect 13024 1996 13032 2162
rect 12884 1786 12894 1956
rect 12894 1786 12928 1956
rect 12928 1786 12936 1956
rect 12884 1776 12936 1786
rect 13172 2162 13224 2176
rect 13172 1996 13182 2162
rect 13182 1996 13216 2162
rect 13216 1996 13224 2162
rect 13076 1786 13086 1956
rect 13086 1786 13120 1956
rect 13120 1786 13128 1956
rect 13076 1776 13128 1786
rect 13364 2162 13416 2176
rect 13364 1996 13374 2162
rect 13374 1996 13408 2162
rect 13408 1996 13416 2162
rect 13268 1786 13278 1956
rect 13278 1786 13312 1956
rect 13312 1786 13320 1956
rect 13268 1776 13320 1786
rect 13460 1786 13470 1956
rect 13470 1786 13504 1956
rect 13504 1786 13512 1956
rect 13460 1776 13512 1786
rect 14020 2162 14072 2176
rect 14020 1996 14030 2162
rect 14030 1996 14064 2162
rect 14064 1996 14072 2162
rect 13924 1786 13934 1956
rect 13934 1786 13968 1956
rect 13968 1786 13976 1956
rect 13924 1776 13976 1786
rect 14212 2162 14264 2176
rect 14212 1996 14222 2162
rect 14222 1996 14256 2162
rect 14256 1996 14264 2162
rect 14116 1786 14126 1956
rect 14126 1786 14160 1956
rect 14160 1786 14168 1956
rect 14116 1776 14168 1786
rect 14404 2162 14456 2176
rect 14404 1996 14414 2162
rect 14414 1996 14448 2162
rect 14448 1996 14456 2162
rect 14308 1786 14318 1956
rect 14318 1786 14352 1956
rect 14352 1786 14360 1956
rect 14308 1776 14360 1786
rect 14500 1786 14510 1956
rect 14510 1786 14544 1956
rect 14544 1786 14552 1956
rect 14500 1776 14552 1786
rect 15060 2162 15112 2176
rect 15060 1996 15070 2162
rect 15070 1996 15104 2162
rect 15104 1996 15112 2162
rect 14964 1786 14974 1956
rect 14974 1786 15008 1956
rect 15008 1786 15016 1956
rect 14964 1776 15016 1786
rect 15252 2162 15304 2176
rect 15252 1996 15262 2162
rect 15262 1996 15296 2162
rect 15296 1996 15304 2162
rect 15156 1786 15166 1956
rect 15166 1786 15200 1956
rect 15200 1786 15208 1956
rect 15156 1776 15208 1786
rect 15444 2162 15496 2176
rect 15444 1996 15454 2162
rect 15454 1996 15488 2162
rect 15488 1996 15496 2162
rect 15348 1786 15358 1956
rect 15358 1786 15392 1956
rect 15392 1786 15400 1956
rect 15348 1776 15400 1786
rect 15540 1786 15550 1956
rect 15550 1786 15584 1956
rect 15584 1786 15592 1956
rect 15540 1776 15592 1786
rect 16100 2162 16152 2176
rect 16100 1996 16110 2162
rect 16110 1996 16144 2162
rect 16144 1996 16152 2162
rect 16004 1786 16014 1956
rect 16014 1786 16048 1956
rect 16048 1786 16056 1956
rect 16004 1776 16056 1786
rect 16292 2162 16344 2176
rect 16292 1996 16302 2162
rect 16302 1996 16336 2162
rect 16336 1996 16344 2162
rect 16196 1786 16206 1956
rect 16206 1786 16240 1956
rect 16240 1786 16248 1956
rect 16196 1776 16248 1786
rect 16484 2162 16536 2176
rect 16484 1996 16494 2162
rect 16494 1996 16528 2162
rect 16528 1996 16536 2162
rect 16388 1786 16398 1956
rect 16398 1786 16432 1956
rect 16432 1786 16440 1956
rect 16388 1776 16440 1786
rect 16580 1786 16590 1956
rect 16590 1786 16624 1956
rect 16624 1786 16632 1956
rect 16580 1776 16632 1786
rect 17140 2162 17192 2176
rect 17140 1996 17150 2162
rect 17150 1996 17184 2162
rect 17184 1996 17192 2162
rect 17044 1786 17054 1956
rect 17054 1786 17088 1956
rect 17088 1786 17096 1956
rect 17044 1776 17096 1786
rect 17332 2162 17384 2176
rect 17332 1996 17342 2162
rect 17342 1996 17376 2162
rect 17376 1996 17384 2162
rect 17236 1786 17246 1956
rect 17246 1786 17280 1956
rect 17280 1786 17288 1956
rect 17236 1776 17288 1786
rect 17524 2162 17576 2176
rect 17524 1996 17534 2162
rect 17534 1996 17568 2162
rect 17568 1996 17576 2162
rect 17428 1786 17438 1956
rect 17438 1786 17472 1956
rect 17472 1786 17480 1956
rect 17428 1776 17480 1786
rect 17620 1786 17630 1956
rect 17630 1786 17664 1956
rect 17664 1786 17672 1956
rect 17620 1776 17672 1786
rect 18180 2162 18232 2176
rect 18180 1996 18190 2162
rect 18190 1996 18224 2162
rect 18224 1996 18232 2162
rect 18084 1786 18094 1956
rect 18094 1786 18128 1956
rect 18128 1786 18136 1956
rect 18084 1776 18136 1786
rect 18372 2162 18424 2176
rect 18372 1996 18382 2162
rect 18382 1996 18416 2162
rect 18416 1996 18424 2162
rect 18276 1786 18286 1956
rect 18286 1786 18320 1956
rect 18320 1786 18328 1956
rect 18276 1776 18328 1786
rect 18564 2162 18616 2176
rect 18564 1996 18574 2162
rect 18574 1996 18608 2162
rect 18608 1996 18616 2162
rect 18468 1786 18478 1956
rect 18478 1786 18512 1956
rect 18512 1786 18520 1956
rect 18468 1776 18520 1786
rect 18660 1786 18670 1956
rect 18670 1786 18704 1956
rect 18704 1786 18712 1956
rect 18660 1776 18712 1786
rect 11964 1358 12016 1372
rect 11964 1192 11972 1358
rect 11972 1192 12006 1358
rect 12006 1192 12016 1358
rect 11844 982 11854 1148
rect 11854 982 11888 1148
rect 11888 982 11896 1148
rect 11844 968 11896 982
rect 12200 1358 12252 1372
rect 12200 1192 12208 1358
rect 12208 1192 12242 1358
rect 12242 1192 12252 1358
rect 12080 982 12090 1148
rect 12090 982 12124 1148
rect 12124 982 12132 1148
rect 12080 968 12132 982
rect 12436 1358 12488 1372
rect 12436 1192 12444 1358
rect 12444 1192 12478 1358
rect 12478 1192 12488 1358
rect 12316 982 12326 1148
rect 12326 982 12360 1148
rect 12360 982 12368 1148
rect 12316 968 12368 982
rect 12552 982 12562 1148
rect 12562 982 12596 1148
rect 12596 982 12604 1148
rect 12552 968 12604 982
rect 13004 1358 13056 1372
rect 13004 1192 13012 1358
rect 13012 1192 13046 1358
rect 13046 1192 13056 1358
rect 12884 982 12894 1148
rect 12894 982 12928 1148
rect 12928 982 12936 1148
rect 12884 968 12936 982
rect 13240 1358 13292 1372
rect 13240 1192 13248 1358
rect 13248 1192 13282 1358
rect 13282 1192 13292 1358
rect 13120 982 13130 1148
rect 13130 982 13164 1148
rect 13164 982 13172 1148
rect 13120 968 13172 982
rect 13476 1358 13528 1372
rect 13476 1192 13484 1358
rect 13484 1192 13518 1358
rect 13518 1192 13528 1358
rect 13356 982 13366 1148
rect 13366 982 13400 1148
rect 13400 982 13408 1148
rect 13356 968 13408 982
rect 13592 982 13602 1148
rect 13602 982 13636 1148
rect 13636 982 13644 1148
rect 13592 968 13644 982
rect 14044 1358 14096 1372
rect 14044 1192 14052 1358
rect 14052 1192 14086 1358
rect 14086 1192 14096 1358
rect 13924 982 13934 1148
rect 13934 982 13968 1148
rect 13968 982 13976 1148
rect 13924 968 13976 982
rect 14280 1358 14332 1372
rect 14280 1192 14288 1358
rect 14288 1192 14322 1358
rect 14322 1192 14332 1358
rect 14160 982 14170 1148
rect 14170 982 14204 1148
rect 14204 982 14212 1148
rect 14160 968 14212 982
rect 14516 1358 14568 1372
rect 14516 1192 14524 1358
rect 14524 1192 14558 1358
rect 14558 1192 14568 1358
rect 14396 982 14406 1148
rect 14406 982 14440 1148
rect 14440 982 14448 1148
rect 14396 968 14448 982
rect 14632 982 14642 1148
rect 14642 982 14676 1148
rect 14676 982 14684 1148
rect 14632 968 14684 982
rect 15084 1358 15136 1372
rect 15084 1192 15092 1358
rect 15092 1192 15126 1358
rect 15126 1192 15136 1358
rect 14964 982 14974 1148
rect 14974 982 15008 1148
rect 15008 982 15016 1148
rect 14964 968 15016 982
rect 15320 1358 15372 1372
rect 15320 1192 15328 1358
rect 15328 1192 15362 1358
rect 15362 1192 15372 1358
rect 15200 982 15210 1148
rect 15210 982 15244 1148
rect 15244 982 15252 1148
rect 15200 968 15252 982
rect 15556 1358 15608 1372
rect 15556 1192 15564 1358
rect 15564 1192 15598 1358
rect 15598 1192 15608 1358
rect 15436 982 15446 1148
rect 15446 982 15480 1148
rect 15480 982 15488 1148
rect 15436 968 15488 982
rect 15672 982 15682 1148
rect 15682 982 15716 1148
rect 15716 982 15724 1148
rect 15672 968 15724 982
rect 16124 1358 16176 1372
rect 16124 1192 16132 1358
rect 16132 1192 16166 1358
rect 16166 1192 16176 1358
rect 16004 982 16014 1148
rect 16014 982 16048 1148
rect 16048 982 16056 1148
rect 16004 968 16056 982
rect 16360 1358 16412 1372
rect 16360 1192 16368 1358
rect 16368 1192 16402 1358
rect 16402 1192 16412 1358
rect 16240 982 16250 1148
rect 16250 982 16284 1148
rect 16284 982 16292 1148
rect 16240 968 16292 982
rect 16596 1358 16648 1372
rect 16596 1192 16604 1358
rect 16604 1192 16638 1358
rect 16638 1192 16648 1358
rect 16476 982 16486 1148
rect 16486 982 16520 1148
rect 16520 982 16528 1148
rect 16476 968 16528 982
rect 16712 982 16722 1148
rect 16722 982 16756 1148
rect 16756 982 16764 1148
rect 16712 968 16764 982
rect 17164 1358 17216 1372
rect 17164 1192 17172 1358
rect 17172 1192 17206 1358
rect 17206 1192 17216 1358
rect 17044 982 17054 1148
rect 17054 982 17088 1148
rect 17088 982 17096 1148
rect 17044 968 17096 982
rect 17400 1358 17452 1372
rect 17400 1192 17408 1358
rect 17408 1192 17442 1358
rect 17442 1192 17452 1358
rect 17280 982 17290 1148
rect 17290 982 17324 1148
rect 17324 982 17332 1148
rect 17280 968 17332 982
rect 17636 1358 17688 1372
rect 17636 1192 17644 1358
rect 17644 1192 17678 1358
rect 17678 1192 17688 1358
rect 17516 982 17526 1148
rect 17526 982 17560 1148
rect 17560 982 17568 1148
rect 17516 968 17568 982
rect 17752 982 17762 1148
rect 17762 982 17796 1148
rect 17796 982 17804 1148
rect 17752 968 17804 982
rect 18204 1358 18256 1372
rect 18204 1192 18212 1358
rect 18212 1192 18246 1358
rect 18246 1192 18256 1358
rect 18084 982 18094 1148
rect 18094 982 18128 1148
rect 18128 982 18136 1148
rect 18084 968 18136 982
rect 18440 1358 18492 1372
rect 18440 1192 18448 1358
rect 18448 1192 18482 1358
rect 18482 1192 18492 1358
rect 18320 982 18330 1148
rect 18330 982 18364 1148
rect 18364 982 18372 1148
rect 18320 968 18372 982
rect 18676 1358 18728 1372
rect 18676 1192 18684 1358
rect 18684 1192 18718 1358
rect 18718 1192 18728 1358
rect 18556 982 18566 1148
rect 18566 982 18600 1148
rect 18600 982 18608 1148
rect 18556 968 18608 982
rect 18792 982 18802 1148
rect 18802 982 18836 1148
rect 18836 982 18844 1148
rect 18792 968 18844 982
rect 11844 540 11896 552
rect 11844 372 11854 540
rect 11854 372 11888 540
rect 11888 372 11896 540
rect 12036 540 12088 552
rect 12036 372 12046 540
rect 12046 372 12080 540
rect 12080 372 12088 540
rect 11940 164 11950 332
rect 11950 164 11984 332
rect 11984 164 11992 332
rect 11940 152 11992 164
rect 12228 540 12280 552
rect 12228 372 12238 540
rect 12238 372 12272 540
rect 12272 372 12280 540
rect 12132 164 12142 332
rect 12142 164 12176 332
rect 12176 164 12184 332
rect 12132 152 12184 164
rect 12420 540 12472 552
rect 12420 372 12430 540
rect 12430 372 12464 540
rect 12464 372 12472 540
rect 12324 164 12334 332
rect 12334 164 12368 332
rect 12368 164 12376 332
rect 12324 152 12376 164
rect 12884 540 12936 552
rect 12884 372 12894 540
rect 12894 372 12928 540
rect 12928 372 12936 540
rect 13076 540 13128 552
rect 13076 372 13086 540
rect 13086 372 13120 540
rect 13120 372 13128 540
rect 12980 164 12990 332
rect 12990 164 13024 332
rect 13024 164 13032 332
rect 12980 152 13032 164
rect 13268 540 13320 552
rect 13268 372 13278 540
rect 13278 372 13312 540
rect 13312 372 13320 540
rect 13172 164 13182 332
rect 13182 164 13216 332
rect 13216 164 13224 332
rect 13172 152 13224 164
rect 13460 540 13512 552
rect 13460 372 13470 540
rect 13470 372 13504 540
rect 13504 372 13512 540
rect 13364 164 13374 332
rect 13374 164 13408 332
rect 13408 164 13416 332
rect 13364 152 13416 164
rect 13924 540 13976 552
rect 13924 372 13934 540
rect 13934 372 13968 540
rect 13968 372 13976 540
rect 14116 540 14168 552
rect 14116 372 14126 540
rect 14126 372 14160 540
rect 14160 372 14168 540
rect 14020 164 14030 332
rect 14030 164 14064 332
rect 14064 164 14072 332
rect 14020 152 14072 164
rect 14308 540 14360 552
rect 14308 372 14318 540
rect 14318 372 14352 540
rect 14352 372 14360 540
rect 14212 164 14222 332
rect 14222 164 14256 332
rect 14256 164 14264 332
rect 14212 152 14264 164
rect 14500 540 14552 552
rect 14500 372 14510 540
rect 14510 372 14544 540
rect 14544 372 14552 540
rect 14404 164 14414 332
rect 14414 164 14448 332
rect 14448 164 14456 332
rect 14404 152 14456 164
rect 14964 540 15016 552
rect 14964 372 14974 540
rect 14974 372 15008 540
rect 15008 372 15016 540
rect 15156 540 15208 552
rect 15156 372 15166 540
rect 15166 372 15200 540
rect 15200 372 15208 540
rect 15060 164 15070 332
rect 15070 164 15104 332
rect 15104 164 15112 332
rect 15060 152 15112 164
rect 15348 540 15400 552
rect 15348 372 15358 540
rect 15358 372 15392 540
rect 15392 372 15400 540
rect 15252 164 15262 332
rect 15262 164 15296 332
rect 15296 164 15304 332
rect 15252 152 15304 164
rect 15540 540 15592 552
rect 15540 372 15550 540
rect 15550 372 15584 540
rect 15584 372 15592 540
rect 15444 164 15454 332
rect 15454 164 15488 332
rect 15488 164 15496 332
rect 15444 152 15496 164
rect 16004 540 16056 552
rect 16004 372 16014 540
rect 16014 372 16048 540
rect 16048 372 16056 540
rect 16196 540 16248 552
rect 16196 372 16206 540
rect 16206 372 16240 540
rect 16240 372 16248 540
rect 16100 164 16110 332
rect 16110 164 16144 332
rect 16144 164 16152 332
rect 16100 152 16152 164
rect 16388 540 16440 552
rect 16388 372 16398 540
rect 16398 372 16432 540
rect 16432 372 16440 540
rect 16292 164 16302 332
rect 16302 164 16336 332
rect 16336 164 16344 332
rect 16292 152 16344 164
rect 16580 540 16632 552
rect 16580 372 16590 540
rect 16590 372 16624 540
rect 16624 372 16632 540
rect 16484 164 16494 332
rect 16494 164 16528 332
rect 16528 164 16536 332
rect 16484 152 16536 164
rect 17044 540 17096 552
rect 17044 372 17054 540
rect 17054 372 17088 540
rect 17088 372 17096 540
rect 17236 540 17288 552
rect 17236 372 17246 540
rect 17246 372 17280 540
rect 17280 372 17288 540
rect 17140 164 17150 332
rect 17150 164 17184 332
rect 17184 164 17192 332
rect 17140 152 17192 164
rect 17428 540 17480 552
rect 17428 372 17438 540
rect 17438 372 17472 540
rect 17472 372 17480 540
rect 17332 164 17342 332
rect 17342 164 17376 332
rect 17376 164 17384 332
rect 17332 152 17384 164
rect 17620 540 17672 552
rect 17620 372 17630 540
rect 17630 372 17664 540
rect 17664 372 17672 540
rect 17524 164 17534 332
rect 17534 164 17568 332
rect 17568 164 17576 332
rect 17524 152 17576 164
rect 18084 540 18136 552
rect 18084 372 18094 540
rect 18094 372 18128 540
rect 18128 372 18136 540
rect 18276 540 18328 552
rect 18276 372 18286 540
rect 18286 372 18320 540
rect 18320 372 18328 540
rect 18180 164 18190 332
rect 18190 164 18224 332
rect 18224 164 18232 332
rect 18180 152 18232 164
rect 18468 540 18520 552
rect 18468 372 18478 540
rect 18478 372 18512 540
rect 18512 372 18520 540
rect 18372 164 18382 332
rect 18382 164 18416 332
rect 18416 164 18424 332
rect 18372 152 18424 164
rect 18660 540 18712 552
rect 18660 372 18670 540
rect 18670 372 18704 540
rect 18704 372 18712 540
rect 18564 164 18574 332
rect 18574 164 18608 332
rect 18608 164 18616 332
rect 18564 152 18616 164
rect 4344 -882 4396 -868
rect 4344 -1048 4352 -882
rect 4352 -1048 4386 -882
rect 4386 -1048 4396 -882
rect 4224 -1258 4234 -1092
rect 4234 -1258 4268 -1092
rect 4268 -1258 4276 -1092
rect 4224 -1272 4276 -1258
rect 4580 -882 4632 -868
rect 4580 -1048 4588 -882
rect 4588 -1048 4622 -882
rect 4622 -1048 4632 -882
rect 4460 -1258 4470 -1092
rect 4470 -1258 4504 -1092
rect 4504 -1258 4512 -1092
rect 4460 -1272 4512 -1258
rect 4816 -882 4868 -868
rect 4816 -1048 4824 -882
rect 4824 -1048 4858 -882
rect 4858 -1048 4868 -882
rect 4696 -1258 4706 -1092
rect 4706 -1258 4740 -1092
rect 4740 -1258 4748 -1092
rect 4696 -1272 4748 -1258
rect 4932 -1258 4942 -1092
rect 4942 -1258 4976 -1092
rect 4976 -1258 4984 -1092
rect 4932 -1272 4984 -1258
rect 5384 -882 5436 -868
rect 5384 -1048 5392 -882
rect 5392 -1048 5426 -882
rect 5426 -1048 5436 -882
rect 5264 -1258 5274 -1092
rect 5274 -1258 5308 -1092
rect 5308 -1258 5316 -1092
rect 5264 -1272 5316 -1258
rect 5620 -882 5672 -868
rect 5620 -1048 5628 -882
rect 5628 -1048 5662 -882
rect 5662 -1048 5672 -882
rect 5500 -1258 5510 -1092
rect 5510 -1258 5544 -1092
rect 5544 -1258 5552 -1092
rect 5500 -1272 5552 -1258
rect 5856 -882 5908 -868
rect 5856 -1048 5864 -882
rect 5864 -1048 5898 -882
rect 5898 -1048 5908 -882
rect 5736 -1258 5746 -1092
rect 5746 -1258 5780 -1092
rect 5780 -1258 5788 -1092
rect 5736 -1272 5788 -1258
rect 5972 -1258 5982 -1092
rect 5982 -1258 6016 -1092
rect 6016 -1258 6024 -1092
rect 5972 -1272 6024 -1258
rect 6424 -882 6476 -868
rect 6424 -1048 6432 -882
rect 6432 -1048 6466 -882
rect 6466 -1048 6476 -882
rect 6304 -1258 6314 -1092
rect 6314 -1258 6348 -1092
rect 6348 -1258 6356 -1092
rect 6304 -1272 6356 -1258
rect 6660 -882 6712 -868
rect 6660 -1048 6668 -882
rect 6668 -1048 6702 -882
rect 6702 -1048 6712 -882
rect 6540 -1258 6550 -1092
rect 6550 -1258 6584 -1092
rect 6584 -1258 6592 -1092
rect 6540 -1272 6592 -1258
rect 6896 -882 6948 -868
rect 6896 -1048 6904 -882
rect 6904 -1048 6938 -882
rect 6938 -1048 6948 -882
rect 6776 -1258 6786 -1092
rect 6786 -1258 6820 -1092
rect 6820 -1258 6828 -1092
rect 6776 -1272 6828 -1258
rect 7012 -1258 7022 -1092
rect 7022 -1258 7056 -1092
rect 7056 -1258 7064 -1092
rect 7012 -1272 7064 -1258
rect 7464 -882 7516 -868
rect 7464 -1048 7472 -882
rect 7472 -1048 7506 -882
rect 7506 -1048 7516 -882
rect 7344 -1258 7354 -1092
rect 7354 -1258 7388 -1092
rect 7388 -1258 7396 -1092
rect 7344 -1272 7396 -1258
rect 7700 -882 7752 -868
rect 7700 -1048 7708 -882
rect 7708 -1048 7742 -882
rect 7742 -1048 7752 -882
rect 7580 -1258 7590 -1092
rect 7590 -1258 7624 -1092
rect 7624 -1258 7632 -1092
rect 7580 -1272 7632 -1258
rect 7936 -882 7988 -868
rect 7936 -1048 7944 -882
rect 7944 -1048 7978 -882
rect 7978 -1048 7988 -882
rect 7816 -1258 7826 -1092
rect 7826 -1258 7860 -1092
rect 7860 -1258 7868 -1092
rect 7816 -1272 7868 -1258
rect 8052 -1258 8062 -1092
rect 8062 -1258 8096 -1092
rect 8096 -1258 8104 -1092
rect 8052 -1272 8104 -1258
rect 8504 -882 8556 -868
rect 8504 -1048 8512 -882
rect 8512 -1048 8546 -882
rect 8546 -1048 8556 -882
rect 8384 -1258 8394 -1092
rect 8394 -1258 8428 -1092
rect 8428 -1258 8436 -1092
rect 8384 -1272 8436 -1258
rect 8740 -882 8792 -868
rect 8740 -1048 8748 -882
rect 8748 -1048 8782 -882
rect 8782 -1048 8792 -882
rect 8620 -1258 8630 -1092
rect 8630 -1258 8664 -1092
rect 8664 -1258 8672 -1092
rect 8620 -1272 8672 -1258
rect 8976 -882 9028 -868
rect 8976 -1048 8984 -882
rect 8984 -1048 9018 -882
rect 9018 -1048 9028 -882
rect 8856 -1258 8866 -1092
rect 8866 -1258 8900 -1092
rect 8900 -1258 8908 -1092
rect 8856 -1272 8908 -1258
rect 9092 -1258 9102 -1092
rect 9102 -1258 9136 -1092
rect 9136 -1258 9144 -1092
rect 9092 -1272 9144 -1258
rect 9544 -882 9596 -868
rect 9544 -1048 9552 -882
rect 9552 -1048 9586 -882
rect 9586 -1048 9596 -882
rect 9424 -1258 9434 -1092
rect 9434 -1258 9468 -1092
rect 9468 -1258 9476 -1092
rect 9424 -1272 9476 -1258
rect 9780 -882 9832 -868
rect 9780 -1048 9788 -882
rect 9788 -1048 9822 -882
rect 9822 -1048 9832 -882
rect 9660 -1258 9670 -1092
rect 9670 -1258 9704 -1092
rect 9704 -1258 9712 -1092
rect 9660 -1272 9712 -1258
rect 10016 -882 10068 -868
rect 10016 -1048 10024 -882
rect 10024 -1048 10058 -882
rect 10058 -1048 10068 -882
rect 9896 -1258 9906 -1092
rect 9906 -1258 9940 -1092
rect 9940 -1258 9948 -1092
rect 9896 -1272 9948 -1258
rect 10132 -1258 10142 -1092
rect 10142 -1258 10176 -1092
rect 10176 -1258 10184 -1092
rect 10132 -1272 10184 -1258
rect 10584 -882 10636 -868
rect 10584 -1048 10592 -882
rect 10592 -1048 10626 -882
rect 10626 -1048 10636 -882
rect 10464 -1258 10474 -1092
rect 10474 -1258 10508 -1092
rect 10508 -1258 10516 -1092
rect 10464 -1272 10516 -1258
rect 10820 -882 10872 -868
rect 10820 -1048 10828 -882
rect 10828 -1048 10862 -882
rect 10862 -1048 10872 -882
rect 10700 -1258 10710 -1092
rect 10710 -1258 10744 -1092
rect 10744 -1258 10752 -1092
rect 10700 -1272 10752 -1258
rect 11056 -882 11108 -868
rect 11056 -1048 11064 -882
rect 11064 -1048 11098 -882
rect 11098 -1048 11108 -882
rect 10936 -1258 10946 -1092
rect 10946 -1258 10980 -1092
rect 10980 -1258 10988 -1092
rect 10936 -1272 10988 -1258
rect 11172 -1258 11182 -1092
rect 11182 -1258 11216 -1092
rect 11216 -1258 11224 -1092
rect 11172 -1272 11224 -1258
rect 4224 -1700 4276 -1688
rect 4224 -1868 4234 -1700
rect 4234 -1868 4268 -1700
rect 4268 -1868 4276 -1700
rect 4416 -1700 4468 -1688
rect 4416 -1868 4426 -1700
rect 4426 -1868 4460 -1700
rect 4460 -1868 4468 -1700
rect 4320 -2076 4330 -1908
rect 4330 -2076 4364 -1908
rect 4364 -2076 4372 -1908
rect 4320 -2088 4372 -2076
rect 4608 -1700 4660 -1688
rect 4608 -1868 4618 -1700
rect 4618 -1868 4652 -1700
rect 4652 -1868 4660 -1700
rect 4512 -2076 4522 -1908
rect 4522 -2076 4556 -1908
rect 4556 -2076 4564 -1908
rect 4512 -2088 4564 -2076
rect 4800 -1700 4852 -1688
rect 4800 -1868 4810 -1700
rect 4810 -1868 4844 -1700
rect 4844 -1868 4852 -1700
rect 4704 -2076 4714 -1908
rect 4714 -2076 4748 -1908
rect 4748 -2076 4756 -1908
rect 4704 -2088 4756 -2076
rect 5264 -1700 5316 -1688
rect 5264 -1868 5274 -1700
rect 5274 -1868 5308 -1700
rect 5308 -1868 5316 -1700
rect 5456 -1700 5508 -1688
rect 5456 -1868 5466 -1700
rect 5466 -1868 5500 -1700
rect 5500 -1868 5508 -1700
rect 5360 -2076 5370 -1908
rect 5370 -2076 5404 -1908
rect 5404 -2076 5412 -1908
rect 5360 -2088 5412 -2076
rect 5648 -1700 5700 -1688
rect 5648 -1868 5658 -1700
rect 5658 -1868 5692 -1700
rect 5692 -1868 5700 -1700
rect 5552 -2076 5562 -1908
rect 5562 -2076 5596 -1908
rect 5596 -2076 5604 -1908
rect 5552 -2088 5604 -2076
rect 5840 -1700 5892 -1688
rect 5840 -1868 5850 -1700
rect 5850 -1868 5884 -1700
rect 5884 -1868 5892 -1700
rect 5744 -2076 5754 -1908
rect 5754 -2076 5788 -1908
rect 5788 -2076 5796 -1908
rect 5744 -2088 5796 -2076
rect 6304 -1700 6356 -1688
rect 6304 -1868 6314 -1700
rect 6314 -1868 6348 -1700
rect 6348 -1868 6356 -1700
rect 6496 -1700 6548 -1688
rect 6496 -1868 6506 -1700
rect 6506 -1868 6540 -1700
rect 6540 -1868 6548 -1700
rect 6400 -2076 6410 -1908
rect 6410 -2076 6444 -1908
rect 6444 -2076 6452 -1908
rect 6400 -2088 6452 -2076
rect 6688 -1700 6740 -1688
rect 6688 -1868 6698 -1700
rect 6698 -1868 6732 -1700
rect 6732 -1868 6740 -1700
rect 6592 -2076 6602 -1908
rect 6602 -2076 6636 -1908
rect 6636 -2076 6644 -1908
rect 6592 -2088 6644 -2076
rect 6880 -1700 6932 -1688
rect 6880 -1868 6890 -1700
rect 6890 -1868 6924 -1700
rect 6924 -1868 6932 -1700
rect 6784 -2076 6794 -1908
rect 6794 -2076 6828 -1908
rect 6828 -2076 6836 -1908
rect 6784 -2088 6836 -2076
rect 7344 -1700 7396 -1688
rect 7344 -1868 7354 -1700
rect 7354 -1868 7388 -1700
rect 7388 -1868 7396 -1700
rect 7536 -1700 7588 -1688
rect 7536 -1868 7546 -1700
rect 7546 -1868 7580 -1700
rect 7580 -1868 7588 -1700
rect 7440 -2076 7450 -1908
rect 7450 -2076 7484 -1908
rect 7484 -2076 7492 -1908
rect 7440 -2088 7492 -2076
rect 7728 -1700 7780 -1688
rect 7728 -1868 7738 -1700
rect 7738 -1868 7772 -1700
rect 7772 -1868 7780 -1700
rect 7632 -2076 7642 -1908
rect 7642 -2076 7676 -1908
rect 7676 -2076 7684 -1908
rect 7632 -2088 7684 -2076
rect 7920 -1700 7972 -1688
rect 7920 -1868 7930 -1700
rect 7930 -1868 7964 -1700
rect 7964 -1868 7972 -1700
rect 7824 -2076 7834 -1908
rect 7834 -2076 7868 -1908
rect 7868 -2076 7876 -1908
rect 7824 -2088 7876 -2076
rect 8384 -1700 8436 -1688
rect 8384 -1868 8394 -1700
rect 8394 -1868 8428 -1700
rect 8428 -1868 8436 -1700
rect 8576 -1700 8628 -1688
rect 8576 -1868 8586 -1700
rect 8586 -1868 8620 -1700
rect 8620 -1868 8628 -1700
rect 8480 -2076 8490 -1908
rect 8490 -2076 8524 -1908
rect 8524 -2076 8532 -1908
rect 8480 -2088 8532 -2076
rect 8768 -1700 8820 -1688
rect 8768 -1868 8778 -1700
rect 8778 -1868 8812 -1700
rect 8812 -1868 8820 -1700
rect 8672 -2076 8682 -1908
rect 8682 -2076 8716 -1908
rect 8716 -2076 8724 -1908
rect 8672 -2088 8724 -2076
rect 8960 -1700 9012 -1688
rect 8960 -1868 8970 -1700
rect 8970 -1868 9004 -1700
rect 9004 -1868 9012 -1700
rect 8864 -2076 8874 -1908
rect 8874 -2076 8908 -1908
rect 8908 -2076 8916 -1908
rect 8864 -2088 8916 -2076
rect 11940 -78 11992 -64
rect 11940 -244 11950 -78
rect 11950 -244 11984 -78
rect 11984 -244 11992 -78
rect 11844 -454 11854 -284
rect 11854 -454 11888 -284
rect 11888 -454 11896 -284
rect 11844 -464 11896 -454
rect 12132 -78 12184 -64
rect 12132 -244 12142 -78
rect 12142 -244 12176 -78
rect 12176 -244 12184 -78
rect 12036 -454 12046 -284
rect 12046 -454 12080 -284
rect 12080 -454 12088 -284
rect 12036 -464 12088 -454
rect 12324 -78 12376 -64
rect 12324 -244 12334 -78
rect 12334 -244 12368 -78
rect 12368 -244 12376 -78
rect 12228 -454 12238 -284
rect 12238 -454 12272 -284
rect 12272 -454 12280 -284
rect 12228 -464 12280 -454
rect 12420 -454 12430 -284
rect 12430 -454 12464 -284
rect 12464 -454 12472 -284
rect 12420 -464 12472 -454
rect 12980 -78 13032 -64
rect 12980 -244 12990 -78
rect 12990 -244 13024 -78
rect 13024 -244 13032 -78
rect 12884 -454 12894 -284
rect 12894 -454 12928 -284
rect 12928 -454 12936 -284
rect 12884 -464 12936 -454
rect 13172 -78 13224 -64
rect 13172 -244 13182 -78
rect 13182 -244 13216 -78
rect 13216 -244 13224 -78
rect 13076 -454 13086 -284
rect 13086 -454 13120 -284
rect 13120 -454 13128 -284
rect 13076 -464 13128 -454
rect 13364 -78 13416 -64
rect 13364 -244 13374 -78
rect 13374 -244 13408 -78
rect 13408 -244 13416 -78
rect 13268 -454 13278 -284
rect 13278 -454 13312 -284
rect 13312 -454 13320 -284
rect 13268 -464 13320 -454
rect 13460 -454 13470 -284
rect 13470 -454 13504 -284
rect 13504 -454 13512 -284
rect 13460 -464 13512 -454
rect 14020 -78 14072 -64
rect 14020 -244 14030 -78
rect 14030 -244 14064 -78
rect 14064 -244 14072 -78
rect 13924 -454 13934 -284
rect 13934 -454 13968 -284
rect 13968 -454 13976 -284
rect 13924 -464 13976 -454
rect 14212 -78 14264 -64
rect 14212 -244 14222 -78
rect 14222 -244 14256 -78
rect 14256 -244 14264 -78
rect 14116 -454 14126 -284
rect 14126 -454 14160 -284
rect 14160 -454 14168 -284
rect 14116 -464 14168 -454
rect 14404 -78 14456 -64
rect 14404 -244 14414 -78
rect 14414 -244 14448 -78
rect 14448 -244 14456 -78
rect 14308 -454 14318 -284
rect 14318 -454 14352 -284
rect 14352 -454 14360 -284
rect 14308 -464 14360 -454
rect 14500 -454 14510 -284
rect 14510 -454 14544 -284
rect 14544 -454 14552 -284
rect 14500 -464 14552 -454
rect 15060 -78 15112 -64
rect 15060 -244 15070 -78
rect 15070 -244 15104 -78
rect 15104 -244 15112 -78
rect 14964 -454 14974 -284
rect 14974 -454 15008 -284
rect 15008 -454 15016 -284
rect 14964 -464 15016 -454
rect 15252 -78 15304 -64
rect 15252 -244 15262 -78
rect 15262 -244 15296 -78
rect 15296 -244 15304 -78
rect 15156 -454 15166 -284
rect 15166 -454 15200 -284
rect 15200 -454 15208 -284
rect 15156 -464 15208 -454
rect 15444 -78 15496 -64
rect 15444 -244 15454 -78
rect 15454 -244 15488 -78
rect 15488 -244 15496 -78
rect 15348 -454 15358 -284
rect 15358 -454 15392 -284
rect 15392 -454 15400 -284
rect 15348 -464 15400 -454
rect 15540 -454 15550 -284
rect 15550 -454 15584 -284
rect 15584 -454 15592 -284
rect 15540 -464 15592 -454
rect 16100 -78 16152 -64
rect 16100 -244 16110 -78
rect 16110 -244 16144 -78
rect 16144 -244 16152 -78
rect 16004 -454 16014 -284
rect 16014 -454 16048 -284
rect 16048 -454 16056 -284
rect 16004 -464 16056 -454
rect 16292 -78 16344 -64
rect 16292 -244 16302 -78
rect 16302 -244 16336 -78
rect 16336 -244 16344 -78
rect 16196 -454 16206 -284
rect 16206 -454 16240 -284
rect 16240 -454 16248 -284
rect 16196 -464 16248 -454
rect 16484 -78 16536 -64
rect 16484 -244 16494 -78
rect 16494 -244 16528 -78
rect 16528 -244 16536 -78
rect 16388 -454 16398 -284
rect 16398 -454 16432 -284
rect 16432 -454 16440 -284
rect 16388 -464 16440 -454
rect 16580 -454 16590 -284
rect 16590 -454 16624 -284
rect 16624 -454 16632 -284
rect 16580 -464 16632 -454
rect 17140 -78 17192 -64
rect 17140 -244 17150 -78
rect 17150 -244 17184 -78
rect 17184 -244 17192 -78
rect 17044 -454 17054 -284
rect 17054 -454 17088 -284
rect 17088 -454 17096 -284
rect 17044 -464 17096 -454
rect 17332 -78 17384 -64
rect 17332 -244 17342 -78
rect 17342 -244 17376 -78
rect 17376 -244 17384 -78
rect 17236 -454 17246 -284
rect 17246 -454 17280 -284
rect 17280 -454 17288 -284
rect 17236 -464 17288 -454
rect 17524 -78 17576 -64
rect 17524 -244 17534 -78
rect 17534 -244 17568 -78
rect 17568 -244 17576 -78
rect 17428 -454 17438 -284
rect 17438 -454 17472 -284
rect 17472 -454 17480 -284
rect 17428 -464 17480 -454
rect 17620 -454 17630 -284
rect 17630 -454 17664 -284
rect 17664 -454 17672 -284
rect 17620 -464 17672 -454
rect 18180 -78 18232 -64
rect 18180 -244 18190 -78
rect 18190 -244 18224 -78
rect 18224 -244 18232 -78
rect 18084 -454 18094 -284
rect 18094 -454 18128 -284
rect 18128 -454 18136 -284
rect 18084 -464 18136 -454
rect 18372 -78 18424 -64
rect 18372 -244 18382 -78
rect 18382 -244 18416 -78
rect 18416 -244 18424 -78
rect 18276 -454 18286 -284
rect 18286 -454 18320 -284
rect 18320 -454 18328 -284
rect 18276 -464 18328 -454
rect 18564 -78 18616 -64
rect 18564 -244 18574 -78
rect 18574 -244 18608 -78
rect 18608 -244 18616 -78
rect 18468 -454 18478 -284
rect 18478 -454 18512 -284
rect 18512 -454 18520 -284
rect 18468 -464 18520 -454
rect 18660 -454 18670 -284
rect 18670 -454 18704 -284
rect 18704 -454 18712 -284
rect 18660 -464 18712 -454
rect 11964 -882 12016 -868
rect 11964 -1048 11972 -882
rect 11972 -1048 12006 -882
rect 12006 -1048 12016 -882
rect 11844 -1258 11854 -1092
rect 11854 -1258 11888 -1092
rect 11888 -1258 11896 -1092
rect 11844 -1272 11896 -1258
rect 12200 -882 12252 -868
rect 12200 -1048 12208 -882
rect 12208 -1048 12242 -882
rect 12242 -1048 12252 -882
rect 12080 -1258 12090 -1092
rect 12090 -1258 12124 -1092
rect 12124 -1258 12132 -1092
rect 12080 -1272 12132 -1258
rect 12436 -882 12488 -868
rect 12436 -1048 12444 -882
rect 12444 -1048 12478 -882
rect 12478 -1048 12488 -882
rect 12316 -1258 12326 -1092
rect 12326 -1258 12360 -1092
rect 12360 -1258 12368 -1092
rect 12316 -1272 12368 -1258
rect 12552 -1258 12562 -1092
rect 12562 -1258 12596 -1092
rect 12596 -1258 12604 -1092
rect 12552 -1272 12604 -1258
rect 13004 -882 13056 -868
rect 13004 -1048 13012 -882
rect 13012 -1048 13046 -882
rect 13046 -1048 13056 -882
rect 12884 -1258 12894 -1092
rect 12894 -1258 12928 -1092
rect 12928 -1258 12936 -1092
rect 12884 -1272 12936 -1258
rect 13240 -882 13292 -868
rect 13240 -1048 13248 -882
rect 13248 -1048 13282 -882
rect 13282 -1048 13292 -882
rect 13120 -1258 13130 -1092
rect 13130 -1258 13164 -1092
rect 13164 -1258 13172 -1092
rect 13120 -1272 13172 -1258
rect 13476 -882 13528 -868
rect 13476 -1048 13484 -882
rect 13484 -1048 13518 -882
rect 13518 -1048 13528 -882
rect 13356 -1258 13366 -1092
rect 13366 -1258 13400 -1092
rect 13400 -1258 13408 -1092
rect 13356 -1272 13408 -1258
rect 13592 -1258 13602 -1092
rect 13602 -1258 13636 -1092
rect 13636 -1258 13644 -1092
rect 13592 -1272 13644 -1258
rect 14044 -882 14096 -868
rect 14044 -1048 14052 -882
rect 14052 -1048 14086 -882
rect 14086 -1048 14096 -882
rect 13924 -1258 13934 -1092
rect 13934 -1258 13968 -1092
rect 13968 -1258 13976 -1092
rect 13924 -1272 13976 -1258
rect 14280 -882 14332 -868
rect 14280 -1048 14288 -882
rect 14288 -1048 14322 -882
rect 14322 -1048 14332 -882
rect 14160 -1258 14170 -1092
rect 14170 -1258 14204 -1092
rect 14204 -1258 14212 -1092
rect 14160 -1272 14212 -1258
rect 14516 -882 14568 -868
rect 14516 -1048 14524 -882
rect 14524 -1048 14558 -882
rect 14558 -1048 14568 -882
rect 14396 -1258 14406 -1092
rect 14406 -1258 14440 -1092
rect 14440 -1258 14448 -1092
rect 14396 -1272 14448 -1258
rect 14632 -1258 14642 -1092
rect 14642 -1258 14676 -1092
rect 14676 -1258 14684 -1092
rect 14632 -1272 14684 -1258
rect 15084 -882 15136 -868
rect 15084 -1048 15092 -882
rect 15092 -1048 15126 -882
rect 15126 -1048 15136 -882
rect 14964 -1258 14974 -1092
rect 14974 -1258 15008 -1092
rect 15008 -1258 15016 -1092
rect 14964 -1272 15016 -1258
rect 15320 -882 15372 -868
rect 15320 -1048 15328 -882
rect 15328 -1048 15362 -882
rect 15362 -1048 15372 -882
rect 15200 -1258 15210 -1092
rect 15210 -1258 15244 -1092
rect 15244 -1258 15252 -1092
rect 15200 -1272 15252 -1258
rect 15556 -882 15608 -868
rect 15556 -1048 15564 -882
rect 15564 -1048 15598 -882
rect 15598 -1048 15608 -882
rect 15436 -1258 15446 -1092
rect 15446 -1258 15480 -1092
rect 15480 -1258 15488 -1092
rect 15436 -1272 15488 -1258
rect 15672 -1258 15682 -1092
rect 15682 -1258 15716 -1092
rect 15716 -1258 15724 -1092
rect 15672 -1272 15724 -1258
rect 16124 -882 16176 -868
rect 16124 -1048 16132 -882
rect 16132 -1048 16166 -882
rect 16166 -1048 16176 -882
rect 16004 -1258 16014 -1092
rect 16014 -1258 16048 -1092
rect 16048 -1258 16056 -1092
rect 16004 -1272 16056 -1258
rect 16360 -882 16412 -868
rect 16360 -1048 16368 -882
rect 16368 -1048 16402 -882
rect 16402 -1048 16412 -882
rect 16240 -1258 16250 -1092
rect 16250 -1258 16284 -1092
rect 16284 -1258 16292 -1092
rect 16240 -1272 16292 -1258
rect 16596 -882 16648 -868
rect 16596 -1048 16604 -882
rect 16604 -1048 16638 -882
rect 16638 -1048 16648 -882
rect 16476 -1258 16486 -1092
rect 16486 -1258 16520 -1092
rect 16520 -1258 16528 -1092
rect 16476 -1272 16528 -1258
rect 16712 -1258 16722 -1092
rect 16722 -1258 16756 -1092
rect 16756 -1258 16764 -1092
rect 16712 -1272 16764 -1258
rect 17164 -882 17216 -868
rect 17164 -1048 17172 -882
rect 17172 -1048 17206 -882
rect 17206 -1048 17216 -882
rect 17044 -1258 17054 -1092
rect 17054 -1258 17088 -1092
rect 17088 -1258 17096 -1092
rect 17044 -1272 17096 -1258
rect 17400 -882 17452 -868
rect 17400 -1048 17408 -882
rect 17408 -1048 17442 -882
rect 17442 -1048 17452 -882
rect 17280 -1258 17290 -1092
rect 17290 -1258 17324 -1092
rect 17324 -1258 17332 -1092
rect 17280 -1272 17332 -1258
rect 17636 -882 17688 -868
rect 17636 -1048 17644 -882
rect 17644 -1048 17678 -882
rect 17678 -1048 17688 -882
rect 17516 -1258 17526 -1092
rect 17526 -1258 17560 -1092
rect 17560 -1258 17568 -1092
rect 17516 -1272 17568 -1258
rect 17752 -1258 17762 -1092
rect 17762 -1258 17796 -1092
rect 17796 -1258 17804 -1092
rect 17752 -1272 17804 -1258
rect 18204 -882 18256 -868
rect 18204 -1048 18212 -882
rect 18212 -1048 18246 -882
rect 18246 -1048 18256 -882
rect 18084 -1258 18094 -1092
rect 18094 -1258 18128 -1092
rect 18128 -1258 18136 -1092
rect 18084 -1272 18136 -1258
rect 18440 -882 18492 -868
rect 18440 -1048 18448 -882
rect 18448 -1048 18482 -882
rect 18482 -1048 18492 -882
rect 18320 -1258 18330 -1092
rect 18330 -1258 18364 -1092
rect 18364 -1258 18372 -1092
rect 18320 -1272 18372 -1258
rect 18676 -882 18728 -868
rect 18676 -1048 18684 -882
rect 18684 -1048 18718 -882
rect 18718 -1048 18728 -882
rect 18556 -1258 18566 -1092
rect 18566 -1258 18600 -1092
rect 18600 -1258 18608 -1092
rect 18556 -1272 18608 -1258
rect 18792 -1258 18802 -1092
rect 18802 -1258 18836 -1092
rect 18836 -1258 18844 -1092
rect 18792 -1272 18844 -1258
rect 11844 -1700 11896 -1688
rect 11844 -1868 11854 -1700
rect 11854 -1868 11888 -1700
rect 11888 -1868 11896 -1700
rect 12036 -1700 12088 -1688
rect 12036 -1868 12046 -1700
rect 12046 -1868 12080 -1700
rect 12080 -1868 12088 -1700
rect 11940 -2076 11950 -1908
rect 11950 -2076 11984 -1908
rect 11984 -2076 11992 -1908
rect 11940 -2088 11992 -2076
rect 12228 -1700 12280 -1688
rect 12228 -1868 12238 -1700
rect 12238 -1868 12272 -1700
rect 12272 -1868 12280 -1700
rect 12132 -2076 12142 -1908
rect 12142 -2076 12176 -1908
rect 12176 -2076 12184 -1908
rect 12132 -2088 12184 -2076
rect 12420 -1700 12472 -1688
rect 12420 -1868 12430 -1700
rect 12430 -1868 12464 -1700
rect 12464 -1868 12472 -1700
rect 12324 -2076 12334 -1908
rect 12334 -2076 12368 -1908
rect 12368 -2076 12376 -1908
rect 12324 -2088 12376 -2076
rect 12884 -1700 12936 -1688
rect 12884 -1868 12894 -1700
rect 12894 -1868 12928 -1700
rect 12928 -1868 12936 -1700
rect 13076 -1700 13128 -1688
rect 13076 -1868 13086 -1700
rect 13086 -1868 13120 -1700
rect 13120 -1868 13128 -1700
rect 12980 -2076 12990 -1908
rect 12990 -2076 13024 -1908
rect 13024 -2076 13032 -1908
rect 12980 -2088 13032 -2076
rect 13268 -1700 13320 -1688
rect 13268 -1868 13278 -1700
rect 13278 -1868 13312 -1700
rect 13312 -1868 13320 -1700
rect 13172 -2076 13182 -1908
rect 13182 -2076 13216 -1908
rect 13216 -2076 13224 -1908
rect 13172 -2088 13224 -2076
rect 13460 -1700 13512 -1688
rect 13460 -1868 13470 -1700
rect 13470 -1868 13504 -1700
rect 13504 -1868 13512 -1700
rect 13364 -2076 13374 -1908
rect 13374 -2076 13408 -1908
rect 13408 -2076 13416 -1908
rect 13364 -2088 13416 -2076
rect 13924 -1700 13976 -1688
rect 13924 -1868 13934 -1700
rect 13934 -1868 13968 -1700
rect 13968 -1868 13976 -1700
rect 14116 -1700 14168 -1688
rect 14116 -1868 14126 -1700
rect 14126 -1868 14160 -1700
rect 14160 -1868 14168 -1700
rect 14020 -2076 14030 -1908
rect 14030 -2076 14064 -1908
rect 14064 -2076 14072 -1908
rect 14020 -2088 14072 -2076
rect 14308 -1700 14360 -1688
rect 14308 -1868 14318 -1700
rect 14318 -1868 14352 -1700
rect 14352 -1868 14360 -1700
rect 14212 -2076 14222 -1908
rect 14222 -2076 14256 -1908
rect 14256 -2076 14264 -1908
rect 14212 -2088 14264 -2076
rect 14500 -1700 14552 -1688
rect 14500 -1868 14510 -1700
rect 14510 -1868 14544 -1700
rect 14544 -1868 14552 -1700
rect 14404 -2076 14414 -1908
rect 14414 -2076 14448 -1908
rect 14448 -2076 14456 -1908
rect 14404 -2088 14456 -2076
rect 14964 -1700 15016 -1688
rect 14964 -1868 14974 -1700
rect 14974 -1868 15008 -1700
rect 15008 -1868 15016 -1700
rect 15156 -1700 15208 -1688
rect 15156 -1868 15166 -1700
rect 15166 -1868 15200 -1700
rect 15200 -1868 15208 -1700
rect 15060 -2076 15070 -1908
rect 15070 -2076 15104 -1908
rect 15104 -2076 15112 -1908
rect 15060 -2088 15112 -2076
rect 15348 -1700 15400 -1688
rect 15348 -1868 15358 -1700
rect 15358 -1868 15392 -1700
rect 15392 -1868 15400 -1700
rect 15252 -2076 15262 -1908
rect 15262 -2076 15296 -1908
rect 15296 -2076 15304 -1908
rect 15252 -2088 15304 -2076
rect 15540 -1700 15592 -1688
rect 15540 -1868 15550 -1700
rect 15550 -1868 15584 -1700
rect 15584 -1868 15592 -1700
rect 15444 -2076 15454 -1908
rect 15454 -2076 15488 -1908
rect 15488 -2076 15496 -1908
rect 15444 -2088 15496 -2076
rect 16004 -1700 16056 -1688
rect 16004 -1868 16014 -1700
rect 16014 -1868 16048 -1700
rect 16048 -1868 16056 -1700
rect 16196 -1700 16248 -1688
rect 16196 -1868 16206 -1700
rect 16206 -1868 16240 -1700
rect 16240 -1868 16248 -1700
rect 16100 -2076 16110 -1908
rect 16110 -2076 16144 -1908
rect 16144 -2076 16152 -1908
rect 16100 -2088 16152 -2076
rect 16388 -1700 16440 -1688
rect 16388 -1868 16398 -1700
rect 16398 -1868 16432 -1700
rect 16432 -1868 16440 -1700
rect 16292 -2076 16302 -1908
rect 16302 -2076 16336 -1908
rect 16336 -2076 16344 -1908
rect 16292 -2088 16344 -2076
rect 16580 -1700 16632 -1688
rect 16580 -1868 16590 -1700
rect 16590 -1868 16624 -1700
rect 16624 -1868 16632 -1700
rect 16484 -2076 16494 -1908
rect 16494 -2076 16528 -1908
rect 16528 -2076 16536 -1908
rect 16484 -2088 16536 -2076
rect -7314 -2520 -7262 -2506
rect -7314 -2686 -7304 -2520
rect -7304 -2686 -7270 -2520
rect -7270 -2686 -7262 -2520
rect -7410 -2896 -7400 -2726
rect -7400 -2896 -7366 -2726
rect -7366 -2896 -7358 -2726
rect -7410 -2906 -7358 -2896
rect -7122 -2520 -7070 -2506
rect -7122 -2686 -7112 -2520
rect -7112 -2686 -7078 -2520
rect -7078 -2686 -7070 -2520
rect -7218 -2896 -7208 -2726
rect -7208 -2896 -7174 -2726
rect -7174 -2896 -7166 -2726
rect -7218 -2906 -7166 -2896
rect -6930 -2520 -6878 -2506
rect -6930 -2686 -6920 -2520
rect -6920 -2686 -6886 -2520
rect -6886 -2686 -6878 -2520
rect -7026 -2896 -7016 -2726
rect -7016 -2896 -6982 -2726
rect -6982 -2896 -6974 -2726
rect -7026 -2906 -6974 -2896
rect -6834 -2896 -6824 -2726
rect -6824 -2896 -6790 -2726
rect -6790 -2896 -6782 -2726
rect -6834 -2906 -6782 -2896
rect 4320 -2318 4372 -2304
rect 4320 -2484 4330 -2318
rect 4330 -2484 4364 -2318
rect 4364 -2484 4372 -2318
rect 4224 -2694 4234 -2524
rect 4234 -2694 4268 -2524
rect 4268 -2694 4276 -2524
rect 4224 -2704 4276 -2694
rect 4512 -2318 4564 -2304
rect 4512 -2484 4522 -2318
rect 4522 -2484 4556 -2318
rect 4556 -2484 4564 -2318
rect 4416 -2694 4426 -2524
rect 4426 -2694 4460 -2524
rect 4460 -2694 4468 -2524
rect 4416 -2704 4468 -2694
rect 4704 -2318 4756 -2304
rect 4704 -2484 4714 -2318
rect 4714 -2484 4748 -2318
rect 4748 -2484 4756 -2318
rect 4608 -2694 4618 -2524
rect 4618 -2694 4652 -2524
rect 4652 -2694 4660 -2524
rect 4608 -2704 4660 -2694
rect 4800 -2694 4810 -2524
rect 4810 -2694 4844 -2524
rect 4844 -2694 4852 -2524
rect 4800 -2704 4852 -2694
rect 5360 -2318 5412 -2304
rect 5360 -2484 5370 -2318
rect 5370 -2484 5404 -2318
rect 5404 -2484 5412 -2318
rect 5264 -2694 5274 -2524
rect 5274 -2694 5308 -2524
rect 5308 -2694 5316 -2524
rect 5264 -2704 5316 -2694
rect 5552 -2318 5604 -2304
rect 5552 -2484 5562 -2318
rect 5562 -2484 5596 -2318
rect 5596 -2484 5604 -2318
rect 5456 -2694 5466 -2524
rect 5466 -2694 5500 -2524
rect 5500 -2694 5508 -2524
rect 5456 -2704 5508 -2694
rect 5744 -2318 5796 -2304
rect 5744 -2484 5754 -2318
rect 5754 -2484 5788 -2318
rect 5788 -2484 5796 -2318
rect 5648 -2694 5658 -2524
rect 5658 -2694 5692 -2524
rect 5692 -2694 5700 -2524
rect 5648 -2704 5700 -2694
rect 5840 -2694 5850 -2524
rect 5850 -2694 5884 -2524
rect 5884 -2694 5892 -2524
rect 5840 -2704 5892 -2694
rect 6400 -2318 6452 -2304
rect 6400 -2484 6410 -2318
rect 6410 -2484 6444 -2318
rect 6444 -2484 6452 -2318
rect 6304 -2694 6314 -2524
rect 6314 -2694 6348 -2524
rect 6348 -2694 6356 -2524
rect 6304 -2704 6356 -2694
rect 6592 -2318 6644 -2304
rect 6592 -2484 6602 -2318
rect 6602 -2484 6636 -2318
rect 6636 -2484 6644 -2318
rect 6496 -2694 6506 -2524
rect 6506 -2694 6540 -2524
rect 6540 -2694 6548 -2524
rect 6496 -2704 6548 -2694
rect 6784 -2318 6836 -2304
rect 6784 -2484 6794 -2318
rect 6794 -2484 6828 -2318
rect 6828 -2484 6836 -2318
rect 6688 -2694 6698 -2524
rect 6698 -2694 6732 -2524
rect 6732 -2694 6740 -2524
rect 6688 -2704 6740 -2694
rect 6880 -2694 6890 -2524
rect 6890 -2694 6924 -2524
rect 6924 -2694 6932 -2524
rect 6880 -2704 6932 -2694
rect 7440 -2318 7492 -2304
rect 7440 -2484 7450 -2318
rect 7450 -2484 7484 -2318
rect 7484 -2484 7492 -2318
rect 7344 -2694 7354 -2524
rect 7354 -2694 7388 -2524
rect 7388 -2694 7396 -2524
rect 7344 -2704 7396 -2694
rect 7632 -2318 7684 -2304
rect 7632 -2484 7642 -2318
rect 7642 -2484 7676 -2318
rect 7676 -2484 7684 -2318
rect 7536 -2694 7546 -2524
rect 7546 -2694 7580 -2524
rect 7580 -2694 7588 -2524
rect 7536 -2704 7588 -2694
rect 7824 -2318 7876 -2304
rect 7824 -2484 7834 -2318
rect 7834 -2484 7868 -2318
rect 7868 -2484 7876 -2318
rect 7728 -2694 7738 -2524
rect 7738 -2694 7772 -2524
rect 7772 -2694 7780 -2524
rect 7728 -2704 7780 -2694
rect 7920 -2694 7930 -2524
rect 7930 -2694 7964 -2524
rect 7964 -2694 7972 -2524
rect 7920 -2704 7972 -2694
rect 8480 -2318 8532 -2304
rect 8480 -2484 8490 -2318
rect 8490 -2484 8524 -2318
rect 8524 -2484 8532 -2318
rect 8384 -2694 8394 -2524
rect 8394 -2694 8428 -2524
rect 8428 -2694 8436 -2524
rect 8384 -2704 8436 -2694
rect 8672 -2318 8724 -2304
rect 8672 -2484 8682 -2318
rect 8682 -2484 8716 -2318
rect 8716 -2484 8724 -2318
rect 8576 -2694 8586 -2524
rect 8586 -2694 8620 -2524
rect 8620 -2694 8628 -2524
rect 8576 -2704 8628 -2694
rect 8864 -2318 8916 -2304
rect 8864 -2484 8874 -2318
rect 8874 -2484 8908 -2318
rect 8908 -2484 8916 -2318
rect 8768 -2694 8778 -2524
rect 8778 -2694 8812 -2524
rect 8812 -2694 8820 -2524
rect 8768 -2704 8820 -2694
rect 8960 -2694 8970 -2524
rect 8970 -2694 9004 -2524
rect 9004 -2694 9012 -2524
rect 8960 -2704 9012 -2694
rect 11940 -2318 11992 -2304
rect 11940 -2484 11950 -2318
rect 11950 -2484 11984 -2318
rect 11984 -2484 11992 -2318
rect 11844 -2694 11854 -2524
rect 11854 -2694 11888 -2524
rect 11888 -2694 11896 -2524
rect 11844 -2704 11896 -2694
rect 12132 -2318 12184 -2304
rect 12132 -2484 12142 -2318
rect 12142 -2484 12176 -2318
rect 12176 -2484 12184 -2318
rect 12036 -2694 12046 -2524
rect 12046 -2694 12080 -2524
rect 12080 -2694 12088 -2524
rect 12036 -2704 12088 -2694
rect 12324 -2318 12376 -2304
rect 12324 -2484 12334 -2318
rect 12334 -2484 12368 -2318
rect 12368 -2484 12376 -2318
rect 12228 -2694 12238 -2524
rect 12238 -2694 12272 -2524
rect 12272 -2694 12280 -2524
rect 12228 -2704 12280 -2694
rect 12420 -2694 12430 -2524
rect 12430 -2694 12464 -2524
rect 12464 -2694 12472 -2524
rect 12420 -2704 12472 -2694
rect 12980 -2318 13032 -2304
rect 12980 -2484 12990 -2318
rect 12990 -2484 13024 -2318
rect 13024 -2484 13032 -2318
rect 12884 -2694 12894 -2524
rect 12894 -2694 12928 -2524
rect 12928 -2694 12936 -2524
rect 12884 -2704 12936 -2694
rect 13172 -2318 13224 -2304
rect 13172 -2484 13182 -2318
rect 13182 -2484 13216 -2318
rect 13216 -2484 13224 -2318
rect 13076 -2694 13086 -2524
rect 13086 -2694 13120 -2524
rect 13120 -2694 13128 -2524
rect 13076 -2704 13128 -2694
rect 13364 -2318 13416 -2304
rect 13364 -2484 13374 -2318
rect 13374 -2484 13408 -2318
rect 13408 -2484 13416 -2318
rect 13268 -2694 13278 -2524
rect 13278 -2694 13312 -2524
rect 13312 -2694 13320 -2524
rect 13268 -2704 13320 -2694
rect 13460 -2694 13470 -2524
rect 13470 -2694 13504 -2524
rect 13504 -2694 13512 -2524
rect 13460 -2704 13512 -2694
rect 14020 -2318 14072 -2304
rect 14020 -2484 14030 -2318
rect 14030 -2484 14064 -2318
rect 14064 -2484 14072 -2318
rect 13924 -2694 13934 -2524
rect 13934 -2694 13968 -2524
rect 13968 -2694 13976 -2524
rect 13924 -2704 13976 -2694
rect 14212 -2318 14264 -2304
rect 14212 -2484 14222 -2318
rect 14222 -2484 14256 -2318
rect 14256 -2484 14264 -2318
rect 14116 -2694 14126 -2524
rect 14126 -2694 14160 -2524
rect 14160 -2694 14168 -2524
rect 14116 -2704 14168 -2694
rect 14404 -2318 14456 -2304
rect 14404 -2484 14414 -2318
rect 14414 -2484 14448 -2318
rect 14448 -2484 14456 -2318
rect 14308 -2694 14318 -2524
rect 14318 -2694 14352 -2524
rect 14352 -2694 14360 -2524
rect 14308 -2704 14360 -2694
rect 14500 -2694 14510 -2524
rect 14510 -2694 14544 -2524
rect 14544 -2694 14552 -2524
rect 14500 -2704 14552 -2694
rect 15060 -2318 15112 -2304
rect 15060 -2484 15070 -2318
rect 15070 -2484 15104 -2318
rect 15104 -2484 15112 -2318
rect 14964 -2694 14974 -2524
rect 14974 -2694 15008 -2524
rect 15008 -2694 15016 -2524
rect 14964 -2704 15016 -2694
rect 15252 -2318 15304 -2304
rect 15252 -2484 15262 -2318
rect 15262 -2484 15296 -2318
rect 15296 -2484 15304 -2318
rect 15156 -2694 15166 -2524
rect 15166 -2694 15200 -2524
rect 15200 -2694 15208 -2524
rect 15156 -2704 15208 -2694
rect 15444 -2318 15496 -2304
rect 15444 -2484 15454 -2318
rect 15454 -2484 15488 -2318
rect 15488 -2484 15496 -2318
rect 15348 -2694 15358 -2524
rect 15358 -2694 15392 -2524
rect 15392 -2694 15400 -2524
rect 15348 -2704 15400 -2694
rect 15540 -2694 15550 -2524
rect 15550 -2694 15584 -2524
rect 15584 -2694 15592 -2524
rect 15540 -2704 15592 -2694
rect 16100 -2318 16152 -2304
rect 16100 -2484 16110 -2318
rect 16110 -2484 16144 -2318
rect 16144 -2484 16152 -2318
rect 16004 -2694 16014 -2524
rect 16014 -2694 16048 -2524
rect 16048 -2694 16056 -2524
rect 16004 -2704 16056 -2694
rect 16292 -2318 16344 -2304
rect 16292 -2484 16302 -2318
rect 16302 -2484 16336 -2318
rect 16336 -2484 16344 -2318
rect 16196 -2694 16206 -2524
rect 16206 -2694 16240 -2524
rect 16240 -2694 16248 -2524
rect 16196 -2704 16248 -2694
rect 16484 -2318 16536 -2304
rect 16484 -2484 16494 -2318
rect 16494 -2484 16528 -2318
rect 16528 -2484 16536 -2318
rect 16388 -2694 16398 -2524
rect 16398 -2694 16432 -2524
rect 16432 -2694 16440 -2524
rect 16388 -2704 16440 -2694
rect 16580 -2694 16590 -2524
rect 16590 -2694 16624 -2524
rect 16624 -2694 16632 -2524
rect 16580 -2704 16632 -2694
rect -7290 -3324 -7238 -3310
rect -7290 -3490 -7282 -3324
rect -7282 -3490 -7248 -3324
rect -7248 -3490 -7238 -3324
rect -7410 -3700 -7400 -3534
rect -7400 -3700 -7366 -3534
rect -7366 -3700 -7358 -3534
rect -7410 -3714 -7358 -3700
rect -7054 -3324 -7002 -3310
rect -7054 -3490 -7046 -3324
rect -7046 -3490 -7012 -3324
rect -7012 -3490 -7002 -3324
rect -7174 -3700 -7164 -3534
rect -7164 -3700 -7130 -3534
rect -7130 -3700 -7122 -3534
rect -7174 -3714 -7122 -3700
rect -6818 -3324 -6766 -3310
rect -6818 -3490 -6810 -3324
rect -6810 -3490 -6776 -3324
rect -6776 -3490 -6766 -3324
rect -6938 -3700 -6928 -3534
rect -6928 -3700 -6894 -3534
rect -6894 -3700 -6886 -3534
rect -6938 -3714 -6886 -3700
rect -6702 -3700 -6692 -3534
rect -6692 -3700 -6658 -3534
rect -6658 -3700 -6650 -3534
rect -6702 -3714 -6650 -3700
rect 4344 -3122 4396 -3108
rect 4344 -3288 4352 -3122
rect 4352 -3288 4386 -3122
rect 4386 -3288 4396 -3122
rect 4224 -3498 4234 -3332
rect 4234 -3498 4268 -3332
rect 4268 -3498 4276 -3332
rect 4224 -3512 4276 -3498
rect 4580 -3122 4632 -3108
rect 4580 -3288 4588 -3122
rect 4588 -3288 4622 -3122
rect 4622 -3288 4632 -3122
rect 4460 -3498 4470 -3332
rect 4470 -3498 4504 -3332
rect 4504 -3498 4512 -3332
rect 4460 -3512 4512 -3498
rect 4816 -3122 4868 -3108
rect 4816 -3288 4824 -3122
rect 4824 -3288 4858 -3122
rect 4858 -3288 4868 -3122
rect 4696 -3498 4706 -3332
rect 4706 -3498 4740 -3332
rect 4740 -3498 4748 -3332
rect 4696 -3512 4748 -3498
rect 4932 -3498 4942 -3332
rect 4942 -3498 4976 -3332
rect 4976 -3498 4984 -3332
rect 4932 -3512 4984 -3498
rect 5384 -3122 5436 -3108
rect 5384 -3288 5392 -3122
rect 5392 -3288 5426 -3122
rect 5426 -3288 5436 -3122
rect 5264 -3498 5274 -3332
rect 5274 -3498 5308 -3332
rect 5308 -3498 5316 -3332
rect 5264 -3512 5316 -3498
rect 5620 -3122 5672 -3108
rect 5620 -3288 5628 -3122
rect 5628 -3288 5662 -3122
rect 5662 -3288 5672 -3122
rect 5500 -3498 5510 -3332
rect 5510 -3498 5544 -3332
rect 5544 -3498 5552 -3332
rect 5500 -3512 5552 -3498
rect 5856 -3122 5908 -3108
rect 5856 -3288 5864 -3122
rect 5864 -3288 5898 -3122
rect 5898 -3288 5908 -3122
rect 5736 -3498 5746 -3332
rect 5746 -3498 5780 -3332
rect 5780 -3498 5788 -3332
rect 5736 -3512 5788 -3498
rect 5972 -3498 5982 -3332
rect 5982 -3498 6016 -3332
rect 6016 -3498 6024 -3332
rect 5972 -3512 6024 -3498
rect 6424 -3122 6476 -3108
rect 6424 -3288 6432 -3122
rect 6432 -3288 6466 -3122
rect 6466 -3288 6476 -3122
rect 6304 -3498 6314 -3332
rect 6314 -3498 6348 -3332
rect 6348 -3498 6356 -3332
rect 6304 -3512 6356 -3498
rect 6660 -3122 6712 -3108
rect 6660 -3288 6668 -3122
rect 6668 -3288 6702 -3122
rect 6702 -3288 6712 -3122
rect 6540 -3498 6550 -3332
rect 6550 -3498 6584 -3332
rect 6584 -3498 6592 -3332
rect 6540 -3512 6592 -3498
rect 6896 -3122 6948 -3108
rect 6896 -3288 6904 -3122
rect 6904 -3288 6938 -3122
rect 6938 -3288 6948 -3122
rect 6776 -3498 6786 -3332
rect 6786 -3498 6820 -3332
rect 6820 -3498 6828 -3332
rect 6776 -3512 6828 -3498
rect 7012 -3498 7022 -3332
rect 7022 -3498 7056 -3332
rect 7056 -3498 7064 -3332
rect 7012 -3512 7064 -3498
rect 7464 -3122 7516 -3108
rect 7464 -3288 7472 -3122
rect 7472 -3288 7506 -3122
rect 7506 -3288 7516 -3122
rect 7344 -3498 7354 -3332
rect 7354 -3498 7388 -3332
rect 7388 -3498 7396 -3332
rect 7344 -3512 7396 -3498
rect 7700 -3122 7752 -3108
rect 7700 -3288 7708 -3122
rect 7708 -3288 7742 -3122
rect 7742 -3288 7752 -3122
rect 7580 -3498 7590 -3332
rect 7590 -3498 7624 -3332
rect 7624 -3498 7632 -3332
rect 7580 -3512 7632 -3498
rect 7936 -3122 7988 -3108
rect 7936 -3288 7944 -3122
rect 7944 -3288 7978 -3122
rect 7978 -3288 7988 -3122
rect 7816 -3498 7826 -3332
rect 7826 -3498 7860 -3332
rect 7860 -3498 7868 -3332
rect 7816 -3512 7868 -3498
rect 8052 -3498 8062 -3332
rect 8062 -3498 8096 -3332
rect 8096 -3498 8104 -3332
rect 8052 -3512 8104 -3498
rect 8504 -3122 8556 -3108
rect 8504 -3288 8512 -3122
rect 8512 -3288 8546 -3122
rect 8546 -3288 8556 -3122
rect 8384 -3498 8394 -3332
rect 8394 -3498 8428 -3332
rect 8428 -3498 8436 -3332
rect 8384 -3512 8436 -3498
rect 8740 -3122 8792 -3108
rect 8740 -3288 8748 -3122
rect 8748 -3288 8782 -3122
rect 8782 -3288 8792 -3122
rect 8620 -3498 8630 -3332
rect 8630 -3498 8664 -3332
rect 8664 -3498 8672 -3332
rect 8620 -3512 8672 -3498
rect 8976 -3122 9028 -3108
rect 8976 -3288 8984 -3122
rect 8984 -3288 9018 -3122
rect 9018 -3288 9028 -3122
rect 8856 -3498 8866 -3332
rect 8866 -3498 8900 -3332
rect 8900 -3498 8908 -3332
rect 8856 -3512 8908 -3498
rect 9092 -3498 9102 -3332
rect 9102 -3498 9136 -3332
rect 9136 -3498 9144 -3332
rect 9092 -3512 9144 -3498
rect 11964 -3122 12016 -3108
rect 11964 -3288 11972 -3122
rect 11972 -3288 12006 -3122
rect 12006 -3288 12016 -3122
rect 11844 -3498 11854 -3332
rect 11854 -3498 11888 -3332
rect 11888 -3498 11896 -3332
rect 11844 -3512 11896 -3498
rect 12200 -3122 12252 -3108
rect 12200 -3288 12208 -3122
rect 12208 -3288 12242 -3122
rect 12242 -3288 12252 -3122
rect 12080 -3498 12090 -3332
rect 12090 -3498 12124 -3332
rect 12124 -3498 12132 -3332
rect 12080 -3512 12132 -3498
rect 12436 -3122 12488 -3108
rect 12436 -3288 12444 -3122
rect 12444 -3288 12478 -3122
rect 12478 -3288 12488 -3122
rect 12316 -3498 12326 -3332
rect 12326 -3498 12360 -3332
rect 12360 -3498 12368 -3332
rect 12316 -3512 12368 -3498
rect 12552 -3498 12562 -3332
rect 12562 -3498 12596 -3332
rect 12596 -3498 12604 -3332
rect 12552 -3512 12604 -3498
rect 13004 -3122 13056 -3108
rect 13004 -3288 13012 -3122
rect 13012 -3288 13046 -3122
rect 13046 -3288 13056 -3122
rect 12884 -3498 12894 -3332
rect 12894 -3498 12928 -3332
rect 12928 -3498 12936 -3332
rect 12884 -3512 12936 -3498
rect 13240 -3122 13292 -3108
rect 13240 -3288 13248 -3122
rect 13248 -3288 13282 -3122
rect 13282 -3288 13292 -3122
rect 13120 -3498 13130 -3332
rect 13130 -3498 13164 -3332
rect 13164 -3498 13172 -3332
rect 13120 -3512 13172 -3498
rect 13476 -3122 13528 -3108
rect 13476 -3288 13484 -3122
rect 13484 -3288 13518 -3122
rect 13518 -3288 13528 -3122
rect 13356 -3498 13366 -3332
rect 13366 -3498 13400 -3332
rect 13400 -3498 13408 -3332
rect 13356 -3512 13408 -3498
rect 13592 -3498 13602 -3332
rect 13602 -3498 13636 -3332
rect 13636 -3498 13644 -3332
rect 13592 -3512 13644 -3498
rect 14044 -3122 14096 -3108
rect 14044 -3288 14052 -3122
rect 14052 -3288 14086 -3122
rect 14086 -3288 14096 -3122
rect 13924 -3498 13934 -3332
rect 13934 -3498 13968 -3332
rect 13968 -3498 13976 -3332
rect 13924 -3512 13976 -3498
rect 14280 -3122 14332 -3108
rect 14280 -3288 14288 -3122
rect 14288 -3288 14322 -3122
rect 14322 -3288 14332 -3122
rect 14160 -3498 14170 -3332
rect 14170 -3498 14204 -3332
rect 14204 -3498 14212 -3332
rect 14160 -3512 14212 -3498
rect 14516 -3122 14568 -3108
rect 14516 -3288 14524 -3122
rect 14524 -3288 14558 -3122
rect 14558 -3288 14568 -3122
rect 14396 -3498 14406 -3332
rect 14406 -3498 14440 -3332
rect 14440 -3498 14448 -3332
rect 14396 -3512 14448 -3498
rect 14632 -3498 14642 -3332
rect 14642 -3498 14676 -3332
rect 14676 -3498 14684 -3332
rect 14632 -3512 14684 -3498
rect 15084 -3122 15136 -3108
rect 15084 -3288 15092 -3122
rect 15092 -3288 15126 -3122
rect 15126 -3288 15136 -3122
rect 14964 -3498 14974 -3332
rect 14974 -3498 15008 -3332
rect 15008 -3498 15016 -3332
rect 14964 -3512 15016 -3498
rect 15320 -3122 15372 -3108
rect 15320 -3288 15328 -3122
rect 15328 -3288 15362 -3122
rect 15362 -3288 15372 -3122
rect 15200 -3498 15210 -3332
rect 15210 -3498 15244 -3332
rect 15244 -3498 15252 -3332
rect 15200 -3512 15252 -3498
rect 15556 -3122 15608 -3108
rect 15556 -3288 15564 -3122
rect 15564 -3288 15598 -3122
rect 15598 -3288 15608 -3122
rect 15436 -3498 15446 -3332
rect 15446 -3498 15480 -3332
rect 15480 -3498 15488 -3332
rect 15436 -3512 15488 -3498
rect 15672 -3498 15682 -3332
rect 15682 -3498 15716 -3332
rect 15716 -3498 15724 -3332
rect 15672 -3512 15724 -3498
rect 16124 -3122 16176 -3108
rect 16124 -3288 16132 -3122
rect 16132 -3288 16166 -3122
rect 16166 -3288 16176 -3122
rect 16004 -3498 16014 -3332
rect 16014 -3498 16048 -3332
rect 16048 -3498 16056 -3332
rect 16004 -3512 16056 -3498
rect 16360 -3122 16412 -3108
rect 16360 -3288 16368 -3122
rect 16368 -3288 16402 -3122
rect 16402 -3288 16412 -3122
rect 16240 -3498 16250 -3332
rect 16250 -3498 16284 -3332
rect 16284 -3498 16292 -3332
rect 16240 -3512 16292 -3498
rect 16596 -3122 16648 -3108
rect 16596 -3288 16604 -3122
rect 16604 -3288 16638 -3122
rect 16638 -3288 16648 -3122
rect 16476 -3498 16486 -3332
rect 16486 -3498 16520 -3332
rect 16520 -3498 16528 -3332
rect 16476 -3512 16528 -3498
rect 16712 -3498 16722 -3332
rect 16722 -3498 16756 -3332
rect 16756 -3498 16764 -3332
rect 16712 -3512 16764 -3498
rect 4924 -3840 5224 -3720
rect 8564 -3840 8864 -3720
rect 12544 -3840 12844 -3720
rect 16184 -3840 16484 -3720
rect -7230 -3982 -6950 -3862
<< metal2 >>
rect -920 6880 15540 7336
rect -1472 6740 -1028 6768
rect -1472 6580 -1440 6740
rect -1080 6580 -1028 6740
rect -1472 6184 -1456 6580
rect -1044 6184 -1028 6580
rect -1472 5212 -1440 6184
rect -1080 5212 -1028 6184
rect -920 5768 -140 6880
rect -52 6720 408 6768
rect -52 6588 0 6720
rect 360 6588 408 6720
rect -52 6192 -28 6588
rect 384 6192 408 6588
rect -1472 4816 -1456 5212
rect -1044 4816 -1028 5212
rect -1472 4804 -1028 4816
rect -944 5744 -124 5768
rect -944 5368 -916 5744
rect -144 5368 -124 5744
rect -944 4372 -124 5368
rect -52 5220 0 6192
rect 360 5220 408 6192
rect -52 4824 -28 5220
rect 384 4824 408 5220
rect -52 4804 408 4824
rect 1328 6740 1772 6768
rect 1328 6580 1360 6740
rect 1720 6580 1772 6740
rect 1328 6184 1344 6580
rect 1756 6184 1772 6580
rect 1328 5212 1360 6184
rect 1720 5212 1772 6184
rect 2748 6720 3208 6768
rect 2748 6588 2800 6720
rect 3160 6588 3208 6720
rect 2748 6192 2772 6588
rect 3184 6192 3208 6588
rect 1328 4816 1344 5212
rect 1756 4816 1772 5212
rect 1328 4804 1772 4816
rect 1856 5744 2676 5768
rect 1856 5368 1884 5744
rect 2656 5368 2676 5744
rect -944 3996 -916 4372
rect -144 3996 -124 4372
rect -944 3608 -124 3996
rect -892 3460 -752 3608
rect -944 3418 -892 3428
rect -700 3460 -560 3608
rect -752 3418 -700 3428
rect -508 3460 -368 3608
rect -560 3418 -508 3428
rect -316 3460 -176 3608
rect -368 3418 -316 3428
rect -176 3418 -124 3428
rect 1856 4372 2676 5368
rect 2748 5220 2800 6192
rect 3160 5220 3208 6192
rect 15080 5780 15540 6880
rect 4520 5550 7260 5560
rect 8160 5550 10900 5560
rect 4520 5540 7324 5550
rect 4520 5468 4864 5540
rect 5264 5468 5884 5540
rect 6284 5468 6924 5540
rect 4572 5292 4712 5468
rect 4520 5274 4572 5284
rect 4764 5320 4864 5468
rect 5264 5320 5288 5468
rect 4764 5292 4904 5320
rect 4712 5274 4764 5284
rect 4956 5292 5096 5320
rect 4904 5274 4956 5284
rect 5148 5292 5288 5320
rect 5096 5274 5148 5284
rect 5340 5292 5480 5468
rect 5288 5274 5340 5284
rect 5532 5292 5672 5468
rect 5480 5274 5532 5284
rect 5724 5292 5864 5468
rect 5672 5274 5724 5284
rect 5916 5292 6056 5320
rect 5864 5274 5916 5284
rect 6108 5292 6248 5320
rect 6056 5274 6108 5284
rect 6300 5292 6440 5468
rect 6248 5274 6300 5284
rect 6492 5292 6632 5468
rect 6440 5274 6492 5284
rect 6684 5292 6824 5468
rect 6632 5274 6684 5284
rect 6876 5320 6924 5468
rect 6876 5292 7016 5320
rect 6824 5274 6876 5284
rect 7068 5292 7208 5320
rect 7016 5274 7068 5284
rect 7260 5310 7324 5320
rect 8004 5540 10900 5550
rect 8404 5468 9024 5540
rect 9424 5468 10044 5540
rect 10444 5468 10900 5540
rect 8004 5310 8160 5320
rect 7208 5274 7260 5284
rect 8212 5292 8352 5320
rect 8160 5274 8212 5284
rect 8404 5292 8544 5468
rect 8352 5274 8404 5284
rect 8596 5292 8736 5468
rect 8544 5274 8596 5284
rect 8788 5292 8928 5468
rect 8736 5274 8788 5284
rect 8980 5320 9024 5468
rect 9424 5320 9504 5468
rect 8980 5292 9120 5320
rect 8928 5274 8980 5284
rect 9172 5292 9312 5320
rect 9120 5274 9172 5284
rect 9364 5292 9504 5320
rect 9312 5274 9364 5284
rect 9556 5292 9696 5468
rect 9504 5274 9556 5284
rect 9748 5292 9888 5468
rect 9696 5274 9748 5284
rect 9940 5320 10044 5468
rect 10444 5320 10464 5468
rect 9940 5292 10080 5320
rect 9888 5274 9940 5284
rect 10132 5292 10272 5320
rect 10080 5274 10132 5284
rect 10324 5292 10464 5320
rect 10272 5274 10324 5284
rect 10516 5292 10656 5468
rect 10464 5274 10516 5284
rect 10708 5292 10848 5468
rect 10656 5274 10708 5284
rect 10848 5274 10900 5284
rect 12140 5550 14880 5560
rect 12140 5540 14944 5550
rect 12140 5468 12484 5540
rect 12884 5468 13504 5540
rect 13904 5468 14544 5540
rect 12192 5292 12332 5468
rect 12140 5274 12192 5284
rect 12384 5320 12484 5468
rect 12884 5320 12908 5468
rect 12384 5292 12524 5320
rect 12332 5274 12384 5284
rect 12576 5292 12716 5320
rect 12524 5274 12576 5284
rect 12768 5292 12908 5320
rect 12716 5274 12768 5284
rect 12960 5292 13100 5468
rect 12908 5274 12960 5284
rect 13152 5292 13292 5468
rect 13100 5274 13152 5284
rect 13344 5292 13484 5468
rect 13292 5274 13344 5284
rect 13536 5292 13676 5320
rect 13484 5274 13536 5284
rect 13728 5292 13868 5320
rect 13676 5274 13728 5284
rect 13920 5292 14060 5468
rect 13868 5274 13920 5284
rect 14112 5292 14252 5468
rect 14060 5274 14112 5284
rect 14304 5292 14444 5468
rect 14252 5274 14304 5284
rect 14496 5320 14544 5468
rect 15780 5550 18520 5560
rect 15080 5410 15540 5420
rect 15624 5540 18520 5550
rect 16024 5468 16644 5540
rect 17044 5468 17664 5540
rect 18064 5468 18520 5540
rect 14496 5292 14636 5320
rect 14444 5274 14496 5284
rect 14688 5292 14828 5320
rect 14636 5274 14688 5284
rect 14880 5310 14944 5320
rect 15624 5310 15780 5320
rect 14828 5274 14880 5284
rect 15832 5292 15972 5320
rect 15780 5274 15832 5284
rect 16024 5292 16164 5468
rect 15972 5274 16024 5284
rect 16216 5292 16356 5468
rect 16164 5274 16216 5284
rect 16408 5292 16548 5468
rect 16356 5274 16408 5284
rect 16600 5320 16644 5468
rect 17044 5320 17124 5468
rect 16600 5292 16740 5320
rect 16548 5274 16600 5284
rect 16792 5292 16932 5320
rect 16740 5274 16792 5284
rect 16984 5292 17124 5320
rect 16932 5274 16984 5284
rect 17176 5292 17316 5468
rect 17124 5274 17176 5284
rect 17368 5292 17508 5468
rect 17316 5274 17368 5284
rect 17560 5320 17664 5468
rect 18064 5320 18084 5468
rect 17560 5292 17700 5320
rect 17508 5274 17560 5284
rect 17752 5292 17892 5320
rect 17700 5274 17752 5284
rect 17944 5292 18084 5320
rect 17892 5274 17944 5284
rect 18136 5292 18276 5468
rect 18084 5274 18136 5284
rect 18328 5292 18468 5468
rect 18276 5274 18328 5284
rect 18468 5274 18520 5284
rect 4424 5248 4476 5258
rect 4420 5230 4424 5240
rect 2748 4824 2772 5220
rect 3184 4824 3208 5220
rect 4304 5220 4424 5230
rect 4616 5248 4668 5258
rect 4476 5220 4616 5240
rect 4808 5248 4860 5258
rect 4668 5220 4808 5240
rect 4744 5064 4808 5220
rect 5000 5248 5052 5258
rect 4860 5064 5000 5240
rect 5192 5248 5244 5258
rect 5052 5064 5192 5240
rect 5384 5248 5436 5258
rect 5244 5064 5384 5240
rect 5576 5248 5628 5258
rect 5436 5200 5576 5240
rect 5768 5248 5820 5258
rect 5628 5200 5768 5240
rect 5960 5248 6012 5258
rect 5820 5064 5960 5240
rect 6152 5248 6204 5258
rect 6012 5064 6152 5240
rect 6344 5248 6396 5258
rect 6204 5064 6344 5240
rect 6536 5248 6588 5258
rect 6396 5200 6536 5240
rect 6728 5248 6780 5258
rect 6588 5200 6728 5240
rect 6920 5248 6972 5258
rect 6780 5200 6920 5240
rect 6396 5064 6424 5200
rect 6824 5064 6920 5200
rect 7112 5248 7164 5258
rect 6972 5064 7112 5240
rect 7304 5248 7356 5258
rect 7164 5064 7304 5240
rect 8064 5248 8116 5258
rect 7356 5200 8064 5240
rect 7356 5064 7464 5200
rect 4744 4980 5384 5064
rect 5784 4980 6424 5064
rect 6824 4980 7464 5064
rect 7864 5064 8064 5200
rect 8256 5248 8308 5258
rect 8116 5064 8256 5240
rect 8448 5248 8500 5258
rect 8308 5064 8448 5240
rect 8640 5248 8692 5258
rect 8500 5220 8640 5240
rect 8832 5248 8884 5258
rect 8692 5220 8832 5240
rect 9024 5248 9076 5258
rect 8884 5220 9024 5240
rect 8500 5064 8504 5220
rect 8904 5064 9024 5220
rect 9216 5248 9268 5258
rect 9076 5064 9216 5240
rect 9408 5248 9460 5258
rect 9268 5064 9408 5240
rect 9600 5248 9652 5258
rect 9460 5220 9600 5240
rect 9792 5248 9844 5258
rect 9652 5220 9792 5240
rect 9984 5248 10036 5258
rect 9844 5220 9984 5240
rect 9460 5064 9544 5220
rect 9944 5064 9984 5220
rect 10176 5248 10228 5258
rect 10036 5064 10176 5240
rect 10368 5248 10420 5258
rect 10228 5064 10368 5240
rect 10560 5248 10612 5258
rect 10420 5064 10560 5240
rect 10752 5248 10804 5258
rect 10612 5220 10752 5240
rect 10944 5248 10996 5258
rect 10804 5220 10944 5240
rect 12044 5248 12096 5258
rect 10996 5064 11004 5240
rect 12040 5230 12044 5240
rect 7864 5000 8504 5064
rect 8904 5000 9544 5064
rect 9944 5000 10584 5064
rect 10984 5000 11004 5064
rect 7864 4980 11004 5000
rect 4304 4972 11004 4980
rect 11924 5220 12044 5230
rect 12236 5248 12288 5258
rect 12096 5220 12236 5240
rect 12428 5248 12480 5258
rect 12288 5220 12428 5240
rect 12364 5064 12428 5220
rect 12620 5248 12672 5258
rect 12480 5064 12620 5240
rect 12812 5248 12864 5258
rect 12672 5064 12812 5240
rect 13004 5248 13056 5258
rect 12864 5064 13004 5240
rect 13196 5248 13248 5258
rect 13056 5200 13196 5240
rect 13388 5248 13440 5258
rect 13248 5200 13388 5240
rect 13580 5248 13632 5258
rect 13440 5064 13580 5240
rect 13772 5248 13824 5258
rect 13632 5064 13772 5240
rect 13964 5248 14016 5258
rect 13824 5064 13964 5240
rect 14156 5248 14208 5258
rect 14016 5200 14156 5240
rect 14348 5248 14400 5258
rect 14208 5200 14348 5240
rect 14540 5248 14592 5258
rect 14400 5200 14540 5240
rect 14016 5064 14044 5200
rect 14444 5064 14540 5200
rect 14732 5248 14784 5258
rect 14592 5064 14732 5240
rect 14924 5248 14976 5258
rect 14784 5064 14924 5240
rect 15684 5248 15736 5258
rect 14976 5200 15684 5240
rect 14976 5064 15084 5200
rect 12364 4980 13004 5064
rect 13404 4980 14044 5064
rect 14444 4980 15084 5064
rect 15484 5064 15684 5200
rect 15876 5248 15928 5258
rect 15736 5064 15876 5240
rect 16068 5248 16120 5258
rect 15928 5064 16068 5240
rect 16260 5248 16312 5258
rect 16120 5220 16260 5240
rect 16452 5248 16504 5258
rect 16312 5220 16452 5240
rect 16644 5248 16696 5258
rect 16504 5220 16644 5240
rect 16120 5064 16124 5220
rect 16524 5064 16644 5220
rect 16836 5248 16888 5258
rect 16696 5064 16836 5240
rect 17028 5248 17080 5258
rect 16888 5064 17028 5240
rect 17220 5248 17272 5258
rect 17080 5220 17220 5240
rect 17412 5248 17464 5258
rect 17272 5220 17412 5240
rect 17604 5248 17656 5258
rect 17464 5220 17604 5240
rect 17080 5064 17164 5220
rect 17564 5064 17604 5220
rect 17796 5248 17848 5258
rect 17656 5064 17796 5240
rect 17988 5248 18040 5258
rect 17848 5064 17988 5240
rect 18180 5248 18232 5258
rect 18040 5064 18180 5240
rect 18372 5248 18424 5258
rect 18232 5220 18372 5240
rect 18564 5248 18616 5258
rect 18424 5220 18564 5240
rect 18616 5064 18624 5240
rect 15484 5000 16124 5064
rect 16524 5000 17164 5064
rect 17564 5000 18204 5064
rect 18604 5000 18624 5064
rect 15484 4980 18624 5000
rect 11924 4972 18624 4980
rect 4304 4970 4744 4972
rect 5384 4970 5784 4972
rect 6424 4970 6824 4972
rect 7464 4970 7864 4972
rect 11924 4970 12364 4972
rect 13004 4970 13404 4972
rect 14044 4970 14444 4972
rect 15084 4970 15484 4972
rect 2748 4804 3208 4824
rect 4520 4930 7260 4940
rect 8160 4930 10900 4940
rect 4520 4920 7324 4930
rect 4520 4848 4864 4920
rect 5264 4848 5884 4920
rect 6284 4848 6924 4920
rect 4572 4672 4712 4848
rect 4520 4654 4572 4664
rect 4764 4700 4864 4848
rect 5264 4700 5288 4848
rect 4764 4672 4904 4700
rect 4712 4654 4764 4664
rect 4956 4672 5096 4700
rect 4904 4654 4956 4664
rect 5148 4672 5288 4700
rect 5096 4654 5148 4664
rect 5340 4672 5480 4848
rect 5288 4654 5340 4664
rect 5532 4672 5672 4848
rect 5480 4654 5532 4664
rect 5724 4672 5864 4848
rect 5672 4654 5724 4664
rect 5916 4672 6056 4700
rect 5864 4654 5916 4664
rect 6108 4672 6248 4700
rect 6056 4654 6108 4664
rect 6300 4672 6440 4848
rect 6248 4654 6300 4664
rect 6492 4672 6632 4848
rect 6440 4654 6492 4664
rect 6684 4672 6824 4848
rect 6632 4654 6684 4664
rect 6876 4700 6924 4848
rect 6876 4672 7016 4700
rect 6824 4654 6876 4664
rect 7068 4672 7208 4700
rect 7016 4654 7068 4664
rect 7260 4690 7324 4700
rect 8004 4920 10900 4930
rect 8404 4848 9024 4920
rect 9424 4848 10044 4920
rect 10444 4848 10900 4920
rect 8004 4690 8160 4700
rect 7208 4654 7260 4664
rect 8212 4672 8352 4700
rect 8160 4654 8212 4664
rect 8404 4672 8544 4848
rect 8352 4654 8404 4664
rect 8596 4672 8736 4848
rect 8544 4654 8596 4664
rect 8788 4672 8928 4848
rect 8736 4654 8788 4664
rect 8980 4700 9024 4848
rect 9424 4700 9504 4848
rect 8980 4672 9120 4700
rect 8928 4654 8980 4664
rect 9172 4672 9312 4700
rect 9120 4654 9172 4664
rect 9364 4672 9504 4700
rect 9312 4654 9364 4664
rect 9556 4672 9696 4848
rect 9504 4654 9556 4664
rect 9748 4672 9888 4848
rect 9696 4654 9748 4664
rect 9940 4700 10044 4848
rect 10444 4700 10464 4848
rect 9940 4672 10080 4700
rect 9888 4654 9940 4664
rect 10132 4672 10272 4700
rect 10080 4654 10132 4664
rect 10324 4672 10464 4700
rect 10272 4654 10324 4664
rect 10516 4672 10656 4848
rect 10464 4654 10516 4664
rect 10708 4672 10848 4848
rect 10656 4654 10708 4664
rect 10848 4654 10900 4664
rect 12140 4930 14880 4940
rect 15780 4930 18520 4940
rect 12140 4920 14944 4930
rect 12140 4848 12484 4920
rect 12884 4848 13504 4920
rect 13904 4848 14544 4920
rect 12192 4672 12332 4848
rect 12140 4654 12192 4664
rect 12384 4700 12484 4848
rect 12884 4700 12908 4848
rect 12384 4672 12524 4700
rect 12332 4654 12384 4664
rect 12576 4672 12716 4700
rect 12524 4654 12576 4664
rect 12768 4672 12908 4700
rect 12716 4654 12768 4664
rect 12960 4672 13100 4848
rect 12908 4654 12960 4664
rect 13152 4672 13292 4848
rect 13100 4654 13152 4664
rect 13344 4672 13484 4848
rect 13292 4654 13344 4664
rect 13536 4672 13676 4700
rect 13484 4654 13536 4664
rect 13728 4672 13868 4700
rect 13676 4654 13728 4664
rect 13920 4672 14060 4848
rect 13868 4654 13920 4664
rect 14112 4672 14252 4848
rect 14060 4654 14112 4664
rect 14304 4672 14444 4848
rect 14252 4654 14304 4664
rect 14496 4700 14544 4848
rect 14496 4672 14636 4700
rect 14444 4654 14496 4664
rect 14688 4672 14828 4700
rect 14636 4654 14688 4664
rect 14880 4690 14944 4700
rect 15624 4920 18520 4930
rect 16024 4848 16644 4920
rect 17044 4848 17664 4920
rect 18064 4848 18520 4920
rect 15624 4690 15780 4700
rect 14828 4654 14880 4664
rect 15832 4672 15972 4700
rect 15780 4654 15832 4664
rect 16024 4672 16164 4848
rect 15972 4654 16024 4664
rect 16216 4672 16356 4848
rect 16164 4654 16216 4664
rect 16408 4672 16548 4848
rect 16356 4654 16408 4664
rect 16600 4700 16644 4848
rect 17044 4700 17124 4848
rect 16600 4672 16740 4700
rect 16548 4654 16600 4664
rect 16792 4672 16932 4700
rect 16740 4654 16792 4664
rect 16984 4672 17124 4700
rect 16932 4654 16984 4664
rect 17176 4672 17316 4848
rect 17124 4654 17176 4664
rect 17368 4672 17508 4848
rect 17316 4654 17368 4664
rect 17560 4700 17664 4848
rect 18064 4700 18084 4848
rect 17560 4672 17700 4700
rect 17508 4654 17560 4664
rect 17752 4672 17892 4700
rect 17700 4654 17752 4664
rect 17944 4672 18084 4700
rect 17892 4654 17944 4664
rect 18136 4672 18276 4848
rect 18084 4654 18136 4664
rect 18328 4672 18468 4848
rect 18276 4654 18328 4664
rect 18468 4654 18520 4664
rect 4424 4628 4476 4638
rect 1856 3996 1884 4372
rect 2656 3996 2676 4372
rect 4304 4600 4424 4610
rect 4616 4628 4668 4638
rect 4476 4600 4616 4620
rect 4808 4628 4860 4638
rect 4668 4600 4808 4620
rect 4744 4444 4808 4600
rect 5000 4628 5052 4638
rect 4860 4444 5000 4620
rect 5192 4628 5244 4638
rect 5052 4444 5192 4620
rect 5384 4628 5436 4638
rect 5244 4444 5384 4620
rect 5576 4628 5628 4638
rect 5436 4600 5576 4620
rect 5768 4628 5820 4638
rect 5628 4600 5768 4620
rect 5960 4628 6012 4638
rect 5820 4444 5960 4620
rect 6152 4628 6204 4638
rect 6012 4444 6152 4620
rect 6344 4628 6396 4638
rect 6204 4444 6344 4620
rect 6536 4628 6588 4638
rect 6396 4600 6536 4620
rect 6728 4628 6780 4638
rect 6588 4600 6728 4620
rect 6920 4628 6972 4638
rect 6780 4600 6920 4620
rect 6396 4444 6424 4600
rect 6824 4444 6920 4600
rect 7112 4628 7164 4638
rect 6972 4444 7112 4620
rect 7304 4628 7356 4638
rect 7164 4444 7304 4620
rect 8064 4628 8116 4638
rect 7356 4600 8064 4620
rect 7356 4444 7464 4600
rect 4744 4380 5384 4444
rect 5784 4380 6424 4444
rect 6824 4380 7464 4444
rect 7864 4444 8064 4600
rect 8256 4628 8308 4638
rect 8116 4444 8256 4620
rect 8448 4628 8500 4638
rect 8308 4444 8448 4620
rect 8640 4628 8692 4638
rect 8500 4600 8640 4620
rect 8832 4628 8884 4638
rect 8692 4600 8832 4620
rect 9024 4628 9076 4638
rect 8884 4600 9024 4620
rect 8500 4444 8504 4600
rect 8904 4444 9024 4600
rect 9216 4628 9268 4638
rect 9076 4444 9216 4620
rect 9408 4628 9460 4638
rect 9268 4444 9408 4620
rect 9600 4628 9652 4638
rect 9460 4600 9600 4620
rect 9792 4628 9844 4638
rect 9652 4600 9792 4620
rect 9984 4628 10036 4638
rect 9844 4600 9984 4620
rect 9460 4444 9544 4600
rect 9944 4444 9984 4600
rect 10176 4628 10228 4638
rect 10036 4444 10176 4620
rect 10368 4628 10420 4638
rect 10228 4444 10368 4620
rect 10560 4628 10612 4638
rect 10420 4444 10560 4620
rect 10752 4628 10804 4638
rect 10612 4600 10752 4620
rect 10944 4628 10996 4638
rect 10804 4600 10944 4620
rect 12044 4628 12096 4638
rect 10996 4444 11004 4620
rect 7864 4380 8504 4444
rect 8904 4380 9544 4444
rect 9944 4380 10584 4444
rect 10984 4380 11004 4444
rect 4304 4370 11004 4380
rect 11924 4600 12044 4610
rect 12236 4628 12288 4638
rect 12096 4600 12236 4620
rect 12428 4628 12480 4638
rect 12288 4600 12428 4620
rect 12364 4444 12428 4600
rect 12620 4628 12672 4638
rect 12480 4444 12620 4620
rect 12812 4628 12864 4638
rect 12672 4444 12812 4620
rect 13004 4628 13056 4638
rect 12864 4444 13004 4620
rect 13196 4628 13248 4638
rect 13056 4600 13196 4620
rect 13388 4628 13440 4638
rect 13248 4600 13388 4620
rect 13580 4628 13632 4638
rect 13440 4444 13580 4620
rect 13772 4628 13824 4638
rect 13632 4444 13772 4620
rect 13964 4628 14016 4638
rect 13824 4444 13964 4620
rect 14156 4628 14208 4638
rect 14016 4600 14156 4620
rect 14348 4628 14400 4638
rect 14208 4600 14348 4620
rect 14540 4628 14592 4638
rect 14400 4600 14540 4620
rect 14016 4444 14044 4600
rect 14444 4444 14540 4600
rect 14732 4628 14784 4638
rect 14592 4444 14732 4620
rect 14924 4628 14976 4638
rect 14784 4444 14924 4620
rect 15684 4628 15736 4638
rect 14976 4600 15684 4620
rect 14976 4444 15084 4600
rect 12364 4380 13004 4444
rect 13404 4380 14044 4444
rect 14444 4380 15084 4444
rect 15484 4444 15684 4600
rect 15876 4628 15928 4638
rect 15736 4444 15876 4620
rect 16068 4628 16120 4638
rect 15928 4444 16068 4620
rect 16260 4628 16312 4638
rect 16120 4600 16260 4620
rect 16452 4628 16504 4638
rect 16312 4600 16452 4620
rect 16644 4628 16696 4638
rect 16504 4600 16644 4620
rect 16120 4444 16124 4600
rect 16524 4444 16644 4600
rect 16836 4628 16888 4638
rect 16696 4444 16836 4620
rect 17028 4628 17080 4638
rect 16888 4444 17028 4620
rect 17220 4628 17272 4638
rect 17080 4600 17220 4620
rect 17412 4628 17464 4638
rect 17272 4600 17412 4620
rect 17604 4628 17656 4638
rect 17464 4600 17604 4620
rect 17080 4444 17164 4600
rect 17564 4444 17604 4600
rect 17796 4628 17848 4638
rect 17656 4444 17796 4620
rect 17988 4628 18040 4638
rect 17848 4444 17988 4620
rect 18180 4628 18232 4638
rect 18040 4444 18180 4620
rect 18372 4628 18424 4638
rect 18232 4600 18372 4620
rect 18564 4628 18616 4638
rect 18424 4600 18564 4620
rect 18616 4444 18624 4620
rect 15484 4380 16124 4444
rect 16524 4380 17164 4444
rect 17564 4380 18204 4444
rect 18604 4380 18624 4444
rect 11924 4370 18624 4380
rect 4424 4352 11004 4370
rect 12044 4352 18624 4370
rect 4520 4310 7260 4324
rect 8160 4310 10900 4324
rect 4520 4300 7324 4310
rect 4520 4232 4864 4300
rect 5264 4232 5884 4300
rect 6284 4232 6924 4300
rect 4572 4056 4712 4232
rect 4520 4038 4572 4048
rect 4764 4080 4864 4232
rect 5264 4080 5288 4232
rect 4764 4056 4904 4080
rect 4712 4038 4764 4048
rect 4956 4056 5096 4080
rect 4904 4038 4956 4048
rect 5148 4056 5288 4080
rect 5096 4038 5148 4048
rect 5340 4056 5480 4232
rect 5288 4038 5340 4048
rect 5532 4056 5672 4232
rect 5480 4038 5532 4048
rect 5724 4056 5864 4232
rect 5672 4038 5724 4048
rect 5916 4056 6056 4080
rect 5864 4038 5916 4048
rect 6108 4056 6248 4080
rect 6056 4038 6108 4048
rect 6300 4056 6440 4232
rect 6248 4038 6300 4048
rect 6492 4056 6632 4232
rect 6440 4038 6492 4048
rect 6684 4056 6824 4232
rect 6632 4038 6684 4048
rect 6876 4080 6924 4232
rect 6876 4056 7016 4080
rect 6824 4038 6876 4048
rect 7068 4056 7208 4080
rect 7016 4038 7068 4048
rect 7260 4070 7324 4080
rect 8004 4300 10900 4310
rect 8404 4232 9024 4300
rect 9424 4232 10044 4300
rect 10444 4232 10900 4300
rect 8004 4070 8160 4080
rect 7208 4038 7260 4048
rect 8212 4056 8352 4080
rect 8160 4038 8212 4048
rect 8404 4056 8544 4232
rect 8352 4038 8404 4048
rect 8596 4056 8736 4232
rect 8544 4038 8596 4048
rect 8788 4056 8928 4232
rect 8736 4038 8788 4048
rect 8980 4080 9024 4232
rect 9424 4080 9504 4232
rect 8980 4056 9120 4080
rect 8928 4038 8980 4048
rect 9172 4056 9312 4080
rect 9120 4038 9172 4048
rect 9364 4056 9504 4080
rect 9312 4038 9364 4048
rect 9556 4056 9696 4232
rect 9504 4038 9556 4048
rect 9748 4056 9888 4232
rect 9696 4038 9748 4048
rect 9940 4080 10044 4232
rect 10444 4080 10464 4232
rect 9940 4056 10080 4080
rect 9888 4038 9940 4048
rect 10132 4056 10272 4080
rect 10080 4038 10132 4048
rect 10324 4056 10464 4080
rect 10272 4038 10324 4048
rect 10516 4056 10656 4232
rect 10464 4038 10516 4048
rect 10708 4056 10848 4232
rect 10656 4038 10708 4048
rect 10848 4038 10900 4048
rect 12140 4310 14880 4324
rect 15780 4310 18520 4324
rect 12140 4300 14944 4310
rect 12140 4232 12484 4300
rect 12884 4232 13504 4300
rect 13904 4232 14544 4300
rect 12192 4056 12332 4232
rect 12140 4038 12192 4048
rect 12384 4080 12484 4232
rect 12884 4080 12908 4232
rect 12384 4056 12524 4080
rect 12332 4038 12384 4048
rect 12576 4056 12716 4080
rect 12524 4038 12576 4048
rect 12768 4056 12908 4080
rect 12716 4038 12768 4048
rect 12960 4056 13100 4232
rect 12908 4038 12960 4048
rect 13152 4056 13292 4232
rect 13100 4038 13152 4048
rect 13344 4056 13484 4232
rect 13292 4038 13344 4048
rect 13536 4056 13676 4080
rect 13484 4038 13536 4048
rect 13728 4056 13868 4080
rect 13676 4038 13728 4048
rect 13920 4056 14060 4232
rect 13868 4038 13920 4048
rect 14112 4056 14252 4232
rect 14060 4038 14112 4048
rect 14304 4056 14444 4232
rect 14252 4038 14304 4048
rect 14496 4080 14544 4232
rect 14496 4056 14636 4080
rect 14444 4038 14496 4048
rect 14688 4056 14828 4080
rect 14636 4038 14688 4048
rect 14880 4070 14944 4080
rect 15624 4300 18520 4310
rect 16024 4232 16644 4300
rect 17044 4232 17664 4300
rect 18064 4232 18520 4300
rect 15624 4070 15780 4080
rect 14828 4038 14880 4048
rect 15832 4056 15972 4080
rect 15780 4038 15832 4048
rect 16024 4056 16164 4232
rect 15972 4038 16024 4048
rect 16216 4056 16356 4232
rect 16164 4038 16216 4048
rect 16408 4056 16548 4232
rect 16356 4038 16408 4048
rect 16600 4080 16644 4232
rect 17044 4080 17124 4232
rect 16600 4056 16740 4080
rect 16548 4038 16600 4048
rect 16792 4056 16932 4080
rect 16740 4038 16792 4048
rect 16984 4056 17124 4080
rect 16932 4038 16984 4048
rect 17176 4056 17316 4232
rect 17124 4038 17176 4048
rect 17368 4056 17508 4232
rect 17316 4038 17368 4048
rect 17560 4080 17664 4232
rect 18064 4080 18084 4232
rect 17560 4056 17700 4080
rect 17508 4038 17560 4048
rect 17752 4056 17892 4080
rect 17700 4038 17752 4048
rect 17944 4056 18084 4080
rect 17892 4038 17944 4048
rect 18136 4056 18276 4232
rect 18084 4038 18136 4048
rect 18328 4056 18468 4232
rect 18276 4038 18328 4048
rect 18468 4038 18520 4048
rect 1856 3608 2676 3996
rect 4424 4012 4476 4022
rect 4304 3980 4424 3990
rect 4616 4012 4668 4022
rect 4476 3980 4616 4008
rect 4808 4012 4860 4022
rect 4668 3980 4808 4008
rect 4744 3828 4808 3980
rect 5000 4012 5052 4022
rect 4860 3828 5000 4008
rect 5192 4012 5244 4022
rect 5052 3828 5192 4008
rect 5384 4012 5436 4022
rect 5244 3828 5384 4008
rect 5576 4012 5628 4022
rect 5436 3980 5576 4008
rect 5768 4012 5820 4022
rect 5628 3980 5768 4008
rect 5960 4012 6012 4022
rect 5820 3828 5960 4008
rect 6152 4012 6204 4022
rect 6012 3828 6152 4008
rect 6344 4012 6396 4022
rect 6204 3828 6344 4008
rect 6536 4012 6588 4022
rect 6396 3980 6536 4008
rect 6728 4012 6780 4022
rect 6588 3980 6728 4008
rect 6920 4012 6972 4022
rect 6780 3980 6920 4008
rect 6396 3828 6424 3980
rect 6824 3828 6920 3980
rect 7112 4012 7164 4022
rect 6972 3828 7112 4008
rect 7304 4012 7356 4022
rect 7164 3828 7304 4008
rect 8064 4012 8116 4022
rect 7356 3980 8064 4008
rect 7356 3828 7464 3980
rect 4744 3760 5384 3828
rect 5784 3760 6424 3828
rect 6824 3760 7464 3828
rect 7864 3828 8064 3980
rect 8256 4012 8308 4022
rect 8116 3828 8256 4008
rect 8448 4012 8500 4022
rect 8308 3828 8448 4008
rect 8640 4012 8692 4022
rect 8500 3980 8640 4008
rect 8832 4012 8884 4022
rect 8692 3980 8832 4008
rect 9024 4012 9076 4022
rect 8884 3980 9024 4008
rect 8500 3828 8504 3980
rect 8904 3828 9024 3980
rect 9216 4012 9268 4022
rect 9076 3828 9216 4008
rect 9408 4012 9460 4022
rect 9268 3828 9408 4008
rect 9600 4012 9652 4022
rect 9460 3980 9600 4008
rect 9792 4012 9844 4022
rect 9652 3980 9792 4008
rect 9984 4012 10036 4022
rect 9844 3980 9984 4008
rect 9460 3828 9544 3980
rect 9944 3828 9984 3980
rect 10176 4012 10228 4022
rect 10036 3828 10176 4008
rect 10368 4012 10420 4022
rect 10228 3828 10368 4008
rect 10560 4012 10612 4022
rect 10420 3828 10560 4008
rect 10752 4012 10804 4022
rect 10612 3980 10752 4008
rect 10944 4012 10996 4022
rect 10804 3980 10944 4008
rect 12044 4012 12096 4022
rect 7864 3760 8504 3828
rect 8904 3760 9544 3828
rect 9944 3760 10584 3828
rect 10984 3760 10996 3828
rect 4304 3750 10996 3760
rect 11924 3980 12044 3990
rect 12236 4012 12288 4022
rect 12096 3980 12236 4008
rect 12428 4012 12480 4022
rect 12288 3980 12428 4008
rect 12364 3828 12428 3980
rect 12620 4012 12672 4022
rect 12480 3828 12620 4008
rect 12812 4012 12864 4022
rect 12672 3828 12812 4008
rect 13004 4012 13056 4022
rect 12864 3828 13004 4008
rect 13196 4012 13248 4022
rect 13056 3980 13196 4008
rect 13388 4012 13440 4022
rect 13248 3980 13388 4008
rect 13580 4012 13632 4022
rect 13440 3828 13580 4008
rect 13772 4012 13824 4022
rect 13632 3828 13772 4008
rect 13964 4012 14016 4022
rect 13824 3828 13964 4008
rect 14156 4012 14208 4022
rect 14016 3980 14156 4008
rect 14348 4012 14400 4022
rect 14208 3980 14348 4008
rect 14540 4012 14592 4022
rect 14400 3980 14540 4008
rect 14016 3828 14044 3980
rect 14444 3828 14540 3980
rect 14732 4012 14784 4022
rect 14592 3828 14732 4008
rect 14924 4012 14976 4022
rect 14784 3828 14924 4008
rect 15684 4012 15736 4022
rect 14976 3980 15684 4008
rect 14976 3828 15084 3980
rect 12364 3760 13004 3828
rect 13404 3760 14044 3828
rect 14444 3760 15084 3828
rect 15484 3828 15684 3980
rect 15876 4012 15928 4022
rect 15736 3828 15876 4008
rect 16068 4012 16120 4022
rect 15928 3828 16068 4008
rect 16260 4012 16312 4022
rect 16120 3980 16260 4008
rect 16452 4012 16504 4022
rect 16312 3980 16452 4008
rect 16644 4012 16696 4022
rect 16504 3980 16644 4008
rect 16120 3828 16124 3980
rect 16524 3828 16644 3980
rect 16836 4012 16888 4022
rect 16696 3828 16836 4008
rect 17028 4012 17080 4022
rect 16888 3828 17028 4008
rect 17220 4012 17272 4022
rect 17080 3980 17220 4008
rect 17412 4012 17464 4022
rect 17272 3980 17412 4008
rect 17604 4012 17656 4022
rect 17464 3980 17604 4008
rect 17080 3828 17164 3980
rect 17564 3828 17604 3980
rect 17796 4012 17848 4022
rect 17656 3828 17796 4008
rect 17988 4012 18040 4022
rect 17848 3828 17988 4008
rect 18180 4012 18232 4022
rect 18040 3828 18180 4008
rect 18372 4012 18424 4022
rect 18232 3980 18372 4008
rect 18564 4012 18616 4022
rect 18424 3980 18564 4008
rect 15484 3760 16124 3828
rect 16524 3760 17164 3828
rect 17564 3760 18204 3828
rect 18604 3760 18616 3828
rect 11924 3750 18616 3760
rect 4424 3740 10996 3750
rect 12044 3740 18616 3750
rect 1908 3460 2048 3608
rect 1856 3418 1908 3428
rect 2100 3460 2240 3608
rect 2048 3418 2100 3428
rect 2292 3460 2432 3608
rect 2240 3418 2292 3428
rect 2484 3460 2624 3608
rect 2432 3418 2484 3428
rect 2624 3418 2676 3428
rect 4520 3690 7260 3704
rect 8160 3690 10900 3704
rect 4520 3680 7324 3690
rect 4520 3612 4864 3680
rect 5264 3612 5884 3680
rect 6284 3612 6924 3680
rect 4572 3436 4712 3612
rect 4520 3418 4572 3428
rect 4764 3460 4864 3612
rect 5264 3460 5288 3612
rect 4764 3436 4904 3460
rect 4712 3418 4764 3428
rect 4956 3436 5096 3460
rect 4904 3418 4956 3428
rect 5148 3436 5288 3460
rect 5096 3418 5148 3428
rect 5340 3436 5480 3612
rect 5288 3418 5340 3428
rect 5532 3436 5672 3612
rect 5480 3418 5532 3428
rect 5724 3436 5864 3612
rect 5672 3418 5724 3428
rect 5916 3436 6056 3460
rect 5864 3418 5916 3428
rect 6108 3436 6248 3460
rect 6056 3418 6108 3428
rect 6300 3436 6440 3612
rect 6248 3418 6300 3428
rect 6492 3436 6632 3612
rect 6440 3418 6492 3428
rect 6684 3436 6824 3612
rect 6632 3418 6684 3428
rect 6876 3460 6924 3612
rect 6876 3436 7016 3460
rect 6824 3418 6876 3428
rect 7068 3436 7208 3460
rect 7016 3418 7068 3428
rect 7260 3450 7324 3460
rect 8004 3680 10900 3690
rect 8404 3612 9024 3680
rect 9424 3612 10044 3680
rect 10444 3612 10900 3680
rect 8004 3450 8160 3460
rect 7208 3418 7260 3428
rect 8212 3436 8352 3460
rect 8160 3418 8212 3428
rect 8404 3436 8544 3612
rect 8352 3418 8404 3428
rect 8596 3436 8736 3612
rect 8544 3418 8596 3428
rect 8788 3436 8928 3612
rect 8736 3418 8788 3428
rect 8980 3460 9024 3612
rect 9424 3460 9504 3612
rect 8980 3436 9120 3460
rect 8928 3418 8980 3428
rect 9172 3436 9312 3460
rect 9120 3418 9172 3428
rect 9364 3436 9504 3460
rect 9312 3418 9364 3428
rect 9556 3436 9696 3612
rect 9504 3418 9556 3428
rect 9748 3436 9888 3612
rect 9696 3418 9748 3428
rect 9940 3460 10044 3612
rect 10444 3460 10464 3612
rect 9940 3436 10080 3460
rect 9888 3418 9940 3428
rect 10132 3436 10272 3460
rect 10080 3418 10132 3428
rect 10324 3436 10464 3460
rect 10272 3418 10324 3428
rect 10516 3436 10656 3612
rect 10464 3418 10516 3428
rect 10708 3436 10848 3612
rect 10656 3418 10708 3428
rect 10848 3418 10900 3428
rect 12140 3690 14880 3704
rect 15780 3690 18520 3704
rect 12140 3680 14944 3690
rect 12140 3612 12484 3680
rect 12884 3612 13504 3680
rect 13904 3612 14544 3680
rect 12192 3436 12332 3612
rect 12140 3418 12192 3428
rect 12384 3460 12484 3612
rect 12884 3460 12908 3612
rect 12384 3436 12524 3460
rect 12332 3418 12384 3428
rect 12576 3436 12716 3460
rect 12524 3418 12576 3428
rect 12768 3436 12908 3460
rect 12716 3418 12768 3428
rect 12960 3436 13100 3612
rect 12908 3418 12960 3428
rect 13152 3436 13292 3612
rect 13100 3418 13152 3428
rect 13344 3436 13484 3612
rect 13292 3418 13344 3428
rect 13536 3436 13676 3460
rect 13484 3418 13536 3428
rect 13728 3436 13868 3460
rect 13676 3418 13728 3428
rect 13920 3436 14060 3612
rect 13868 3418 13920 3428
rect 14112 3436 14252 3612
rect 14060 3418 14112 3428
rect 14304 3436 14444 3612
rect 14252 3418 14304 3428
rect 14496 3460 14544 3612
rect 14496 3436 14636 3460
rect 14444 3418 14496 3428
rect 14688 3436 14828 3460
rect 14636 3418 14688 3428
rect 14880 3450 14944 3460
rect 15624 3680 18520 3690
rect 16024 3612 16644 3680
rect 17044 3612 17664 3680
rect 18064 3612 18520 3680
rect 15624 3450 15780 3460
rect 14828 3418 14880 3428
rect 15832 3436 15972 3460
rect 15780 3418 15832 3428
rect 16024 3436 16164 3612
rect 15972 3418 16024 3428
rect 16216 3436 16356 3612
rect 16164 3418 16216 3428
rect 16408 3436 16548 3612
rect 16356 3418 16408 3428
rect 16600 3460 16644 3612
rect 17044 3460 17124 3612
rect 16600 3436 16740 3460
rect 16548 3418 16600 3428
rect 16792 3436 16932 3460
rect 16740 3418 16792 3428
rect 16984 3436 17124 3460
rect 16932 3418 16984 3428
rect 17176 3436 17316 3612
rect 17124 3418 17176 3428
rect 17368 3436 17508 3612
rect 17316 3418 17368 3428
rect 17560 3460 17664 3612
rect 18064 3460 18084 3612
rect 17560 3436 17700 3460
rect 17508 3418 17560 3428
rect 17752 3436 17892 3460
rect 17700 3418 17752 3428
rect 17944 3436 18084 3460
rect 17892 3418 17944 3428
rect 18136 3436 18276 3612
rect 18084 3418 18136 3428
rect 18328 3436 18468 3612
rect 18276 3418 18328 3428
rect 18468 3418 18520 3428
rect -1040 3392 -988 3402
rect -1100 3290 -1040 3320
rect -1140 3280 -1040 3290
rect -848 3392 -796 3402
rect -988 3280 -848 3364
rect -656 3392 -604 3402
rect -796 3280 -656 3364
rect -464 3392 -412 3402
rect -604 3280 -464 3364
rect -272 3392 -220 3402
rect -412 3280 -272 3364
rect -80 3392 -28 3402
rect -220 3280 -80 3364
rect 1760 3392 1812 3402
rect -28 3280 120 3320
rect 60 2980 120 3280
rect 1620 3280 1760 3320
rect 1952 3392 2004 3402
rect 1812 3280 1952 3364
rect 2144 3392 2196 3402
rect 2004 3280 2144 3364
rect 2336 3392 2388 3402
rect 2196 3280 2336 3364
rect 2528 3392 2580 3402
rect 2388 3280 2528 3364
rect 2720 3392 2772 3402
rect 2580 3280 2720 3364
rect 4424 3392 4476 3402
rect 4304 3360 4424 3370
rect 4616 3392 4668 3402
rect 4476 3360 4616 3384
rect 4808 3392 4860 3402
rect 4668 3360 4808 3384
rect 2772 3280 2860 3320
rect 1620 2980 1660 3280
rect -1140 2770 60 2780
rect 4744 3208 4808 3360
rect 5000 3392 5052 3402
rect 4860 3208 5000 3384
rect 5192 3392 5244 3402
rect 5052 3208 5192 3384
rect 5384 3392 5436 3402
rect 5244 3208 5384 3384
rect 5576 3392 5628 3402
rect 5436 3360 5576 3384
rect 5768 3392 5820 3402
rect 5628 3360 5768 3384
rect 5960 3392 6012 3402
rect 5820 3208 5960 3384
rect 6152 3392 6204 3402
rect 6012 3208 6152 3384
rect 6344 3392 6396 3402
rect 6204 3208 6344 3384
rect 6536 3392 6588 3402
rect 6396 3360 6536 3384
rect 6728 3392 6780 3402
rect 6588 3360 6728 3384
rect 6920 3392 6972 3402
rect 6780 3360 6920 3384
rect 6396 3208 6424 3360
rect 6824 3208 6920 3360
rect 7112 3392 7164 3402
rect 6972 3208 7112 3384
rect 7304 3392 7356 3402
rect 7164 3208 7304 3384
rect 8064 3392 8116 3402
rect 7356 3360 8064 3384
rect 7356 3208 7464 3360
rect 4744 3140 5384 3208
rect 5784 3140 6424 3208
rect 6824 3140 7464 3208
rect 7864 3208 8064 3360
rect 8256 3392 8308 3402
rect 8116 3208 8256 3384
rect 8448 3392 8500 3402
rect 8308 3208 8448 3384
rect 8640 3392 8692 3402
rect 8500 3360 8640 3384
rect 8832 3392 8884 3402
rect 8692 3360 8832 3384
rect 9024 3392 9076 3402
rect 8884 3360 9024 3384
rect 8500 3208 8504 3360
rect 8904 3208 9024 3360
rect 9216 3392 9268 3402
rect 9076 3208 9216 3384
rect 9408 3392 9460 3402
rect 9268 3208 9408 3384
rect 9600 3392 9652 3402
rect 9460 3360 9600 3384
rect 9792 3392 9844 3402
rect 9652 3360 9792 3384
rect 9984 3392 10036 3402
rect 9844 3360 9984 3384
rect 9460 3208 9544 3360
rect 9944 3208 9984 3360
rect 10176 3392 10228 3402
rect 10036 3208 10176 3384
rect 10368 3392 10420 3402
rect 10228 3208 10368 3384
rect 10560 3392 10612 3402
rect 10420 3208 10560 3384
rect 10752 3392 10804 3402
rect 10612 3360 10752 3384
rect 10944 3392 10996 3402
rect 10804 3360 10944 3384
rect 12044 3392 12096 3402
rect 10996 3208 11000 3384
rect 7864 3140 8504 3208
rect 8904 3140 9544 3208
rect 9944 3140 10584 3208
rect 10984 3140 11000 3208
rect 4304 3130 11000 3140
rect 11924 3360 12044 3370
rect 12236 3392 12288 3402
rect 12096 3360 12236 3384
rect 12428 3392 12480 3402
rect 12288 3360 12428 3384
rect 12364 3208 12428 3360
rect 12620 3392 12672 3402
rect 12480 3208 12620 3384
rect 12812 3392 12864 3402
rect 12672 3208 12812 3384
rect 13004 3392 13056 3402
rect 12864 3208 13004 3384
rect 13196 3392 13248 3402
rect 13056 3360 13196 3384
rect 13388 3392 13440 3402
rect 13248 3360 13388 3384
rect 13580 3392 13632 3402
rect 13440 3208 13580 3384
rect 13772 3392 13824 3402
rect 13632 3208 13772 3384
rect 13964 3392 14016 3402
rect 13824 3208 13964 3384
rect 14156 3392 14208 3402
rect 14016 3360 14156 3384
rect 14348 3392 14400 3402
rect 14208 3360 14348 3384
rect 14540 3392 14592 3402
rect 14400 3360 14540 3384
rect 14016 3208 14044 3360
rect 14444 3208 14540 3360
rect 14732 3392 14784 3402
rect 14592 3208 14732 3384
rect 14924 3392 14976 3402
rect 14784 3208 14924 3384
rect 15684 3392 15736 3402
rect 14976 3360 15684 3384
rect 14976 3208 15084 3360
rect 12364 3140 13004 3208
rect 13404 3140 14044 3208
rect 14444 3140 15084 3208
rect 15484 3208 15684 3360
rect 15876 3392 15928 3402
rect 15736 3208 15876 3384
rect 16068 3392 16120 3402
rect 15928 3208 16068 3384
rect 16260 3392 16312 3402
rect 16120 3360 16260 3384
rect 16452 3392 16504 3402
rect 16312 3360 16452 3384
rect 16644 3392 16696 3402
rect 16504 3360 16644 3384
rect 16120 3208 16124 3360
rect 16524 3208 16644 3360
rect 16836 3392 16888 3402
rect 16696 3208 16836 3384
rect 17028 3392 17080 3402
rect 16888 3208 17028 3384
rect 17220 3392 17272 3402
rect 17080 3360 17220 3384
rect 17412 3392 17464 3402
rect 17272 3360 17412 3384
rect 17604 3392 17656 3402
rect 17464 3360 17604 3384
rect 17080 3208 17164 3360
rect 17564 3208 17604 3360
rect 17796 3392 17848 3402
rect 17656 3208 17796 3384
rect 17988 3392 18040 3402
rect 17848 3208 17988 3384
rect 18180 3392 18232 3402
rect 18040 3208 18180 3384
rect 18372 3392 18424 3402
rect 18232 3360 18372 3384
rect 18564 3392 18616 3402
rect 18424 3360 18564 3384
rect 18616 3208 18620 3384
rect 15484 3140 16124 3208
rect 16524 3140 17164 3208
rect 17564 3140 18204 3208
rect 18604 3140 18620 3208
rect 11924 3130 18620 3140
rect 4424 3116 11000 3130
rect 12044 3116 18620 3130
rect 1660 2770 2860 2780
rect 4084 2792 4984 2844
rect -1720 2632 -820 2684
rect -1720 2452 -1580 2632
rect -1528 2460 -1388 2632
rect -1720 2442 -1528 2452
rect -1336 2460 -1196 2632
rect -1388 2442 -1336 2452
rect -1144 2460 -1004 2632
rect -1196 2442 -1144 2452
rect -1012 2452 -1004 2460
rect -952 2452 -820 2632
rect -1720 1804 -1540 2442
rect -1012 2432 -820 2452
rect -1484 2412 -1432 2422
rect -1292 2412 -1240 2422
rect -1432 2372 -1292 2404
rect -1100 2412 -1048 2422
rect -1240 2372 -1100 2404
rect -1092 2016 -1048 2232
rect -1432 1844 -1292 1880
rect -1484 1826 -1432 1836
rect -1240 1844 -1100 1880
rect -1292 1826 -1240 1836
rect -1000 1844 -820 2432
rect -1100 1826 -1048 1836
rect -1720 1796 -1528 1804
rect -1720 1616 -1580 1796
rect -1388 1796 -1336 1806
rect -1528 1616 -1388 1788
rect -1196 1796 -1144 1806
rect -1336 1616 -1196 1788
rect -1012 1796 -820 1844
rect -1012 1788 -1004 1796
rect -1144 1616 -1004 1788
rect -952 1660 -820 1796
rect -680 2632 220 2684
rect -680 2452 -540 2632
rect -488 2460 -348 2632
rect -680 2442 -488 2452
rect -296 2460 -156 2632
rect -348 2442 -296 2452
rect -104 2460 36 2632
rect -156 2442 -104 2452
rect 28 2452 36 2460
rect 88 2452 220 2632
rect -680 1804 -500 2442
rect 28 2432 220 2452
rect -444 2412 -392 2422
rect -252 2412 -200 2422
rect -392 2380 -252 2404
rect -60 2412 -8 2422
rect -200 2380 -60 2404
rect -444 2016 -440 2232
rect -48 2016 -8 2232
rect -392 1844 -252 1888
rect -444 1826 -392 1836
rect -200 1844 -60 1888
rect -252 1826 -200 1836
rect 40 1844 220 2432
rect -60 1826 -8 1836
rect -680 1796 -488 1804
rect -680 1660 -540 1796
rect -952 1616 -540 1660
rect -348 1796 -296 1806
rect -488 1616 -348 1788
rect -156 1796 -104 1806
rect -296 1616 -156 1788
rect 28 1796 220 1844
rect 28 1788 36 1796
rect -104 1616 36 1788
rect 88 1660 220 1796
rect 360 2632 1260 2684
rect 360 2452 500 2632
rect 552 2460 692 2632
rect 360 2442 552 2452
rect 744 2460 884 2632
rect 692 2442 744 2452
rect 936 2460 1076 2632
rect 884 2442 936 2452
rect 1068 2452 1076 2460
rect 1128 2452 1260 2632
rect 360 1804 540 2442
rect 1068 2432 1260 2452
rect 596 2412 648 2422
rect 788 2412 840 2422
rect 648 2376 788 2404
rect 980 2412 1032 2422
rect 840 2376 980 2404
rect 596 2016 604 2232
rect 996 2016 1032 2232
rect 648 1844 788 1884
rect 596 1826 648 1836
rect 840 1844 980 1884
rect 788 1826 840 1836
rect 1080 1844 1260 2432
rect 980 1826 1032 1836
rect 360 1796 552 1804
rect 360 1660 500 1796
rect 88 1616 500 1660
rect 692 1796 744 1806
rect 552 1616 692 1788
rect 884 1796 936 1806
rect 744 1616 884 1788
rect 1068 1796 1260 1844
rect 1068 1788 1076 1796
rect 936 1616 1076 1788
rect 1128 1660 1260 1796
rect 1400 2632 2300 2684
rect 1400 2452 1540 2632
rect 1592 2460 1732 2632
rect 1400 2442 1592 2452
rect 1784 2460 1924 2632
rect 1732 2442 1784 2452
rect 1976 2460 2116 2632
rect 1924 2442 1976 2452
rect 2108 2452 2116 2460
rect 2168 2452 2300 2632
rect 1400 1804 1580 2442
rect 2108 2432 2300 2452
rect 1636 2412 1688 2422
rect 1828 2412 1880 2422
rect 1688 2372 1828 2404
rect 2020 2412 2072 2422
rect 1880 2372 2020 2404
rect 1636 2016 1648 2232
rect 2040 2016 2072 2232
rect 1688 1844 1828 1880
rect 1636 1826 1688 1836
rect 1880 1844 2020 1880
rect 1828 1826 1880 1836
rect 2120 1844 2300 2432
rect 2020 1826 2072 1836
rect 1400 1796 1592 1804
rect 1400 1660 1540 1796
rect 1128 1616 1540 1660
rect 1732 1796 1784 1806
rect 1592 1616 1732 1788
rect 1924 1796 1976 1806
rect 1784 1616 1924 1788
rect 2108 1796 2300 1844
rect 2108 1788 2116 1796
rect 1976 1616 2116 1788
rect 2168 1660 2300 1796
rect 2440 2632 3340 2684
rect 2440 2452 2580 2632
rect 2632 2460 2772 2632
rect 2440 2442 2632 2452
rect 2824 2460 2964 2632
rect 2772 2442 2824 2452
rect 3016 2460 3156 2632
rect 2964 2442 3016 2452
rect 3148 2452 3156 2460
rect 3208 2452 3340 2632
rect 2440 1804 2620 2442
rect 3148 2432 3340 2452
rect 2676 2412 2728 2422
rect 2868 2412 2920 2422
rect 2728 2372 2868 2404
rect 3060 2412 3112 2422
rect 2920 2372 3060 2404
rect 2676 2016 2704 2232
rect 3096 2016 3112 2232
rect 2728 1844 2868 1880
rect 2676 1826 2728 1836
rect 2920 1844 3060 1880
rect 2868 1826 2920 1836
rect 3160 1844 3340 2432
rect 3060 1826 3112 1836
rect 2440 1796 2632 1804
rect 2440 1660 2580 1796
rect 2168 1616 2580 1660
rect 2772 1796 2824 1806
rect 2632 1616 2772 1788
rect 2964 1796 3016 1806
rect 2824 1616 2964 1788
rect 3148 1796 3340 1844
rect 4084 2612 4224 2792
rect 4276 2620 4416 2792
rect 4084 2602 4276 2612
rect 4468 2620 4608 2792
rect 4416 2602 4468 2612
rect 4660 2620 4800 2792
rect 4608 2602 4660 2612
rect 4792 2612 4800 2620
rect 4852 2612 4984 2792
rect 4084 1964 4264 2602
rect 4792 2592 4984 2612
rect 4320 2572 4372 2582
rect 4512 2572 4564 2582
rect 4372 2550 4512 2564
rect 4704 2572 4756 2582
rect 4564 2550 4704 2564
rect 4320 2176 4328 2392
rect 4748 2176 4756 2392
rect 4372 2004 4512 2016
rect 4320 1986 4372 1996
rect 4564 2004 4704 2016
rect 4512 1986 4564 1996
rect 4804 2004 4984 2592
rect 4704 1986 4756 1996
rect 4084 1956 4276 1964
rect 4084 1808 4224 1956
rect 3148 1788 3156 1796
rect 3016 1616 3156 1788
rect 3208 1616 3340 1796
rect -1720 1504 3340 1616
rect 4000 1776 4224 1808
rect 4416 1956 4468 1966
rect 4276 1776 4416 1948
rect 4608 1956 4660 1966
rect 4468 1776 4608 1948
rect 4792 1956 4984 2004
rect 4792 1948 4800 1956
rect 4660 1776 4800 1948
rect 4852 1808 4984 1956
rect 5124 2792 6024 2844
rect 5124 2612 5264 2792
rect 5316 2620 5456 2792
rect 5124 2602 5316 2612
rect 5508 2620 5648 2792
rect 5456 2602 5508 2612
rect 5700 2620 5840 2792
rect 5648 2602 5700 2612
rect 5832 2612 5840 2620
rect 5892 2612 6024 2792
rect 5124 1964 5304 2602
rect 5832 2592 6024 2612
rect 5360 2572 5412 2582
rect 5552 2572 5604 2582
rect 5412 2550 5552 2564
rect 5744 2572 5796 2582
rect 5604 2550 5744 2564
rect 5360 2176 5368 2392
rect 5788 2176 5796 2392
rect 5412 2004 5552 2016
rect 5360 1986 5412 1996
rect 5604 2004 5744 2016
rect 5552 1986 5604 1996
rect 5844 2004 6024 2592
rect 5744 1986 5796 1996
rect 5124 1956 5316 1964
rect 5124 1808 5264 1956
rect 4852 1776 5264 1808
rect 5456 1956 5508 1966
rect 5316 1776 5456 1948
rect 5648 1956 5700 1966
rect 5508 1776 5648 1948
rect 5832 1956 6024 2004
rect 5832 1948 5840 1956
rect 5700 1776 5840 1948
rect 5892 1808 6024 1956
rect 6164 2792 7064 2844
rect 6164 2612 6304 2792
rect 6356 2620 6496 2792
rect 6164 2602 6356 2612
rect 6548 2620 6688 2792
rect 6496 2602 6548 2612
rect 6740 2620 6880 2792
rect 6688 2602 6740 2612
rect 6872 2612 6880 2620
rect 6932 2612 7064 2792
rect 6164 1964 6344 2602
rect 6872 2592 7064 2612
rect 6400 2572 6452 2582
rect 6592 2572 6644 2582
rect 6452 2550 6592 2564
rect 6784 2572 6836 2582
rect 6644 2550 6784 2564
rect 6400 2176 6408 2392
rect 6828 2176 6836 2392
rect 6452 2004 6592 2016
rect 6400 1986 6452 1996
rect 6644 2004 6784 2016
rect 6592 1986 6644 1996
rect 6884 2004 7064 2592
rect 6784 1986 6836 1996
rect 6164 1956 6356 1964
rect 6164 1808 6304 1956
rect 5892 1776 6304 1808
rect 6496 1956 6548 1966
rect 6356 1776 6496 1948
rect 6688 1956 6740 1966
rect 6548 1776 6688 1948
rect 6872 1956 7064 2004
rect 6872 1948 6880 1956
rect 6740 1776 6880 1948
rect 6932 1808 7064 1956
rect 7204 2792 8104 2844
rect 7204 2612 7344 2792
rect 7396 2620 7536 2792
rect 7204 2602 7396 2612
rect 7588 2620 7728 2792
rect 7536 2602 7588 2612
rect 7780 2620 7920 2792
rect 7728 2602 7780 2612
rect 7912 2612 7920 2620
rect 7972 2612 8104 2792
rect 7204 1964 7384 2602
rect 7912 2592 8104 2612
rect 7440 2572 7492 2582
rect 7632 2572 7684 2582
rect 7492 2550 7632 2564
rect 7824 2572 7876 2582
rect 7684 2550 7824 2564
rect 7440 2176 7448 2392
rect 7868 2176 7876 2392
rect 7492 2004 7632 2016
rect 7440 1986 7492 1996
rect 7684 2004 7824 2016
rect 7632 1986 7684 1996
rect 7924 2004 8104 2592
rect 7824 1986 7876 1996
rect 7204 1956 7396 1964
rect 7204 1808 7344 1956
rect 6932 1776 7344 1808
rect 7536 1956 7588 1966
rect 7396 1776 7536 1948
rect 7728 1956 7780 1966
rect 7588 1776 7728 1948
rect 7912 1956 8104 2004
rect 7912 1948 7920 1956
rect 7780 1776 7920 1948
rect 7972 1808 8104 1956
rect 8244 2792 9144 2844
rect 8244 2612 8384 2792
rect 8436 2620 8576 2792
rect 8244 2602 8436 2612
rect 8628 2620 8768 2792
rect 8576 2602 8628 2612
rect 8820 2620 8960 2792
rect 8768 2602 8820 2612
rect 8952 2612 8960 2620
rect 9012 2612 9144 2792
rect 8244 1964 8424 2602
rect 8952 2592 9144 2612
rect 8480 2572 8532 2582
rect 8672 2572 8724 2582
rect 8532 2546 8672 2564
rect 8864 2572 8916 2582
rect 8724 2546 8864 2564
rect 8480 2176 8488 2392
rect 8908 2176 8916 2392
rect 8532 2002 8672 2012
rect 8480 1986 8532 1996
rect 8724 2002 8864 2012
rect 8672 1986 8724 1996
rect 8964 2004 9144 2592
rect 8864 1986 8916 1996
rect 8244 1956 8436 1964
rect 8244 1808 8384 1956
rect 7972 1776 8384 1808
rect 8576 1956 8628 1966
rect 8436 1776 8576 1948
rect 8768 1956 8820 1966
rect 8628 1776 8768 1948
rect 8952 1956 9144 2004
rect 8952 1948 8960 1956
rect 8820 1776 8960 1948
rect 9012 1808 9144 1956
rect 9284 2792 10184 2844
rect 9284 2612 9424 2792
rect 9476 2620 9616 2792
rect 9284 2602 9476 2612
rect 9668 2620 9808 2792
rect 9616 2602 9668 2612
rect 9860 2620 10000 2792
rect 9808 2602 9860 2612
rect 9992 2612 10000 2620
rect 10052 2612 10184 2792
rect 9284 1964 9464 2602
rect 9992 2592 10184 2612
rect 9520 2572 9572 2582
rect 9712 2572 9764 2582
rect 9572 2550 9712 2564
rect 9904 2572 9956 2582
rect 9764 2550 9904 2564
rect 9520 2176 9528 2392
rect 9948 2176 9956 2392
rect 9572 2004 9712 2016
rect 9520 1986 9572 1996
rect 9764 2004 9904 2016
rect 9712 1986 9764 1996
rect 10004 2004 10184 2592
rect 9904 1986 9956 1996
rect 9284 1956 9476 1964
rect 9284 1808 9424 1956
rect 9012 1776 9424 1808
rect 9616 1956 9668 1966
rect 9476 1776 9616 1948
rect 9808 1956 9860 1966
rect 9668 1776 9808 1948
rect 9992 1956 10184 2004
rect 9992 1948 10000 1956
rect 9860 1776 10000 1948
rect 10052 1808 10184 1956
rect 10324 2792 11224 2844
rect 10324 2612 10464 2792
rect 10516 2620 10656 2792
rect 10324 2602 10516 2612
rect 10708 2620 10848 2792
rect 10656 2602 10708 2612
rect 10900 2620 11040 2792
rect 10848 2602 10900 2612
rect 11032 2612 11040 2620
rect 11092 2612 11224 2792
rect 10324 1964 10504 2602
rect 11032 2592 11224 2612
rect 10560 2572 10612 2582
rect 10752 2572 10804 2582
rect 10612 2546 10752 2564
rect 10944 2572 10996 2582
rect 10804 2546 10944 2564
rect 10560 2176 10568 2392
rect 10988 2176 10996 2392
rect 10612 2002 10752 2012
rect 10560 1986 10612 1996
rect 10804 2002 10944 2012
rect 10752 1986 10804 1996
rect 11044 2004 11224 2592
rect 10944 1986 10996 1996
rect 10324 1956 10516 1964
rect 10324 1808 10464 1956
rect 10052 1776 10464 1808
rect 10656 1956 10708 1966
rect 10516 1776 10656 1948
rect 10848 1956 10900 1966
rect 10708 1776 10848 1948
rect 11032 1956 11224 2004
rect 11032 1948 11040 1956
rect 10900 1776 11040 1948
rect 11092 1808 11224 1956
rect 11704 2792 12604 2844
rect 11704 2612 11844 2792
rect 11896 2620 12036 2792
rect 11704 2602 11896 2612
rect 12088 2620 12228 2792
rect 12036 2602 12088 2612
rect 12280 2620 12420 2792
rect 12228 2602 12280 2612
rect 12412 2612 12420 2620
rect 12472 2612 12604 2792
rect 11704 1964 11884 2602
rect 12412 2592 12604 2612
rect 11940 2572 11992 2582
rect 12132 2572 12184 2582
rect 11992 2550 12132 2564
rect 12324 2572 12376 2582
rect 12184 2550 12324 2564
rect 11940 2176 11948 2392
rect 12368 2176 12376 2392
rect 11992 2004 12132 2016
rect 11940 1986 11992 1996
rect 12184 2004 12324 2016
rect 12132 1986 12184 1996
rect 12424 2004 12604 2592
rect 12324 1986 12376 1996
rect 11704 1956 11896 1964
rect 11704 1808 11844 1956
rect 11092 1776 11316 1808
rect 4000 1664 11316 1776
rect 11620 1776 11844 1808
rect 12036 1956 12088 1966
rect 11896 1776 12036 1948
rect 12228 1956 12280 1966
rect 12088 1776 12228 1948
rect 12412 1956 12604 2004
rect 12412 1948 12420 1956
rect 12280 1776 12420 1948
rect 12472 1808 12604 1956
rect 12744 2792 13644 2844
rect 12744 2612 12884 2792
rect 12936 2620 13076 2792
rect 12744 2602 12936 2612
rect 13128 2620 13268 2792
rect 13076 2602 13128 2612
rect 13320 2620 13460 2792
rect 13268 2602 13320 2612
rect 13452 2612 13460 2620
rect 13512 2612 13644 2792
rect 12744 1964 12924 2602
rect 13452 2592 13644 2612
rect 12980 2572 13032 2582
rect 13172 2572 13224 2582
rect 13032 2550 13172 2564
rect 13364 2572 13416 2582
rect 13224 2550 13364 2564
rect 12980 2176 12988 2392
rect 13408 2176 13416 2392
rect 13032 2004 13172 2016
rect 12980 1986 13032 1996
rect 13224 2004 13364 2016
rect 13172 1986 13224 1996
rect 13464 2004 13644 2592
rect 13364 1986 13416 1996
rect 12744 1956 12936 1964
rect 12744 1808 12884 1956
rect 12472 1776 12884 1808
rect 13076 1956 13128 1966
rect 12936 1776 13076 1948
rect 13268 1956 13320 1966
rect 13128 1776 13268 1948
rect 13452 1956 13644 2004
rect 13452 1948 13460 1956
rect 13320 1776 13460 1948
rect 13512 1808 13644 1956
rect 13784 2792 14684 2844
rect 13784 2612 13924 2792
rect 13976 2620 14116 2792
rect 13784 2602 13976 2612
rect 14168 2620 14308 2792
rect 14116 2602 14168 2612
rect 14360 2620 14500 2792
rect 14308 2602 14360 2612
rect 14492 2612 14500 2620
rect 14552 2612 14684 2792
rect 13784 1964 13964 2602
rect 14492 2592 14684 2612
rect 14020 2572 14072 2582
rect 14212 2572 14264 2582
rect 14072 2550 14212 2564
rect 14404 2572 14456 2582
rect 14264 2550 14404 2564
rect 14020 2176 14028 2392
rect 14448 2176 14456 2392
rect 14072 2004 14212 2016
rect 14020 1986 14072 1996
rect 14264 2004 14404 2016
rect 14212 1986 14264 1996
rect 14504 2004 14684 2592
rect 14404 1986 14456 1996
rect 13784 1956 13976 1964
rect 13784 1808 13924 1956
rect 13512 1776 13924 1808
rect 14116 1956 14168 1966
rect 13976 1776 14116 1948
rect 14308 1956 14360 1966
rect 14168 1776 14308 1948
rect 14492 1956 14684 2004
rect 14492 1948 14500 1956
rect 14360 1776 14500 1948
rect 14552 1808 14684 1956
rect 14824 2792 15724 2844
rect 14824 2612 14964 2792
rect 15016 2620 15156 2792
rect 14824 2602 15016 2612
rect 15208 2620 15348 2792
rect 15156 2602 15208 2612
rect 15400 2620 15540 2792
rect 15348 2602 15400 2612
rect 15532 2612 15540 2620
rect 15592 2612 15724 2792
rect 14824 1964 15004 2602
rect 15532 2592 15724 2612
rect 15060 2572 15112 2582
rect 15252 2572 15304 2582
rect 15112 2550 15252 2564
rect 15444 2572 15496 2582
rect 15304 2550 15444 2564
rect 15060 2176 15068 2392
rect 15488 2176 15496 2392
rect 15112 2004 15252 2016
rect 15060 1986 15112 1996
rect 15304 2004 15444 2016
rect 15252 1986 15304 1996
rect 15544 2004 15724 2592
rect 15444 1986 15496 1996
rect 14824 1956 15016 1964
rect 14824 1808 14964 1956
rect 14552 1776 14964 1808
rect 15156 1956 15208 1966
rect 15016 1776 15156 1948
rect 15348 1956 15400 1966
rect 15208 1776 15348 1948
rect 15532 1956 15724 2004
rect 15532 1948 15540 1956
rect 15400 1776 15540 1948
rect 15592 1808 15724 1956
rect 15864 2792 16764 2844
rect 15864 2612 16004 2792
rect 16056 2620 16196 2792
rect 15864 2602 16056 2612
rect 16248 2620 16388 2792
rect 16196 2602 16248 2612
rect 16440 2620 16580 2792
rect 16388 2602 16440 2612
rect 16572 2612 16580 2620
rect 16632 2612 16764 2792
rect 15864 1964 16044 2602
rect 16572 2592 16764 2612
rect 16100 2572 16152 2582
rect 16292 2572 16344 2582
rect 16152 2546 16292 2564
rect 16484 2572 16536 2582
rect 16344 2546 16484 2564
rect 16100 2176 16108 2392
rect 16528 2176 16536 2392
rect 16152 2002 16292 2012
rect 16100 1986 16152 1996
rect 16344 2002 16484 2012
rect 16292 1986 16344 1996
rect 16584 2004 16764 2592
rect 16484 1986 16536 1996
rect 15864 1956 16056 1964
rect 15864 1808 16004 1956
rect 15592 1776 16004 1808
rect 16196 1956 16248 1966
rect 16056 1776 16196 1948
rect 16388 1956 16440 1966
rect 16248 1776 16388 1948
rect 16572 1956 16764 2004
rect 16572 1948 16580 1956
rect 16440 1776 16580 1948
rect 16632 1808 16764 1956
rect 16904 2792 17804 2844
rect 16904 2612 17044 2792
rect 17096 2620 17236 2792
rect 16904 2602 17096 2612
rect 17288 2620 17428 2792
rect 17236 2602 17288 2612
rect 17480 2620 17620 2792
rect 17428 2602 17480 2612
rect 17612 2612 17620 2620
rect 17672 2612 17804 2792
rect 16904 1964 17084 2602
rect 17612 2592 17804 2612
rect 17140 2572 17192 2582
rect 17332 2572 17384 2582
rect 17192 2550 17332 2564
rect 17524 2572 17576 2582
rect 17384 2550 17524 2564
rect 17140 2176 17148 2392
rect 17568 2176 17576 2392
rect 17192 2004 17332 2016
rect 17140 1986 17192 1996
rect 17384 2004 17524 2016
rect 17332 1986 17384 1996
rect 17624 2004 17804 2592
rect 17524 1986 17576 1996
rect 16904 1956 17096 1964
rect 16904 1808 17044 1956
rect 16632 1776 17044 1808
rect 17236 1956 17288 1966
rect 17096 1776 17236 1948
rect 17428 1956 17480 1966
rect 17288 1776 17428 1948
rect 17612 1956 17804 2004
rect 17612 1948 17620 1956
rect 17480 1776 17620 1948
rect 17672 1808 17804 1956
rect 17944 2792 18844 2844
rect 17944 2612 18084 2792
rect 18136 2620 18276 2792
rect 17944 2602 18136 2612
rect 18328 2620 18468 2792
rect 18276 2602 18328 2612
rect 18520 2620 18660 2792
rect 18468 2602 18520 2612
rect 18652 2612 18660 2620
rect 18712 2612 18844 2792
rect 17944 1964 18124 2602
rect 18652 2592 18844 2612
rect 18180 2572 18232 2582
rect 18372 2572 18424 2582
rect 18232 2546 18372 2564
rect 18564 2572 18616 2582
rect 18424 2546 18564 2564
rect 18180 2176 18188 2392
rect 18608 2176 18616 2392
rect 18232 2002 18372 2012
rect 18180 1986 18232 1996
rect 18424 2002 18564 2012
rect 18372 1986 18424 1996
rect 18664 2004 18844 2592
rect 18564 1986 18616 1996
rect 17944 1956 18136 1964
rect 17944 1808 18084 1956
rect 17672 1776 18084 1808
rect 18276 1956 18328 1966
rect 18136 1776 18276 1948
rect 18468 1956 18520 1966
rect 18328 1776 18468 1948
rect 18652 1956 18844 2004
rect 18652 1948 18660 1956
rect 18520 1776 18660 1948
rect 18712 1808 18844 1956
rect 18712 1776 18936 1808
rect 11620 1664 18936 1776
rect -1460 1500 2540 1504
rect -1460 1212 -920 1500
rect -1408 1044 -1224 1212
rect -1460 1022 -1408 1032
rect -1172 1044 -988 1212
rect -1224 1022 -1172 1032
rect -936 1044 -920 1212
rect -420 1212 120 1500
rect -988 1022 -936 1032
rect -368 1044 -184 1212
rect -420 1022 -368 1032
rect -132 1044 52 1212
rect -184 1022 -132 1032
rect 104 1044 120 1212
rect 620 1212 1160 1500
rect 52 1022 104 1032
rect 672 1044 856 1212
rect 620 1022 672 1032
rect 908 1044 1092 1212
rect 856 1022 908 1032
rect 1144 1044 1160 1212
rect 1660 1212 2200 1500
rect 1092 1022 1144 1032
rect 1712 1044 1896 1212
rect 1660 1022 1712 1032
rect 1948 1044 2132 1212
rect 1896 1022 1948 1032
rect 2184 1044 2200 1212
rect 2700 1212 3240 1504
rect 2132 1022 2184 1032
rect 2752 1044 2936 1212
rect 2700 1022 2752 1032
rect 2988 1044 3172 1212
rect 2936 1022 2988 1032
rect 3224 1044 3240 1212
rect 3172 1022 3224 1032
rect -1580 988 -1528 998
rect -1344 988 -1292 998
rect -1528 920 -1344 980
rect -1108 988 -1056 998
rect -1292 920 -1108 980
rect -872 988 -820 998
rect -1056 920 -872 980
rect -1580 440 -1540 808
rect -860 440 -820 808
rect -5998 406 -5802 416
rect -1580 412 -1308 440
rect -1128 412 -820 440
rect -1580 400 -820 412
rect -540 988 -488 998
rect -304 988 -252 998
rect -488 920 -304 980
rect -68 988 -16 998
rect -252 920 -68 980
rect 168 988 220 998
rect -16 920 168 980
rect -540 440 -500 808
rect 180 440 220 808
rect -540 400 220 440
rect 500 988 552 998
rect 736 988 788 998
rect 552 920 736 980
rect 972 988 1024 998
rect 788 920 972 980
rect 1208 988 1260 998
rect 1024 920 1208 980
rect 500 440 540 808
rect 1220 440 1260 808
rect 500 400 1260 440
rect 1540 988 1592 998
rect 1776 988 1828 998
rect 1592 920 1776 980
rect 2012 988 2064 998
rect 1828 920 2012 980
rect 2248 988 2300 998
rect 2064 920 2248 980
rect 1540 440 1580 808
rect 2260 440 2300 808
rect 1540 400 2300 440
rect 2580 988 2632 998
rect 2816 988 2868 998
rect 2632 920 2816 980
rect 3052 988 3104 998
rect 2868 920 3052 980
rect 3288 988 3340 998
rect 3104 920 3288 980
rect 2580 440 2620 808
rect 3300 440 3340 808
rect 2580 408 2800 440
rect 3068 408 3340 440
rect 2580 400 3340 408
rect 4000 604 4156 1664
rect 4344 1372 4884 1664
rect 4396 1204 4580 1372
rect 4344 1182 4396 1192
rect 4632 1204 4816 1372
rect 4580 1182 4632 1192
rect 4868 1204 4884 1372
rect 5384 1372 5924 1664
rect 4816 1182 4868 1192
rect 5436 1204 5620 1372
rect 5384 1182 5436 1192
rect 5672 1204 5856 1372
rect 5620 1182 5672 1192
rect 5908 1204 5924 1372
rect 6424 1372 6964 1664
rect 5856 1182 5908 1192
rect 6476 1204 6660 1372
rect 6424 1182 6476 1192
rect 6712 1204 6896 1372
rect 6660 1182 6712 1192
rect 6948 1204 6964 1372
rect 7464 1372 8004 1664
rect 6896 1182 6948 1192
rect 7516 1204 7700 1372
rect 7464 1182 7516 1192
rect 7752 1204 7936 1372
rect 7700 1182 7752 1192
rect 7988 1204 8004 1372
rect 8504 1372 9044 1664
rect 7936 1182 7988 1192
rect 8556 1204 8740 1372
rect 8504 1182 8556 1192
rect 8792 1204 8976 1372
rect 8740 1182 8792 1192
rect 9028 1204 9044 1372
rect 9544 1372 10084 1664
rect 8976 1182 9028 1192
rect 9596 1204 9780 1372
rect 9544 1182 9596 1192
rect 9832 1204 10016 1372
rect 9780 1182 9832 1192
rect 10068 1204 10084 1372
rect 10584 1372 11124 1664
rect 10016 1182 10068 1192
rect 10636 1204 10820 1372
rect 10584 1182 10636 1192
rect 10872 1204 11056 1372
rect 10820 1182 10872 1192
rect 11108 1204 11124 1372
rect 11056 1182 11108 1192
rect 4224 1148 4276 1158
rect 4460 1148 4512 1158
rect 4276 968 4460 1140
rect 4696 1148 4748 1158
rect 4512 968 4696 1140
rect 4932 1148 4984 1158
rect 4748 1120 4932 1140
rect 5264 1148 5316 1158
rect 4984 1120 5264 1130
rect 4748 968 4864 1120
rect 5500 1148 5552 1158
rect 5316 968 5500 1140
rect 5736 1148 5788 1158
rect 5552 968 5736 1140
rect 5972 1148 6024 1158
rect 5788 1120 5972 1140
rect 6304 1148 6356 1158
rect 6024 1120 6304 1130
rect 6540 1148 6592 1158
rect 5788 968 5904 1120
rect 6356 968 6540 1140
rect 6776 1148 6828 1158
rect 6592 968 6776 1140
rect 7012 1148 7064 1158
rect 6828 1120 7012 1140
rect 7344 1148 7396 1158
rect 7064 1120 7344 1130
rect 6828 968 6924 1120
rect 7580 1148 7632 1158
rect 7396 968 7580 1140
rect 7816 1148 7868 1158
rect 7632 968 7816 1140
rect 8052 1148 8104 1158
rect 7868 1120 8052 1140
rect 8384 1148 8436 1158
rect 8104 1120 8384 1130
rect 8620 1148 8672 1158
rect 7868 968 7984 1120
rect 8436 968 8620 1140
rect 8856 1148 8908 1158
rect 8672 968 8856 1140
rect 9092 1148 9144 1158
rect 8908 1120 9092 1140
rect 9424 1148 9476 1158
rect 9144 1120 9424 1130
rect 9660 1148 9712 1158
rect 8908 968 9024 1120
rect 9476 968 9660 1140
rect 9896 1148 9948 1158
rect 9712 968 9896 1140
rect 10132 1148 10184 1158
rect 9948 1120 10132 1140
rect 10464 1148 10516 1158
rect 10184 1120 10464 1130
rect 9948 968 10044 1120
rect 10700 1148 10752 1158
rect 10516 968 10700 1140
rect 10936 1148 10988 1158
rect 10752 968 10936 1140
rect 11172 1148 11224 1158
rect 10988 968 11172 1140
rect 4224 868 4864 968
rect 5264 868 5904 968
rect 5264 790 5284 868
rect 6324 868 6924 968
rect 5904 790 6324 800
rect 7344 868 7984 968
rect 6924 790 7344 800
rect 8404 868 9024 968
rect 7984 790 8404 800
rect 9444 868 10044 968
rect 9024 790 9444 800
rect 10464 868 11224 968
rect 10044 790 10464 800
rect 4864 770 5264 780
rect 11620 604 11776 1664
rect 11964 1372 12504 1664
rect 12016 1204 12200 1372
rect 11964 1182 12016 1192
rect 12252 1204 12436 1372
rect 12200 1182 12252 1192
rect 12488 1204 12504 1372
rect 13004 1372 13544 1664
rect 12436 1182 12488 1192
rect 13056 1204 13240 1372
rect 13004 1182 13056 1192
rect 13292 1204 13476 1372
rect 13240 1182 13292 1192
rect 13528 1204 13544 1372
rect 14044 1372 14584 1664
rect 13476 1182 13528 1192
rect 14096 1204 14280 1372
rect 14044 1182 14096 1192
rect 14332 1204 14516 1372
rect 14280 1182 14332 1192
rect 14568 1204 14584 1372
rect 15084 1372 15624 1664
rect 14516 1182 14568 1192
rect 15136 1204 15320 1372
rect 15084 1182 15136 1192
rect 15372 1204 15556 1372
rect 15320 1182 15372 1192
rect 15608 1204 15624 1372
rect 16124 1372 16664 1664
rect 15556 1182 15608 1192
rect 16176 1204 16360 1372
rect 16124 1182 16176 1192
rect 16412 1204 16596 1372
rect 16360 1182 16412 1192
rect 16648 1204 16664 1372
rect 17164 1372 17704 1664
rect 16596 1182 16648 1192
rect 17216 1204 17400 1372
rect 17164 1182 17216 1192
rect 17452 1204 17636 1372
rect 17400 1182 17452 1192
rect 17688 1204 17704 1372
rect 18204 1372 18744 1664
rect 17636 1182 17688 1192
rect 18256 1204 18440 1372
rect 18204 1182 18256 1192
rect 18492 1204 18676 1372
rect 18440 1182 18492 1192
rect 18728 1204 18744 1372
rect 18676 1182 18728 1192
rect 11844 1148 11896 1158
rect 12080 1148 12132 1158
rect 11896 968 12080 1140
rect 12316 1148 12368 1158
rect 12132 968 12316 1140
rect 12552 1148 12604 1158
rect 12368 1120 12552 1140
rect 12884 1148 12936 1158
rect 12604 1120 12884 1130
rect 12368 968 12484 1120
rect 13120 1148 13172 1158
rect 12936 968 13120 1140
rect 13356 1148 13408 1158
rect 13172 968 13356 1140
rect 13592 1148 13644 1158
rect 13408 1120 13592 1140
rect 13924 1148 13976 1158
rect 13644 1120 13924 1130
rect 14160 1148 14212 1158
rect 13408 968 13524 1120
rect 13976 968 14160 1140
rect 14396 1148 14448 1158
rect 14212 968 14396 1140
rect 14632 1148 14684 1158
rect 14448 1120 14632 1140
rect 14964 1148 15016 1158
rect 14684 1120 14964 1130
rect 14448 968 14544 1120
rect 15200 1148 15252 1158
rect 15016 968 15200 1140
rect 15436 1148 15488 1158
rect 15252 968 15436 1140
rect 15672 1148 15724 1158
rect 15488 1120 15672 1140
rect 16004 1148 16056 1158
rect 15724 1120 16004 1130
rect 16240 1148 16292 1158
rect 15488 968 15604 1120
rect 16056 968 16240 1140
rect 16476 1148 16528 1158
rect 16292 968 16476 1140
rect 16712 1148 16764 1158
rect 16528 1120 16712 1140
rect 17044 1148 17096 1158
rect 16764 1120 17044 1130
rect 17280 1148 17332 1158
rect 16528 968 16644 1120
rect 17096 968 17280 1140
rect 17516 1148 17568 1158
rect 17332 968 17516 1140
rect 17752 1148 17804 1158
rect 17568 1120 17752 1140
rect 18084 1148 18136 1158
rect 17804 1120 18084 1130
rect 17568 968 17664 1120
rect 18320 1148 18372 1158
rect 18136 968 18320 1140
rect 18556 1148 18608 1158
rect 18372 968 18556 1140
rect 18792 1148 18844 1158
rect 18608 968 18792 1140
rect 11844 868 12484 968
rect 12884 868 13524 968
rect 12884 790 12904 868
rect 13944 868 14544 968
rect 13524 790 13944 800
rect 14964 868 15604 968
rect 14544 790 14964 800
rect 16024 868 16644 968
rect 15604 790 16024 800
rect 17064 868 17664 968
rect 16644 790 17064 800
rect 18084 868 18844 968
rect 17664 790 18084 800
rect 12484 770 12884 780
rect 4000 552 4984 604
rect 2800 398 3068 400
rect -5998 144 -5802 154
rect 4000 372 4224 552
rect 4276 380 4416 552
rect 4000 362 4276 372
rect 4468 380 4608 552
rect 4416 362 4468 372
rect 4660 380 4800 552
rect 4608 362 4660 372
rect 4792 372 4800 380
rect 4852 372 4984 552
rect 3712 76 3912 86
rect -7314 22 -6490 38
rect -7314 -54 -7030 22
rect -6698 -54 -6490 22
rect -7262 -222 -7122 -54
rect -7314 -244 -7262 -234
rect -7070 -210 -7030 -54
rect -7070 -222 -6930 -210
rect -7122 -244 -7070 -234
rect -6878 -222 -6738 -210
rect -6930 -244 -6878 -234
rect -6686 -222 -6546 -54
rect -6738 -244 -6686 -234
rect -6494 -222 -6490 -54
rect 3712 -150 3912 -140
rect -6546 -244 -6494 -234
rect -7410 -274 -7358 -264
rect -7478 -294 -7410 -284
rect -7218 -274 -7166 -264
rect -7358 -294 -7218 -282
rect -7026 -274 -6974 -264
rect -7166 -294 -7026 -282
rect -7146 -454 -7026 -294
rect -6834 -274 -6782 -264
rect -6974 -454 -6834 -282
rect -6642 -274 -6590 -264
rect -6782 -454 -6642 -282
rect -6450 -274 -6398 -264
rect -6590 -454 -6450 -282
rect -7146 -526 -6398 -454
rect -7478 -536 -6398 -526
rect -7410 -542 -6398 -536
rect 4000 -276 4264 362
rect 4792 352 4984 372
rect 4320 332 4372 342
rect 4512 332 4564 342
rect 4372 310 4512 324
rect 4704 332 4756 342
rect 4564 310 4704 324
rect 4320 -64 4332 152
rect 4752 -64 4756 152
rect 4372 -236 4512 -224
rect 4320 -254 4372 -244
rect 4564 -236 4704 -224
rect 4512 -254 4564 -244
rect 4804 -236 4984 352
rect 4704 -254 4756 -244
rect 4000 -284 4276 -276
rect 4000 -464 4224 -284
rect 4416 -284 4468 -274
rect 4276 -464 4416 -292
rect 4608 -284 4660 -274
rect 4468 -464 4608 -292
rect 4792 -284 4984 -236
rect 4792 -292 4800 -284
rect 4660 -464 4800 -292
rect 4852 -432 4984 -284
rect 5124 552 6024 604
rect 5124 372 5264 552
rect 5316 380 5456 552
rect 5124 362 5316 372
rect 5508 380 5648 552
rect 5456 362 5508 372
rect 5700 380 5840 552
rect 5648 362 5700 372
rect 5832 372 5840 380
rect 5892 372 6024 552
rect 5124 -276 5304 362
rect 5832 352 6024 372
rect 5360 332 5412 342
rect 5552 332 5604 342
rect 5412 310 5552 324
rect 5744 332 5796 342
rect 5604 310 5744 324
rect 5360 -64 5376 152
rect 5412 -236 5552 -224
rect 5360 -254 5412 -244
rect 5604 -236 5744 -224
rect 5552 -254 5604 -244
rect 5844 -236 6024 352
rect 5744 -254 5796 -244
rect 5124 -284 5316 -276
rect 5124 -432 5264 -284
rect 4852 -464 5264 -432
rect 5456 -284 5508 -274
rect 5316 -464 5456 -292
rect 5648 -284 5700 -274
rect 5508 -464 5648 -292
rect 5832 -284 6024 -236
rect 5832 -292 5840 -284
rect 5700 -464 5840 -292
rect 5892 -432 6024 -284
rect 6164 552 7064 604
rect 6164 372 6304 552
rect 6356 380 6496 552
rect 6164 362 6356 372
rect 6548 380 6688 552
rect 6496 362 6548 372
rect 6740 380 6880 552
rect 6688 362 6740 372
rect 6872 372 6880 380
rect 6932 372 7064 552
rect 6164 -276 6344 362
rect 6872 352 7064 372
rect 6400 332 6452 342
rect 6592 332 6644 342
rect 6452 310 6592 324
rect 6784 332 6836 342
rect 6644 310 6784 324
rect 6400 -64 6412 152
rect 6832 -64 6836 152
rect 6452 -236 6592 -224
rect 6400 -254 6452 -244
rect 6644 -236 6784 -224
rect 6592 -254 6644 -244
rect 6884 -236 7064 352
rect 6784 -254 6836 -244
rect 6164 -284 6356 -276
rect 6164 -432 6304 -284
rect 5892 -464 6304 -432
rect 6496 -284 6548 -274
rect 6356 -464 6496 -292
rect 6688 -284 6740 -274
rect 6548 -464 6688 -292
rect 6872 -284 7064 -236
rect 6872 -292 6880 -284
rect 6740 -464 6880 -292
rect 6932 -432 7064 -284
rect 7204 552 8104 604
rect 7204 372 7344 552
rect 7396 380 7536 552
rect 7204 362 7396 372
rect 7588 380 7728 552
rect 7536 362 7588 372
rect 7780 380 7920 552
rect 7728 362 7780 372
rect 7912 372 7920 380
rect 7972 372 8104 552
rect 7204 -276 7384 362
rect 7912 352 8104 372
rect 7440 332 7492 342
rect 7632 332 7684 342
rect 7492 310 7632 324
rect 7824 332 7876 342
rect 7684 310 7824 324
rect 7440 -64 7452 152
rect 7872 -64 7876 152
rect 7492 -236 7632 -224
rect 7440 -254 7492 -244
rect 7684 -236 7824 -224
rect 7632 -254 7684 -244
rect 7924 -236 8104 352
rect 7824 -254 7876 -244
rect 7204 -284 7396 -276
rect 7204 -432 7344 -284
rect 6932 -464 7344 -432
rect 7536 -284 7588 -274
rect 7396 -464 7536 -292
rect 7728 -284 7780 -274
rect 7588 -464 7728 -292
rect 7912 -284 8104 -236
rect 7912 -292 7920 -284
rect 7780 -464 7920 -292
rect 7972 -432 8104 -284
rect 8244 552 9144 604
rect 8244 372 8384 552
rect 8436 380 8576 552
rect 8244 362 8436 372
rect 8628 380 8768 552
rect 8576 362 8628 372
rect 8820 380 8960 552
rect 8768 362 8820 372
rect 8952 372 8960 380
rect 9012 372 9144 552
rect 8244 -276 8424 362
rect 8952 352 9144 372
rect 8480 332 8532 342
rect 8672 332 8724 342
rect 8532 310 8672 324
rect 8864 332 8916 342
rect 8724 310 8864 324
rect 8480 -64 8488 152
rect 8908 -64 8916 152
rect 8532 -236 8672 -224
rect 8480 -254 8532 -244
rect 8724 -236 8864 -224
rect 8672 -254 8724 -244
rect 8964 -236 9144 352
rect 8864 -254 8916 -244
rect 8244 -284 8436 -276
rect 8244 -432 8384 -284
rect 7972 -464 8384 -432
rect 8576 -284 8628 -274
rect 8436 -464 8576 -292
rect 8768 -284 8820 -274
rect 8628 -464 8768 -292
rect 8952 -284 9144 -236
rect 8952 -292 8960 -284
rect 8820 -464 8960 -292
rect 9012 -432 9144 -284
rect 9284 552 10184 604
rect 9284 372 9424 552
rect 9476 380 9616 552
rect 9284 362 9476 372
rect 9668 380 9808 552
rect 9616 362 9668 372
rect 9860 380 10000 552
rect 9808 362 9860 372
rect 9992 372 10000 380
rect 10052 372 10184 552
rect 9284 -276 9464 362
rect 9992 352 10184 372
rect 9520 332 9572 342
rect 9712 332 9764 342
rect 9572 310 9712 324
rect 9904 332 9956 342
rect 9764 310 9904 324
rect 9940 -64 9956 152
rect 9572 -236 9712 -224
rect 9520 -254 9572 -244
rect 9764 -236 9904 -224
rect 9712 -254 9764 -244
rect 10004 -236 10184 352
rect 9904 -254 9956 -244
rect 9284 -284 9476 -276
rect 9284 -432 9424 -284
rect 9012 -464 9424 -432
rect 9616 -284 9668 -274
rect 9476 -464 9616 -292
rect 9808 -284 9860 -274
rect 9668 -464 9808 -292
rect 9992 -284 10184 -236
rect 9992 -292 10000 -284
rect 9860 -464 10000 -292
rect 10052 -432 10184 -284
rect 10324 552 11224 604
rect 10324 372 10464 552
rect 10516 380 10656 552
rect 10324 362 10516 372
rect 10708 380 10848 552
rect 10656 362 10708 372
rect 10900 380 11040 552
rect 10848 362 10900 372
rect 11032 372 11040 380
rect 11092 372 11224 552
rect 10324 -276 10504 362
rect 11032 352 11224 372
rect 10560 332 10612 342
rect 10752 332 10804 342
rect 10612 310 10752 324
rect 10944 332 10996 342
rect 10804 310 10944 324
rect 10980 -64 10996 152
rect 10612 -236 10752 -224
rect 10560 -254 10612 -244
rect 10804 -236 10944 -224
rect 10752 -254 10804 -244
rect 11044 -236 11224 352
rect 10944 -254 10996 -244
rect 10324 -284 10516 -276
rect 10324 -432 10464 -284
rect 10052 -464 10464 -432
rect 10656 -284 10708 -274
rect 10516 -464 10656 -292
rect 10848 -284 10900 -274
rect 10708 -464 10848 -292
rect 11032 -284 11224 -236
rect 11032 -292 11040 -284
rect 10900 -464 11040 -292
rect 11092 -464 11224 -284
rect 4000 -576 11224 -464
rect 11620 552 12604 604
rect 11620 372 11844 552
rect 11896 380 12036 552
rect 11620 362 11896 372
rect 12088 380 12228 552
rect 12036 362 12088 372
rect 12280 380 12420 552
rect 12228 362 12280 372
rect 12412 372 12420 380
rect 12472 372 12604 552
rect 11620 -276 11884 362
rect 12412 352 12604 372
rect 11940 332 11992 342
rect 12132 332 12184 342
rect 11992 310 12132 324
rect 12324 332 12376 342
rect 12184 310 12324 324
rect 11940 -64 11952 152
rect 12372 -64 12376 152
rect 11992 -236 12132 -224
rect 11940 -254 11992 -244
rect 12184 -236 12324 -224
rect 12132 -254 12184 -244
rect 12424 -236 12604 352
rect 12324 -254 12376 -244
rect 11620 -284 11896 -276
rect 11620 -464 11844 -284
rect 12036 -284 12088 -274
rect 11896 -464 12036 -292
rect 12228 -284 12280 -274
rect 12088 -464 12228 -292
rect 12412 -284 12604 -236
rect 12412 -292 12420 -284
rect 12280 -464 12420 -292
rect 12472 -432 12604 -284
rect 12744 552 13644 604
rect 12744 372 12884 552
rect 12936 380 13076 552
rect 12744 362 12936 372
rect 13128 380 13268 552
rect 13076 362 13128 372
rect 13320 380 13460 552
rect 13268 362 13320 372
rect 13452 372 13460 380
rect 13512 372 13644 552
rect 12744 -276 12924 362
rect 13452 352 13644 372
rect 12980 332 13032 342
rect 13172 332 13224 342
rect 13032 310 13172 324
rect 13364 332 13416 342
rect 13224 310 13364 324
rect 12980 -64 12996 152
rect 13032 -236 13172 -224
rect 12980 -254 13032 -244
rect 13224 -236 13364 -224
rect 13172 -254 13224 -244
rect 13464 -236 13644 352
rect 13364 -254 13416 -244
rect 12744 -284 12936 -276
rect 12744 -432 12884 -284
rect 12472 -464 12884 -432
rect 13076 -284 13128 -274
rect 12936 -464 13076 -292
rect 13268 -284 13320 -274
rect 13128 -464 13268 -292
rect 13452 -284 13644 -236
rect 13452 -292 13460 -284
rect 13320 -464 13460 -292
rect 13512 -432 13644 -284
rect 13784 552 14684 604
rect 13784 372 13924 552
rect 13976 380 14116 552
rect 13784 362 13976 372
rect 14168 380 14308 552
rect 14116 362 14168 372
rect 14360 380 14500 552
rect 14308 362 14360 372
rect 14492 372 14500 380
rect 14552 372 14684 552
rect 13784 -276 13964 362
rect 14492 352 14684 372
rect 14020 332 14072 342
rect 14212 332 14264 342
rect 14072 310 14212 324
rect 14404 332 14456 342
rect 14264 310 14404 324
rect 14020 -64 14032 152
rect 14452 -64 14456 152
rect 14072 -236 14212 -224
rect 14020 -254 14072 -244
rect 14264 -236 14404 -224
rect 14212 -254 14264 -244
rect 14504 -236 14684 352
rect 14404 -254 14456 -244
rect 13784 -284 13976 -276
rect 13784 -432 13924 -284
rect 13512 -464 13924 -432
rect 14116 -284 14168 -274
rect 13976 -464 14116 -292
rect 14308 -284 14360 -274
rect 14168 -464 14308 -292
rect 14492 -284 14684 -236
rect 14492 -292 14500 -284
rect 14360 -464 14500 -292
rect 14552 -432 14684 -284
rect 14824 552 15724 604
rect 14824 372 14964 552
rect 15016 380 15156 552
rect 14824 362 15016 372
rect 15208 380 15348 552
rect 15156 362 15208 372
rect 15400 380 15540 552
rect 15348 362 15400 372
rect 15532 372 15540 380
rect 15592 372 15724 552
rect 14824 -276 15004 362
rect 15532 352 15724 372
rect 15060 332 15112 342
rect 15252 332 15304 342
rect 15112 310 15252 324
rect 15444 332 15496 342
rect 15304 310 15444 324
rect 15060 -64 15072 152
rect 15492 -64 15496 152
rect 15112 -236 15252 -224
rect 15060 -254 15112 -244
rect 15304 -236 15444 -224
rect 15252 -254 15304 -244
rect 15544 -236 15724 352
rect 15444 -254 15496 -244
rect 14824 -284 15016 -276
rect 14824 -432 14964 -284
rect 14552 -464 14964 -432
rect 15156 -284 15208 -274
rect 15016 -464 15156 -292
rect 15348 -284 15400 -274
rect 15208 -464 15348 -292
rect 15532 -284 15724 -236
rect 15532 -292 15540 -284
rect 15400 -464 15540 -292
rect 15592 -432 15724 -284
rect 15864 552 16764 604
rect 15864 372 16004 552
rect 16056 380 16196 552
rect 15864 362 16056 372
rect 16248 380 16388 552
rect 16196 362 16248 372
rect 16440 380 16580 552
rect 16388 362 16440 372
rect 16572 372 16580 380
rect 16632 372 16764 552
rect 15864 -276 16044 362
rect 16572 352 16764 372
rect 16100 332 16152 342
rect 16292 332 16344 342
rect 16152 310 16292 324
rect 16484 332 16536 342
rect 16344 310 16484 324
rect 16100 -64 16108 152
rect 16528 -64 16536 152
rect 16152 -236 16292 -224
rect 16100 -254 16152 -244
rect 16344 -236 16484 -224
rect 16292 -254 16344 -244
rect 16584 -236 16764 352
rect 16484 -254 16536 -244
rect 15864 -284 16056 -276
rect 15864 -432 16004 -284
rect 15592 -464 16004 -432
rect 16196 -284 16248 -274
rect 16056 -464 16196 -292
rect 16388 -284 16440 -274
rect 16248 -464 16388 -292
rect 16572 -284 16764 -236
rect 16572 -292 16580 -284
rect 16440 -464 16580 -292
rect 16632 -432 16764 -284
rect 16904 552 17804 604
rect 16904 372 17044 552
rect 17096 380 17236 552
rect 16904 362 17096 372
rect 17288 380 17428 552
rect 17236 362 17288 372
rect 17480 380 17620 552
rect 17428 362 17480 372
rect 17612 372 17620 380
rect 17672 372 17804 552
rect 16904 -276 17084 362
rect 17612 352 17804 372
rect 17140 332 17192 342
rect 17332 332 17384 342
rect 17192 310 17332 324
rect 17524 332 17576 342
rect 17384 310 17524 324
rect 17560 -64 17576 152
rect 17192 -236 17332 -224
rect 17140 -254 17192 -244
rect 17384 -236 17524 -224
rect 17332 -254 17384 -244
rect 17624 -236 17804 352
rect 17524 -254 17576 -244
rect 16904 -284 17096 -276
rect 16904 -432 17044 -284
rect 16632 -464 17044 -432
rect 17236 -284 17288 -274
rect 17096 -464 17236 -292
rect 17428 -284 17480 -274
rect 17288 -464 17428 -292
rect 17612 -284 17804 -236
rect 17612 -292 17620 -284
rect 17480 -464 17620 -292
rect 17672 -432 17804 -284
rect 17944 552 18844 604
rect 17944 372 18084 552
rect 18136 380 18276 552
rect 17944 362 18136 372
rect 18328 380 18468 552
rect 18276 362 18328 372
rect 18520 380 18660 552
rect 18468 362 18520 372
rect 18652 372 18660 380
rect 18712 372 18844 552
rect 17944 -276 18124 362
rect 18652 352 18844 372
rect 18180 332 18232 342
rect 18372 332 18424 342
rect 18232 310 18372 324
rect 18564 332 18616 342
rect 18424 310 18564 324
rect 18600 -64 18616 152
rect 18232 -236 18372 -224
rect 18180 -254 18232 -244
rect 18424 -236 18564 -224
rect 18372 -254 18424 -244
rect 18664 -236 18844 352
rect 18564 -254 18616 -244
rect 17944 -284 18136 -276
rect 17944 -432 18084 -284
rect 17672 -464 18084 -432
rect 18276 -284 18328 -274
rect 18136 -464 18276 -292
rect 18468 -284 18520 -274
rect 18328 -464 18468 -292
rect 18652 -284 18844 -236
rect 18652 -292 18660 -284
rect 18520 -464 18660 -292
rect 18712 -464 18844 -284
rect 11620 -576 18844 -464
rect -7314 -598 -6494 -582
rect -7314 -670 -7030 -598
rect -6698 -670 -6494 -598
rect -7262 -842 -7122 -670
rect -7314 -860 -7262 -850
rect -7070 -830 -7030 -670
rect -7070 -842 -6930 -830
rect -7122 -860 -7070 -850
rect -6878 -842 -6738 -830
rect -6930 -860 -6878 -850
rect -6686 -842 -6546 -670
rect -6738 -860 -6686 -850
rect -6546 -860 -6494 -850
rect -7410 -894 -7358 -884
rect -7478 -918 -7410 -908
rect -7218 -894 -7166 -884
rect -7358 -918 -7218 -902
rect -7026 -894 -6974 -884
rect -7166 -918 -7026 -902
rect -7146 -1074 -7026 -918
rect -6834 -894 -6782 -884
rect -6974 -1074 -6834 -902
rect -6642 -894 -6590 -884
rect -6782 -1074 -6642 -902
rect -6450 -894 -6398 -884
rect -6590 -1074 -6450 -902
rect -7146 -1150 -6398 -1074
rect -7478 -1160 -6398 -1150
rect -7410 -1162 -6398 -1160
rect 4000 -1636 4156 -576
rect 4344 -868 4884 -576
rect 4396 -1036 4580 -868
rect 4344 -1058 4396 -1048
rect 4632 -1036 4816 -868
rect 4580 -1058 4632 -1048
rect 4868 -1036 4884 -868
rect 5384 -868 5924 -576
rect 4816 -1058 4868 -1048
rect 5436 -1036 5620 -868
rect 5384 -1058 5436 -1048
rect 5672 -1036 5856 -868
rect 5620 -1058 5672 -1048
rect 5908 -1036 5924 -868
rect 6424 -868 6964 -576
rect 5856 -1058 5908 -1048
rect 6476 -1036 6660 -868
rect 6424 -1058 6476 -1048
rect 6712 -1036 6896 -868
rect 6660 -1058 6712 -1048
rect 6948 -1036 6964 -868
rect 7464 -868 8004 -576
rect 6896 -1058 6948 -1048
rect 7516 -1036 7700 -868
rect 7464 -1058 7516 -1048
rect 7752 -1036 7936 -868
rect 7700 -1058 7752 -1048
rect 7988 -1036 8004 -868
rect 8504 -868 9044 -576
rect 7936 -1058 7988 -1048
rect 8556 -1036 8740 -868
rect 8504 -1058 8556 -1048
rect 8792 -1036 8976 -868
rect 8740 -1058 8792 -1048
rect 9028 -1036 9044 -868
rect 9544 -868 10084 -576
rect 8976 -1058 9028 -1048
rect 9596 -1036 9780 -868
rect 9544 -1058 9596 -1048
rect 9832 -1036 10016 -868
rect 9780 -1058 9832 -1048
rect 10068 -1036 10084 -868
rect 10584 -868 11124 -576
rect 10016 -1058 10068 -1048
rect 10636 -1036 10820 -868
rect 10584 -1058 10636 -1048
rect 10872 -1036 11056 -868
rect 10820 -1058 10872 -1048
rect 11108 -1036 11124 -868
rect 11056 -1058 11108 -1048
rect 4224 -1092 4276 -1082
rect 4460 -1092 4512 -1082
rect 4276 -1272 4460 -1100
rect 4696 -1092 4748 -1082
rect 4512 -1272 4696 -1100
rect 4932 -1092 4984 -1082
rect 4748 -1120 4932 -1100
rect 5264 -1092 5316 -1082
rect 4984 -1120 5264 -1110
rect 4748 -1272 4844 -1120
rect 5500 -1092 5552 -1082
rect 5316 -1272 5500 -1100
rect 5736 -1092 5788 -1082
rect 5552 -1272 5736 -1100
rect 5972 -1092 6024 -1082
rect 5788 -1120 5972 -1100
rect 6304 -1092 6356 -1082
rect 6024 -1120 6304 -1110
rect 6540 -1092 6592 -1082
rect 5788 -1272 5904 -1120
rect 6356 -1272 6540 -1100
rect 6776 -1092 6828 -1082
rect 6592 -1272 6776 -1100
rect 7012 -1092 7064 -1082
rect 6828 -1120 7012 -1100
rect 7344 -1092 7396 -1082
rect 7064 -1120 7344 -1110
rect 6828 -1272 6924 -1120
rect 7580 -1092 7632 -1082
rect 7396 -1272 7580 -1100
rect 7816 -1092 7868 -1082
rect 7632 -1272 7816 -1100
rect 8052 -1092 8104 -1082
rect 7868 -1120 8052 -1100
rect 8384 -1092 8436 -1082
rect 8104 -1120 8384 -1110
rect 8620 -1092 8672 -1082
rect 7868 -1272 7984 -1120
rect 8436 -1272 8620 -1100
rect 8856 -1092 8908 -1082
rect 8672 -1272 8856 -1100
rect 9092 -1092 9144 -1082
rect 8908 -1120 9092 -1100
rect 9424 -1092 9476 -1082
rect 9144 -1120 9424 -1110
rect 8908 -1272 9004 -1120
rect 9660 -1092 9712 -1082
rect 9476 -1272 9660 -1100
rect 9896 -1092 9948 -1082
rect 9712 -1272 9896 -1100
rect 10132 -1092 10184 -1082
rect 9948 -1120 10132 -1100
rect 10464 -1092 10516 -1082
rect 10184 -1120 10464 -1110
rect 9948 -1272 10044 -1120
rect 10700 -1092 10752 -1082
rect 10516 -1272 10700 -1100
rect 10936 -1092 10988 -1082
rect 10752 -1272 10936 -1100
rect 11172 -1092 11224 -1082
rect 10988 -1272 11172 -1100
rect 4224 -1372 4844 -1272
rect 5264 -1372 5904 -1272
rect 4844 -1450 5264 -1440
rect 6324 -1372 6924 -1272
rect 5904 -1450 6324 -1440
rect 7344 -1372 7984 -1272
rect 6924 -1450 7344 -1440
rect 8404 -1372 9004 -1272
rect 7984 -1450 8404 -1440
rect 9424 -1372 10044 -1272
rect 9004 -1450 9424 -1440
rect 10464 -1372 11224 -1272
rect 10044 -1450 10464 -1440
rect 11620 -1636 11776 -576
rect 11964 -868 12504 -576
rect 12016 -1036 12200 -868
rect 11964 -1058 12016 -1048
rect 12252 -1036 12436 -868
rect 12200 -1058 12252 -1048
rect 12488 -1036 12504 -868
rect 13004 -868 13544 -576
rect 12436 -1058 12488 -1048
rect 13056 -1036 13240 -868
rect 13004 -1058 13056 -1048
rect 13292 -1036 13476 -868
rect 13240 -1058 13292 -1048
rect 13528 -1036 13544 -868
rect 14044 -868 14584 -576
rect 13476 -1058 13528 -1048
rect 14096 -1036 14280 -868
rect 14044 -1058 14096 -1048
rect 14332 -1036 14516 -868
rect 14280 -1058 14332 -1048
rect 14568 -1036 14584 -868
rect 15084 -868 15624 -576
rect 14516 -1058 14568 -1048
rect 15136 -1036 15320 -868
rect 15084 -1058 15136 -1048
rect 15372 -1036 15556 -868
rect 15320 -1058 15372 -1048
rect 15608 -1036 15624 -868
rect 16124 -868 16664 -576
rect 15556 -1058 15608 -1048
rect 16176 -1036 16360 -868
rect 16124 -1058 16176 -1048
rect 16412 -1036 16596 -868
rect 16360 -1058 16412 -1048
rect 16648 -1036 16664 -868
rect 17164 -868 17704 -576
rect 16596 -1058 16648 -1048
rect 17216 -1036 17400 -868
rect 17164 -1058 17216 -1048
rect 17452 -1036 17636 -868
rect 17400 -1058 17452 -1048
rect 17688 -1036 17704 -868
rect 18204 -868 18744 -576
rect 17636 -1058 17688 -1048
rect 18256 -1036 18440 -868
rect 18204 -1058 18256 -1048
rect 18492 -1036 18676 -868
rect 18440 -1058 18492 -1048
rect 18728 -1036 18744 -868
rect 18676 -1058 18728 -1048
rect 11844 -1092 11896 -1082
rect 12080 -1092 12132 -1082
rect 11896 -1272 12080 -1100
rect 12316 -1092 12368 -1082
rect 12132 -1272 12316 -1100
rect 12552 -1092 12604 -1082
rect 12368 -1120 12552 -1100
rect 12884 -1092 12936 -1082
rect 12604 -1120 12884 -1110
rect 12368 -1272 12464 -1120
rect 13120 -1092 13172 -1082
rect 12936 -1272 13120 -1100
rect 13356 -1092 13408 -1082
rect 13172 -1272 13356 -1100
rect 13592 -1092 13644 -1082
rect 13408 -1120 13592 -1100
rect 13924 -1092 13976 -1082
rect 13644 -1120 13924 -1110
rect 14160 -1092 14212 -1082
rect 13408 -1272 13524 -1120
rect 13976 -1272 14160 -1100
rect 14396 -1092 14448 -1082
rect 14212 -1272 14396 -1100
rect 14632 -1092 14684 -1082
rect 14448 -1120 14632 -1100
rect 14964 -1092 15016 -1082
rect 14684 -1120 14964 -1110
rect 14448 -1272 14544 -1120
rect 15200 -1092 15252 -1082
rect 15016 -1272 15200 -1100
rect 15436 -1092 15488 -1082
rect 15252 -1272 15436 -1100
rect 15672 -1092 15724 -1082
rect 15488 -1120 15672 -1100
rect 16004 -1092 16056 -1082
rect 15724 -1120 16004 -1110
rect 16240 -1092 16292 -1082
rect 15488 -1272 15604 -1120
rect 16056 -1272 16240 -1100
rect 16476 -1092 16528 -1082
rect 16292 -1272 16476 -1100
rect 16712 -1092 16764 -1082
rect 16528 -1120 16712 -1100
rect 17044 -1092 17096 -1082
rect 16764 -1120 17044 -1110
rect 16528 -1272 16624 -1120
rect 17280 -1092 17332 -1082
rect 17096 -1272 17280 -1100
rect 17516 -1092 17568 -1082
rect 17332 -1272 17516 -1100
rect 17752 -1092 17804 -1082
rect 17568 -1120 17752 -1100
rect 18084 -1092 18136 -1082
rect 17804 -1120 18084 -1110
rect 17568 -1272 17664 -1120
rect 18320 -1092 18372 -1082
rect 18136 -1272 18320 -1100
rect 18556 -1092 18608 -1082
rect 18372 -1272 18556 -1100
rect 18792 -1092 18844 -1082
rect 18608 -1272 18792 -1100
rect 11844 -1372 12464 -1272
rect 12884 -1372 13524 -1272
rect 12464 -1450 12884 -1440
rect 13944 -1372 14544 -1272
rect 13524 -1450 13944 -1440
rect 14964 -1372 15604 -1272
rect 14544 -1450 14964 -1440
rect 16024 -1372 16624 -1272
rect 15604 -1450 16024 -1440
rect 17044 -1372 17664 -1272
rect 16624 -1450 17044 -1440
rect 18084 -1372 18844 -1272
rect 17664 -1450 18084 -1440
rect 4000 -1688 4984 -1636
rect -7550 -1890 -6650 -1838
rect -7550 -2070 -7410 -1890
rect -7358 -2062 -7218 -1890
rect -7550 -2080 -7358 -2070
rect -7166 -2062 -7026 -1890
rect -7218 -2080 -7166 -2070
rect -6974 -2062 -6834 -1890
rect -7026 -2080 -6974 -2070
rect -6842 -2070 -6834 -2062
rect -6782 -2070 -6650 -1890
rect -7550 -2718 -7370 -2080
rect -6842 -2090 -6650 -2070
rect -7314 -2110 -7262 -2100
rect -7122 -2110 -7070 -2100
rect -7262 -2154 -7122 -2118
rect -6930 -2110 -6878 -2100
rect -7070 -2154 -6930 -2118
rect -7314 -2506 -7298 -2290
rect -6910 -2506 -6878 -2290
rect -7262 -2678 -7122 -2646
rect -7314 -2696 -7262 -2686
rect -7070 -2678 -6930 -2646
rect -7122 -2696 -7070 -2686
rect -6830 -2678 -6650 -2090
rect -6930 -2696 -6878 -2686
rect -7550 -2726 -7358 -2718
rect -7550 -2906 -7410 -2726
rect -7218 -2726 -7166 -2716
rect -7358 -2906 -7218 -2734
rect -7026 -2726 -6974 -2716
rect -7166 -2906 -7026 -2734
rect -6842 -2726 -6650 -2678
rect -6842 -2734 -6834 -2726
rect -6974 -2906 -6834 -2734
rect -6782 -2906 -6650 -2726
rect 4000 -1868 4224 -1688
rect 4276 -1860 4416 -1688
rect 4000 -1878 4276 -1868
rect 4468 -1860 4608 -1688
rect 4416 -1878 4468 -1868
rect 4660 -1860 4800 -1688
rect 4608 -1878 4660 -1868
rect 4792 -1868 4800 -1860
rect 4852 -1868 4984 -1688
rect 4000 -2516 4264 -1878
rect 4792 -1888 4984 -1868
rect 4320 -1908 4372 -1898
rect 4512 -1908 4564 -1898
rect 4372 -1936 4512 -1916
rect 4704 -1908 4756 -1898
rect 4564 -1936 4704 -1916
rect 4320 -2304 4332 -2088
rect 4732 -2304 4756 -2088
rect 4372 -2476 4512 -2460
rect 4320 -2494 4372 -2484
rect 4564 -2476 4704 -2460
rect 4512 -2494 4564 -2484
rect 4804 -2476 4984 -1888
rect 4704 -2494 4756 -2484
rect 4000 -2524 4276 -2516
rect 4000 -2704 4224 -2524
rect 4416 -2524 4468 -2514
rect 4276 -2704 4416 -2532
rect 4608 -2524 4660 -2514
rect 4468 -2704 4608 -2532
rect 4792 -2524 4984 -2476
rect 4792 -2532 4800 -2524
rect 4660 -2704 4800 -2532
rect 4852 -2672 4984 -2524
rect 5124 -1688 6024 -1636
rect 5124 -1868 5264 -1688
rect 5316 -1860 5456 -1688
rect 5124 -1878 5316 -1868
rect 5508 -1860 5648 -1688
rect 5456 -1878 5508 -1868
rect 5700 -1860 5840 -1688
rect 5648 -1878 5700 -1868
rect 5832 -1868 5840 -1860
rect 5892 -1868 6024 -1688
rect 5124 -2516 5304 -1878
rect 5832 -1888 6024 -1868
rect 5360 -1908 5412 -1898
rect 5552 -1908 5604 -1898
rect 5412 -1936 5552 -1916
rect 5744 -1908 5796 -1898
rect 5604 -1936 5744 -1916
rect 5360 -2304 5372 -2088
rect 5772 -2304 5796 -2088
rect 5412 -2476 5552 -2460
rect 5360 -2494 5412 -2484
rect 5604 -2476 5744 -2460
rect 5552 -2494 5604 -2484
rect 5844 -2476 6024 -1888
rect 5744 -2494 5796 -2484
rect 5124 -2524 5316 -2516
rect 5124 -2672 5264 -2524
rect 4852 -2704 5264 -2672
rect 5456 -2524 5508 -2514
rect 5316 -2704 5456 -2532
rect 5648 -2524 5700 -2514
rect 5508 -2704 5648 -2532
rect 5832 -2524 6024 -2476
rect 5832 -2532 5840 -2524
rect 5700 -2704 5840 -2532
rect 5892 -2672 6024 -2524
rect 6164 -1688 7064 -1636
rect 6164 -1868 6304 -1688
rect 6356 -1860 6496 -1688
rect 6164 -1878 6356 -1868
rect 6548 -1860 6688 -1688
rect 6496 -1878 6548 -1868
rect 6740 -1860 6880 -1688
rect 6688 -1878 6740 -1868
rect 6872 -1868 6880 -1860
rect 6932 -1868 7064 -1688
rect 6164 -2516 6344 -1878
rect 6872 -1888 7064 -1868
rect 6400 -1908 6452 -1898
rect 6592 -1908 6644 -1898
rect 6452 -1936 6592 -1916
rect 6784 -1908 6836 -1898
rect 6644 -1936 6784 -1916
rect 6400 -2304 6412 -2088
rect 6812 -2304 6836 -2088
rect 6452 -2476 6592 -2460
rect 6400 -2494 6452 -2484
rect 6644 -2476 6784 -2460
rect 6592 -2494 6644 -2484
rect 6884 -2476 7064 -1888
rect 6784 -2494 6836 -2484
rect 6164 -2524 6356 -2516
rect 6164 -2672 6304 -2524
rect 5892 -2704 6304 -2672
rect 6496 -2524 6548 -2514
rect 6356 -2704 6496 -2532
rect 6688 -2524 6740 -2514
rect 6548 -2704 6688 -2532
rect 6872 -2524 7064 -2476
rect 6872 -2532 6880 -2524
rect 6740 -2704 6880 -2532
rect 6932 -2672 7064 -2524
rect 7204 -1688 8104 -1636
rect 7204 -1868 7344 -1688
rect 7396 -1860 7536 -1688
rect 7204 -1878 7396 -1868
rect 7588 -1860 7728 -1688
rect 7536 -1878 7588 -1868
rect 7780 -1860 7920 -1688
rect 7728 -1878 7780 -1868
rect 7912 -1868 7920 -1860
rect 7972 -1868 8104 -1688
rect 7204 -2516 7384 -1878
rect 7912 -1888 8104 -1868
rect 7440 -1908 7492 -1898
rect 7632 -1908 7684 -1898
rect 7492 -1936 7632 -1916
rect 7824 -1908 7876 -1898
rect 7684 -1936 7824 -1916
rect 7440 -2304 7452 -2088
rect 7852 -2304 7876 -2088
rect 7492 -2476 7632 -2460
rect 7440 -2494 7492 -2484
rect 7684 -2476 7824 -2460
rect 7632 -2494 7684 -2484
rect 7924 -2476 8104 -1888
rect 7824 -2494 7876 -2484
rect 7204 -2524 7396 -2516
rect 7204 -2672 7344 -2524
rect 6932 -2704 7344 -2672
rect 7536 -2524 7588 -2514
rect 7396 -2704 7536 -2532
rect 7728 -2524 7780 -2514
rect 7588 -2704 7728 -2532
rect 7912 -2524 8104 -2476
rect 7912 -2532 7920 -2524
rect 7780 -2704 7920 -2532
rect 7972 -2672 8104 -2524
rect 8244 -1688 9144 -1636
rect 8244 -1868 8384 -1688
rect 8436 -1860 8576 -1688
rect 8244 -1878 8436 -1868
rect 8628 -1860 8768 -1688
rect 8576 -1878 8628 -1868
rect 8820 -1860 8960 -1688
rect 8768 -1878 8820 -1868
rect 8952 -1868 8960 -1860
rect 9012 -1868 9144 -1688
rect 8244 -2516 8424 -1878
rect 8952 -1888 9144 -1868
rect 8480 -1908 8532 -1898
rect 8672 -1908 8724 -1898
rect 8532 -1936 8672 -1916
rect 8864 -1908 8916 -1898
rect 8724 -1936 8864 -1916
rect 8480 -2304 8488 -2088
rect 8888 -2304 8916 -2088
rect 8532 -2476 8672 -2460
rect 8480 -2494 8532 -2484
rect 8724 -2476 8864 -2460
rect 8672 -2494 8724 -2484
rect 8964 -2476 9144 -1888
rect 8864 -2494 8916 -2484
rect 8244 -2524 8436 -2516
rect 8244 -2672 8384 -2524
rect 7972 -2704 8384 -2672
rect 8576 -2524 8628 -2514
rect 8436 -2704 8576 -2532
rect 8768 -2524 8820 -2514
rect 8628 -2704 8768 -2532
rect 8952 -2524 9144 -2476
rect 8952 -2532 8960 -2524
rect 8820 -2704 8960 -2532
rect 9012 -2704 9144 -2524
rect 4000 -2816 9144 -2704
rect 11620 -1688 12604 -1636
rect 11620 -1868 11844 -1688
rect 11896 -1860 12036 -1688
rect 11620 -1878 11896 -1868
rect 12088 -1860 12228 -1688
rect 12036 -1878 12088 -1868
rect 12280 -1860 12420 -1688
rect 12228 -1878 12280 -1868
rect 12412 -1868 12420 -1860
rect 12472 -1868 12604 -1688
rect 11620 -2516 11884 -1878
rect 12412 -1888 12604 -1868
rect 11940 -1908 11992 -1898
rect 12132 -1908 12184 -1898
rect 11992 -1936 12132 -1916
rect 12324 -1908 12376 -1898
rect 12184 -1936 12324 -1916
rect 11940 -2304 11952 -2088
rect 12352 -2304 12376 -2088
rect 11992 -2476 12132 -2460
rect 11940 -2494 11992 -2484
rect 12184 -2476 12324 -2460
rect 12132 -2494 12184 -2484
rect 12424 -2476 12604 -1888
rect 12324 -2494 12376 -2484
rect 11620 -2524 11896 -2516
rect 11620 -2704 11844 -2524
rect 12036 -2524 12088 -2514
rect 11896 -2704 12036 -2532
rect 12228 -2524 12280 -2514
rect 12088 -2704 12228 -2532
rect 12412 -2524 12604 -2476
rect 12412 -2532 12420 -2524
rect 12280 -2704 12420 -2532
rect 12472 -2672 12604 -2524
rect 12744 -1688 13644 -1636
rect 12744 -1868 12884 -1688
rect 12936 -1860 13076 -1688
rect 12744 -1878 12936 -1868
rect 13128 -1860 13268 -1688
rect 13076 -1878 13128 -1868
rect 13320 -1860 13460 -1688
rect 13268 -1878 13320 -1868
rect 13452 -1868 13460 -1860
rect 13512 -1868 13644 -1688
rect 12744 -2516 12924 -1878
rect 13452 -1888 13644 -1868
rect 12980 -1908 13032 -1898
rect 13172 -1908 13224 -1898
rect 13032 -1936 13172 -1916
rect 13364 -1908 13416 -1898
rect 13224 -1936 13364 -1916
rect 12980 -2304 12992 -2088
rect 13392 -2304 13416 -2088
rect 13032 -2476 13172 -2460
rect 12980 -2494 13032 -2484
rect 13224 -2476 13364 -2460
rect 13172 -2494 13224 -2484
rect 13464 -2476 13644 -1888
rect 13364 -2494 13416 -2484
rect 12744 -2524 12936 -2516
rect 12744 -2672 12884 -2524
rect 12472 -2704 12884 -2672
rect 13076 -2524 13128 -2514
rect 12936 -2704 13076 -2532
rect 13268 -2524 13320 -2514
rect 13128 -2704 13268 -2532
rect 13452 -2524 13644 -2476
rect 13452 -2532 13460 -2524
rect 13320 -2704 13460 -2532
rect 13512 -2672 13644 -2524
rect 13784 -1688 14684 -1636
rect 13784 -1868 13924 -1688
rect 13976 -1860 14116 -1688
rect 13784 -1878 13976 -1868
rect 14168 -1860 14308 -1688
rect 14116 -1878 14168 -1868
rect 14360 -1860 14500 -1688
rect 14308 -1878 14360 -1868
rect 14492 -1868 14500 -1860
rect 14552 -1868 14684 -1688
rect 13784 -2516 13964 -1878
rect 14492 -1888 14684 -1868
rect 14020 -1908 14072 -1898
rect 14212 -1908 14264 -1898
rect 14072 -1936 14212 -1916
rect 14404 -1908 14456 -1898
rect 14264 -1936 14404 -1916
rect 14020 -2304 14032 -2088
rect 14432 -2304 14456 -2088
rect 14072 -2476 14212 -2460
rect 14020 -2494 14072 -2484
rect 14264 -2476 14404 -2460
rect 14212 -2494 14264 -2484
rect 14504 -2476 14684 -1888
rect 14404 -2494 14456 -2484
rect 13784 -2524 13976 -2516
rect 13784 -2672 13924 -2524
rect 13512 -2704 13924 -2672
rect 14116 -2524 14168 -2514
rect 13976 -2704 14116 -2532
rect 14308 -2524 14360 -2514
rect 14168 -2704 14308 -2532
rect 14492 -2524 14684 -2476
rect 14492 -2532 14500 -2524
rect 14360 -2704 14500 -2532
rect 14552 -2672 14684 -2524
rect 14824 -1688 15724 -1636
rect 14824 -1868 14964 -1688
rect 15016 -1860 15156 -1688
rect 14824 -1878 15016 -1868
rect 15208 -1860 15348 -1688
rect 15156 -1878 15208 -1868
rect 15400 -1860 15540 -1688
rect 15348 -1878 15400 -1868
rect 15532 -1868 15540 -1860
rect 15592 -1868 15724 -1688
rect 14824 -2516 15004 -1878
rect 15532 -1888 15724 -1868
rect 15060 -1908 15112 -1898
rect 15252 -1908 15304 -1898
rect 15112 -1936 15252 -1916
rect 15444 -1908 15496 -1898
rect 15304 -1936 15444 -1916
rect 15060 -2304 15072 -2088
rect 15472 -2304 15496 -2088
rect 15112 -2476 15252 -2460
rect 15060 -2494 15112 -2484
rect 15304 -2476 15444 -2460
rect 15252 -2494 15304 -2484
rect 15544 -2476 15724 -1888
rect 15444 -2494 15496 -2484
rect 14824 -2524 15016 -2516
rect 14824 -2672 14964 -2524
rect 14552 -2704 14964 -2672
rect 15156 -2524 15208 -2514
rect 15016 -2704 15156 -2532
rect 15348 -2524 15400 -2514
rect 15208 -2704 15348 -2532
rect 15532 -2524 15724 -2476
rect 15532 -2532 15540 -2524
rect 15400 -2704 15540 -2532
rect 15592 -2672 15724 -2524
rect 15864 -1688 16764 -1636
rect 15864 -1868 16004 -1688
rect 16056 -1860 16196 -1688
rect 15864 -1878 16056 -1868
rect 16248 -1860 16388 -1688
rect 16196 -1878 16248 -1868
rect 16440 -1860 16580 -1688
rect 16388 -1878 16440 -1868
rect 16572 -1868 16580 -1860
rect 16632 -1868 16764 -1688
rect 15864 -2516 16044 -1878
rect 16572 -1888 16764 -1868
rect 16100 -1908 16152 -1898
rect 16292 -1908 16344 -1898
rect 16152 -1936 16292 -1916
rect 16484 -1908 16536 -1898
rect 16344 -1936 16484 -1916
rect 16100 -2304 16108 -2088
rect 16508 -2304 16536 -2088
rect 16152 -2476 16292 -2460
rect 16100 -2494 16152 -2484
rect 16344 -2476 16484 -2460
rect 16292 -2494 16344 -2484
rect 16584 -2476 16764 -1888
rect 16484 -2494 16536 -2484
rect 15864 -2524 16056 -2516
rect 15864 -2672 16004 -2524
rect 15592 -2704 16004 -2672
rect 16196 -2524 16248 -2514
rect 16056 -2704 16196 -2532
rect 16388 -2524 16440 -2514
rect 16248 -2704 16388 -2532
rect 16572 -2524 16764 -2476
rect 16572 -2532 16580 -2524
rect 16440 -2704 16580 -2532
rect 16632 -2704 16764 -2524
rect 11620 -2816 16764 -2704
rect -7550 -3018 -6650 -2906
rect -7290 -3310 -6750 -3018
rect 4344 -3108 4884 -2816
rect 4396 -3276 4580 -3108
rect 4344 -3298 4396 -3288
rect 4632 -3276 4816 -3108
rect 4580 -3298 4632 -3288
rect 4868 -3276 4884 -3108
rect 5384 -3108 5924 -2816
rect 4816 -3298 4868 -3288
rect 5436 -3276 5620 -3108
rect 5384 -3298 5436 -3288
rect 5672 -3276 5856 -3108
rect 5620 -3298 5672 -3288
rect 5908 -3276 5924 -3108
rect 6424 -3108 6964 -2816
rect 5856 -3298 5908 -3288
rect 6476 -3276 6660 -3108
rect 6424 -3298 6476 -3288
rect 6712 -3276 6896 -3108
rect 6660 -3298 6712 -3288
rect 6948 -3276 6964 -3108
rect 7464 -3108 8004 -2816
rect 6896 -3298 6948 -3288
rect 7516 -3276 7700 -3108
rect 7464 -3298 7516 -3288
rect 7752 -3276 7936 -3108
rect 7700 -3298 7752 -3288
rect 7988 -3276 8004 -3108
rect 8504 -3108 9044 -2816
rect 7936 -3298 7988 -3288
rect 8556 -3276 8740 -3108
rect 8504 -3298 8556 -3288
rect 8792 -3276 8976 -3108
rect 8740 -3298 8792 -3288
rect 9028 -3276 9044 -3108
rect 11964 -3108 12504 -2816
rect 8976 -3298 9028 -3288
rect 12016 -3276 12200 -3108
rect 11964 -3298 12016 -3288
rect 12252 -3276 12436 -3108
rect 12200 -3298 12252 -3288
rect 12488 -3276 12504 -3108
rect 13004 -3108 13544 -2816
rect 12436 -3298 12488 -3288
rect 13056 -3276 13240 -3108
rect 13004 -3298 13056 -3288
rect 13292 -3276 13476 -3108
rect 13240 -3298 13292 -3288
rect 13528 -3276 13544 -3108
rect 14044 -3108 14584 -2816
rect 13476 -3298 13528 -3288
rect 14096 -3276 14280 -3108
rect 14044 -3298 14096 -3288
rect 14332 -3276 14516 -3108
rect 14280 -3298 14332 -3288
rect 14568 -3276 14584 -3108
rect 15084 -3108 15624 -2816
rect 14516 -3298 14568 -3288
rect 15136 -3276 15320 -3108
rect 15084 -3298 15136 -3288
rect 15372 -3276 15556 -3108
rect 15320 -3298 15372 -3288
rect 15608 -3276 15624 -3108
rect 16124 -3108 16664 -2816
rect 15556 -3298 15608 -3288
rect 16176 -3276 16360 -3108
rect 16124 -3298 16176 -3288
rect 16412 -3276 16596 -3108
rect 16360 -3298 16412 -3288
rect 16648 -3276 16664 -3108
rect 16596 -3298 16648 -3288
rect -7238 -3478 -7054 -3310
rect -7290 -3500 -7238 -3490
rect -7002 -3478 -6818 -3310
rect -7054 -3500 -7002 -3490
rect -6766 -3478 -6750 -3310
rect 4224 -3332 4276 -3322
rect -6818 -3500 -6766 -3490
rect 4460 -3332 4512 -3322
rect 4276 -3512 4460 -3340
rect 4696 -3332 4748 -3322
rect 4512 -3512 4696 -3340
rect 4932 -3332 4984 -3322
rect 4748 -3360 4932 -3340
rect 5264 -3332 5316 -3322
rect 4984 -3360 5264 -3350
rect 5500 -3332 5552 -3322
rect 4748 -3512 4844 -3360
rect 5316 -3512 5500 -3340
rect 5736 -3332 5788 -3322
rect 5552 -3512 5736 -3340
rect 5972 -3332 6024 -3322
rect 5788 -3380 5972 -3340
rect 6304 -3332 6356 -3322
rect 6024 -3380 6304 -3350
rect 5788 -3512 5904 -3380
rect 6540 -3332 6592 -3322
rect 6356 -3512 6540 -3340
rect 6776 -3332 6828 -3322
rect 6592 -3512 6776 -3340
rect 7012 -3332 7064 -3322
rect 6828 -3380 7012 -3340
rect 7344 -3332 7396 -3322
rect 7064 -3380 7344 -3370
rect 6828 -3512 6924 -3380
rect 7580 -3332 7632 -3322
rect 7396 -3512 7580 -3340
rect 7816 -3332 7868 -3322
rect 7632 -3512 7816 -3340
rect 8052 -3332 8104 -3322
rect 7868 -3380 8052 -3340
rect 8384 -3332 8436 -3322
rect 8104 -3380 8384 -3370
rect 8620 -3332 8672 -3322
rect 7868 -3512 7984 -3380
rect 8436 -3512 8620 -3340
rect 8856 -3332 8908 -3322
rect 8672 -3512 8856 -3340
rect 9092 -3332 9144 -3322
rect 8908 -3380 9092 -3340
rect 11844 -3332 11896 -3322
rect 9144 -3380 9424 -3370
rect 8908 -3512 9004 -3380
rect -7410 -3534 -7358 -3524
rect -7420 -3580 -7410 -3570
rect -7174 -3534 -7122 -3524
rect -7358 -3580 -7174 -3542
rect -6938 -3534 -6886 -3524
rect -7122 -3580 -6938 -3542
rect -6702 -3534 -6650 -3524
rect -6886 -3580 -6702 -3542
rect -6650 -3580 -6620 -3570
rect 4224 -3612 4844 -3512
rect 5284 -3612 5904 -3512
rect 4844 -3630 5284 -3620
rect 5884 -3630 5904 -3612
rect 6304 -3612 6924 -3512
rect 6304 -3630 6324 -3612
rect 5904 -3710 6304 -3700
rect 7344 -3612 7984 -3512
rect 6924 -3710 7344 -3700
rect 8404 -3612 9004 -3512
rect 7984 -3710 8404 -3700
rect 12080 -3332 12132 -3322
rect 11896 -3512 12080 -3340
rect 12316 -3332 12368 -3322
rect 12132 -3512 12316 -3340
rect 12552 -3332 12604 -3322
rect 12368 -3360 12552 -3340
rect 12884 -3332 12936 -3322
rect 12604 -3360 12884 -3350
rect 13120 -3332 13172 -3322
rect 12368 -3512 12464 -3360
rect 12936 -3512 13120 -3340
rect 13356 -3332 13408 -3322
rect 13172 -3512 13356 -3340
rect 13592 -3332 13644 -3322
rect 13408 -3380 13592 -3340
rect 13924 -3332 13976 -3322
rect 13644 -3380 13924 -3350
rect 13408 -3512 13524 -3380
rect 14160 -3332 14212 -3322
rect 13976 -3512 14160 -3340
rect 14396 -3332 14448 -3322
rect 14212 -3512 14396 -3340
rect 14632 -3332 14684 -3322
rect 14448 -3380 14632 -3340
rect 14964 -3332 15016 -3322
rect 14684 -3380 14964 -3370
rect 14448 -3512 14544 -3380
rect 15200 -3332 15252 -3322
rect 15016 -3512 15200 -3340
rect 15436 -3332 15488 -3322
rect 15252 -3512 15436 -3340
rect 15672 -3332 15724 -3322
rect 15488 -3380 15672 -3340
rect 16004 -3332 16056 -3322
rect 15724 -3380 16004 -3370
rect 16240 -3332 16292 -3322
rect 15488 -3512 15604 -3380
rect 16056 -3512 16240 -3340
rect 16476 -3332 16528 -3322
rect 16292 -3512 16476 -3340
rect 16712 -3332 16764 -3322
rect 16528 -3380 16712 -3340
rect 16764 -3380 17044 -3370
rect 16528 -3512 16624 -3380
rect 11844 -3612 12464 -3512
rect 12904 -3612 13524 -3512
rect 12464 -3630 12904 -3620
rect 13504 -3630 13524 -3612
rect 9004 -3710 9424 -3700
rect 13924 -3612 14544 -3512
rect 13924 -3630 13944 -3612
rect 13524 -3710 13924 -3700
rect 14964 -3612 15604 -3512
rect 14544 -3710 14964 -3700
rect 16024 -3612 16624 -3512
rect 15604 -3710 16024 -3700
rect 16624 -3710 17044 -3700
rect 4924 -3720 5224 -3710
rect 4924 -3850 5224 -3840
rect 8564 -3720 8864 -3710
rect 8564 -3850 8864 -3840
rect 12544 -3720 12844 -3710
rect 12544 -3850 12844 -3840
rect 16184 -3720 16484 -3710
rect 16184 -3850 16484 -3840
rect -7420 -3970 -7230 -3960
rect -6950 -3970 -6620 -3960
rect -7230 -3992 -6950 -3982
<< via2 >>
rect -1440 6580 -1080 6740
rect -1440 6184 -1080 6580
rect -1440 5212 -1080 6184
rect 0 6588 360 6720
rect 0 6192 360 6588
rect -1440 4860 -1080 5212
rect 0 5220 360 6192
rect 0 4840 360 5220
rect 1360 6580 1720 6740
rect 1360 6184 1720 6580
rect 1360 5212 1720 6184
rect 2800 6588 3160 6720
rect 2800 6192 3160 6588
rect 1360 4860 1720 5212
rect 2800 5220 3160 6192
rect 4864 5468 5264 5540
rect 5884 5468 6284 5540
rect 6924 5468 7324 5540
rect 4864 5320 4904 5468
rect 4904 5320 4956 5468
rect 4956 5320 5096 5468
rect 5096 5320 5148 5468
rect 5148 5320 5264 5468
rect 5884 5320 5916 5468
rect 5916 5320 6056 5468
rect 6056 5320 6108 5468
rect 6108 5320 6248 5468
rect 6248 5320 6284 5468
rect 6924 5320 7016 5468
rect 7016 5320 7068 5468
rect 7068 5320 7208 5468
rect 7208 5320 7260 5468
rect 7260 5320 7324 5468
rect 8004 5468 8404 5540
rect 9024 5468 9424 5540
rect 10044 5468 10444 5540
rect 8004 5320 8160 5468
rect 8160 5320 8212 5468
rect 8212 5320 8352 5468
rect 8352 5320 8404 5468
rect 9024 5320 9120 5468
rect 9120 5320 9172 5468
rect 9172 5320 9312 5468
rect 9312 5320 9364 5468
rect 9364 5320 9424 5468
rect 10044 5320 10080 5468
rect 10080 5320 10132 5468
rect 10132 5320 10272 5468
rect 10272 5320 10324 5468
rect 10324 5320 10444 5468
rect 12484 5468 12884 5540
rect 13504 5468 13904 5540
rect 14544 5468 14944 5540
rect 12484 5320 12524 5468
rect 12524 5320 12576 5468
rect 12576 5320 12716 5468
rect 12716 5320 12768 5468
rect 12768 5320 12884 5468
rect 13504 5320 13536 5468
rect 13536 5320 13676 5468
rect 13676 5320 13728 5468
rect 13728 5320 13868 5468
rect 13868 5320 13904 5468
rect 14544 5320 14636 5468
rect 14636 5320 14688 5468
rect 14688 5320 14828 5468
rect 14828 5320 14880 5468
rect 14880 5320 14944 5468
rect 15624 5468 16024 5540
rect 16644 5468 17044 5540
rect 17664 5468 18064 5540
rect 15624 5320 15780 5468
rect 15780 5320 15832 5468
rect 15832 5320 15972 5468
rect 15972 5320 16024 5468
rect 16644 5320 16740 5468
rect 16740 5320 16792 5468
rect 16792 5320 16932 5468
rect 16932 5320 16984 5468
rect 16984 5320 17044 5468
rect 17664 5320 17700 5468
rect 17700 5320 17752 5468
rect 17752 5320 17892 5468
rect 17892 5320 17944 5468
rect 17944 5320 18064 5468
rect 2800 4840 3160 5220
rect 4304 5064 4424 5220
rect 4424 5064 4476 5220
rect 4476 5064 4616 5220
rect 4616 5064 4668 5220
rect 4668 5064 4744 5220
rect 5384 5064 5436 5200
rect 5436 5064 5576 5200
rect 5576 5064 5628 5200
rect 5628 5064 5768 5200
rect 5768 5064 5784 5200
rect 6424 5064 6536 5200
rect 6536 5064 6588 5200
rect 6588 5064 6728 5200
rect 6728 5064 6780 5200
rect 6780 5064 6824 5200
rect 4304 4980 4744 5064
rect 5384 4980 5784 5064
rect 6424 4980 6824 5064
rect 7464 4980 7864 5200
rect 8504 5064 8640 5220
rect 8640 5064 8692 5220
rect 8692 5064 8832 5220
rect 8832 5064 8884 5220
rect 8884 5064 8904 5220
rect 9544 5064 9600 5220
rect 9600 5064 9652 5220
rect 9652 5064 9792 5220
rect 9792 5064 9844 5220
rect 9844 5064 9944 5220
rect 10584 5064 10612 5220
rect 10612 5064 10752 5220
rect 10752 5064 10804 5220
rect 10804 5064 10944 5220
rect 10944 5064 10984 5220
rect 8504 5000 8904 5064
rect 9544 5000 9944 5064
rect 10584 5000 10984 5064
rect 11924 5064 12044 5220
rect 12044 5064 12096 5220
rect 12096 5064 12236 5220
rect 12236 5064 12288 5220
rect 12288 5064 12364 5220
rect 13004 5064 13056 5200
rect 13056 5064 13196 5200
rect 13196 5064 13248 5200
rect 13248 5064 13388 5200
rect 13388 5064 13404 5200
rect 14044 5064 14156 5200
rect 14156 5064 14208 5200
rect 14208 5064 14348 5200
rect 14348 5064 14400 5200
rect 14400 5064 14444 5200
rect 11924 4980 12364 5064
rect 13004 4980 13404 5064
rect 14044 4980 14444 5064
rect 15084 4980 15484 5200
rect 16124 5064 16260 5220
rect 16260 5064 16312 5220
rect 16312 5064 16452 5220
rect 16452 5064 16504 5220
rect 16504 5064 16524 5220
rect 17164 5064 17220 5220
rect 17220 5064 17272 5220
rect 17272 5064 17412 5220
rect 17412 5064 17464 5220
rect 17464 5064 17564 5220
rect 18204 5064 18232 5220
rect 18232 5064 18372 5220
rect 18372 5064 18424 5220
rect 18424 5064 18564 5220
rect 18564 5064 18604 5220
rect 16124 5000 16524 5064
rect 17164 5000 17564 5064
rect 18204 5000 18604 5064
rect 4864 4848 5264 4920
rect 5884 4848 6284 4920
rect 6924 4848 7324 4920
rect 4864 4700 4904 4848
rect 4904 4700 4956 4848
rect 4956 4700 5096 4848
rect 5096 4700 5148 4848
rect 5148 4700 5264 4848
rect 5884 4700 5916 4848
rect 5916 4700 6056 4848
rect 6056 4700 6108 4848
rect 6108 4700 6248 4848
rect 6248 4700 6284 4848
rect 6924 4700 7016 4848
rect 7016 4700 7068 4848
rect 7068 4700 7208 4848
rect 7208 4700 7260 4848
rect 7260 4700 7324 4848
rect 8004 4848 8404 4920
rect 9024 4848 9424 4920
rect 10044 4848 10444 4920
rect 8004 4700 8160 4848
rect 8160 4700 8212 4848
rect 8212 4700 8352 4848
rect 8352 4700 8404 4848
rect 9024 4700 9120 4848
rect 9120 4700 9172 4848
rect 9172 4700 9312 4848
rect 9312 4700 9364 4848
rect 9364 4700 9424 4848
rect 10044 4700 10080 4848
rect 10080 4700 10132 4848
rect 10132 4700 10272 4848
rect 10272 4700 10324 4848
rect 10324 4700 10444 4848
rect 12484 4848 12884 4920
rect 13504 4848 13904 4920
rect 14544 4848 14944 4920
rect 12484 4700 12524 4848
rect 12524 4700 12576 4848
rect 12576 4700 12716 4848
rect 12716 4700 12768 4848
rect 12768 4700 12884 4848
rect 13504 4700 13536 4848
rect 13536 4700 13676 4848
rect 13676 4700 13728 4848
rect 13728 4700 13868 4848
rect 13868 4700 13904 4848
rect 14544 4700 14636 4848
rect 14636 4700 14688 4848
rect 14688 4700 14828 4848
rect 14828 4700 14880 4848
rect 14880 4700 14944 4848
rect 15624 4848 16024 4920
rect 16644 4848 17044 4920
rect 17664 4848 18064 4920
rect 15624 4700 15780 4848
rect 15780 4700 15832 4848
rect 15832 4700 15972 4848
rect 15972 4700 16024 4848
rect 16644 4700 16740 4848
rect 16740 4700 16792 4848
rect 16792 4700 16932 4848
rect 16932 4700 16984 4848
rect 16984 4700 17044 4848
rect 17664 4700 17700 4848
rect 17700 4700 17752 4848
rect 17752 4700 17892 4848
rect 17892 4700 17944 4848
rect 17944 4700 18064 4848
rect 4304 4444 4424 4600
rect 4424 4444 4476 4600
rect 4476 4444 4616 4600
rect 4616 4444 4668 4600
rect 4668 4444 4744 4600
rect 5384 4444 5436 4600
rect 5436 4444 5576 4600
rect 5576 4444 5628 4600
rect 5628 4444 5768 4600
rect 5768 4444 5784 4600
rect 6424 4444 6536 4600
rect 6536 4444 6588 4600
rect 6588 4444 6728 4600
rect 6728 4444 6780 4600
rect 6780 4444 6824 4600
rect 4304 4380 4744 4444
rect 5384 4380 5784 4444
rect 6424 4380 6824 4444
rect 7464 4380 7864 4600
rect 8504 4444 8640 4600
rect 8640 4444 8692 4600
rect 8692 4444 8832 4600
rect 8832 4444 8884 4600
rect 8884 4444 8904 4600
rect 9544 4444 9600 4600
rect 9600 4444 9652 4600
rect 9652 4444 9792 4600
rect 9792 4444 9844 4600
rect 9844 4444 9944 4600
rect 10584 4444 10612 4600
rect 10612 4444 10752 4600
rect 10752 4444 10804 4600
rect 10804 4444 10944 4600
rect 10944 4444 10984 4600
rect 8504 4380 8904 4444
rect 9544 4380 9944 4444
rect 10584 4380 10984 4444
rect 11924 4444 12044 4600
rect 12044 4444 12096 4600
rect 12096 4444 12236 4600
rect 12236 4444 12288 4600
rect 12288 4444 12364 4600
rect 13004 4444 13056 4600
rect 13056 4444 13196 4600
rect 13196 4444 13248 4600
rect 13248 4444 13388 4600
rect 13388 4444 13404 4600
rect 14044 4444 14156 4600
rect 14156 4444 14208 4600
rect 14208 4444 14348 4600
rect 14348 4444 14400 4600
rect 14400 4444 14444 4600
rect 11924 4380 12364 4444
rect 13004 4380 13404 4444
rect 14044 4380 14444 4444
rect 15084 4380 15484 4600
rect 16124 4444 16260 4600
rect 16260 4444 16312 4600
rect 16312 4444 16452 4600
rect 16452 4444 16504 4600
rect 16504 4444 16524 4600
rect 17164 4444 17220 4600
rect 17220 4444 17272 4600
rect 17272 4444 17412 4600
rect 17412 4444 17464 4600
rect 17464 4444 17564 4600
rect 18204 4444 18232 4600
rect 18232 4444 18372 4600
rect 18372 4444 18424 4600
rect 18424 4444 18564 4600
rect 18564 4444 18604 4600
rect 16124 4380 16524 4444
rect 17164 4380 17564 4444
rect 18204 4380 18604 4444
rect 4864 4232 5264 4300
rect 5884 4232 6284 4300
rect 6924 4232 7324 4300
rect 4864 4080 4904 4232
rect 4904 4080 4956 4232
rect 4956 4080 5096 4232
rect 5096 4080 5148 4232
rect 5148 4080 5264 4232
rect 5884 4080 5916 4232
rect 5916 4080 6056 4232
rect 6056 4080 6108 4232
rect 6108 4080 6248 4232
rect 6248 4080 6284 4232
rect 6924 4080 7016 4232
rect 7016 4080 7068 4232
rect 7068 4080 7208 4232
rect 7208 4080 7260 4232
rect 7260 4080 7324 4232
rect 8004 4232 8404 4300
rect 9024 4232 9424 4300
rect 10044 4232 10444 4300
rect 8004 4080 8160 4232
rect 8160 4080 8212 4232
rect 8212 4080 8352 4232
rect 8352 4080 8404 4232
rect 9024 4080 9120 4232
rect 9120 4080 9172 4232
rect 9172 4080 9312 4232
rect 9312 4080 9364 4232
rect 9364 4080 9424 4232
rect 10044 4080 10080 4232
rect 10080 4080 10132 4232
rect 10132 4080 10272 4232
rect 10272 4080 10324 4232
rect 10324 4080 10444 4232
rect 12484 4232 12884 4300
rect 13504 4232 13904 4300
rect 14544 4232 14944 4300
rect 12484 4080 12524 4232
rect 12524 4080 12576 4232
rect 12576 4080 12716 4232
rect 12716 4080 12768 4232
rect 12768 4080 12884 4232
rect 13504 4080 13536 4232
rect 13536 4080 13676 4232
rect 13676 4080 13728 4232
rect 13728 4080 13868 4232
rect 13868 4080 13904 4232
rect 14544 4080 14636 4232
rect 14636 4080 14688 4232
rect 14688 4080 14828 4232
rect 14828 4080 14880 4232
rect 14880 4080 14944 4232
rect 15624 4232 16024 4300
rect 16644 4232 17044 4300
rect 17664 4232 18064 4300
rect 15624 4080 15780 4232
rect 15780 4080 15832 4232
rect 15832 4080 15972 4232
rect 15972 4080 16024 4232
rect 16644 4080 16740 4232
rect 16740 4080 16792 4232
rect 16792 4080 16932 4232
rect 16932 4080 16984 4232
rect 16984 4080 17044 4232
rect 17664 4080 17700 4232
rect 17700 4080 17752 4232
rect 17752 4080 17892 4232
rect 17892 4080 17944 4232
rect 17944 4080 18064 4232
rect 4304 3828 4424 3980
rect 4424 3828 4476 3980
rect 4476 3828 4616 3980
rect 4616 3828 4668 3980
rect 4668 3828 4744 3980
rect 5384 3828 5436 3980
rect 5436 3828 5576 3980
rect 5576 3828 5628 3980
rect 5628 3828 5768 3980
rect 5768 3828 5784 3980
rect 6424 3828 6536 3980
rect 6536 3828 6588 3980
rect 6588 3828 6728 3980
rect 6728 3828 6780 3980
rect 6780 3828 6824 3980
rect 4304 3760 4744 3828
rect 5384 3760 5784 3828
rect 6424 3760 6824 3828
rect 7464 3760 7864 3980
rect 8504 3828 8640 3980
rect 8640 3828 8692 3980
rect 8692 3828 8832 3980
rect 8832 3828 8884 3980
rect 8884 3828 8904 3980
rect 9544 3828 9600 3980
rect 9600 3828 9652 3980
rect 9652 3828 9792 3980
rect 9792 3828 9844 3980
rect 9844 3828 9944 3980
rect 10584 3828 10612 3980
rect 10612 3828 10752 3980
rect 10752 3828 10804 3980
rect 10804 3828 10944 3980
rect 10944 3828 10984 3980
rect 8504 3760 8904 3828
rect 9544 3760 9944 3828
rect 10584 3760 10984 3828
rect 11924 3828 12044 3980
rect 12044 3828 12096 3980
rect 12096 3828 12236 3980
rect 12236 3828 12288 3980
rect 12288 3828 12364 3980
rect 13004 3828 13056 3980
rect 13056 3828 13196 3980
rect 13196 3828 13248 3980
rect 13248 3828 13388 3980
rect 13388 3828 13404 3980
rect 14044 3828 14156 3980
rect 14156 3828 14208 3980
rect 14208 3828 14348 3980
rect 14348 3828 14400 3980
rect 14400 3828 14444 3980
rect 11924 3760 12364 3828
rect 13004 3760 13404 3828
rect 14044 3760 14444 3828
rect 15084 3760 15484 3980
rect 16124 3828 16260 3980
rect 16260 3828 16312 3980
rect 16312 3828 16452 3980
rect 16452 3828 16504 3980
rect 16504 3828 16524 3980
rect 17164 3828 17220 3980
rect 17220 3828 17272 3980
rect 17272 3828 17412 3980
rect 17412 3828 17464 3980
rect 17464 3828 17564 3980
rect 18204 3828 18232 3980
rect 18232 3828 18372 3980
rect 18372 3828 18424 3980
rect 18424 3828 18564 3980
rect 18564 3828 18604 3980
rect 16124 3760 16524 3828
rect 17164 3760 17564 3828
rect 18204 3760 18604 3828
rect 4864 3612 5264 3680
rect 5884 3612 6284 3680
rect 6924 3612 7324 3680
rect 4864 3460 4904 3612
rect 4904 3460 4956 3612
rect 4956 3460 5096 3612
rect 5096 3460 5148 3612
rect 5148 3460 5264 3612
rect 5884 3460 5916 3612
rect 5916 3460 6056 3612
rect 6056 3460 6108 3612
rect 6108 3460 6248 3612
rect 6248 3460 6284 3612
rect 6924 3460 7016 3612
rect 7016 3460 7068 3612
rect 7068 3460 7208 3612
rect 7208 3460 7260 3612
rect 7260 3460 7324 3612
rect 8004 3612 8404 3680
rect 9024 3612 9424 3680
rect 10044 3612 10444 3680
rect 8004 3460 8160 3612
rect 8160 3460 8212 3612
rect 8212 3460 8352 3612
rect 8352 3460 8404 3612
rect 9024 3460 9120 3612
rect 9120 3460 9172 3612
rect 9172 3460 9312 3612
rect 9312 3460 9364 3612
rect 9364 3460 9424 3612
rect 10044 3460 10080 3612
rect 10080 3460 10132 3612
rect 10132 3460 10272 3612
rect 10272 3460 10324 3612
rect 10324 3460 10444 3612
rect 12484 3612 12884 3680
rect 13504 3612 13904 3680
rect 14544 3612 14944 3680
rect 12484 3460 12524 3612
rect 12524 3460 12576 3612
rect 12576 3460 12716 3612
rect 12716 3460 12768 3612
rect 12768 3460 12884 3612
rect 13504 3460 13536 3612
rect 13536 3460 13676 3612
rect 13676 3460 13728 3612
rect 13728 3460 13868 3612
rect 13868 3460 13904 3612
rect 14544 3460 14636 3612
rect 14636 3460 14688 3612
rect 14688 3460 14828 3612
rect 14828 3460 14880 3612
rect 14880 3460 14944 3612
rect 15624 3612 16024 3680
rect 16644 3612 17044 3680
rect 17664 3612 18064 3680
rect 15624 3460 15780 3612
rect 15780 3460 15832 3612
rect 15832 3460 15972 3612
rect 15972 3460 16024 3612
rect 16644 3460 16740 3612
rect 16740 3460 16792 3612
rect 16792 3460 16932 3612
rect 16932 3460 16984 3612
rect 16984 3460 17044 3612
rect 17664 3460 17700 3612
rect 17700 3460 17752 3612
rect 17752 3460 17892 3612
rect 17892 3460 17944 3612
rect 17944 3460 18064 3612
rect -1140 3212 -1040 3280
rect -1040 3212 -988 3280
rect -988 3212 -848 3280
rect -848 3212 -796 3280
rect -796 3212 -656 3280
rect -656 3212 -604 3280
rect -604 3212 -464 3280
rect -464 3212 -412 3280
rect -412 3212 -272 3280
rect -272 3212 -220 3280
rect -220 3212 -80 3280
rect -80 3212 -28 3280
rect -28 3212 60 3280
rect -1140 2780 60 3212
rect 1660 3212 1760 3280
rect 1760 3212 1812 3280
rect 1812 3212 1952 3280
rect 1952 3212 2004 3280
rect 2004 3212 2144 3280
rect 2144 3212 2196 3280
rect 2196 3212 2336 3280
rect 2336 3212 2388 3280
rect 2388 3212 2528 3280
rect 2528 3212 2580 3280
rect 2580 3212 2720 3280
rect 2720 3212 2772 3280
rect 2772 3212 2860 3280
rect 1660 2780 2860 3212
rect 4304 3208 4424 3360
rect 4424 3208 4476 3360
rect 4476 3208 4616 3360
rect 4616 3208 4668 3360
rect 4668 3208 4744 3360
rect 5384 3208 5436 3360
rect 5436 3208 5576 3360
rect 5576 3208 5628 3360
rect 5628 3208 5768 3360
rect 5768 3208 5784 3360
rect 6424 3208 6536 3360
rect 6536 3208 6588 3360
rect 6588 3208 6728 3360
rect 6728 3208 6780 3360
rect 6780 3208 6824 3360
rect 4304 3140 4744 3208
rect 5384 3140 5784 3208
rect 6424 3140 6824 3208
rect 7464 3140 7864 3360
rect 8504 3208 8640 3360
rect 8640 3208 8692 3360
rect 8692 3208 8832 3360
rect 8832 3208 8884 3360
rect 8884 3208 8904 3360
rect 9544 3208 9600 3360
rect 9600 3208 9652 3360
rect 9652 3208 9792 3360
rect 9792 3208 9844 3360
rect 9844 3208 9944 3360
rect 10584 3208 10612 3360
rect 10612 3208 10752 3360
rect 10752 3208 10804 3360
rect 10804 3208 10944 3360
rect 10944 3208 10984 3360
rect 8504 3140 8904 3208
rect 9544 3140 9944 3208
rect 10584 3140 10984 3208
rect 11924 3208 12044 3360
rect 12044 3208 12096 3360
rect 12096 3208 12236 3360
rect 12236 3208 12288 3360
rect 12288 3208 12364 3360
rect 13004 3208 13056 3360
rect 13056 3208 13196 3360
rect 13196 3208 13248 3360
rect 13248 3208 13388 3360
rect 13388 3208 13404 3360
rect 14044 3208 14156 3360
rect 14156 3208 14208 3360
rect 14208 3208 14348 3360
rect 14348 3208 14400 3360
rect 14400 3208 14444 3360
rect 11924 3140 12364 3208
rect 13004 3140 13404 3208
rect 14044 3140 14444 3208
rect 15084 3140 15484 3360
rect 16124 3208 16260 3360
rect 16260 3208 16312 3360
rect 16312 3208 16452 3360
rect 16452 3208 16504 3360
rect 16504 3208 16524 3360
rect 17164 3208 17220 3360
rect 17220 3208 17272 3360
rect 17272 3208 17412 3360
rect 17412 3208 17464 3360
rect 17464 3208 17564 3360
rect 18204 3208 18232 3360
rect 18232 3208 18372 3360
rect 18372 3208 18424 3360
rect 18424 3208 18564 3360
rect 18564 3208 18604 3360
rect 16124 3140 16524 3208
rect 17164 3140 17564 3208
rect 18204 3140 18604 3208
rect -1484 2232 -1432 2372
rect -1432 2232 -1292 2372
rect -1292 2232 -1240 2372
rect -1240 2232 -1100 2372
rect -1100 2232 -1092 2372
rect -1484 2016 -1092 2232
rect -1484 1880 -1432 2016
rect -1432 1880 -1292 2016
rect -1292 1880 -1240 2016
rect -1240 1880 -1100 2016
rect -1100 1880 -1092 2016
rect -440 2232 -392 2380
rect -392 2232 -252 2380
rect -252 2232 -200 2380
rect -200 2232 -60 2380
rect -60 2232 -48 2380
rect -440 2016 -48 2232
rect -440 1888 -392 2016
rect -392 1888 -252 2016
rect -252 1888 -200 2016
rect -200 1888 -60 2016
rect -60 1888 -48 2016
rect 604 2232 648 2376
rect 648 2232 788 2376
rect 788 2232 840 2376
rect 840 2232 980 2376
rect 980 2232 996 2376
rect 604 2016 996 2232
rect 604 1884 648 2016
rect 648 1884 788 2016
rect 788 1884 840 2016
rect 840 1884 980 2016
rect 980 1884 996 2016
rect 1648 2232 1688 2372
rect 1688 2232 1828 2372
rect 1828 2232 1880 2372
rect 1880 2232 2020 2372
rect 2020 2232 2040 2372
rect 1648 2016 2040 2232
rect 1648 1880 1688 2016
rect 1688 1880 1828 2016
rect 1828 1880 1880 2016
rect 1880 1880 2020 2016
rect 2020 1880 2040 2016
rect 2704 2232 2728 2372
rect 2728 2232 2868 2372
rect 2868 2232 2920 2372
rect 2920 2232 3060 2372
rect 3060 2232 3096 2372
rect 2704 2016 3096 2232
rect 2704 1880 2728 2016
rect 2728 1880 2868 2016
rect 2868 1880 2920 2016
rect 2920 1880 3060 2016
rect 3060 1880 3096 2016
rect 4328 2392 4372 2550
rect 4372 2392 4512 2550
rect 4512 2392 4564 2550
rect 4564 2392 4704 2550
rect 4704 2392 4748 2550
rect 4328 2176 4748 2392
rect 4328 2016 4372 2176
rect 4372 2016 4512 2176
rect 4512 2016 4564 2176
rect 4564 2016 4704 2176
rect 4704 2016 4748 2176
rect 5368 2392 5412 2550
rect 5412 2392 5552 2550
rect 5552 2392 5604 2550
rect 5604 2392 5744 2550
rect 5744 2392 5788 2550
rect 5368 2176 5788 2392
rect 5368 2016 5412 2176
rect 5412 2016 5552 2176
rect 5552 2016 5604 2176
rect 5604 2016 5744 2176
rect 5744 2016 5788 2176
rect 6408 2392 6452 2550
rect 6452 2392 6592 2550
rect 6592 2392 6644 2550
rect 6644 2392 6784 2550
rect 6784 2392 6828 2550
rect 6408 2176 6828 2392
rect 6408 2016 6452 2176
rect 6452 2016 6592 2176
rect 6592 2016 6644 2176
rect 6644 2016 6784 2176
rect 6784 2016 6828 2176
rect 7448 2392 7492 2550
rect 7492 2392 7632 2550
rect 7632 2392 7684 2550
rect 7684 2392 7824 2550
rect 7824 2392 7868 2550
rect 7448 2176 7868 2392
rect 7448 2016 7492 2176
rect 7492 2016 7632 2176
rect 7632 2016 7684 2176
rect 7684 2016 7824 2176
rect 7824 2016 7868 2176
rect 8488 2392 8532 2546
rect 8532 2392 8672 2546
rect 8672 2392 8724 2546
rect 8724 2392 8864 2546
rect 8864 2392 8908 2546
rect 8488 2176 8908 2392
rect 8488 2012 8532 2176
rect 8532 2012 8672 2176
rect 8672 2012 8724 2176
rect 8724 2012 8864 2176
rect 8864 2012 8908 2176
rect 9528 2392 9572 2550
rect 9572 2392 9712 2550
rect 9712 2392 9764 2550
rect 9764 2392 9904 2550
rect 9904 2392 9948 2550
rect 9528 2176 9948 2392
rect 9528 2016 9572 2176
rect 9572 2016 9712 2176
rect 9712 2016 9764 2176
rect 9764 2016 9904 2176
rect 9904 2016 9948 2176
rect 10568 2392 10612 2546
rect 10612 2392 10752 2546
rect 10752 2392 10804 2546
rect 10804 2392 10944 2546
rect 10944 2392 10988 2546
rect 10568 2176 10988 2392
rect 10568 2012 10612 2176
rect 10612 2012 10752 2176
rect 10752 2012 10804 2176
rect 10804 2012 10944 2176
rect 10944 2012 10988 2176
rect 11948 2392 11992 2550
rect 11992 2392 12132 2550
rect 12132 2392 12184 2550
rect 12184 2392 12324 2550
rect 12324 2392 12368 2550
rect 11948 2176 12368 2392
rect 11948 2016 11992 2176
rect 11992 2016 12132 2176
rect 12132 2016 12184 2176
rect 12184 2016 12324 2176
rect 12324 2016 12368 2176
rect 12988 2392 13032 2550
rect 13032 2392 13172 2550
rect 13172 2392 13224 2550
rect 13224 2392 13364 2550
rect 13364 2392 13408 2550
rect 12988 2176 13408 2392
rect 12988 2016 13032 2176
rect 13032 2016 13172 2176
rect 13172 2016 13224 2176
rect 13224 2016 13364 2176
rect 13364 2016 13408 2176
rect 14028 2392 14072 2550
rect 14072 2392 14212 2550
rect 14212 2392 14264 2550
rect 14264 2392 14404 2550
rect 14404 2392 14448 2550
rect 14028 2176 14448 2392
rect 14028 2016 14072 2176
rect 14072 2016 14212 2176
rect 14212 2016 14264 2176
rect 14264 2016 14404 2176
rect 14404 2016 14448 2176
rect 15068 2392 15112 2550
rect 15112 2392 15252 2550
rect 15252 2392 15304 2550
rect 15304 2392 15444 2550
rect 15444 2392 15488 2550
rect 15068 2176 15488 2392
rect 15068 2016 15112 2176
rect 15112 2016 15252 2176
rect 15252 2016 15304 2176
rect 15304 2016 15444 2176
rect 15444 2016 15488 2176
rect 16108 2392 16152 2546
rect 16152 2392 16292 2546
rect 16292 2392 16344 2546
rect 16344 2392 16484 2546
rect 16484 2392 16528 2546
rect 16108 2176 16528 2392
rect 16108 2012 16152 2176
rect 16152 2012 16292 2176
rect 16292 2012 16344 2176
rect 16344 2012 16484 2176
rect 16484 2012 16528 2176
rect 17148 2392 17192 2550
rect 17192 2392 17332 2550
rect 17332 2392 17384 2550
rect 17384 2392 17524 2550
rect 17524 2392 17568 2550
rect 17148 2176 17568 2392
rect 17148 2016 17192 2176
rect 17192 2016 17332 2176
rect 17332 2016 17384 2176
rect 17384 2016 17524 2176
rect 17524 2016 17568 2176
rect 18188 2392 18232 2546
rect 18232 2392 18372 2546
rect 18372 2392 18424 2546
rect 18424 2392 18564 2546
rect 18564 2392 18608 2546
rect 18188 2176 18608 2392
rect 18188 2012 18232 2176
rect 18232 2012 18372 2176
rect 18372 2012 18424 2176
rect 18424 2012 18564 2176
rect 18564 2012 18608 2176
rect -1540 808 -1528 920
rect -1528 808 -1344 920
rect -1344 808 -1292 920
rect -1292 808 -1108 920
rect -1108 808 -1056 920
rect -1056 808 -872 920
rect -872 808 -860 920
rect -1540 476 -860 808
rect -1540 440 -1308 476
rect -1308 440 -1128 476
rect -1128 440 -860 476
rect -5998 154 -5802 406
rect -500 808 -488 920
rect -488 808 -304 920
rect -304 808 -252 920
rect -252 808 -68 920
rect -68 808 -16 920
rect -16 808 168 920
rect 168 808 180 920
rect -500 440 180 808
rect 540 808 552 920
rect 552 808 736 920
rect 736 808 788 920
rect 788 808 972 920
rect 972 808 1024 920
rect 1024 808 1208 920
rect 1208 808 1220 920
rect 540 440 1220 808
rect 1580 808 1592 920
rect 1592 808 1776 920
rect 1776 808 1828 920
rect 1828 808 2012 920
rect 2012 808 2064 920
rect 2064 808 2248 920
rect 2248 808 2260 920
rect 1580 440 2260 808
rect 2620 808 2632 920
rect 2632 808 2816 920
rect 2816 808 2868 920
rect 2868 808 3052 920
rect 3052 808 3104 920
rect 3104 808 3288 920
rect 3288 808 3300 920
rect 2620 492 3300 808
rect 2620 440 2800 492
rect 2800 440 3068 492
rect 3068 440 3300 492
rect 4864 968 4932 1120
rect 4932 968 4984 1120
rect 4984 968 5264 1120
rect 5904 968 5972 1120
rect 5972 968 6024 1120
rect 6024 968 6304 1120
rect 6304 968 6324 1120
rect 6924 968 7012 1120
rect 7012 968 7064 1120
rect 7064 968 7344 1120
rect 7984 968 8052 1120
rect 8052 968 8104 1120
rect 8104 968 8384 1120
rect 8384 968 8404 1120
rect 9024 968 9092 1120
rect 9092 968 9144 1120
rect 9144 968 9424 1120
rect 9424 968 9444 1120
rect 10044 968 10132 1120
rect 10132 968 10184 1120
rect 10184 968 10464 1120
rect 4864 780 5264 968
rect 5904 800 6324 968
rect 6924 800 7344 968
rect 7984 800 8404 968
rect 9024 800 9444 968
rect 10044 800 10464 968
rect 12484 968 12552 1120
rect 12552 968 12604 1120
rect 12604 968 12884 1120
rect 13524 968 13592 1120
rect 13592 968 13644 1120
rect 13644 968 13924 1120
rect 13924 968 13944 1120
rect 14544 968 14632 1120
rect 14632 968 14684 1120
rect 14684 968 14964 1120
rect 15604 968 15672 1120
rect 15672 968 15724 1120
rect 15724 968 16004 1120
rect 16004 968 16024 1120
rect 16644 968 16712 1120
rect 16712 968 16764 1120
rect 16764 968 17044 1120
rect 17044 968 17064 1120
rect 17664 968 17752 1120
rect 17752 968 17804 1120
rect 17804 968 18084 1120
rect 12484 780 12884 968
rect 13524 800 13944 968
rect 14544 800 14964 968
rect 15604 800 16024 968
rect 16644 800 17064 968
rect 17664 800 18084 968
rect -7030 -54 -6698 22
rect -7030 -210 -6930 -54
rect -6930 -210 -6878 -54
rect -6878 -210 -6738 -54
rect -6738 -210 -6698 -54
rect 3712 -140 3912 76
rect -7478 -454 -7410 -294
rect -7410 -454 -7358 -294
rect -7358 -454 -7218 -294
rect -7218 -454 -7166 -294
rect -7166 -454 -7146 -294
rect -7478 -526 -7146 -454
rect 4332 152 4372 310
rect 4372 152 4512 310
rect 4512 152 4564 310
rect 4564 152 4704 310
rect 4704 152 4752 310
rect 4332 -64 4752 152
rect 4332 -224 4372 -64
rect 4372 -224 4512 -64
rect 4512 -224 4564 -64
rect 4564 -224 4704 -64
rect 4704 -224 4752 -64
rect 5376 152 5412 310
rect 5412 152 5552 310
rect 5552 152 5604 310
rect 5604 152 5744 310
rect 5744 152 5796 310
rect 5376 -64 5796 152
rect 5376 -224 5412 -64
rect 5412 -224 5552 -64
rect 5552 -224 5604 -64
rect 5604 -224 5744 -64
rect 5744 -224 5796 -64
rect 6412 152 6452 310
rect 6452 152 6592 310
rect 6592 152 6644 310
rect 6644 152 6784 310
rect 6784 152 6832 310
rect 6412 -64 6832 152
rect 6412 -224 6452 -64
rect 6452 -224 6592 -64
rect 6592 -224 6644 -64
rect 6644 -224 6784 -64
rect 6784 -224 6832 -64
rect 7452 152 7492 310
rect 7492 152 7632 310
rect 7632 152 7684 310
rect 7684 152 7824 310
rect 7824 152 7872 310
rect 7452 -64 7872 152
rect 7452 -224 7492 -64
rect 7492 -224 7632 -64
rect 7632 -224 7684 -64
rect 7684 -224 7824 -64
rect 7824 -224 7872 -64
rect 8488 152 8532 310
rect 8532 152 8672 310
rect 8672 152 8724 310
rect 8724 152 8864 310
rect 8864 152 8908 310
rect 8488 -64 8908 152
rect 8488 -224 8532 -64
rect 8532 -224 8672 -64
rect 8672 -224 8724 -64
rect 8724 -224 8864 -64
rect 8864 -224 8908 -64
rect 9520 152 9572 310
rect 9572 152 9712 310
rect 9712 152 9764 310
rect 9764 152 9904 310
rect 9904 152 9940 310
rect 9520 -64 9940 152
rect 9520 -224 9572 -64
rect 9572 -224 9712 -64
rect 9712 -224 9764 -64
rect 9764 -224 9904 -64
rect 9904 -224 9940 -64
rect 10560 152 10612 310
rect 10612 152 10752 310
rect 10752 152 10804 310
rect 10804 152 10944 310
rect 10944 152 10980 310
rect 10560 -64 10980 152
rect 10560 -224 10612 -64
rect 10612 -224 10752 -64
rect 10752 -224 10804 -64
rect 10804 -224 10944 -64
rect 10944 -224 10980 -64
rect 11952 152 11992 310
rect 11992 152 12132 310
rect 12132 152 12184 310
rect 12184 152 12324 310
rect 12324 152 12372 310
rect 11952 -64 12372 152
rect 11952 -224 11992 -64
rect 11992 -224 12132 -64
rect 12132 -224 12184 -64
rect 12184 -224 12324 -64
rect 12324 -224 12372 -64
rect 12996 152 13032 310
rect 13032 152 13172 310
rect 13172 152 13224 310
rect 13224 152 13364 310
rect 13364 152 13416 310
rect 12996 -64 13416 152
rect 12996 -224 13032 -64
rect 13032 -224 13172 -64
rect 13172 -224 13224 -64
rect 13224 -224 13364 -64
rect 13364 -224 13416 -64
rect 14032 152 14072 310
rect 14072 152 14212 310
rect 14212 152 14264 310
rect 14264 152 14404 310
rect 14404 152 14452 310
rect 14032 -64 14452 152
rect 14032 -224 14072 -64
rect 14072 -224 14212 -64
rect 14212 -224 14264 -64
rect 14264 -224 14404 -64
rect 14404 -224 14452 -64
rect 15072 152 15112 310
rect 15112 152 15252 310
rect 15252 152 15304 310
rect 15304 152 15444 310
rect 15444 152 15492 310
rect 15072 -64 15492 152
rect 15072 -224 15112 -64
rect 15112 -224 15252 -64
rect 15252 -224 15304 -64
rect 15304 -224 15444 -64
rect 15444 -224 15492 -64
rect 16108 152 16152 310
rect 16152 152 16292 310
rect 16292 152 16344 310
rect 16344 152 16484 310
rect 16484 152 16528 310
rect 16108 -64 16528 152
rect 16108 -224 16152 -64
rect 16152 -224 16292 -64
rect 16292 -224 16344 -64
rect 16344 -224 16484 -64
rect 16484 -224 16528 -64
rect 17140 152 17192 310
rect 17192 152 17332 310
rect 17332 152 17384 310
rect 17384 152 17524 310
rect 17524 152 17560 310
rect 17140 -64 17560 152
rect 17140 -224 17192 -64
rect 17192 -224 17332 -64
rect 17332 -224 17384 -64
rect 17384 -224 17524 -64
rect 17524 -224 17560 -64
rect 18180 152 18232 310
rect 18232 152 18372 310
rect 18372 152 18424 310
rect 18424 152 18564 310
rect 18564 152 18600 310
rect 18180 -64 18600 152
rect 18180 -224 18232 -64
rect 18232 -224 18372 -64
rect 18372 -224 18424 -64
rect 18424 -224 18564 -64
rect 18564 -224 18600 -64
rect -7030 -670 -6698 -598
rect -7030 -830 -6930 -670
rect -6930 -830 -6878 -670
rect -6878 -830 -6738 -670
rect -6738 -830 -6698 -670
rect -7478 -1074 -7410 -918
rect -7410 -1074 -7358 -918
rect -7358 -1074 -7218 -918
rect -7218 -1074 -7166 -918
rect -7166 -1074 -7146 -918
rect -7478 -1150 -7146 -1074
rect 4844 -1272 4932 -1120
rect 4932 -1272 4984 -1120
rect 4984 -1272 5264 -1120
rect 5904 -1272 5972 -1120
rect 5972 -1272 6024 -1120
rect 6024 -1272 6304 -1120
rect 6304 -1272 6324 -1120
rect 6924 -1272 7012 -1120
rect 7012 -1272 7064 -1120
rect 7064 -1272 7344 -1120
rect 7984 -1272 8052 -1120
rect 8052 -1272 8104 -1120
rect 8104 -1272 8384 -1120
rect 8384 -1272 8404 -1120
rect 9004 -1272 9092 -1120
rect 9092 -1272 9144 -1120
rect 9144 -1272 9424 -1120
rect 10044 -1272 10132 -1120
rect 10132 -1272 10184 -1120
rect 10184 -1272 10464 -1120
rect 4844 -1440 5264 -1272
rect 5904 -1440 6324 -1272
rect 6924 -1440 7344 -1272
rect 7984 -1440 8404 -1272
rect 9004 -1440 9424 -1272
rect 10044 -1440 10464 -1272
rect 12464 -1272 12552 -1120
rect 12552 -1272 12604 -1120
rect 12604 -1272 12884 -1120
rect 13524 -1272 13592 -1120
rect 13592 -1272 13644 -1120
rect 13644 -1272 13924 -1120
rect 13924 -1272 13944 -1120
rect 14544 -1272 14632 -1120
rect 14632 -1272 14684 -1120
rect 14684 -1272 14964 -1120
rect 15604 -1272 15672 -1120
rect 15672 -1272 15724 -1120
rect 15724 -1272 16004 -1120
rect 16004 -1272 16024 -1120
rect 16624 -1272 16712 -1120
rect 16712 -1272 16764 -1120
rect 16764 -1272 17044 -1120
rect 17664 -1272 17752 -1120
rect 17752 -1272 17804 -1120
rect 17804 -1272 18084 -1120
rect 12464 -1440 12884 -1272
rect 13524 -1440 13944 -1272
rect 14544 -1440 14964 -1272
rect 15604 -1440 16024 -1272
rect 16624 -1440 17044 -1272
rect 17664 -1440 18084 -1272
rect -7298 -2290 -7262 -2154
rect -7262 -2290 -7122 -2154
rect -7122 -2290 -7070 -2154
rect -7070 -2290 -6930 -2154
rect -6930 -2290 -6910 -2154
rect -7298 -2506 -6910 -2290
rect -7298 -2646 -7262 -2506
rect -7262 -2646 -7122 -2506
rect -7122 -2646 -7070 -2506
rect -7070 -2646 -6930 -2506
rect -6930 -2646 -6910 -2506
rect 4332 -2088 4372 -1936
rect 4372 -2088 4512 -1936
rect 4512 -2088 4564 -1936
rect 4564 -2088 4704 -1936
rect 4704 -2088 4732 -1936
rect 4332 -2304 4732 -2088
rect 4332 -2460 4372 -2304
rect 4372 -2460 4512 -2304
rect 4512 -2460 4564 -2304
rect 4564 -2460 4704 -2304
rect 4704 -2460 4732 -2304
rect 5372 -2088 5412 -1936
rect 5412 -2088 5552 -1936
rect 5552 -2088 5604 -1936
rect 5604 -2088 5744 -1936
rect 5744 -2088 5772 -1936
rect 5372 -2304 5772 -2088
rect 5372 -2460 5412 -2304
rect 5412 -2460 5552 -2304
rect 5552 -2460 5604 -2304
rect 5604 -2460 5744 -2304
rect 5744 -2460 5772 -2304
rect 6412 -2088 6452 -1936
rect 6452 -2088 6592 -1936
rect 6592 -2088 6644 -1936
rect 6644 -2088 6784 -1936
rect 6784 -2088 6812 -1936
rect 6412 -2304 6812 -2088
rect 6412 -2460 6452 -2304
rect 6452 -2460 6592 -2304
rect 6592 -2460 6644 -2304
rect 6644 -2460 6784 -2304
rect 6784 -2460 6812 -2304
rect 7452 -2088 7492 -1936
rect 7492 -2088 7632 -1936
rect 7632 -2088 7684 -1936
rect 7684 -2088 7824 -1936
rect 7824 -2088 7852 -1936
rect 7452 -2304 7852 -2088
rect 7452 -2460 7492 -2304
rect 7492 -2460 7632 -2304
rect 7632 -2460 7684 -2304
rect 7684 -2460 7824 -2304
rect 7824 -2460 7852 -2304
rect 8488 -2088 8532 -1936
rect 8532 -2088 8672 -1936
rect 8672 -2088 8724 -1936
rect 8724 -2088 8864 -1936
rect 8864 -2088 8888 -1936
rect 8488 -2304 8888 -2088
rect 8488 -2460 8532 -2304
rect 8532 -2460 8672 -2304
rect 8672 -2460 8724 -2304
rect 8724 -2460 8864 -2304
rect 8864 -2460 8888 -2304
rect 11952 -2088 11992 -1936
rect 11992 -2088 12132 -1936
rect 12132 -2088 12184 -1936
rect 12184 -2088 12324 -1936
rect 12324 -2088 12352 -1936
rect 11952 -2304 12352 -2088
rect 11952 -2460 11992 -2304
rect 11992 -2460 12132 -2304
rect 12132 -2460 12184 -2304
rect 12184 -2460 12324 -2304
rect 12324 -2460 12352 -2304
rect 12992 -2088 13032 -1936
rect 13032 -2088 13172 -1936
rect 13172 -2088 13224 -1936
rect 13224 -2088 13364 -1936
rect 13364 -2088 13392 -1936
rect 12992 -2304 13392 -2088
rect 12992 -2460 13032 -2304
rect 13032 -2460 13172 -2304
rect 13172 -2460 13224 -2304
rect 13224 -2460 13364 -2304
rect 13364 -2460 13392 -2304
rect 14032 -2088 14072 -1936
rect 14072 -2088 14212 -1936
rect 14212 -2088 14264 -1936
rect 14264 -2088 14404 -1936
rect 14404 -2088 14432 -1936
rect 14032 -2304 14432 -2088
rect 14032 -2460 14072 -2304
rect 14072 -2460 14212 -2304
rect 14212 -2460 14264 -2304
rect 14264 -2460 14404 -2304
rect 14404 -2460 14432 -2304
rect 15072 -2088 15112 -1936
rect 15112 -2088 15252 -1936
rect 15252 -2088 15304 -1936
rect 15304 -2088 15444 -1936
rect 15444 -2088 15472 -1936
rect 15072 -2304 15472 -2088
rect 15072 -2460 15112 -2304
rect 15112 -2460 15252 -2304
rect 15252 -2460 15304 -2304
rect 15304 -2460 15444 -2304
rect 15444 -2460 15472 -2304
rect 16108 -2088 16152 -1936
rect 16152 -2088 16292 -1936
rect 16292 -2088 16344 -1936
rect 16344 -2088 16484 -1936
rect 16484 -2088 16508 -1936
rect 16108 -2304 16508 -2088
rect 16108 -2460 16152 -2304
rect 16152 -2460 16292 -2304
rect 16292 -2460 16344 -2304
rect 16344 -2460 16484 -2304
rect 16484 -2460 16508 -2304
rect 4844 -3512 4932 -3360
rect 4932 -3512 4984 -3360
rect 4984 -3512 5264 -3360
rect 5264 -3512 5284 -3360
rect 5904 -3512 5972 -3380
rect 5972 -3512 6024 -3380
rect 6024 -3512 6304 -3380
rect 6924 -3512 7012 -3380
rect 7012 -3512 7064 -3380
rect 7064 -3512 7344 -3380
rect 7984 -3512 8052 -3380
rect 8052 -3512 8104 -3380
rect 8104 -3512 8384 -3380
rect 8384 -3512 8404 -3380
rect 9004 -3512 9092 -3380
rect 9092 -3512 9144 -3380
rect 9144 -3512 9424 -3380
rect -7420 -3714 -7410 -3580
rect -7410 -3714 -7358 -3580
rect -7358 -3714 -7174 -3580
rect -7174 -3714 -7122 -3580
rect -7122 -3714 -6938 -3580
rect -6938 -3714 -6886 -3580
rect -6886 -3714 -6702 -3580
rect -6702 -3714 -6650 -3580
rect -6650 -3714 -6620 -3580
rect 4844 -3620 5284 -3512
rect 5904 -3700 6304 -3512
rect 6924 -3700 7344 -3512
rect 7984 -3700 8404 -3512
rect 9004 -3700 9424 -3512
rect 12464 -3512 12552 -3360
rect 12552 -3512 12604 -3360
rect 12604 -3512 12884 -3360
rect 12884 -3512 12904 -3360
rect 13524 -3512 13592 -3380
rect 13592 -3512 13644 -3380
rect 13644 -3512 13924 -3380
rect 14544 -3512 14632 -3380
rect 14632 -3512 14684 -3380
rect 14684 -3512 14964 -3380
rect 15604 -3512 15672 -3380
rect 15672 -3512 15724 -3380
rect 15724 -3512 16004 -3380
rect 16004 -3512 16024 -3380
rect 16624 -3512 16712 -3380
rect 16712 -3512 16764 -3380
rect 16764 -3512 17044 -3380
rect 12464 -3620 12904 -3512
rect 13524 -3700 13924 -3512
rect 14544 -3700 14964 -3512
rect 15604 -3700 16024 -3512
rect 16624 -3700 17044 -3512
rect -7420 -3862 -6620 -3714
rect 4924 -3840 5224 -3720
rect 8564 -3840 8864 -3720
rect 12544 -3840 12844 -3720
rect 16184 -3840 16484 -3720
rect -7420 -3960 -7230 -3862
rect -7230 -3960 -6950 -3862
rect -6950 -3960 -6620 -3862
<< metal3 >>
rect -10420 6740 18720 8900
rect -10420 6580 -1440 6740
rect -10420 6300 -9020 6580
rect -3140 6300 -1440 6580
rect -10420 6042 -1440 6300
rect -10420 5978 -10328 6042
rect -6304 5978 -6008 6042
rect -1984 5978 -1440 6042
rect -10420 5300 -1440 5978
rect -10356 1690 -6276 5300
rect -6036 1690 -1956 5300
rect -1672 4860 -1440 5300
rect -1080 6720 1360 6740
rect -1080 4860 0 6720
rect -1672 4840 0 4860
rect 360 4860 1360 6720
rect 1720 6720 18720 6740
rect 1720 4860 2800 6720
rect 360 4840 2800 4860
rect 3160 5660 18720 6720
rect 3160 4840 3420 5660
rect 4844 5540 5284 5660
rect 4844 5320 4864 5540
rect 5264 5320 5284 5540
rect 4324 5225 4764 5240
rect 4294 5220 4764 5225
rect 4294 4980 4304 5220
rect 4744 4980 4764 5220
rect 4294 4975 4764 4980
rect -1672 4180 3420 4840
rect 4324 4605 4764 4975
rect 4294 4600 4764 4605
rect 4294 4380 4304 4600
rect 4744 4380 4764 4600
rect 4294 4375 4764 4380
rect 4324 3985 4764 4375
rect 4294 3980 4764 3985
rect 4294 3760 4304 3980
rect 4744 3760 4764 3980
rect 4294 3755 4320 3760
rect 4310 3365 4320 3755
rect 4294 3360 4320 3365
rect 4740 3360 4764 3760
rect 4844 4920 5284 5320
rect 5864 5540 6304 5660
rect 5864 5320 5884 5540
rect 6284 5320 6304 5540
rect 4844 4700 4864 4920
rect 5264 4700 5284 4920
rect 4844 4300 5284 4700
rect 4844 4080 4864 4300
rect 5264 4080 5284 4300
rect 4844 3680 5284 4080
rect 4844 3460 4864 3680
rect 5264 3460 5284 3680
rect 4844 3440 5284 3460
rect 5364 5200 5804 5240
rect 5364 4980 5384 5200
rect 5784 4980 5804 5200
rect 5364 4600 5804 4980
rect 5364 4380 5384 4600
rect 5784 4380 5804 4600
rect 5364 3980 5804 4380
rect -1644 3280 3112 3320
rect -1644 2780 -1140 3280
rect 60 2780 1660 3280
rect 2860 2780 3112 3280
rect 4294 3140 4304 3360
rect 4744 3140 4764 3360
rect 5364 3336 5380 3980
rect 5784 3760 5804 3980
rect 5780 3360 5804 3760
rect 5864 4920 6304 5320
rect 6904 5540 7344 5660
rect 6904 5320 6924 5540
rect 7324 5320 7344 5540
rect 5864 4700 5884 4920
rect 6284 4700 6304 4920
rect 5864 4300 6304 4700
rect 5864 4080 5884 4300
rect 6284 4080 6304 4300
rect 5864 3680 6304 4080
rect 5864 3460 5884 3680
rect 6284 3460 6304 3680
rect 5864 3440 6304 3460
rect 6404 5200 6844 5240
rect 6404 4980 6424 5200
rect 6824 4980 6844 5200
rect 6404 4600 6844 4980
rect 6404 4380 6424 4600
rect 6824 4380 6844 4600
rect 6404 3980 6844 4380
rect 4294 3135 4764 3140
rect -1644 2552 3112 2780
rect 4316 2980 4764 3135
rect 5360 3140 5380 3336
rect 5784 3140 5804 3360
rect 6404 3336 6420 3980
rect 6824 3760 6844 3980
rect 6820 3360 6844 3760
rect 6904 4920 7344 5320
rect 7984 5540 8424 5660
rect 7984 5320 8004 5540
rect 8404 5320 8424 5540
rect 6904 4700 6924 4920
rect 7324 4700 7344 4920
rect 6904 4300 7344 4700
rect 6904 4080 6924 4300
rect 7324 4080 7344 4300
rect 6904 3680 7344 4080
rect 6904 3460 6924 3680
rect 7324 3460 7344 3680
rect 6904 3440 7344 3460
rect 7444 5200 7884 5240
rect 7444 4980 7464 5200
rect 7864 4980 7884 5200
rect 7444 4600 7884 4980
rect 7444 4380 7464 4600
rect 7864 4380 7884 4600
rect 7444 3980 7884 4380
rect -1488 2377 -1084 2552
rect -444 2385 -40 2552
rect -450 2380 -38 2385
rect 596 2381 1000 2552
rect -1494 2372 -1082 2377
rect -1494 1880 -1484 2372
rect -1092 1880 -1082 2372
rect -450 1888 -440 2380
rect -48 1888 -38 2380
rect -450 1883 -38 1888
rect 594 2376 1006 2381
rect 1644 2377 2048 2552
rect 2700 2377 3104 2552
rect 4316 2550 4760 2980
rect 5360 2555 5804 3140
rect 594 1884 604 2376
rect 996 1884 1006 2376
rect -1494 1875 -1082 1880
rect 594 1879 1006 1884
rect 1638 2372 2050 2377
rect 1638 1880 1648 2372
rect 2040 1880 2050 2372
rect 1638 1875 2050 1880
rect 2694 2372 3106 2377
rect 2694 1880 2704 2372
rect 3096 1880 3106 2372
rect 2694 1875 3106 1880
rect 4316 2016 4328 2550
rect 4748 2016 4760 2550
rect 1644 1872 2048 1875
rect -1580 1040 3340 1080
rect -1580 920 420 1040
rect 1380 920 3340 1040
rect -7040 202 -6680 520
rect -5510 454 -5330 458
rect -6018 406 -5330 454
rect -7042 22 -6674 202
rect -6018 154 -5998 406
rect -5802 158 -5330 406
rect -1580 440 -1540 920
rect -860 440 -500 920
rect 180 440 420 920
rect 1380 440 1580 920
rect 2260 440 2620 920
rect 3300 440 3340 920
rect -1580 400 3340 440
rect 4316 315 4760 2016
rect 5358 2550 5804 2555
rect 5358 2016 5368 2550
rect 5788 2016 5804 2550
rect 5358 2011 5804 2016
rect 4844 1120 5284 1140
rect 4844 780 4864 1120
rect 5264 780 5284 1120
rect 4316 310 4762 315
rect -5802 154 3474 158
rect -6018 146 3474 154
rect -7042 -210 -7030 22
rect -6698 -210 -6674 22
rect -7494 -294 -7130 -282
rect -7494 -526 -7478 -294
rect -7146 -526 -7130 -294
rect -7494 -918 -7130 -526
rect -7042 -598 -6674 -210
rect -7042 -830 -7030 -598
rect -6698 -830 -6674 -598
rect -7042 -846 -6674 -830
rect -5510 130 3474 146
rect -7494 -1150 -7478 -918
rect -7146 -1150 -7130 -918
rect -7494 -2149 -7130 -1150
rect -7494 -2154 -6900 -2149
rect -7494 -2646 -7298 -2154
rect -6910 -2646 -6900 -2154
rect -7494 -2650 -6900 -2646
rect -7308 -2651 -6900 -2650
rect -7430 -3580 -6610 -3575
rect -7430 -3960 -7420 -3580
rect -6620 -3960 -6610 -3580
rect -5510 -3894 -1222 130
rect -1158 -222 3390 130
rect -1158 -3894 -1138 -222
rect -5510 -3922 -1138 -3894
rect -898 -3894 3390 -222
rect 3454 100 3474 130
rect 3454 76 3932 100
rect 3454 -140 3712 76
rect 3912 -140 3932 76
rect 3454 -160 3932 -140
rect 3454 -3894 3474 -160
rect 4316 -224 4332 310
rect 4752 -224 4762 310
rect 4844 -120 5284 780
rect 4316 -229 4762 -224
rect 4316 -1936 4760 -229
rect 4316 -2460 4332 -1936
rect 4732 -2460 4760 -1936
rect 4316 -2480 4760 -2460
rect 4824 -1120 5284 -120
rect 4824 -1440 4844 -1120
rect 5264 -1440 5284 -1120
rect -898 -3922 3474 -3894
rect 4824 -3300 5284 -1440
rect 5360 315 5804 2011
rect 6396 3140 6420 3336
rect 6824 3140 6844 3360
rect 6396 2980 6844 3140
rect 7444 3140 7460 3980
rect 7864 3760 7884 3980
rect 7860 3360 7884 3760
rect 7984 4920 8424 5320
rect 9004 5540 9444 5660
rect 9004 5320 9024 5540
rect 9424 5320 9444 5540
rect 7984 4700 8004 4920
rect 8404 4700 8424 4920
rect 7984 4300 8424 4700
rect 7984 4080 8004 4300
rect 8404 4080 8424 4300
rect 7984 3680 8424 4080
rect 7984 3460 8004 3680
rect 8404 3460 8424 3680
rect 7984 3440 8424 3460
rect 8484 5220 8924 5240
rect 8484 5000 8504 5220
rect 8904 5000 8924 5220
rect 8484 4600 8924 5000
rect 8484 4380 8504 4600
rect 8904 4380 8924 4600
rect 8484 3980 8924 4380
rect 7864 3336 7884 3360
rect 8484 3336 8500 3980
rect 8904 3760 8924 3980
rect 8900 3360 8924 3760
rect 9004 4920 9444 5320
rect 10024 5540 10464 5660
rect 10024 5320 10044 5540
rect 10444 5320 10464 5540
rect 9004 4700 9024 4920
rect 9424 4700 9444 4920
rect 9004 4300 9444 4700
rect 9004 4080 9024 4300
rect 9424 4080 9444 4300
rect 9004 3680 9444 4080
rect 9004 3460 9024 3680
rect 9424 3460 9444 3680
rect 9004 3440 9444 3460
rect 9524 5220 9964 5240
rect 9524 5000 9544 5220
rect 9944 5000 9964 5220
rect 9524 4600 9964 5000
rect 9524 4380 9544 4600
rect 9944 4380 9964 4600
rect 9524 3980 9964 4380
rect 7864 3140 7888 3336
rect 6396 2550 6840 2980
rect 7444 2555 7888 3140
rect 6396 2016 6408 2550
rect 6828 2016 6840 2550
rect 5884 1125 6324 1140
rect 5884 1120 6334 1125
rect 5884 800 5904 1120
rect 6324 800 6334 1120
rect 5884 795 6334 800
rect 5360 310 5806 315
rect 5360 -224 5376 310
rect 5796 -224 5806 310
rect 5360 -229 5806 -224
rect 5360 -1936 5804 -229
rect 5884 -660 6324 795
rect 5864 -940 6324 -660
rect 5360 -2460 5372 -1936
rect 5772 -2460 5804 -1936
rect 5360 -2480 5804 -2460
rect 5884 -1115 6324 -940
rect 6396 315 6840 2016
rect 7438 2550 7888 2555
rect 7438 2016 7448 2550
rect 7868 2016 7888 2550
rect 7438 2011 7888 2016
rect 6904 1125 7344 1140
rect 6904 1120 7354 1125
rect 6904 800 6924 1120
rect 7344 800 7354 1120
rect 6904 795 7354 800
rect 6396 310 6842 315
rect 6396 -224 6412 310
rect 6832 -224 6842 310
rect 6396 -229 6842 -224
rect 6904 -120 7344 795
rect 7444 315 7888 2011
rect 8476 3140 8500 3336
rect 8904 3140 8924 3360
rect 9524 3336 9540 3980
rect 9944 3760 9964 3980
rect 9940 3360 9964 3760
rect 10024 4920 10464 5320
rect 12464 5540 12904 5660
rect 12464 5320 12484 5540
rect 12884 5320 12904 5540
rect 10024 4700 10044 4920
rect 10444 4700 10464 4920
rect 10024 4300 10464 4700
rect 10024 4080 10044 4300
rect 10444 4080 10464 4300
rect 10024 3680 10464 4080
rect 10024 3460 10044 3680
rect 10444 3460 10464 3680
rect 10024 3440 10464 3460
rect 10564 5220 11004 5240
rect 11944 5225 12384 5240
rect 10564 5000 10584 5220
rect 10984 5000 11004 5220
rect 10564 4600 11004 5000
rect 11914 5220 12384 5225
rect 11914 4980 11924 5220
rect 12364 4980 12384 5220
rect 11914 4975 12384 4980
rect 11944 4605 12384 4975
rect 10564 4380 10584 4600
rect 10984 4380 11004 4600
rect 10564 3980 11004 4380
rect 11914 4600 12384 4605
rect 11914 4380 11924 4600
rect 12364 4380 12384 4600
rect 11914 4375 12384 4380
rect 11944 3985 12384 4375
rect 8476 2980 8924 3140
rect 9520 3140 9540 3336
rect 9944 3140 9964 3360
rect 8476 2546 8920 2980
rect 9520 2555 9964 3140
rect 8476 2012 8488 2546
rect 8908 2012 8920 2546
rect 7442 310 7888 315
rect 5884 -1120 6334 -1115
rect 5884 -1440 5904 -1120
rect 6324 -1440 6334 -1120
rect 5884 -1445 6334 -1440
rect 5884 -3300 6324 -1445
rect 6396 -1936 6840 -229
rect 6396 -2460 6412 -1936
rect 6812 -2460 6840 -1936
rect 6396 -2480 6840 -2460
rect 6904 -1120 7364 -120
rect 7442 -224 7452 310
rect 7872 -224 7888 310
rect 7442 -229 7888 -224
rect 6904 -1440 6924 -1120
rect 7344 -1440 7364 -1120
rect 6904 -3300 7364 -1440
rect 7444 -1931 7888 -229
rect 7442 -1936 7888 -1931
rect 7442 -2460 7452 -1936
rect 7852 -2460 7888 -1936
rect 7442 -2465 7888 -2460
rect 7444 -2480 7888 -2465
rect 7964 1125 8404 1140
rect 7964 1120 8414 1125
rect 7964 800 7984 1120
rect 8404 800 8414 1120
rect 7964 795 8414 800
rect 7964 -1115 8404 795
rect 8476 310 8920 2012
rect 9518 2550 9964 2555
rect 10564 3140 10580 3980
rect 10984 3760 11004 3980
rect 10980 3360 11004 3760
rect 11914 3980 12384 3985
rect 11914 3760 11924 3980
rect 12364 3760 12384 3980
rect 11914 3755 12384 3760
rect 11944 3365 12384 3755
rect 12464 4920 12904 5320
rect 13484 5540 13924 5660
rect 13484 5320 13504 5540
rect 13904 5320 13924 5540
rect 12464 4700 12484 4920
rect 12884 4700 12904 4920
rect 12464 4300 12904 4700
rect 12464 4080 12484 4300
rect 12884 4080 12904 4300
rect 12464 3680 12904 4080
rect 12464 3460 12484 3680
rect 12884 3460 12904 3680
rect 12464 3440 12904 3460
rect 12984 5200 13424 5240
rect 12984 4980 13004 5200
rect 13404 4980 13424 5200
rect 12984 4600 13424 4980
rect 12984 4380 13004 4600
rect 13404 4380 13424 4600
rect 12984 3980 13424 4380
rect 12984 3760 13004 3980
rect 13404 3760 13424 3980
rect 10984 3336 11004 3360
rect 11914 3360 12384 3365
rect 10984 3140 11008 3336
rect 10564 2551 11008 3140
rect 11914 3140 11924 3360
rect 12364 3140 12384 3360
rect 12984 3360 13424 3760
rect 13484 4920 13924 5320
rect 14524 5540 14964 5660
rect 14524 5320 14544 5540
rect 14944 5320 14964 5540
rect 13484 4700 13504 4920
rect 13904 4700 13924 4920
rect 13484 4300 13924 4700
rect 13484 4080 13504 4300
rect 13904 4080 13924 4300
rect 13484 3680 13924 4080
rect 13484 3460 13504 3680
rect 13904 3460 13924 3680
rect 13484 3440 13924 3460
rect 14024 5200 14464 5240
rect 14024 4980 14044 5200
rect 14444 4980 14464 5200
rect 14024 4600 14464 4980
rect 14024 4380 14044 4600
rect 14444 4380 14464 4600
rect 14024 3980 14464 4380
rect 14024 3760 14044 3980
rect 14444 3760 14464 3980
rect 12984 3336 13004 3360
rect 11914 3135 12384 3140
rect 9518 2016 9528 2550
rect 9948 2016 9964 2550
rect 9518 2011 9964 2016
rect 8476 -224 8488 310
rect 8908 -224 8920 310
rect 9004 1125 9444 1140
rect 9004 1120 9454 1125
rect 9004 800 9024 1120
rect 9444 800 9454 1120
rect 9004 795 9454 800
rect 9004 -120 9444 795
rect 9520 315 9964 2011
rect 10558 2546 11008 2551
rect 10558 2012 10568 2546
rect 10988 2012 11008 2546
rect 10558 2007 11008 2012
rect 7964 -1120 8414 -1115
rect 7964 -1440 7984 -1120
rect 8404 -1440 8414 -1120
rect 7964 -1445 8414 -1440
rect 7964 -2720 8404 -1445
rect 8476 -1936 8920 -224
rect 8476 -2460 8488 -1936
rect 8888 -2460 8920 -1936
rect 8476 -2480 8920 -2460
rect 8984 -1120 9444 -120
rect 9510 310 9964 315
rect 9510 -224 9520 310
rect 9940 -224 9964 310
rect 9510 -229 9964 -224
rect 9520 -244 9964 -229
rect 10024 1120 10484 1140
rect 10024 800 10044 1120
rect 10464 800 10484 1120
rect 8984 -1440 9004 -1120
rect 9424 -1440 9444 -1120
rect 8984 -2720 9444 -1440
rect 7964 -3300 9444 -2720
rect 10024 -1120 10484 800
rect 10564 315 11008 2007
rect 10550 310 11008 315
rect 10550 -224 10560 310
rect 10980 -224 11008 310
rect 10550 -229 11008 -224
rect 10564 -244 11008 -229
rect 11936 2980 12384 3135
rect 12980 3140 13004 3336
rect 13404 3140 13424 3360
rect 14024 3360 14464 3760
rect 14524 4920 14964 5320
rect 15604 5540 16044 5660
rect 15604 5320 15624 5540
rect 16024 5320 16044 5540
rect 14524 4700 14544 4920
rect 14944 4700 14964 4920
rect 14524 4300 14964 4700
rect 14524 4080 14544 4300
rect 14944 4080 14964 4300
rect 14524 3680 14964 4080
rect 14524 3460 14544 3680
rect 14944 3460 14964 3680
rect 14524 3440 14964 3460
rect 15064 5200 15504 5240
rect 15064 4980 15084 5200
rect 15484 4980 15504 5200
rect 15064 4600 15504 4980
rect 15064 4380 15084 4600
rect 15484 4380 15504 4600
rect 15064 3980 15504 4380
rect 15064 3760 15084 3980
rect 15484 3760 15504 3980
rect 14024 3336 14044 3360
rect 11936 2550 12380 2980
rect 12980 2555 13424 3140
rect 11936 2016 11948 2550
rect 12368 2016 12380 2550
rect 11936 940 12380 2016
rect 12978 2550 13424 2555
rect 12978 2016 12988 2550
rect 13408 2016 13424 2550
rect 12978 2011 13424 2016
rect 11936 310 11960 940
rect 12360 315 12380 940
rect 12464 1120 12904 1140
rect 12464 780 12484 1120
rect 12884 780 12904 1120
rect 12360 310 12382 315
rect 11936 -224 11952 310
rect 12372 -224 12382 310
rect 12464 -120 12904 780
rect 11936 -229 12382 -224
rect 10024 -1440 10044 -1120
rect 10464 -1440 10484 -1120
rect 10024 -3300 10484 -1440
rect 11936 -1936 12380 -229
rect 11936 -2460 11952 -1936
rect 12352 -2460 12380 -1936
rect 11936 -2480 12380 -2460
rect 12444 -1120 12904 -120
rect 12444 -1440 12464 -1120
rect 12884 -1440 12904 -1120
rect 4824 -3360 10484 -3300
rect 4824 -3620 4844 -3360
rect 5284 -3380 10484 -3360
rect 5284 -3620 5904 -3380
rect 4824 -3880 4880 -3620
rect 5240 -3700 5904 -3620
rect 6304 -3700 6924 -3380
rect 7344 -3700 7984 -3380
rect 8404 -3700 9004 -3380
rect 9424 -3400 10484 -3380
rect 9424 -3700 10060 -3400
rect 5240 -3880 5940 -3700
rect 6300 -3880 6960 -3700
rect 7320 -3880 8020 -3700
rect 8380 -3720 9020 -3700
rect 8380 -3840 8564 -3720
rect 8864 -3840 9020 -3720
rect 8380 -3880 9020 -3840
rect 9380 -3880 10060 -3700
rect 10420 -3880 10484 -3400
rect 4824 -3920 10484 -3880
rect 12444 -3300 12904 -1440
rect 12980 940 13424 2011
rect 14016 3140 14044 3336
rect 14444 3140 14464 3360
rect 14016 2980 14464 3140
rect 15064 3360 15504 3760
rect 15604 4920 16044 5320
rect 16624 5540 17064 5660
rect 16624 5320 16644 5540
rect 17044 5320 17064 5540
rect 15604 4700 15624 4920
rect 16024 4700 16044 4920
rect 15604 4300 16044 4700
rect 15604 4080 15624 4300
rect 16024 4080 16044 4300
rect 15604 3680 16044 4080
rect 15604 3460 15624 3680
rect 16024 3460 16044 3680
rect 15604 3440 16044 3460
rect 16104 5220 16544 5240
rect 16104 5000 16124 5220
rect 16524 5000 16544 5220
rect 16104 4600 16544 5000
rect 16104 4380 16124 4600
rect 16524 4380 16544 4600
rect 16104 3980 16544 4380
rect 16104 3760 16124 3980
rect 16524 3760 16544 3980
rect 15064 3140 15084 3360
rect 15484 3336 15504 3360
rect 16104 3360 16544 3760
rect 16624 4920 17064 5320
rect 17644 5540 18084 5660
rect 17644 5320 17664 5540
rect 18064 5320 18084 5540
rect 16624 4700 16644 4920
rect 17044 4700 17064 4920
rect 16624 4300 17064 4700
rect 16624 4080 16644 4300
rect 17044 4080 17064 4300
rect 16624 3680 17064 4080
rect 16624 3460 16644 3680
rect 17044 3460 17064 3680
rect 16624 3440 17064 3460
rect 17144 5220 17584 5240
rect 17144 5000 17164 5220
rect 17564 5000 17584 5220
rect 17144 4600 17584 5000
rect 17144 4380 17164 4600
rect 17564 4380 17584 4600
rect 17144 3980 17584 4380
rect 17144 3760 17164 3980
rect 17564 3760 17584 3980
rect 16104 3336 16124 3360
rect 15484 3140 15508 3336
rect 14016 2550 14460 2980
rect 15064 2555 15508 3140
rect 14016 2016 14028 2550
rect 14448 2016 14460 2550
rect 12980 310 13000 940
rect 13400 315 13424 940
rect 13504 1125 13944 1140
rect 13504 1120 13954 1125
rect 13504 800 13524 1120
rect 13944 800 13954 1120
rect 13504 795 13954 800
rect 14016 940 14460 2016
rect 15058 2550 15508 2555
rect 15058 2016 15068 2550
rect 15488 2016 15508 2550
rect 15058 2011 15508 2016
rect 13400 310 13426 315
rect 12980 -224 12996 310
rect 13416 -224 13426 310
rect 12980 -229 13426 -224
rect 12980 -1936 13424 -229
rect 13504 -660 13944 795
rect 13484 -940 13944 -660
rect 12980 -2460 12992 -1936
rect 13392 -2460 13424 -1936
rect 12980 -2480 13424 -2460
rect 13504 -1115 13944 -940
rect 14016 310 14040 940
rect 14440 315 14460 940
rect 14524 1125 14964 1140
rect 14524 1120 14974 1125
rect 14524 800 14544 1120
rect 14964 800 14974 1120
rect 14524 795 14974 800
rect 15064 940 15508 2011
rect 16096 3140 16124 3336
rect 16524 3140 16544 3360
rect 17144 3360 17584 3760
rect 17644 4920 18084 5320
rect 17644 4700 17664 4920
rect 18064 4700 18084 4920
rect 17644 4300 18084 4700
rect 17644 4080 17664 4300
rect 18064 4080 18084 4300
rect 17644 3680 18084 4080
rect 17644 3460 17664 3680
rect 18064 3460 18084 3680
rect 17644 3440 18084 3460
rect 18184 5220 18624 5240
rect 18184 5000 18204 5220
rect 18604 5000 18624 5220
rect 18184 4600 18624 5000
rect 18184 4380 18204 4600
rect 18604 4380 18624 4600
rect 18184 3980 18624 4380
rect 18184 3760 18204 3980
rect 18604 3760 18624 3980
rect 17144 3336 17164 3360
rect 16096 2980 16544 3140
rect 17140 3140 17164 3336
rect 17564 3140 17584 3360
rect 16096 2546 16540 2980
rect 17140 2555 17584 3140
rect 16096 2012 16108 2546
rect 16528 2012 16540 2546
rect 14440 310 14462 315
rect 14016 -224 14032 310
rect 14452 -224 14462 310
rect 14016 -229 14462 -224
rect 14524 -120 14964 795
rect 15064 315 15080 940
rect 15062 310 15080 315
rect 15480 310 15508 940
rect 13504 -1120 13954 -1115
rect 13504 -1440 13524 -1120
rect 13944 -1440 13954 -1120
rect 13504 -1445 13954 -1440
rect 13504 -3300 13944 -1445
rect 14016 -1936 14460 -229
rect 14016 -2460 14032 -1936
rect 14432 -2460 14460 -1936
rect 14016 -2480 14460 -2460
rect 14524 -1120 14984 -120
rect 15062 -224 15072 310
rect 15492 -224 15508 310
rect 15062 -229 15508 -224
rect 14524 -1440 14544 -1120
rect 14964 -1440 14984 -1120
rect 14524 -3300 14984 -1440
rect 15064 -1931 15508 -229
rect 15062 -1936 15508 -1931
rect 15062 -2460 15072 -1936
rect 15472 -2460 15508 -1936
rect 15062 -2465 15508 -2460
rect 15064 -2480 15508 -2465
rect 15584 1125 16024 1140
rect 15584 1120 16034 1125
rect 15584 800 15604 1120
rect 16024 800 16034 1120
rect 15584 795 16034 800
rect 16096 940 16540 2012
rect 17138 2550 17584 2555
rect 18184 3360 18624 3760
rect 18184 3140 18204 3360
rect 18604 3336 18624 3360
rect 18604 3140 18628 3336
rect 18184 2551 18628 3140
rect 17138 2016 17148 2550
rect 17568 2016 17584 2550
rect 17138 2011 17584 2016
rect 15584 -1115 16024 795
rect 16096 310 16120 940
rect 16520 310 16540 940
rect 16096 -224 16108 310
rect 16528 -224 16540 310
rect 16624 1125 17064 1140
rect 16624 1120 17074 1125
rect 16624 800 16644 1120
rect 17064 800 17074 1120
rect 16624 795 17074 800
rect 17140 940 17584 2011
rect 18178 2546 18628 2551
rect 18178 2012 18188 2546
rect 18608 2012 18628 2546
rect 18178 2007 18628 2012
rect 16624 -120 17064 795
rect 17140 315 17160 940
rect 15584 -1120 16034 -1115
rect 15584 -1440 15604 -1120
rect 16024 -1440 16034 -1120
rect 15584 -1445 16034 -1440
rect 15584 -2720 16024 -1445
rect 16096 -1936 16540 -224
rect 16096 -2460 16108 -1936
rect 16508 -2460 16540 -1936
rect 16096 -2480 16540 -2460
rect 16604 -1120 17064 -120
rect 17130 310 17160 315
rect 17130 -224 17140 310
rect 17560 -224 17584 940
rect 17130 -229 17584 -224
rect 17140 -244 17584 -229
rect 17644 1120 18104 1140
rect 17644 800 17664 1120
rect 18084 800 18104 1120
rect 16604 -1440 16624 -1120
rect 17044 -1440 17064 -1120
rect 16604 -2720 17064 -1440
rect 15584 -3300 17064 -2720
rect 17644 -1120 18104 800
rect 18184 940 18628 2007
rect 18184 315 18200 940
rect 18170 310 18200 315
rect 18170 -224 18180 310
rect 18600 -224 18628 940
rect 18170 -229 18628 -224
rect 18184 -244 18628 -229
rect 17644 -1440 17664 -1120
rect 18084 -1440 18104 -1120
rect 17644 -3300 18104 -1440
rect 12444 -3360 18104 -3300
rect 12444 -3620 12464 -3360
rect 12904 -3380 18104 -3360
rect 12904 -3620 13524 -3380
rect 12444 -3880 12500 -3620
rect 12860 -3700 13524 -3620
rect 13924 -3700 14544 -3380
rect 14964 -3700 15604 -3380
rect 16024 -3700 16624 -3380
rect 17044 -3400 18104 -3380
rect 17044 -3700 17700 -3400
rect 12860 -3880 13560 -3700
rect 13920 -3880 14580 -3700
rect 14940 -3880 15640 -3700
rect 16000 -3720 16660 -3700
rect 16000 -3840 16184 -3720
rect 16484 -3840 16660 -3720
rect 16000 -3880 16660 -3840
rect 17020 -3880 17700 -3700
rect 18060 -3880 18104 -3400
rect 12444 -3920 18104 -3880
rect -7430 -3965 -6610 -3960
<< via3 >>
rect -10328 5978 -6304 6042
rect -6008 5978 -1984 6042
rect 4320 3760 4740 3980
rect 4320 3360 4740 3760
rect 4320 3140 4740 3360
rect 5380 3760 5384 3980
rect 5384 3760 5780 3980
rect 5380 3360 5780 3760
rect 5380 3140 5384 3360
rect 5384 3140 5780 3360
rect 6420 3760 6424 3980
rect 6424 3760 6820 3980
rect 6420 3360 6820 3760
rect 420 920 1380 1040
rect 420 440 540 920
rect 540 440 1220 920
rect 1220 440 1380 920
rect -7420 -3960 -6620 -3580
rect -1222 -3894 -1158 130
rect 3390 -3894 3454 130
rect 6420 3140 6424 3360
rect 6424 3140 6820 3360
rect 7460 3760 7464 3980
rect 7464 3760 7860 3980
rect 7460 3360 7860 3760
rect 7460 3140 7464 3360
rect 7464 3140 7860 3360
rect 8500 3760 8504 3980
rect 8504 3760 8900 3980
rect 8500 3360 8900 3760
rect 8500 3140 8504 3360
rect 8504 3140 8900 3360
rect 9540 3760 9544 3980
rect 9544 3760 9940 3980
rect 9540 3360 9940 3760
rect 9540 3140 9544 3360
rect 9544 3140 9940 3360
rect 10580 3760 10584 3980
rect 10584 3760 10980 3980
rect 10580 3360 10980 3760
rect 10580 3140 10584 3360
rect 10584 3140 10980 3360
rect 11960 310 12360 940
rect 11960 100 12360 310
rect 4880 -3620 5240 -3400
rect 4880 -3720 5240 -3620
rect 5940 -3700 6300 -3400
rect 6960 -3700 7320 -3400
rect 8020 -3700 8380 -3400
rect 9020 -3700 9380 -3400
rect 4880 -3840 4924 -3720
rect 4924 -3840 5224 -3720
rect 5224 -3840 5240 -3720
rect 4880 -3880 5240 -3840
rect 5940 -3880 6300 -3700
rect 6960 -3880 7320 -3700
rect 8020 -3880 8380 -3700
rect 9020 -3880 9380 -3700
rect 10060 -3880 10420 -3400
rect 13000 310 13400 940
rect 13000 100 13400 310
rect 14040 310 14440 940
rect 14040 100 14440 310
rect 15080 310 15480 940
rect 15080 100 15480 310
rect 16120 310 16520 940
rect 16120 100 16520 310
rect 17160 310 17560 940
rect 17160 100 17560 310
rect 18200 310 18600 940
rect 18200 100 18600 310
rect 12500 -3620 12860 -3400
rect 12500 -3720 12860 -3620
rect 13560 -3700 13920 -3400
rect 14580 -3700 14940 -3400
rect 15640 -3700 16000 -3400
rect 16660 -3700 17020 -3400
rect 12500 -3840 12544 -3720
rect 12544 -3840 12844 -3720
rect 12844 -3840 12860 -3720
rect 12500 -3880 12860 -3840
rect 13560 -3880 13920 -3700
rect 14580 -3880 14940 -3700
rect 15640 -3880 16000 -3700
rect 16660 -3880 17020 -3700
rect 17700 -3880 18060 -3400
<< mimcap >>
rect -10316 5690 -6316 5730
rect -10316 1770 -10276 5690
rect -6356 1770 -6316 5690
rect -10316 1730 -6316 1770
rect -5996 5690 -1996 5730
rect -5996 1770 -5956 5690
rect -2036 1770 -1996 5690
rect -5996 1730 -1996 1770
rect -5470 78 -1470 118
rect -5470 -3842 -5430 78
rect -1510 -3842 -1470 78
rect -5470 -3882 -1470 -3842
rect -858 78 3142 118
rect -858 -3842 -818 78
rect 3102 -3842 3142 78
rect -858 -3882 3142 -3842
<< mimcapcontact >>
rect -10276 1770 -6356 5690
rect -5956 1770 -2036 5690
rect -5430 -3842 -1510 78
rect -818 -3842 3102 78
<< metal4 >>
rect -10344 6042 -6288 6058
rect -10344 5978 -10328 6042
rect -6304 5978 -6288 6042
rect -10344 5962 -6288 5978
rect -6024 6042 -1968 6058
rect -6024 5978 -6008 6042
rect -1984 5978 -1968 6042
rect -6024 5962 -1968 5978
rect -10277 5690 -6355 5691
rect -10277 1770 -10276 5690
rect -6356 2798 -6355 5690
rect -5957 5690 -2035 5691
rect -5957 2798 -5956 5690
rect -6356 1814 -5956 2798
rect -6356 1770 -6355 1814
rect -10277 1769 -6355 1770
rect -5957 1770 -5956 1814
rect -2036 1770 -2035 5690
rect 4400 3981 19800 4400
rect 4319 3980 19800 3981
rect 4319 3140 4320 3980
rect 4740 3140 5380 3980
rect 5780 3140 6420 3980
rect 6820 3140 7460 3980
rect 7860 3140 8500 3980
rect 8900 3140 9540 3980
rect 9940 3140 10580 3980
rect 10980 3140 19800 3980
rect 4319 3139 19800 3140
rect 4400 2400 19800 3139
rect -5957 1769 -2035 1770
rect -10084 -4200 -8316 1769
rect 380 1040 1420 1080
rect 380 440 420 1040
rect 1380 440 1420 1040
rect -1238 130 -1142 146
rect -5431 78 -1509 79
rect -7421 -3580 -6619 -3579
rect -7421 -3960 -7420 -3580
rect -6620 -3960 -6619 -3580
rect -5431 -3842 -5430 78
rect -1510 -3842 -1509 78
rect -5431 -3843 -1509 -3842
rect -7421 -3961 -6619 -3960
rect -7420 -4200 -6620 -3961
rect -4000 -4200 -2800 -3843
rect -1238 -3894 -1222 130
rect -1158 -3894 -1142 130
rect 380 79 1420 440
rect 11540 940 19800 1600
rect 3374 130 3470 146
rect -819 78 3103 79
rect -819 -3842 -818 78
rect 3102 -3842 3103 78
rect -819 -3843 3103 -3842
rect -1238 -3910 -1142 -3894
rect 0 -4200 1200 -3843
rect 3374 -3894 3390 130
rect 3454 -3894 3470 130
rect 11540 100 11960 940
rect 12360 100 13000 940
rect 13400 100 14040 940
rect 14440 100 15080 940
rect 15480 100 16120 940
rect 16520 100 17160 940
rect 17560 100 18200 940
rect 18600 100 19800 940
rect 11540 -400 19800 100
rect 3374 -3910 3470 -3894
rect 4840 -3400 5280 -3360
rect 4840 -3880 4880 -3400
rect 5240 -3880 5280 -3400
rect 3512 -4196 4488 -4188
rect 3132 -4200 4632 -4196
rect 4840 -4200 5280 -3880
rect 5900 -3400 6340 -3360
rect 5900 -3880 5940 -3400
rect 6300 -3880 6340 -3400
rect 5900 -4200 6340 -3880
rect 6920 -3400 7360 -3360
rect 6920 -3880 6960 -3400
rect 7320 -3880 7360 -3400
rect 6920 -4200 7360 -3880
rect 7980 -3400 8420 -3360
rect 7980 -3880 8020 -3400
rect 8380 -3880 8420 -3400
rect 7980 -4200 8420 -3880
rect 8980 -3400 9420 -3360
rect 8980 -3880 9020 -3400
rect 9380 -3880 9420 -3400
rect 8980 -4200 9420 -3880
rect 10020 -3400 10460 -3360
rect 10020 -3880 10060 -3400
rect 10420 -3880 10460 -3400
rect 10020 -4200 10460 -3880
rect 12460 -3400 12900 -3360
rect 12460 -3880 12500 -3400
rect 12860 -3880 12900 -3400
rect 12460 -4200 12900 -3880
rect 13520 -3400 13960 -3360
rect 13520 -3880 13560 -3400
rect 13920 -3880 13960 -3400
rect 13520 -4200 13960 -3880
rect 14540 -3400 14980 -3360
rect 14540 -3880 14580 -3400
rect 14940 -3880 14980 -3400
rect 14540 -4200 14980 -3880
rect 15600 -3400 16040 -3360
rect 15600 -3880 15640 -3400
rect 16000 -3880 16040 -3400
rect 15600 -4200 16040 -3880
rect 16620 -3400 17060 -3360
rect 16620 -3880 16660 -3400
rect 17020 -3880 17060 -3400
rect 16620 -4200 17060 -3880
rect 17660 -3400 18100 -3360
rect 17660 -3880 17700 -3400
rect 18060 -3880 18100 -3400
rect 17660 -4200 18100 -3880
rect -10200 -5288 19800 -4200
rect -10200 -6528 -8052 -5288
rect -7024 -6528 19800 -5288
rect -10200 -7796 19800 -6528
rect -10200 -7800 3680 -7796
rect 4300 -7800 19800 -7796
<< res1p41 >>
rect -1436 5768 -1150 6172
rect -1058 5768 -772 6172
rect -680 5768 -394 6172
rect -302 5768 -16 6172
rect 76 5768 362 6172
rect 1364 5768 1650 6172
rect 1742 5768 2028 6172
rect 2120 5768 2406 6172
rect 2498 5768 2784 6172
rect 2876 5768 3162 6172
rect -1436 4400 -1150 4804
rect -1058 4400 -772 4804
rect -680 4400 -394 4804
rect -302 4400 -16 4804
rect 76 4400 362 4804
rect 1364 4400 1650 4804
rect 1742 4400 2028 4804
rect 2120 4400 2406 4804
rect 2498 4400 2784 4804
rect 2876 4400 3162 4804
<< labels >>
rlabel metal1 1400 3500 1600 3700 1 InputSignal
port 1 n
rlabel metal1 140 3480 300 3700 1 InputRef
port 2 n
rlabel metal3 -7020 280 -6700 500 1 I_Bias
port 3 n
rlabel metal4 -9960 -6980 -9240 -4660 1 VN
port 4 n
rlabel metal3 -10200 6280 -9760 6680 1 VP
port 5 n
rlabel metal4 19140 2800 19560 3740 1 OutP
port 6 n
rlabel metal4 19200 220 19620 1160 1 OutN
port 7 n
<< end >>
