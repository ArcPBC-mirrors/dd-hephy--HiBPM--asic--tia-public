magic
tech sky130A
magscale 1 2
timestamp 1683714046
<< error_p >>
rect -845 2744 -787 2750
rect -653 2744 -595 2750
rect -461 2744 -403 2750
rect -269 2744 -211 2750
rect -77 2744 -19 2750
rect 115 2744 173 2750
rect 307 2744 365 2750
rect 499 2744 557 2750
rect 691 2744 749 2750
rect 883 2744 941 2750
rect -845 2710 -833 2744
rect -653 2710 -641 2744
rect -461 2710 -449 2744
rect -269 2710 -257 2744
rect -77 2710 -65 2744
rect 115 2710 127 2744
rect 307 2710 319 2744
rect 499 2710 511 2744
rect 691 2710 703 2744
rect 883 2710 895 2744
rect -845 2704 -787 2710
rect -653 2704 -595 2710
rect -461 2704 -403 2710
rect -269 2704 -211 2710
rect -77 2704 -19 2710
rect 115 2704 173 2710
rect 307 2704 365 2710
rect 499 2704 557 2710
rect 691 2704 749 2710
rect 883 2704 941 2710
rect -941 2234 -883 2240
rect -749 2234 -691 2240
rect -557 2234 -499 2240
rect -365 2234 -307 2240
rect -173 2234 -115 2240
rect 19 2234 77 2240
rect 211 2234 269 2240
rect 403 2234 461 2240
rect 595 2234 653 2240
rect 787 2234 845 2240
rect -941 2200 -929 2234
rect -749 2200 -737 2234
rect -557 2200 -545 2234
rect -365 2200 -353 2234
rect -173 2200 -161 2234
rect 19 2200 31 2234
rect 211 2200 223 2234
rect 403 2200 415 2234
rect 595 2200 607 2234
rect 787 2200 799 2234
rect -941 2194 -883 2200
rect -749 2194 -691 2200
rect -557 2194 -499 2200
rect -365 2194 -307 2200
rect -173 2194 -115 2200
rect 19 2194 77 2200
rect 211 2194 269 2200
rect 403 2194 461 2200
rect 595 2194 653 2200
rect 787 2194 845 2200
rect -941 2126 -883 2132
rect -749 2126 -691 2132
rect -557 2126 -499 2132
rect -365 2126 -307 2132
rect -173 2126 -115 2132
rect 19 2126 77 2132
rect 211 2126 269 2132
rect 403 2126 461 2132
rect 595 2126 653 2132
rect 787 2126 845 2132
rect -941 2092 -929 2126
rect -749 2092 -737 2126
rect -557 2092 -545 2126
rect -365 2092 -353 2126
rect -173 2092 -161 2126
rect 19 2092 31 2126
rect 211 2092 223 2126
rect 403 2092 415 2126
rect 595 2092 607 2126
rect 787 2092 799 2126
rect -941 2086 -883 2092
rect -749 2086 -691 2092
rect -557 2086 -499 2092
rect -365 2086 -307 2092
rect -173 2086 -115 2092
rect 19 2086 77 2092
rect 211 2086 269 2092
rect 403 2086 461 2092
rect 595 2086 653 2092
rect 787 2086 845 2092
rect -845 1616 -787 1622
rect -653 1616 -595 1622
rect -461 1616 -403 1622
rect -269 1616 -211 1622
rect -77 1616 -19 1622
rect 115 1616 173 1622
rect 307 1616 365 1622
rect 499 1616 557 1622
rect 691 1616 749 1622
rect 883 1616 941 1622
rect -845 1582 -833 1616
rect -653 1582 -641 1616
rect -461 1582 -449 1616
rect -269 1582 -257 1616
rect -77 1582 -65 1616
rect 115 1582 127 1616
rect 307 1582 319 1616
rect 499 1582 511 1616
rect 691 1582 703 1616
rect 883 1582 895 1616
rect -845 1576 -787 1582
rect -653 1576 -595 1582
rect -461 1576 -403 1582
rect -269 1576 -211 1582
rect -77 1576 -19 1582
rect 115 1576 173 1582
rect 307 1576 365 1582
rect 499 1576 557 1582
rect 691 1576 749 1582
rect 883 1576 941 1582
rect -845 1508 -787 1514
rect -653 1508 -595 1514
rect -461 1508 -403 1514
rect -269 1508 -211 1514
rect -77 1508 -19 1514
rect 115 1508 173 1514
rect 307 1508 365 1514
rect 499 1508 557 1514
rect 691 1508 749 1514
rect 883 1508 941 1514
rect -845 1474 -833 1508
rect -653 1474 -641 1508
rect -461 1474 -449 1508
rect -269 1474 -257 1508
rect -77 1474 -65 1508
rect 115 1474 127 1508
rect 307 1474 319 1508
rect 499 1474 511 1508
rect 691 1474 703 1508
rect 883 1474 895 1508
rect -845 1468 -787 1474
rect -653 1468 -595 1474
rect -461 1468 -403 1474
rect -269 1468 -211 1474
rect -77 1468 -19 1474
rect 115 1468 173 1474
rect 307 1468 365 1474
rect 499 1468 557 1474
rect 691 1468 749 1474
rect 883 1468 941 1474
rect -941 998 -883 1004
rect -749 998 -691 1004
rect -557 998 -499 1004
rect -365 998 -307 1004
rect -173 998 -115 1004
rect 19 998 77 1004
rect 211 998 269 1004
rect 403 998 461 1004
rect 595 998 653 1004
rect 787 998 845 1004
rect -941 964 -929 998
rect -749 964 -737 998
rect -557 964 -545 998
rect -365 964 -353 998
rect -173 964 -161 998
rect 19 964 31 998
rect 211 964 223 998
rect 403 964 415 998
rect 595 964 607 998
rect 787 964 799 998
rect -941 958 -883 964
rect -749 958 -691 964
rect -557 958 -499 964
rect -365 958 -307 964
rect -173 958 -115 964
rect 19 958 77 964
rect 211 958 269 964
rect 403 958 461 964
rect 595 958 653 964
rect 787 958 845 964
rect -941 890 -883 896
rect -749 890 -691 896
rect -557 890 -499 896
rect -365 890 -307 896
rect -173 890 -115 896
rect 19 890 77 896
rect 211 890 269 896
rect 403 890 461 896
rect 595 890 653 896
rect 787 890 845 896
rect -941 856 -929 890
rect -749 856 -737 890
rect -557 856 -545 890
rect -365 856 -353 890
rect -173 856 -161 890
rect 19 856 31 890
rect 211 856 223 890
rect 403 856 415 890
rect 595 856 607 890
rect 787 856 799 890
rect -941 850 -883 856
rect -749 850 -691 856
rect -557 850 -499 856
rect -365 850 -307 856
rect -173 850 -115 856
rect 19 850 77 856
rect 211 850 269 856
rect 403 850 461 856
rect 595 850 653 856
rect 787 850 845 856
rect -845 380 -787 386
rect -653 380 -595 386
rect -461 380 -403 386
rect -269 380 -211 386
rect -77 380 -19 386
rect 115 380 173 386
rect 307 380 365 386
rect 499 380 557 386
rect 691 380 749 386
rect 883 380 941 386
rect -845 346 -833 380
rect -653 346 -641 380
rect -461 346 -449 380
rect -269 346 -257 380
rect -77 346 -65 380
rect 115 346 127 380
rect 307 346 319 380
rect 499 346 511 380
rect 691 346 703 380
rect 883 346 895 380
rect -845 340 -787 346
rect -653 340 -595 346
rect -461 340 -403 346
rect -269 340 -211 346
rect -77 340 -19 346
rect 115 340 173 346
rect 307 340 365 346
rect 499 340 557 346
rect 691 340 749 346
rect 883 340 941 346
rect -845 272 -787 278
rect -653 272 -595 278
rect -461 272 -403 278
rect -269 272 -211 278
rect -77 272 -19 278
rect 115 272 173 278
rect 307 272 365 278
rect 499 272 557 278
rect 691 272 749 278
rect 883 272 941 278
rect -845 238 -833 272
rect -653 238 -641 272
rect -461 238 -449 272
rect -269 238 -257 272
rect -77 238 -65 272
rect 115 238 127 272
rect 307 238 319 272
rect 499 238 511 272
rect 691 238 703 272
rect 883 238 895 272
rect -845 232 -787 238
rect -653 232 -595 238
rect -461 232 -403 238
rect -269 232 -211 238
rect -77 232 -19 238
rect 115 232 173 238
rect 307 232 365 238
rect 499 232 557 238
rect 691 232 749 238
rect 883 232 941 238
rect -941 -238 -883 -232
rect -749 -238 -691 -232
rect -557 -238 -499 -232
rect -365 -238 -307 -232
rect -173 -238 -115 -232
rect 19 -238 77 -232
rect 211 -238 269 -232
rect 403 -238 461 -232
rect 595 -238 653 -232
rect 787 -238 845 -232
rect -941 -272 -929 -238
rect -749 -272 -737 -238
rect -557 -272 -545 -238
rect -365 -272 -353 -238
rect -173 -272 -161 -238
rect 19 -272 31 -238
rect 211 -272 223 -238
rect 403 -272 415 -238
rect 595 -272 607 -238
rect 787 -272 799 -238
rect -941 -278 -883 -272
rect -749 -278 -691 -272
rect -557 -278 -499 -272
rect -365 -278 -307 -272
rect -173 -278 -115 -272
rect 19 -278 77 -272
rect 211 -278 269 -272
rect 403 -278 461 -272
rect 595 -278 653 -272
rect 787 -278 845 -272
rect -941 -346 -883 -340
rect -749 -346 -691 -340
rect -557 -346 -499 -340
rect -365 -346 -307 -340
rect -173 -346 -115 -340
rect 19 -346 77 -340
rect 211 -346 269 -340
rect 403 -346 461 -340
rect 595 -346 653 -340
rect 787 -346 845 -340
rect -941 -380 -929 -346
rect -749 -380 -737 -346
rect -557 -380 -545 -346
rect -365 -380 -353 -346
rect -173 -380 -161 -346
rect 19 -380 31 -346
rect 211 -380 223 -346
rect 403 -380 415 -346
rect 595 -380 607 -346
rect 787 -380 799 -346
rect -941 -386 -883 -380
rect -749 -386 -691 -380
rect -557 -386 -499 -380
rect -365 -386 -307 -380
rect -173 -386 -115 -380
rect 19 -386 77 -380
rect 211 -386 269 -380
rect 403 -386 461 -380
rect 595 -386 653 -380
rect 787 -386 845 -380
rect -845 -856 -787 -850
rect -653 -856 -595 -850
rect -461 -856 -403 -850
rect -269 -856 -211 -850
rect -77 -856 -19 -850
rect 115 -856 173 -850
rect 307 -856 365 -850
rect 499 -856 557 -850
rect 691 -856 749 -850
rect 883 -856 941 -850
rect -845 -890 -833 -856
rect -653 -890 -641 -856
rect -461 -890 -449 -856
rect -269 -890 -257 -856
rect -77 -890 -65 -856
rect 115 -890 127 -856
rect 307 -890 319 -856
rect 499 -890 511 -856
rect 691 -890 703 -856
rect 883 -890 895 -856
rect -845 -896 -787 -890
rect -653 -896 -595 -890
rect -461 -896 -403 -890
rect -269 -896 -211 -890
rect -77 -896 -19 -890
rect 115 -896 173 -890
rect 307 -896 365 -890
rect 499 -896 557 -890
rect 691 -896 749 -890
rect 883 -896 941 -890
rect -845 -964 -787 -958
rect -653 -964 -595 -958
rect -461 -964 -403 -958
rect -269 -964 -211 -958
rect -77 -964 -19 -958
rect 115 -964 173 -958
rect 307 -964 365 -958
rect 499 -964 557 -958
rect 691 -964 749 -958
rect 883 -964 941 -958
rect -845 -998 -833 -964
rect -653 -998 -641 -964
rect -461 -998 -449 -964
rect -269 -998 -257 -964
rect -77 -998 -65 -964
rect 115 -998 127 -964
rect 307 -998 319 -964
rect 499 -998 511 -964
rect 691 -998 703 -964
rect 883 -998 895 -964
rect -845 -1004 -787 -998
rect -653 -1004 -595 -998
rect -461 -1004 -403 -998
rect -269 -1004 -211 -998
rect -77 -1004 -19 -998
rect 115 -1004 173 -998
rect 307 -1004 365 -998
rect 499 -1004 557 -998
rect 691 -1004 749 -998
rect 883 -1004 941 -998
rect -941 -1474 -883 -1468
rect -749 -1474 -691 -1468
rect -557 -1474 -499 -1468
rect -365 -1474 -307 -1468
rect -173 -1474 -115 -1468
rect 19 -1474 77 -1468
rect 211 -1474 269 -1468
rect 403 -1474 461 -1468
rect 595 -1474 653 -1468
rect 787 -1474 845 -1468
rect -941 -1508 -929 -1474
rect -749 -1508 -737 -1474
rect -557 -1508 -545 -1474
rect -365 -1508 -353 -1474
rect -173 -1508 -161 -1474
rect 19 -1508 31 -1474
rect 211 -1508 223 -1474
rect 403 -1508 415 -1474
rect 595 -1508 607 -1474
rect 787 -1508 799 -1474
rect -941 -1514 -883 -1508
rect -749 -1514 -691 -1508
rect -557 -1514 -499 -1508
rect -365 -1514 -307 -1508
rect -173 -1514 -115 -1508
rect 19 -1514 77 -1508
rect 211 -1514 269 -1508
rect 403 -1514 461 -1508
rect 595 -1514 653 -1508
rect 787 -1514 845 -1508
rect -941 -1582 -883 -1576
rect -749 -1582 -691 -1576
rect -557 -1582 -499 -1576
rect -365 -1582 -307 -1576
rect -173 -1582 -115 -1576
rect 19 -1582 77 -1576
rect 211 -1582 269 -1576
rect 403 -1582 461 -1576
rect 595 -1582 653 -1576
rect 787 -1582 845 -1576
rect -941 -1616 -929 -1582
rect -749 -1616 -737 -1582
rect -557 -1616 -545 -1582
rect -365 -1616 -353 -1582
rect -173 -1616 -161 -1582
rect 19 -1616 31 -1582
rect 211 -1616 223 -1582
rect 403 -1616 415 -1582
rect 595 -1616 607 -1582
rect 787 -1616 799 -1582
rect -941 -1622 -883 -1616
rect -749 -1622 -691 -1616
rect -557 -1622 -499 -1616
rect -365 -1622 -307 -1616
rect -173 -1622 -115 -1616
rect 19 -1622 77 -1616
rect 211 -1622 269 -1616
rect 403 -1622 461 -1616
rect 595 -1622 653 -1616
rect 787 -1622 845 -1616
rect -845 -2092 -787 -2086
rect -653 -2092 -595 -2086
rect -461 -2092 -403 -2086
rect -269 -2092 -211 -2086
rect -77 -2092 -19 -2086
rect 115 -2092 173 -2086
rect 307 -2092 365 -2086
rect 499 -2092 557 -2086
rect 691 -2092 749 -2086
rect 883 -2092 941 -2086
rect -845 -2126 -833 -2092
rect -653 -2126 -641 -2092
rect -461 -2126 -449 -2092
rect -269 -2126 -257 -2092
rect -77 -2126 -65 -2092
rect 115 -2126 127 -2092
rect 307 -2126 319 -2092
rect 499 -2126 511 -2092
rect 691 -2126 703 -2092
rect 883 -2126 895 -2092
rect -845 -2132 -787 -2126
rect -653 -2132 -595 -2126
rect -461 -2132 -403 -2126
rect -269 -2132 -211 -2126
rect -77 -2132 -19 -2126
rect 115 -2132 173 -2126
rect 307 -2132 365 -2126
rect 499 -2132 557 -2126
rect 691 -2132 749 -2126
rect 883 -2132 941 -2126
rect -845 -2200 -787 -2194
rect -653 -2200 -595 -2194
rect -461 -2200 -403 -2194
rect -269 -2200 -211 -2194
rect -77 -2200 -19 -2194
rect 115 -2200 173 -2194
rect 307 -2200 365 -2194
rect 499 -2200 557 -2194
rect 691 -2200 749 -2194
rect 883 -2200 941 -2194
rect -845 -2234 -833 -2200
rect -653 -2234 -641 -2200
rect -461 -2234 -449 -2200
rect -269 -2234 -257 -2200
rect -77 -2234 -65 -2200
rect 115 -2234 127 -2200
rect 307 -2234 319 -2200
rect 499 -2234 511 -2200
rect 691 -2234 703 -2200
rect 883 -2234 895 -2200
rect -845 -2240 -787 -2234
rect -653 -2240 -595 -2234
rect -461 -2240 -403 -2234
rect -269 -2240 -211 -2234
rect -77 -2240 -19 -2234
rect 115 -2240 173 -2234
rect 307 -2240 365 -2234
rect 499 -2240 557 -2234
rect 691 -2240 749 -2234
rect 883 -2240 941 -2234
rect -941 -2710 -883 -2704
rect -749 -2710 -691 -2704
rect -557 -2710 -499 -2704
rect -365 -2710 -307 -2704
rect -173 -2710 -115 -2704
rect 19 -2710 77 -2704
rect 211 -2710 269 -2704
rect 403 -2710 461 -2704
rect 595 -2710 653 -2704
rect 787 -2710 845 -2704
rect -941 -2744 -929 -2710
rect -749 -2744 -737 -2710
rect -557 -2744 -545 -2710
rect -365 -2744 -353 -2710
rect -173 -2744 -161 -2710
rect 19 -2744 31 -2710
rect 211 -2744 223 -2710
rect 403 -2744 415 -2710
rect 595 -2744 607 -2710
rect 787 -2744 799 -2710
rect -941 -2750 -883 -2744
rect -749 -2750 -691 -2744
rect -557 -2750 -499 -2744
rect -365 -2750 -307 -2744
rect -173 -2750 -115 -2744
rect 19 -2750 77 -2744
rect 211 -2750 269 -2744
rect 403 -2750 461 -2744
rect 595 -2750 653 -2744
rect 787 -2750 845 -2744
<< pwell >>
rect -1127 -2882 1127 2882
<< nmoslvt >>
rect -927 2272 -897 2672
rect -831 2272 -801 2672
rect -735 2272 -705 2672
rect -639 2272 -609 2672
rect -543 2272 -513 2672
rect -447 2272 -417 2672
rect -351 2272 -321 2672
rect -255 2272 -225 2672
rect -159 2272 -129 2672
rect -63 2272 -33 2672
rect 33 2272 63 2672
rect 129 2272 159 2672
rect 225 2272 255 2672
rect 321 2272 351 2672
rect 417 2272 447 2672
rect 513 2272 543 2672
rect 609 2272 639 2672
rect 705 2272 735 2672
rect 801 2272 831 2672
rect 897 2272 927 2672
rect -927 1654 -897 2054
rect -831 1654 -801 2054
rect -735 1654 -705 2054
rect -639 1654 -609 2054
rect -543 1654 -513 2054
rect -447 1654 -417 2054
rect -351 1654 -321 2054
rect -255 1654 -225 2054
rect -159 1654 -129 2054
rect -63 1654 -33 2054
rect 33 1654 63 2054
rect 129 1654 159 2054
rect 225 1654 255 2054
rect 321 1654 351 2054
rect 417 1654 447 2054
rect 513 1654 543 2054
rect 609 1654 639 2054
rect 705 1654 735 2054
rect 801 1654 831 2054
rect 897 1654 927 2054
rect -927 1036 -897 1436
rect -831 1036 -801 1436
rect -735 1036 -705 1436
rect -639 1036 -609 1436
rect -543 1036 -513 1436
rect -447 1036 -417 1436
rect -351 1036 -321 1436
rect -255 1036 -225 1436
rect -159 1036 -129 1436
rect -63 1036 -33 1436
rect 33 1036 63 1436
rect 129 1036 159 1436
rect 225 1036 255 1436
rect 321 1036 351 1436
rect 417 1036 447 1436
rect 513 1036 543 1436
rect 609 1036 639 1436
rect 705 1036 735 1436
rect 801 1036 831 1436
rect 897 1036 927 1436
rect -927 418 -897 818
rect -831 418 -801 818
rect -735 418 -705 818
rect -639 418 -609 818
rect -543 418 -513 818
rect -447 418 -417 818
rect -351 418 -321 818
rect -255 418 -225 818
rect -159 418 -129 818
rect -63 418 -33 818
rect 33 418 63 818
rect 129 418 159 818
rect 225 418 255 818
rect 321 418 351 818
rect 417 418 447 818
rect 513 418 543 818
rect 609 418 639 818
rect 705 418 735 818
rect 801 418 831 818
rect 897 418 927 818
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
rect -927 -818 -897 -418
rect -831 -818 -801 -418
rect -735 -818 -705 -418
rect -639 -818 -609 -418
rect -543 -818 -513 -418
rect -447 -818 -417 -418
rect -351 -818 -321 -418
rect -255 -818 -225 -418
rect -159 -818 -129 -418
rect -63 -818 -33 -418
rect 33 -818 63 -418
rect 129 -818 159 -418
rect 225 -818 255 -418
rect 321 -818 351 -418
rect 417 -818 447 -418
rect 513 -818 543 -418
rect 609 -818 639 -418
rect 705 -818 735 -418
rect 801 -818 831 -418
rect 897 -818 927 -418
rect -927 -1436 -897 -1036
rect -831 -1436 -801 -1036
rect -735 -1436 -705 -1036
rect -639 -1436 -609 -1036
rect -543 -1436 -513 -1036
rect -447 -1436 -417 -1036
rect -351 -1436 -321 -1036
rect -255 -1436 -225 -1036
rect -159 -1436 -129 -1036
rect -63 -1436 -33 -1036
rect 33 -1436 63 -1036
rect 129 -1436 159 -1036
rect 225 -1436 255 -1036
rect 321 -1436 351 -1036
rect 417 -1436 447 -1036
rect 513 -1436 543 -1036
rect 609 -1436 639 -1036
rect 705 -1436 735 -1036
rect 801 -1436 831 -1036
rect 897 -1436 927 -1036
rect -927 -2054 -897 -1654
rect -831 -2054 -801 -1654
rect -735 -2054 -705 -1654
rect -639 -2054 -609 -1654
rect -543 -2054 -513 -1654
rect -447 -2054 -417 -1654
rect -351 -2054 -321 -1654
rect -255 -2054 -225 -1654
rect -159 -2054 -129 -1654
rect -63 -2054 -33 -1654
rect 33 -2054 63 -1654
rect 129 -2054 159 -1654
rect 225 -2054 255 -1654
rect 321 -2054 351 -1654
rect 417 -2054 447 -1654
rect 513 -2054 543 -1654
rect 609 -2054 639 -1654
rect 705 -2054 735 -1654
rect 801 -2054 831 -1654
rect 897 -2054 927 -1654
rect -927 -2672 -897 -2272
rect -831 -2672 -801 -2272
rect -735 -2672 -705 -2272
rect -639 -2672 -609 -2272
rect -543 -2672 -513 -2272
rect -447 -2672 -417 -2272
rect -351 -2672 -321 -2272
rect -255 -2672 -225 -2272
rect -159 -2672 -129 -2272
rect -63 -2672 -33 -2272
rect 33 -2672 63 -2272
rect 129 -2672 159 -2272
rect 225 -2672 255 -2272
rect 321 -2672 351 -2272
rect 417 -2672 447 -2272
rect 513 -2672 543 -2272
rect 609 -2672 639 -2272
rect 705 -2672 735 -2272
rect 801 -2672 831 -2272
rect 897 -2672 927 -2272
<< ndiff >>
rect -989 2660 -927 2672
rect -989 2284 -977 2660
rect -943 2284 -927 2660
rect -989 2272 -927 2284
rect -897 2660 -831 2672
rect -897 2284 -881 2660
rect -847 2284 -831 2660
rect -897 2272 -831 2284
rect -801 2660 -735 2672
rect -801 2284 -785 2660
rect -751 2284 -735 2660
rect -801 2272 -735 2284
rect -705 2660 -639 2672
rect -705 2284 -689 2660
rect -655 2284 -639 2660
rect -705 2272 -639 2284
rect -609 2660 -543 2672
rect -609 2284 -593 2660
rect -559 2284 -543 2660
rect -609 2272 -543 2284
rect -513 2660 -447 2672
rect -513 2284 -497 2660
rect -463 2284 -447 2660
rect -513 2272 -447 2284
rect -417 2660 -351 2672
rect -417 2284 -401 2660
rect -367 2284 -351 2660
rect -417 2272 -351 2284
rect -321 2660 -255 2672
rect -321 2284 -305 2660
rect -271 2284 -255 2660
rect -321 2272 -255 2284
rect -225 2660 -159 2672
rect -225 2284 -209 2660
rect -175 2284 -159 2660
rect -225 2272 -159 2284
rect -129 2660 -63 2672
rect -129 2284 -113 2660
rect -79 2284 -63 2660
rect -129 2272 -63 2284
rect -33 2660 33 2672
rect -33 2284 -17 2660
rect 17 2284 33 2660
rect -33 2272 33 2284
rect 63 2660 129 2672
rect 63 2284 79 2660
rect 113 2284 129 2660
rect 63 2272 129 2284
rect 159 2660 225 2672
rect 159 2284 175 2660
rect 209 2284 225 2660
rect 159 2272 225 2284
rect 255 2660 321 2672
rect 255 2284 271 2660
rect 305 2284 321 2660
rect 255 2272 321 2284
rect 351 2660 417 2672
rect 351 2284 367 2660
rect 401 2284 417 2660
rect 351 2272 417 2284
rect 447 2660 513 2672
rect 447 2284 463 2660
rect 497 2284 513 2660
rect 447 2272 513 2284
rect 543 2660 609 2672
rect 543 2284 559 2660
rect 593 2284 609 2660
rect 543 2272 609 2284
rect 639 2660 705 2672
rect 639 2284 655 2660
rect 689 2284 705 2660
rect 639 2272 705 2284
rect 735 2660 801 2672
rect 735 2284 751 2660
rect 785 2284 801 2660
rect 735 2272 801 2284
rect 831 2660 897 2672
rect 831 2284 847 2660
rect 881 2284 897 2660
rect 831 2272 897 2284
rect 927 2660 989 2672
rect 927 2284 943 2660
rect 977 2284 989 2660
rect 927 2272 989 2284
rect -989 2042 -927 2054
rect -989 1666 -977 2042
rect -943 1666 -927 2042
rect -989 1654 -927 1666
rect -897 2042 -831 2054
rect -897 1666 -881 2042
rect -847 1666 -831 2042
rect -897 1654 -831 1666
rect -801 2042 -735 2054
rect -801 1666 -785 2042
rect -751 1666 -735 2042
rect -801 1654 -735 1666
rect -705 2042 -639 2054
rect -705 1666 -689 2042
rect -655 1666 -639 2042
rect -705 1654 -639 1666
rect -609 2042 -543 2054
rect -609 1666 -593 2042
rect -559 1666 -543 2042
rect -609 1654 -543 1666
rect -513 2042 -447 2054
rect -513 1666 -497 2042
rect -463 1666 -447 2042
rect -513 1654 -447 1666
rect -417 2042 -351 2054
rect -417 1666 -401 2042
rect -367 1666 -351 2042
rect -417 1654 -351 1666
rect -321 2042 -255 2054
rect -321 1666 -305 2042
rect -271 1666 -255 2042
rect -321 1654 -255 1666
rect -225 2042 -159 2054
rect -225 1666 -209 2042
rect -175 1666 -159 2042
rect -225 1654 -159 1666
rect -129 2042 -63 2054
rect -129 1666 -113 2042
rect -79 1666 -63 2042
rect -129 1654 -63 1666
rect -33 2042 33 2054
rect -33 1666 -17 2042
rect 17 1666 33 2042
rect -33 1654 33 1666
rect 63 2042 129 2054
rect 63 1666 79 2042
rect 113 1666 129 2042
rect 63 1654 129 1666
rect 159 2042 225 2054
rect 159 1666 175 2042
rect 209 1666 225 2042
rect 159 1654 225 1666
rect 255 2042 321 2054
rect 255 1666 271 2042
rect 305 1666 321 2042
rect 255 1654 321 1666
rect 351 2042 417 2054
rect 351 1666 367 2042
rect 401 1666 417 2042
rect 351 1654 417 1666
rect 447 2042 513 2054
rect 447 1666 463 2042
rect 497 1666 513 2042
rect 447 1654 513 1666
rect 543 2042 609 2054
rect 543 1666 559 2042
rect 593 1666 609 2042
rect 543 1654 609 1666
rect 639 2042 705 2054
rect 639 1666 655 2042
rect 689 1666 705 2042
rect 639 1654 705 1666
rect 735 2042 801 2054
rect 735 1666 751 2042
rect 785 1666 801 2042
rect 735 1654 801 1666
rect 831 2042 897 2054
rect 831 1666 847 2042
rect 881 1666 897 2042
rect 831 1654 897 1666
rect 927 2042 989 2054
rect 927 1666 943 2042
rect 977 1666 989 2042
rect 927 1654 989 1666
rect -989 1424 -927 1436
rect -989 1048 -977 1424
rect -943 1048 -927 1424
rect -989 1036 -927 1048
rect -897 1424 -831 1436
rect -897 1048 -881 1424
rect -847 1048 -831 1424
rect -897 1036 -831 1048
rect -801 1424 -735 1436
rect -801 1048 -785 1424
rect -751 1048 -735 1424
rect -801 1036 -735 1048
rect -705 1424 -639 1436
rect -705 1048 -689 1424
rect -655 1048 -639 1424
rect -705 1036 -639 1048
rect -609 1424 -543 1436
rect -609 1048 -593 1424
rect -559 1048 -543 1424
rect -609 1036 -543 1048
rect -513 1424 -447 1436
rect -513 1048 -497 1424
rect -463 1048 -447 1424
rect -513 1036 -447 1048
rect -417 1424 -351 1436
rect -417 1048 -401 1424
rect -367 1048 -351 1424
rect -417 1036 -351 1048
rect -321 1424 -255 1436
rect -321 1048 -305 1424
rect -271 1048 -255 1424
rect -321 1036 -255 1048
rect -225 1424 -159 1436
rect -225 1048 -209 1424
rect -175 1048 -159 1424
rect -225 1036 -159 1048
rect -129 1424 -63 1436
rect -129 1048 -113 1424
rect -79 1048 -63 1424
rect -129 1036 -63 1048
rect -33 1424 33 1436
rect -33 1048 -17 1424
rect 17 1048 33 1424
rect -33 1036 33 1048
rect 63 1424 129 1436
rect 63 1048 79 1424
rect 113 1048 129 1424
rect 63 1036 129 1048
rect 159 1424 225 1436
rect 159 1048 175 1424
rect 209 1048 225 1424
rect 159 1036 225 1048
rect 255 1424 321 1436
rect 255 1048 271 1424
rect 305 1048 321 1424
rect 255 1036 321 1048
rect 351 1424 417 1436
rect 351 1048 367 1424
rect 401 1048 417 1424
rect 351 1036 417 1048
rect 447 1424 513 1436
rect 447 1048 463 1424
rect 497 1048 513 1424
rect 447 1036 513 1048
rect 543 1424 609 1436
rect 543 1048 559 1424
rect 593 1048 609 1424
rect 543 1036 609 1048
rect 639 1424 705 1436
rect 639 1048 655 1424
rect 689 1048 705 1424
rect 639 1036 705 1048
rect 735 1424 801 1436
rect 735 1048 751 1424
rect 785 1048 801 1424
rect 735 1036 801 1048
rect 831 1424 897 1436
rect 831 1048 847 1424
rect 881 1048 897 1424
rect 831 1036 897 1048
rect 927 1424 989 1436
rect 927 1048 943 1424
rect 977 1048 989 1424
rect 927 1036 989 1048
rect -989 806 -927 818
rect -989 430 -977 806
rect -943 430 -927 806
rect -989 418 -927 430
rect -897 806 -831 818
rect -897 430 -881 806
rect -847 430 -831 806
rect -897 418 -831 430
rect -801 806 -735 818
rect -801 430 -785 806
rect -751 430 -735 806
rect -801 418 -735 430
rect -705 806 -639 818
rect -705 430 -689 806
rect -655 430 -639 806
rect -705 418 -639 430
rect -609 806 -543 818
rect -609 430 -593 806
rect -559 430 -543 806
rect -609 418 -543 430
rect -513 806 -447 818
rect -513 430 -497 806
rect -463 430 -447 806
rect -513 418 -447 430
rect -417 806 -351 818
rect -417 430 -401 806
rect -367 430 -351 806
rect -417 418 -351 430
rect -321 806 -255 818
rect -321 430 -305 806
rect -271 430 -255 806
rect -321 418 -255 430
rect -225 806 -159 818
rect -225 430 -209 806
rect -175 430 -159 806
rect -225 418 -159 430
rect -129 806 -63 818
rect -129 430 -113 806
rect -79 430 -63 806
rect -129 418 -63 430
rect -33 806 33 818
rect -33 430 -17 806
rect 17 430 33 806
rect -33 418 33 430
rect 63 806 129 818
rect 63 430 79 806
rect 113 430 129 806
rect 63 418 129 430
rect 159 806 225 818
rect 159 430 175 806
rect 209 430 225 806
rect 159 418 225 430
rect 255 806 321 818
rect 255 430 271 806
rect 305 430 321 806
rect 255 418 321 430
rect 351 806 417 818
rect 351 430 367 806
rect 401 430 417 806
rect 351 418 417 430
rect 447 806 513 818
rect 447 430 463 806
rect 497 430 513 806
rect 447 418 513 430
rect 543 806 609 818
rect 543 430 559 806
rect 593 430 609 806
rect 543 418 609 430
rect 639 806 705 818
rect 639 430 655 806
rect 689 430 705 806
rect 639 418 705 430
rect 735 806 801 818
rect 735 430 751 806
rect 785 430 801 806
rect 735 418 801 430
rect 831 806 897 818
rect 831 430 847 806
rect 881 430 897 806
rect 831 418 897 430
rect 927 806 989 818
rect 927 430 943 806
rect 977 430 989 806
rect 927 418 989 430
rect -989 188 -927 200
rect -989 -188 -977 188
rect -943 -188 -927 188
rect -989 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 989 200
rect 927 -188 943 188
rect 977 -188 989 188
rect 927 -200 989 -188
rect -989 -430 -927 -418
rect -989 -806 -977 -430
rect -943 -806 -927 -430
rect -989 -818 -927 -806
rect -897 -430 -831 -418
rect -897 -806 -881 -430
rect -847 -806 -831 -430
rect -897 -818 -831 -806
rect -801 -430 -735 -418
rect -801 -806 -785 -430
rect -751 -806 -735 -430
rect -801 -818 -735 -806
rect -705 -430 -639 -418
rect -705 -806 -689 -430
rect -655 -806 -639 -430
rect -705 -818 -639 -806
rect -609 -430 -543 -418
rect -609 -806 -593 -430
rect -559 -806 -543 -430
rect -609 -818 -543 -806
rect -513 -430 -447 -418
rect -513 -806 -497 -430
rect -463 -806 -447 -430
rect -513 -818 -447 -806
rect -417 -430 -351 -418
rect -417 -806 -401 -430
rect -367 -806 -351 -430
rect -417 -818 -351 -806
rect -321 -430 -255 -418
rect -321 -806 -305 -430
rect -271 -806 -255 -430
rect -321 -818 -255 -806
rect -225 -430 -159 -418
rect -225 -806 -209 -430
rect -175 -806 -159 -430
rect -225 -818 -159 -806
rect -129 -430 -63 -418
rect -129 -806 -113 -430
rect -79 -806 -63 -430
rect -129 -818 -63 -806
rect -33 -430 33 -418
rect -33 -806 -17 -430
rect 17 -806 33 -430
rect -33 -818 33 -806
rect 63 -430 129 -418
rect 63 -806 79 -430
rect 113 -806 129 -430
rect 63 -818 129 -806
rect 159 -430 225 -418
rect 159 -806 175 -430
rect 209 -806 225 -430
rect 159 -818 225 -806
rect 255 -430 321 -418
rect 255 -806 271 -430
rect 305 -806 321 -430
rect 255 -818 321 -806
rect 351 -430 417 -418
rect 351 -806 367 -430
rect 401 -806 417 -430
rect 351 -818 417 -806
rect 447 -430 513 -418
rect 447 -806 463 -430
rect 497 -806 513 -430
rect 447 -818 513 -806
rect 543 -430 609 -418
rect 543 -806 559 -430
rect 593 -806 609 -430
rect 543 -818 609 -806
rect 639 -430 705 -418
rect 639 -806 655 -430
rect 689 -806 705 -430
rect 639 -818 705 -806
rect 735 -430 801 -418
rect 735 -806 751 -430
rect 785 -806 801 -430
rect 735 -818 801 -806
rect 831 -430 897 -418
rect 831 -806 847 -430
rect 881 -806 897 -430
rect 831 -818 897 -806
rect 927 -430 989 -418
rect 927 -806 943 -430
rect 977 -806 989 -430
rect 927 -818 989 -806
rect -989 -1048 -927 -1036
rect -989 -1424 -977 -1048
rect -943 -1424 -927 -1048
rect -989 -1436 -927 -1424
rect -897 -1048 -831 -1036
rect -897 -1424 -881 -1048
rect -847 -1424 -831 -1048
rect -897 -1436 -831 -1424
rect -801 -1048 -735 -1036
rect -801 -1424 -785 -1048
rect -751 -1424 -735 -1048
rect -801 -1436 -735 -1424
rect -705 -1048 -639 -1036
rect -705 -1424 -689 -1048
rect -655 -1424 -639 -1048
rect -705 -1436 -639 -1424
rect -609 -1048 -543 -1036
rect -609 -1424 -593 -1048
rect -559 -1424 -543 -1048
rect -609 -1436 -543 -1424
rect -513 -1048 -447 -1036
rect -513 -1424 -497 -1048
rect -463 -1424 -447 -1048
rect -513 -1436 -447 -1424
rect -417 -1048 -351 -1036
rect -417 -1424 -401 -1048
rect -367 -1424 -351 -1048
rect -417 -1436 -351 -1424
rect -321 -1048 -255 -1036
rect -321 -1424 -305 -1048
rect -271 -1424 -255 -1048
rect -321 -1436 -255 -1424
rect -225 -1048 -159 -1036
rect -225 -1424 -209 -1048
rect -175 -1424 -159 -1048
rect -225 -1436 -159 -1424
rect -129 -1048 -63 -1036
rect -129 -1424 -113 -1048
rect -79 -1424 -63 -1048
rect -129 -1436 -63 -1424
rect -33 -1048 33 -1036
rect -33 -1424 -17 -1048
rect 17 -1424 33 -1048
rect -33 -1436 33 -1424
rect 63 -1048 129 -1036
rect 63 -1424 79 -1048
rect 113 -1424 129 -1048
rect 63 -1436 129 -1424
rect 159 -1048 225 -1036
rect 159 -1424 175 -1048
rect 209 -1424 225 -1048
rect 159 -1436 225 -1424
rect 255 -1048 321 -1036
rect 255 -1424 271 -1048
rect 305 -1424 321 -1048
rect 255 -1436 321 -1424
rect 351 -1048 417 -1036
rect 351 -1424 367 -1048
rect 401 -1424 417 -1048
rect 351 -1436 417 -1424
rect 447 -1048 513 -1036
rect 447 -1424 463 -1048
rect 497 -1424 513 -1048
rect 447 -1436 513 -1424
rect 543 -1048 609 -1036
rect 543 -1424 559 -1048
rect 593 -1424 609 -1048
rect 543 -1436 609 -1424
rect 639 -1048 705 -1036
rect 639 -1424 655 -1048
rect 689 -1424 705 -1048
rect 639 -1436 705 -1424
rect 735 -1048 801 -1036
rect 735 -1424 751 -1048
rect 785 -1424 801 -1048
rect 735 -1436 801 -1424
rect 831 -1048 897 -1036
rect 831 -1424 847 -1048
rect 881 -1424 897 -1048
rect 831 -1436 897 -1424
rect 927 -1048 989 -1036
rect 927 -1424 943 -1048
rect 977 -1424 989 -1048
rect 927 -1436 989 -1424
rect -989 -1666 -927 -1654
rect -989 -2042 -977 -1666
rect -943 -2042 -927 -1666
rect -989 -2054 -927 -2042
rect -897 -1666 -831 -1654
rect -897 -2042 -881 -1666
rect -847 -2042 -831 -1666
rect -897 -2054 -831 -2042
rect -801 -1666 -735 -1654
rect -801 -2042 -785 -1666
rect -751 -2042 -735 -1666
rect -801 -2054 -735 -2042
rect -705 -1666 -639 -1654
rect -705 -2042 -689 -1666
rect -655 -2042 -639 -1666
rect -705 -2054 -639 -2042
rect -609 -1666 -543 -1654
rect -609 -2042 -593 -1666
rect -559 -2042 -543 -1666
rect -609 -2054 -543 -2042
rect -513 -1666 -447 -1654
rect -513 -2042 -497 -1666
rect -463 -2042 -447 -1666
rect -513 -2054 -447 -2042
rect -417 -1666 -351 -1654
rect -417 -2042 -401 -1666
rect -367 -2042 -351 -1666
rect -417 -2054 -351 -2042
rect -321 -1666 -255 -1654
rect -321 -2042 -305 -1666
rect -271 -2042 -255 -1666
rect -321 -2054 -255 -2042
rect -225 -1666 -159 -1654
rect -225 -2042 -209 -1666
rect -175 -2042 -159 -1666
rect -225 -2054 -159 -2042
rect -129 -1666 -63 -1654
rect -129 -2042 -113 -1666
rect -79 -2042 -63 -1666
rect -129 -2054 -63 -2042
rect -33 -1666 33 -1654
rect -33 -2042 -17 -1666
rect 17 -2042 33 -1666
rect -33 -2054 33 -2042
rect 63 -1666 129 -1654
rect 63 -2042 79 -1666
rect 113 -2042 129 -1666
rect 63 -2054 129 -2042
rect 159 -1666 225 -1654
rect 159 -2042 175 -1666
rect 209 -2042 225 -1666
rect 159 -2054 225 -2042
rect 255 -1666 321 -1654
rect 255 -2042 271 -1666
rect 305 -2042 321 -1666
rect 255 -2054 321 -2042
rect 351 -1666 417 -1654
rect 351 -2042 367 -1666
rect 401 -2042 417 -1666
rect 351 -2054 417 -2042
rect 447 -1666 513 -1654
rect 447 -2042 463 -1666
rect 497 -2042 513 -1666
rect 447 -2054 513 -2042
rect 543 -1666 609 -1654
rect 543 -2042 559 -1666
rect 593 -2042 609 -1666
rect 543 -2054 609 -2042
rect 639 -1666 705 -1654
rect 639 -2042 655 -1666
rect 689 -2042 705 -1666
rect 639 -2054 705 -2042
rect 735 -1666 801 -1654
rect 735 -2042 751 -1666
rect 785 -2042 801 -1666
rect 735 -2054 801 -2042
rect 831 -1666 897 -1654
rect 831 -2042 847 -1666
rect 881 -2042 897 -1666
rect 831 -2054 897 -2042
rect 927 -1666 989 -1654
rect 927 -2042 943 -1666
rect 977 -2042 989 -1666
rect 927 -2054 989 -2042
rect -989 -2284 -927 -2272
rect -989 -2660 -977 -2284
rect -943 -2660 -927 -2284
rect -989 -2672 -927 -2660
rect -897 -2284 -831 -2272
rect -897 -2660 -881 -2284
rect -847 -2660 -831 -2284
rect -897 -2672 -831 -2660
rect -801 -2284 -735 -2272
rect -801 -2660 -785 -2284
rect -751 -2660 -735 -2284
rect -801 -2672 -735 -2660
rect -705 -2284 -639 -2272
rect -705 -2660 -689 -2284
rect -655 -2660 -639 -2284
rect -705 -2672 -639 -2660
rect -609 -2284 -543 -2272
rect -609 -2660 -593 -2284
rect -559 -2660 -543 -2284
rect -609 -2672 -543 -2660
rect -513 -2284 -447 -2272
rect -513 -2660 -497 -2284
rect -463 -2660 -447 -2284
rect -513 -2672 -447 -2660
rect -417 -2284 -351 -2272
rect -417 -2660 -401 -2284
rect -367 -2660 -351 -2284
rect -417 -2672 -351 -2660
rect -321 -2284 -255 -2272
rect -321 -2660 -305 -2284
rect -271 -2660 -255 -2284
rect -321 -2672 -255 -2660
rect -225 -2284 -159 -2272
rect -225 -2660 -209 -2284
rect -175 -2660 -159 -2284
rect -225 -2672 -159 -2660
rect -129 -2284 -63 -2272
rect -129 -2660 -113 -2284
rect -79 -2660 -63 -2284
rect -129 -2672 -63 -2660
rect -33 -2284 33 -2272
rect -33 -2660 -17 -2284
rect 17 -2660 33 -2284
rect -33 -2672 33 -2660
rect 63 -2284 129 -2272
rect 63 -2660 79 -2284
rect 113 -2660 129 -2284
rect 63 -2672 129 -2660
rect 159 -2284 225 -2272
rect 159 -2660 175 -2284
rect 209 -2660 225 -2284
rect 159 -2672 225 -2660
rect 255 -2284 321 -2272
rect 255 -2660 271 -2284
rect 305 -2660 321 -2284
rect 255 -2672 321 -2660
rect 351 -2284 417 -2272
rect 351 -2660 367 -2284
rect 401 -2660 417 -2284
rect 351 -2672 417 -2660
rect 447 -2284 513 -2272
rect 447 -2660 463 -2284
rect 497 -2660 513 -2284
rect 447 -2672 513 -2660
rect 543 -2284 609 -2272
rect 543 -2660 559 -2284
rect 593 -2660 609 -2284
rect 543 -2672 609 -2660
rect 639 -2284 705 -2272
rect 639 -2660 655 -2284
rect 689 -2660 705 -2284
rect 639 -2672 705 -2660
rect 735 -2284 801 -2272
rect 735 -2660 751 -2284
rect 785 -2660 801 -2284
rect 735 -2672 801 -2660
rect 831 -2284 897 -2272
rect 831 -2660 847 -2284
rect 881 -2660 897 -2284
rect 831 -2672 897 -2660
rect 927 -2284 989 -2272
rect 927 -2660 943 -2284
rect 977 -2660 989 -2284
rect 927 -2672 989 -2660
<< ndiffc >>
rect -977 2284 -943 2660
rect -881 2284 -847 2660
rect -785 2284 -751 2660
rect -689 2284 -655 2660
rect -593 2284 -559 2660
rect -497 2284 -463 2660
rect -401 2284 -367 2660
rect -305 2284 -271 2660
rect -209 2284 -175 2660
rect -113 2284 -79 2660
rect -17 2284 17 2660
rect 79 2284 113 2660
rect 175 2284 209 2660
rect 271 2284 305 2660
rect 367 2284 401 2660
rect 463 2284 497 2660
rect 559 2284 593 2660
rect 655 2284 689 2660
rect 751 2284 785 2660
rect 847 2284 881 2660
rect 943 2284 977 2660
rect -977 1666 -943 2042
rect -881 1666 -847 2042
rect -785 1666 -751 2042
rect -689 1666 -655 2042
rect -593 1666 -559 2042
rect -497 1666 -463 2042
rect -401 1666 -367 2042
rect -305 1666 -271 2042
rect -209 1666 -175 2042
rect -113 1666 -79 2042
rect -17 1666 17 2042
rect 79 1666 113 2042
rect 175 1666 209 2042
rect 271 1666 305 2042
rect 367 1666 401 2042
rect 463 1666 497 2042
rect 559 1666 593 2042
rect 655 1666 689 2042
rect 751 1666 785 2042
rect 847 1666 881 2042
rect 943 1666 977 2042
rect -977 1048 -943 1424
rect -881 1048 -847 1424
rect -785 1048 -751 1424
rect -689 1048 -655 1424
rect -593 1048 -559 1424
rect -497 1048 -463 1424
rect -401 1048 -367 1424
rect -305 1048 -271 1424
rect -209 1048 -175 1424
rect -113 1048 -79 1424
rect -17 1048 17 1424
rect 79 1048 113 1424
rect 175 1048 209 1424
rect 271 1048 305 1424
rect 367 1048 401 1424
rect 463 1048 497 1424
rect 559 1048 593 1424
rect 655 1048 689 1424
rect 751 1048 785 1424
rect 847 1048 881 1424
rect 943 1048 977 1424
rect -977 430 -943 806
rect -881 430 -847 806
rect -785 430 -751 806
rect -689 430 -655 806
rect -593 430 -559 806
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect 559 430 593 806
rect 655 430 689 806
rect 751 430 785 806
rect 847 430 881 806
rect 943 430 977 806
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect -977 -806 -943 -430
rect -881 -806 -847 -430
rect -785 -806 -751 -430
rect -689 -806 -655 -430
rect -593 -806 -559 -430
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect 559 -806 593 -430
rect 655 -806 689 -430
rect 751 -806 785 -430
rect 847 -806 881 -430
rect 943 -806 977 -430
rect -977 -1424 -943 -1048
rect -881 -1424 -847 -1048
rect -785 -1424 -751 -1048
rect -689 -1424 -655 -1048
rect -593 -1424 -559 -1048
rect -497 -1424 -463 -1048
rect -401 -1424 -367 -1048
rect -305 -1424 -271 -1048
rect -209 -1424 -175 -1048
rect -113 -1424 -79 -1048
rect -17 -1424 17 -1048
rect 79 -1424 113 -1048
rect 175 -1424 209 -1048
rect 271 -1424 305 -1048
rect 367 -1424 401 -1048
rect 463 -1424 497 -1048
rect 559 -1424 593 -1048
rect 655 -1424 689 -1048
rect 751 -1424 785 -1048
rect 847 -1424 881 -1048
rect 943 -1424 977 -1048
rect -977 -2042 -943 -1666
rect -881 -2042 -847 -1666
rect -785 -2042 -751 -1666
rect -689 -2042 -655 -1666
rect -593 -2042 -559 -1666
rect -497 -2042 -463 -1666
rect -401 -2042 -367 -1666
rect -305 -2042 -271 -1666
rect -209 -2042 -175 -1666
rect -113 -2042 -79 -1666
rect -17 -2042 17 -1666
rect 79 -2042 113 -1666
rect 175 -2042 209 -1666
rect 271 -2042 305 -1666
rect 367 -2042 401 -1666
rect 463 -2042 497 -1666
rect 559 -2042 593 -1666
rect 655 -2042 689 -1666
rect 751 -2042 785 -1666
rect 847 -2042 881 -1666
rect 943 -2042 977 -1666
rect -977 -2660 -943 -2284
rect -881 -2660 -847 -2284
rect -785 -2660 -751 -2284
rect -689 -2660 -655 -2284
rect -593 -2660 -559 -2284
rect -497 -2660 -463 -2284
rect -401 -2660 -367 -2284
rect -305 -2660 -271 -2284
rect -209 -2660 -175 -2284
rect -113 -2660 -79 -2284
rect -17 -2660 17 -2284
rect 79 -2660 113 -2284
rect 175 -2660 209 -2284
rect 271 -2660 305 -2284
rect 367 -2660 401 -2284
rect 463 -2660 497 -2284
rect 559 -2660 593 -2284
rect 655 -2660 689 -2284
rect 751 -2660 785 -2284
rect 847 -2660 881 -2284
rect 943 -2660 977 -2284
<< psubdiff >>
rect -1091 2812 -995 2846
rect 995 2812 1091 2846
rect -1091 2750 -1057 2812
rect 1057 2750 1091 2812
rect -1091 -2812 -1057 -2750
rect 1057 -2812 1091 -2750
rect -1091 -2846 -995 -2812
rect 995 -2846 1091 -2812
<< psubdiffcont >>
rect -995 2812 995 2846
rect -1091 -2750 -1057 2750
rect 1057 -2750 1091 2750
rect -995 -2846 995 -2812
<< poly >>
rect -849 2744 -783 2760
rect -849 2710 -833 2744
rect -799 2710 -783 2744
rect -927 2672 -897 2698
rect -849 2694 -783 2710
rect -657 2744 -591 2760
rect -657 2710 -641 2744
rect -607 2710 -591 2744
rect -831 2672 -801 2694
rect -735 2672 -705 2698
rect -657 2694 -591 2710
rect -465 2744 -399 2760
rect -465 2710 -449 2744
rect -415 2710 -399 2744
rect -639 2672 -609 2694
rect -543 2672 -513 2698
rect -465 2694 -399 2710
rect -273 2744 -207 2760
rect -273 2710 -257 2744
rect -223 2710 -207 2744
rect -447 2672 -417 2694
rect -351 2672 -321 2698
rect -273 2694 -207 2710
rect -81 2744 -15 2760
rect -81 2710 -65 2744
rect -31 2710 -15 2744
rect -255 2672 -225 2694
rect -159 2672 -129 2698
rect -81 2694 -15 2710
rect 111 2744 177 2760
rect 111 2710 127 2744
rect 161 2710 177 2744
rect -63 2672 -33 2694
rect 33 2672 63 2698
rect 111 2694 177 2710
rect 303 2744 369 2760
rect 303 2710 319 2744
rect 353 2710 369 2744
rect 129 2672 159 2694
rect 225 2672 255 2698
rect 303 2694 369 2710
rect 495 2744 561 2760
rect 495 2710 511 2744
rect 545 2710 561 2744
rect 321 2672 351 2694
rect 417 2672 447 2698
rect 495 2694 561 2710
rect 687 2744 753 2760
rect 687 2710 703 2744
rect 737 2710 753 2744
rect 513 2672 543 2694
rect 609 2672 639 2698
rect 687 2694 753 2710
rect 879 2744 945 2760
rect 879 2710 895 2744
rect 929 2710 945 2744
rect 705 2672 735 2694
rect 801 2672 831 2698
rect 879 2694 945 2710
rect 897 2672 927 2694
rect -927 2250 -897 2272
rect -945 2234 -879 2250
rect -831 2246 -801 2272
rect -735 2250 -705 2272
rect -945 2200 -929 2234
rect -895 2200 -879 2234
rect -945 2184 -879 2200
rect -753 2234 -687 2250
rect -639 2246 -609 2272
rect -543 2250 -513 2272
rect -753 2200 -737 2234
rect -703 2200 -687 2234
rect -753 2184 -687 2200
rect -561 2234 -495 2250
rect -447 2246 -417 2272
rect -351 2250 -321 2272
rect -561 2200 -545 2234
rect -511 2200 -495 2234
rect -561 2184 -495 2200
rect -369 2234 -303 2250
rect -255 2246 -225 2272
rect -159 2250 -129 2272
rect -369 2200 -353 2234
rect -319 2200 -303 2234
rect -369 2184 -303 2200
rect -177 2234 -111 2250
rect -63 2246 -33 2272
rect 33 2250 63 2272
rect -177 2200 -161 2234
rect -127 2200 -111 2234
rect -177 2184 -111 2200
rect 15 2234 81 2250
rect 129 2246 159 2272
rect 225 2250 255 2272
rect 15 2200 31 2234
rect 65 2200 81 2234
rect 15 2184 81 2200
rect 207 2234 273 2250
rect 321 2246 351 2272
rect 417 2250 447 2272
rect 207 2200 223 2234
rect 257 2200 273 2234
rect 207 2184 273 2200
rect 399 2234 465 2250
rect 513 2246 543 2272
rect 609 2250 639 2272
rect 399 2200 415 2234
rect 449 2200 465 2234
rect 399 2184 465 2200
rect 591 2234 657 2250
rect 705 2246 735 2272
rect 801 2250 831 2272
rect 591 2200 607 2234
rect 641 2200 657 2234
rect 591 2184 657 2200
rect 783 2234 849 2250
rect 897 2246 927 2272
rect 783 2200 799 2234
rect 833 2200 849 2234
rect 783 2184 849 2200
rect -945 2126 -879 2142
rect -945 2092 -929 2126
rect -895 2092 -879 2126
rect -945 2076 -879 2092
rect -753 2126 -687 2142
rect -753 2092 -737 2126
rect -703 2092 -687 2126
rect -927 2054 -897 2076
rect -831 2054 -801 2080
rect -753 2076 -687 2092
rect -561 2126 -495 2142
rect -561 2092 -545 2126
rect -511 2092 -495 2126
rect -735 2054 -705 2076
rect -639 2054 -609 2080
rect -561 2076 -495 2092
rect -369 2126 -303 2142
rect -369 2092 -353 2126
rect -319 2092 -303 2126
rect -543 2054 -513 2076
rect -447 2054 -417 2080
rect -369 2076 -303 2092
rect -177 2126 -111 2142
rect -177 2092 -161 2126
rect -127 2092 -111 2126
rect -351 2054 -321 2076
rect -255 2054 -225 2080
rect -177 2076 -111 2092
rect 15 2126 81 2142
rect 15 2092 31 2126
rect 65 2092 81 2126
rect -159 2054 -129 2076
rect -63 2054 -33 2080
rect 15 2076 81 2092
rect 207 2126 273 2142
rect 207 2092 223 2126
rect 257 2092 273 2126
rect 33 2054 63 2076
rect 129 2054 159 2080
rect 207 2076 273 2092
rect 399 2126 465 2142
rect 399 2092 415 2126
rect 449 2092 465 2126
rect 225 2054 255 2076
rect 321 2054 351 2080
rect 399 2076 465 2092
rect 591 2126 657 2142
rect 591 2092 607 2126
rect 641 2092 657 2126
rect 417 2054 447 2076
rect 513 2054 543 2080
rect 591 2076 657 2092
rect 783 2126 849 2142
rect 783 2092 799 2126
rect 833 2092 849 2126
rect 609 2054 639 2076
rect 705 2054 735 2080
rect 783 2076 849 2092
rect 801 2054 831 2076
rect 897 2054 927 2080
rect -927 1628 -897 1654
rect -831 1632 -801 1654
rect -849 1616 -783 1632
rect -735 1628 -705 1654
rect -639 1632 -609 1654
rect -849 1582 -833 1616
rect -799 1582 -783 1616
rect -849 1566 -783 1582
rect -657 1616 -591 1632
rect -543 1628 -513 1654
rect -447 1632 -417 1654
rect -657 1582 -641 1616
rect -607 1582 -591 1616
rect -657 1566 -591 1582
rect -465 1616 -399 1632
rect -351 1628 -321 1654
rect -255 1632 -225 1654
rect -465 1582 -449 1616
rect -415 1582 -399 1616
rect -465 1566 -399 1582
rect -273 1616 -207 1632
rect -159 1628 -129 1654
rect -63 1632 -33 1654
rect -273 1582 -257 1616
rect -223 1582 -207 1616
rect -273 1566 -207 1582
rect -81 1616 -15 1632
rect 33 1628 63 1654
rect 129 1632 159 1654
rect -81 1582 -65 1616
rect -31 1582 -15 1616
rect -81 1566 -15 1582
rect 111 1616 177 1632
rect 225 1628 255 1654
rect 321 1632 351 1654
rect 111 1582 127 1616
rect 161 1582 177 1616
rect 111 1566 177 1582
rect 303 1616 369 1632
rect 417 1628 447 1654
rect 513 1632 543 1654
rect 303 1582 319 1616
rect 353 1582 369 1616
rect 303 1566 369 1582
rect 495 1616 561 1632
rect 609 1628 639 1654
rect 705 1632 735 1654
rect 495 1582 511 1616
rect 545 1582 561 1616
rect 495 1566 561 1582
rect 687 1616 753 1632
rect 801 1628 831 1654
rect 897 1632 927 1654
rect 687 1582 703 1616
rect 737 1582 753 1616
rect 687 1566 753 1582
rect 879 1616 945 1632
rect 879 1582 895 1616
rect 929 1582 945 1616
rect 879 1566 945 1582
rect -849 1508 -783 1524
rect -849 1474 -833 1508
rect -799 1474 -783 1508
rect -927 1436 -897 1462
rect -849 1458 -783 1474
rect -657 1508 -591 1524
rect -657 1474 -641 1508
rect -607 1474 -591 1508
rect -831 1436 -801 1458
rect -735 1436 -705 1462
rect -657 1458 -591 1474
rect -465 1508 -399 1524
rect -465 1474 -449 1508
rect -415 1474 -399 1508
rect -639 1436 -609 1458
rect -543 1436 -513 1462
rect -465 1458 -399 1474
rect -273 1508 -207 1524
rect -273 1474 -257 1508
rect -223 1474 -207 1508
rect -447 1436 -417 1458
rect -351 1436 -321 1462
rect -273 1458 -207 1474
rect -81 1508 -15 1524
rect -81 1474 -65 1508
rect -31 1474 -15 1508
rect -255 1436 -225 1458
rect -159 1436 -129 1462
rect -81 1458 -15 1474
rect 111 1508 177 1524
rect 111 1474 127 1508
rect 161 1474 177 1508
rect -63 1436 -33 1458
rect 33 1436 63 1462
rect 111 1458 177 1474
rect 303 1508 369 1524
rect 303 1474 319 1508
rect 353 1474 369 1508
rect 129 1436 159 1458
rect 225 1436 255 1462
rect 303 1458 369 1474
rect 495 1508 561 1524
rect 495 1474 511 1508
rect 545 1474 561 1508
rect 321 1436 351 1458
rect 417 1436 447 1462
rect 495 1458 561 1474
rect 687 1508 753 1524
rect 687 1474 703 1508
rect 737 1474 753 1508
rect 513 1436 543 1458
rect 609 1436 639 1462
rect 687 1458 753 1474
rect 879 1508 945 1524
rect 879 1474 895 1508
rect 929 1474 945 1508
rect 705 1436 735 1458
rect 801 1436 831 1462
rect 879 1458 945 1474
rect 897 1436 927 1458
rect -927 1014 -897 1036
rect -945 998 -879 1014
rect -831 1010 -801 1036
rect -735 1014 -705 1036
rect -945 964 -929 998
rect -895 964 -879 998
rect -945 948 -879 964
rect -753 998 -687 1014
rect -639 1010 -609 1036
rect -543 1014 -513 1036
rect -753 964 -737 998
rect -703 964 -687 998
rect -753 948 -687 964
rect -561 998 -495 1014
rect -447 1010 -417 1036
rect -351 1014 -321 1036
rect -561 964 -545 998
rect -511 964 -495 998
rect -561 948 -495 964
rect -369 998 -303 1014
rect -255 1010 -225 1036
rect -159 1014 -129 1036
rect -369 964 -353 998
rect -319 964 -303 998
rect -369 948 -303 964
rect -177 998 -111 1014
rect -63 1010 -33 1036
rect 33 1014 63 1036
rect -177 964 -161 998
rect -127 964 -111 998
rect -177 948 -111 964
rect 15 998 81 1014
rect 129 1010 159 1036
rect 225 1014 255 1036
rect 15 964 31 998
rect 65 964 81 998
rect 15 948 81 964
rect 207 998 273 1014
rect 321 1010 351 1036
rect 417 1014 447 1036
rect 207 964 223 998
rect 257 964 273 998
rect 207 948 273 964
rect 399 998 465 1014
rect 513 1010 543 1036
rect 609 1014 639 1036
rect 399 964 415 998
rect 449 964 465 998
rect 399 948 465 964
rect 591 998 657 1014
rect 705 1010 735 1036
rect 801 1014 831 1036
rect 591 964 607 998
rect 641 964 657 998
rect 591 948 657 964
rect 783 998 849 1014
rect 897 1010 927 1036
rect 783 964 799 998
rect 833 964 849 998
rect 783 948 849 964
rect -945 890 -879 906
rect -945 856 -929 890
rect -895 856 -879 890
rect -945 840 -879 856
rect -753 890 -687 906
rect -753 856 -737 890
rect -703 856 -687 890
rect -927 818 -897 840
rect -831 818 -801 844
rect -753 840 -687 856
rect -561 890 -495 906
rect -561 856 -545 890
rect -511 856 -495 890
rect -735 818 -705 840
rect -639 818 -609 844
rect -561 840 -495 856
rect -369 890 -303 906
rect -369 856 -353 890
rect -319 856 -303 890
rect -543 818 -513 840
rect -447 818 -417 844
rect -369 840 -303 856
rect -177 890 -111 906
rect -177 856 -161 890
rect -127 856 -111 890
rect -351 818 -321 840
rect -255 818 -225 844
rect -177 840 -111 856
rect 15 890 81 906
rect 15 856 31 890
rect 65 856 81 890
rect -159 818 -129 840
rect -63 818 -33 844
rect 15 840 81 856
rect 207 890 273 906
rect 207 856 223 890
rect 257 856 273 890
rect 33 818 63 840
rect 129 818 159 844
rect 207 840 273 856
rect 399 890 465 906
rect 399 856 415 890
rect 449 856 465 890
rect 225 818 255 840
rect 321 818 351 844
rect 399 840 465 856
rect 591 890 657 906
rect 591 856 607 890
rect 641 856 657 890
rect 417 818 447 840
rect 513 818 543 844
rect 591 840 657 856
rect 783 890 849 906
rect 783 856 799 890
rect 833 856 849 890
rect 609 818 639 840
rect 705 818 735 844
rect 783 840 849 856
rect 801 818 831 840
rect 897 818 927 844
rect -927 392 -897 418
rect -831 396 -801 418
rect -849 380 -783 396
rect -735 392 -705 418
rect -639 396 -609 418
rect -849 346 -833 380
rect -799 346 -783 380
rect -849 330 -783 346
rect -657 380 -591 396
rect -543 392 -513 418
rect -447 396 -417 418
rect -657 346 -641 380
rect -607 346 -591 380
rect -657 330 -591 346
rect -465 380 -399 396
rect -351 392 -321 418
rect -255 396 -225 418
rect -465 346 -449 380
rect -415 346 -399 380
rect -465 330 -399 346
rect -273 380 -207 396
rect -159 392 -129 418
rect -63 396 -33 418
rect -273 346 -257 380
rect -223 346 -207 380
rect -273 330 -207 346
rect -81 380 -15 396
rect 33 392 63 418
rect 129 396 159 418
rect -81 346 -65 380
rect -31 346 -15 380
rect -81 330 -15 346
rect 111 380 177 396
rect 225 392 255 418
rect 321 396 351 418
rect 111 346 127 380
rect 161 346 177 380
rect 111 330 177 346
rect 303 380 369 396
rect 417 392 447 418
rect 513 396 543 418
rect 303 346 319 380
rect 353 346 369 380
rect 303 330 369 346
rect 495 380 561 396
rect 609 392 639 418
rect 705 396 735 418
rect 495 346 511 380
rect 545 346 561 380
rect 495 330 561 346
rect 687 380 753 396
rect 801 392 831 418
rect 897 396 927 418
rect 687 346 703 380
rect 737 346 753 380
rect 687 330 753 346
rect 879 380 945 396
rect 879 346 895 380
rect 929 346 945 380
rect 879 330 945 346
rect -849 272 -783 288
rect -849 238 -833 272
rect -799 238 -783 272
rect -927 200 -897 226
rect -849 222 -783 238
rect -657 272 -591 288
rect -657 238 -641 272
rect -607 238 -591 272
rect -831 200 -801 222
rect -735 200 -705 226
rect -657 222 -591 238
rect -465 272 -399 288
rect -465 238 -449 272
rect -415 238 -399 272
rect -639 200 -609 222
rect -543 200 -513 226
rect -465 222 -399 238
rect -273 272 -207 288
rect -273 238 -257 272
rect -223 238 -207 272
rect -447 200 -417 222
rect -351 200 -321 226
rect -273 222 -207 238
rect -81 272 -15 288
rect -81 238 -65 272
rect -31 238 -15 272
rect -255 200 -225 222
rect -159 200 -129 226
rect -81 222 -15 238
rect 111 272 177 288
rect 111 238 127 272
rect 161 238 177 272
rect -63 200 -33 222
rect 33 200 63 226
rect 111 222 177 238
rect 303 272 369 288
rect 303 238 319 272
rect 353 238 369 272
rect 129 200 159 222
rect 225 200 255 226
rect 303 222 369 238
rect 495 272 561 288
rect 495 238 511 272
rect 545 238 561 272
rect 321 200 351 222
rect 417 200 447 226
rect 495 222 561 238
rect 687 272 753 288
rect 687 238 703 272
rect 737 238 753 272
rect 513 200 543 222
rect 609 200 639 226
rect 687 222 753 238
rect 879 272 945 288
rect 879 238 895 272
rect 929 238 945 272
rect 705 200 735 222
rect 801 200 831 226
rect 879 222 945 238
rect 897 200 927 222
rect -927 -222 -897 -200
rect -945 -238 -879 -222
rect -831 -226 -801 -200
rect -735 -222 -705 -200
rect -945 -272 -929 -238
rect -895 -272 -879 -238
rect -945 -288 -879 -272
rect -753 -238 -687 -222
rect -639 -226 -609 -200
rect -543 -222 -513 -200
rect -753 -272 -737 -238
rect -703 -272 -687 -238
rect -753 -288 -687 -272
rect -561 -238 -495 -222
rect -447 -226 -417 -200
rect -351 -222 -321 -200
rect -561 -272 -545 -238
rect -511 -272 -495 -238
rect -561 -288 -495 -272
rect -369 -238 -303 -222
rect -255 -226 -225 -200
rect -159 -222 -129 -200
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -369 -288 -303 -272
rect -177 -238 -111 -222
rect -63 -226 -33 -200
rect 33 -222 63 -200
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect -177 -288 -111 -272
rect 15 -238 81 -222
rect 129 -226 159 -200
rect 225 -222 255 -200
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 15 -288 81 -272
rect 207 -238 273 -222
rect 321 -226 351 -200
rect 417 -222 447 -200
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 207 -288 273 -272
rect 399 -238 465 -222
rect 513 -226 543 -200
rect 609 -222 639 -200
rect 399 -272 415 -238
rect 449 -272 465 -238
rect 399 -288 465 -272
rect 591 -238 657 -222
rect 705 -226 735 -200
rect 801 -222 831 -200
rect 591 -272 607 -238
rect 641 -272 657 -238
rect 591 -288 657 -272
rect 783 -238 849 -222
rect 897 -226 927 -200
rect 783 -272 799 -238
rect 833 -272 849 -238
rect 783 -288 849 -272
rect -945 -346 -879 -330
rect -945 -380 -929 -346
rect -895 -380 -879 -346
rect -945 -396 -879 -380
rect -753 -346 -687 -330
rect -753 -380 -737 -346
rect -703 -380 -687 -346
rect -927 -418 -897 -396
rect -831 -418 -801 -392
rect -753 -396 -687 -380
rect -561 -346 -495 -330
rect -561 -380 -545 -346
rect -511 -380 -495 -346
rect -735 -418 -705 -396
rect -639 -418 -609 -392
rect -561 -396 -495 -380
rect -369 -346 -303 -330
rect -369 -380 -353 -346
rect -319 -380 -303 -346
rect -543 -418 -513 -396
rect -447 -418 -417 -392
rect -369 -396 -303 -380
rect -177 -346 -111 -330
rect -177 -380 -161 -346
rect -127 -380 -111 -346
rect -351 -418 -321 -396
rect -255 -418 -225 -392
rect -177 -396 -111 -380
rect 15 -346 81 -330
rect 15 -380 31 -346
rect 65 -380 81 -346
rect -159 -418 -129 -396
rect -63 -418 -33 -392
rect 15 -396 81 -380
rect 207 -346 273 -330
rect 207 -380 223 -346
rect 257 -380 273 -346
rect 33 -418 63 -396
rect 129 -418 159 -392
rect 207 -396 273 -380
rect 399 -346 465 -330
rect 399 -380 415 -346
rect 449 -380 465 -346
rect 225 -418 255 -396
rect 321 -418 351 -392
rect 399 -396 465 -380
rect 591 -346 657 -330
rect 591 -380 607 -346
rect 641 -380 657 -346
rect 417 -418 447 -396
rect 513 -418 543 -392
rect 591 -396 657 -380
rect 783 -346 849 -330
rect 783 -380 799 -346
rect 833 -380 849 -346
rect 609 -418 639 -396
rect 705 -418 735 -392
rect 783 -396 849 -380
rect 801 -418 831 -396
rect 897 -418 927 -392
rect -927 -844 -897 -818
rect -831 -840 -801 -818
rect -849 -856 -783 -840
rect -735 -844 -705 -818
rect -639 -840 -609 -818
rect -849 -890 -833 -856
rect -799 -890 -783 -856
rect -849 -906 -783 -890
rect -657 -856 -591 -840
rect -543 -844 -513 -818
rect -447 -840 -417 -818
rect -657 -890 -641 -856
rect -607 -890 -591 -856
rect -657 -906 -591 -890
rect -465 -856 -399 -840
rect -351 -844 -321 -818
rect -255 -840 -225 -818
rect -465 -890 -449 -856
rect -415 -890 -399 -856
rect -465 -906 -399 -890
rect -273 -856 -207 -840
rect -159 -844 -129 -818
rect -63 -840 -33 -818
rect -273 -890 -257 -856
rect -223 -890 -207 -856
rect -273 -906 -207 -890
rect -81 -856 -15 -840
rect 33 -844 63 -818
rect 129 -840 159 -818
rect -81 -890 -65 -856
rect -31 -890 -15 -856
rect -81 -906 -15 -890
rect 111 -856 177 -840
rect 225 -844 255 -818
rect 321 -840 351 -818
rect 111 -890 127 -856
rect 161 -890 177 -856
rect 111 -906 177 -890
rect 303 -856 369 -840
rect 417 -844 447 -818
rect 513 -840 543 -818
rect 303 -890 319 -856
rect 353 -890 369 -856
rect 303 -906 369 -890
rect 495 -856 561 -840
rect 609 -844 639 -818
rect 705 -840 735 -818
rect 495 -890 511 -856
rect 545 -890 561 -856
rect 495 -906 561 -890
rect 687 -856 753 -840
rect 801 -844 831 -818
rect 897 -840 927 -818
rect 687 -890 703 -856
rect 737 -890 753 -856
rect 687 -906 753 -890
rect 879 -856 945 -840
rect 879 -890 895 -856
rect 929 -890 945 -856
rect 879 -906 945 -890
rect -849 -964 -783 -948
rect -849 -998 -833 -964
rect -799 -998 -783 -964
rect -927 -1036 -897 -1010
rect -849 -1014 -783 -998
rect -657 -964 -591 -948
rect -657 -998 -641 -964
rect -607 -998 -591 -964
rect -831 -1036 -801 -1014
rect -735 -1036 -705 -1010
rect -657 -1014 -591 -998
rect -465 -964 -399 -948
rect -465 -998 -449 -964
rect -415 -998 -399 -964
rect -639 -1036 -609 -1014
rect -543 -1036 -513 -1010
rect -465 -1014 -399 -998
rect -273 -964 -207 -948
rect -273 -998 -257 -964
rect -223 -998 -207 -964
rect -447 -1036 -417 -1014
rect -351 -1036 -321 -1010
rect -273 -1014 -207 -998
rect -81 -964 -15 -948
rect -81 -998 -65 -964
rect -31 -998 -15 -964
rect -255 -1036 -225 -1014
rect -159 -1036 -129 -1010
rect -81 -1014 -15 -998
rect 111 -964 177 -948
rect 111 -998 127 -964
rect 161 -998 177 -964
rect -63 -1036 -33 -1014
rect 33 -1036 63 -1010
rect 111 -1014 177 -998
rect 303 -964 369 -948
rect 303 -998 319 -964
rect 353 -998 369 -964
rect 129 -1036 159 -1014
rect 225 -1036 255 -1010
rect 303 -1014 369 -998
rect 495 -964 561 -948
rect 495 -998 511 -964
rect 545 -998 561 -964
rect 321 -1036 351 -1014
rect 417 -1036 447 -1010
rect 495 -1014 561 -998
rect 687 -964 753 -948
rect 687 -998 703 -964
rect 737 -998 753 -964
rect 513 -1036 543 -1014
rect 609 -1036 639 -1010
rect 687 -1014 753 -998
rect 879 -964 945 -948
rect 879 -998 895 -964
rect 929 -998 945 -964
rect 705 -1036 735 -1014
rect 801 -1036 831 -1010
rect 879 -1014 945 -998
rect 897 -1036 927 -1014
rect -927 -1458 -897 -1436
rect -945 -1474 -879 -1458
rect -831 -1462 -801 -1436
rect -735 -1458 -705 -1436
rect -945 -1508 -929 -1474
rect -895 -1508 -879 -1474
rect -945 -1524 -879 -1508
rect -753 -1474 -687 -1458
rect -639 -1462 -609 -1436
rect -543 -1458 -513 -1436
rect -753 -1508 -737 -1474
rect -703 -1508 -687 -1474
rect -753 -1524 -687 -1508
rect -561 -1474 -495 -1458
rect -447 -1462 -417 -1436
rect -351 -1458 -321 -1436
rect -561 -1508 -545 -1474
rect -511 -1508 -495 -1474
rect -561 -1524 -495 -1508
rect -369 -1474 -303 -1458
rect -255 -1462 -225 -1436
rect -159 -1458 -129 -1436
rect -369 -1508 -353 -1474
rect -319 -1508 -303 -1474
rect -369 -1524 -303 -1508
rect -177 -1474 -111 -1458
rect -63 -1462 -33 -1436
rect 33 -1458 63 -1436
rect -177 -1508 -161 -1474
rect -127 -1508 -111 -1474
rect -177 -1524 -111 -1508
rect 15 -1474 81 -1458
rect 129 -1462 159 -1436
rect 225 -1458 255 -1436
rect 15 -1508 31 -1474
rect 65 -1508 81 -1474
rect 15 -1524 81 -1508
rect 207 -1474 273 -1458
rect 321 -1462 351 -1436
rect 417 -1458 447 -1436
rect 207 -1508 223 -1474
rect 257 -1508 273 -1474
rect 207 -1524 273 -1508
rect 399 -1474 465 -1458
rect 513 -1462 543 -1436
rect 609 -1458 639 -1436
rect 399 -1508 415 -1474
rect 449 -1508 465 -1474
rect 399 -1524 465 -1508
rect 591 -1474 657 -1458
rect 705 -1462 735 -1436
rect 801 -1458 831 -1436
rect 591 -1508 607 -1474
rect 641 -1508 657 -1474
rect 591 -1524 657 -1508
rect 783 -1474 849 -1458
rect 897 -1462 927 -1436
rect 783 -1508 799 -1474
rect 833 -1508 849 -1474
rect 783 -1524 849 -1508
rect -945 -1582 -879 -1566
rect -945 -1616 -929 -1582
rect -895 -1616 -879 -1582
rect -945 -1632 -879 -1616
rect -753 -1582 -687 -1566
rect -753 -1616 -737 -1582
rect -703 -1616 -687 -1582
rect -927 -1654 -897 -1632
rect -831 -1654 -801 -1628
rect -753 -1632 -687 -1616
rect -561 -1582 -495 -1566
rect -561 -1616 -545 -1582
rect -511 -1616 -495 -1582
rect -735 -1654 -705 -1632
rect -639 -1654 -609 -1628
rect -561 -1632 -495 -1616
rect -369 -1582 -303 -1566
rect -369 -1616 -353 -1582
rect -319 -1616 -303 -1582
rect -543 -1654 -513 -1632
rect -447 -1654 -417 -1628
rect -369 -1632 -303 -1616
rect -177 -1582 -111 -1566
rect -177 -1616 -161 -1582
rect -127 -1616 -111 -1582
rect -351 -1654 -321 -1632
rect -255 -1654 -225 -1628
rect -177 -1632 -111 -1616
rect 15 -1582 81 -1566
rect 15 -1616 31 -1582
rect 65 -1616 81 -1582
rect -159 -1654 -129 -1632
rect -63 -1654 -33 -1628
rect 15 -1632 81 -1616
rect 207 -1582 273 -1566
rect 207 -1616 223 -1582
rect 257 -1616 273 -1582
rect 33 -1654 63 -1632
rect 129 -1654 159 -1628
rect 207 -1632 273 -1616
rect 399 -1582 465 -1566
rect 399 -1616 415 -1582
rect 449 -1616 465 -1582
rect 225 -1654 255 -1632
rect 321 -1654 351 -1628
rect 399 -1632 465 -1616
rect 591 -1582 657 -1566
rect 591 -1616 607 -1582
rect 641 -1616 657 -1582
rect 417 -1654 447 -1632
rect 513 -1654 543 -1628
rect 591 -1632 657 -1616
rect 783 -1582 849 -1566
rect 783 -1616 799 -1582
rect 833 -1616 849 -1582
rect 609 -1654 639 -1632
rect 705 -1654 735 -1628
rect 783 -1632 849 -1616
rect 801 -1654 831 -1632
rect 897 -1654 927 -1628
rect -927 -2080 -897 -2054
rect -831 -2076 -801 -2054
rect -849 -2092 -783 -2076
rect -735 -2080 -705 -2054
rect -639 -2076 -609 -2054
rect -849 -2126 -833 -2092
rect -799 -2126 -783 -2092
rect -849 -2142 -783 -2126
rect -657 -2092 -591 -2076
rect -543 -2080 -513 -2054
rect -447 -2076 -417 -2054
rect -657 -2126 -641 -2092
rect -607 -2126 -591 -2092
rect -657 -2142 -591 -2126
rect -465 -2092 -399 -2076
rect -351 -2080 -321 -2054
rect -255 -2076 -225 -2054
rect -465 -2126 -449 -2092
rect -415 -2126 -399 -2092
rect -465 -2142 -399 -2126
rect -273 -2092 -207 -2076
rect -159 -2080 -129 -2054
rect -63 -2076 -33 -2054
rect -273 -2126 -257 -2092
rect -223 -2126 -207 -2092
rect -273 -2142 -207 -2126
rect -81 -2092 -15 -2076
rect 33 -2080 63 -2054
rect 129 -2076 159 -2054
rect -81 -2126 -65 -2092
rect -31 -2126 -15 -2092
rect -81 -2142 -15 -2126
rect 111 -2092 177 -2076
rect 225 -2080 255 -2054
rect 321 -2076 351 -2054
rect 111 -2126 127 -2092
rect 161 -2126 177 -2092
rect 111 -2142 177 -2126
rect 303 -2092 369 -2076
rect 417 -2080 447 -2054
rect 513 -2076 543 -2054
rect 303 -2126 319 -2092
rect 353 -2126 369 -2092
rect 303 -2142 369 -2126
rect 495 -2092 561 -2076
rect 609 -2080 639 -2054
rect 705 -2076 735 -2054
rect 495 -2126 511 -2092
rect 545 -2126 561 -2092
rect 495 -2142 561 -2126
rect 687 -2092 753 -2076
rect 801 -2080 831 -2054
rect 897 -2076 927 -2054
rect 687 -2126 703 -2092
rect 737 -2126 753 -2092
rect 687 -2142 753 -2126
rect 879 -2092 945 -2076
rect 879 -2126 895 -2092
rect 929 -2126 945 -2092
rect 879 -2142 945 -2126
rect -849 -2200 -783 -2184
rect -849 -2234 -833 -2200
rect -799 -2234 -783 -2200
rect -927 -2272 -897 -2246
rect -849 -2250 -783 -2234
rect -657 -2200 -591 -2184
rect -657 -2234 -641 -2200
rect -607 -2234 -591 -2200
rect -831 -2272 -801 -2250
rect -735 -2272 -705 -2246
rect -657 -2250 -591 -2234
rect -465 -2200 -399 -2184
rect -465 -2234 -449 -2200
rect -415 -2234 -399 -2200
rect -639 -2272 -609 -2250
rect -543 -2272 -513 -2246
rect -465 -2250 -399 -2234
rect -273 -2200 -207 -2184
rect -273 -2234 -257 -2200
rect -223 -2234 -207 -2200
rect -447 -2272 -417 -2250
rect -351 -2272 -321 -2246
rect -273 -2250 -207 -2234
rect -81 -2200 -15 -2184
rect -81 -2234 -65 -2200
rect -31 -2234 -15 -2200
rect -255 -2272 -225 -2250
rect -159 -2272 -129 -2246
rect -81 -2250 -15 -2234
rect 111 -2200 177 -2184
rect 111 -2234 127 -2200
rect 161 -2234 177 -2200
rect -63 -2272 -33 -2250
rect 33 -2272 63 -2246
rect 111 -2250 177 -2234
rect 303 -2200 369 -2184
rect 303 -2234 319 -2200
rect 353 -2234 369 -2200
rect 129 -2272 159 -2250
rect 225 -2272 255 -2246
rect 303 -2250 369 -2234
rect 495 -2200 561 -2184
rect 495 -2234 511 -2200
rect 545 -2234 561 -2200
rect 321 -2272 351 -2250
rect 417 -2272 447 -2246
rect 495 -2250 561 -2234
rect 687 -2200 753 -2184
rect 687 -2234 703 -2200
rect 737 -2234 753 -2200
rect 513 -2272 543 -2250
rect 609 -2272 639 -2246
rect 687 -2250 753 -2234
rect 879 -2200 945 -2184
rect 879 -2234 895 -2200
rect 929 -2234 945 -2200
rect 705 -2272 735 -2250
rect 801 -2272 831 -2246
rect 879 -2250 945 -2234
rect 897 -2272 927 -2250
rect -927 -2694 -897 -2672
rect -945 -2710 -879 -2694
rect -831 -2698 -801 -2672
rect -735 -2694 -705 -2672
rect -945 -2744 -929 -2710
rect -895 -2744 -879 -2710
rect -945 -2760 -879 -2744
rect -753 -2710 -687 -2694
rect -639 -2698 -609 -2672
rect -543 -2694 -513 -2672
rect -753 -2744 -737 -2710
rect -703 -2744 -687 -2710
rect -753 -2760 -687 -2744
rect -561 -2710 -495 -2694
rect -447 -2698 -417 -2672
rect -351 -2694 -321 -2672
rect -561 -2744 -545 -2710
rect -511 -2744 -495 -2710
rect -561 -2760 -495 -2744
rect -369 -2710 -303 -2694
rect -255 -2698 -225 -2672
rect -159 -2694 -129 -2672
rect -369 -2744 -353 -2710
rect -319 -2744 -303 -2710
rect -369 -2760 -303 -2744
rect -177 -2710 -111 -2694
rect -63 -2698 -33 -2672
rect 33 -2694 63 -2672
rect -177 -2744 -161 -2710
rect -127 -2744 -111 -2710
rect -177 -2760 -111 -2744
rect 15 -2710 81 -2694
rect 129 -2698 159 -2672
rect 225 -2694 255 -2672
rect 15 -2744 31 -2710
rect 65 -2744 81 -2710
rect 15 -2760 81 -2744
rect 207 -2710 273 -2694
rect 321 -2698 351 -2672
rect 417 -2694 447 -2672
rect 207 -2744 223 -2710
rect 257 -2744 273 -2710
rect 207 -2760 273 -2744
rect 399 -2710 465 -2694
rect 513 -2698 543 -2672
rect 609 -2694 639 -2672
rect 399 -2744 415 -2710
rect 449 -2744 465 -2710
rect 399 -2760 465 -2744
rect 591 -2710 657 -2694
rect 705 -2698 735 -2672
rect 801 -2694 831 -2672
rect 591 -2744 607 -2710
rect 641 -2744 657 -2710
rect 591 -2760 657 -2744
rect 783 -2710 849 -2694
rect 897 -2698 927 -2672
rect 783 -2744 799 -2710
rect 833 -2744 849 -2710
rect 783 -2760 849 -2744
<< polycont >>
rect -833 2710 -799 2744
rect -641 2710 -607 2744
rect -449 2710 -415 2744
rect -257 2710 -223 2744
rect -65 2710 -31 2744
rect 127 2710 161 2744
rect 319 2710 353 2744
rect 511 2710 545 2744
rect 703 2710 737 2744
rect 895 2710 929 2744
rect -929 2200 -895 2234
rect -737 2200 -703 2234
rect -545 2200 -511 2234
rect -353 2200 -319 2234
rect -161 2200 -127 2234
rect 31 2200 65 2234
rect 223 2200 257 2234
rect 415 2200 449 2234
rect 607 2200 641 2234
rect 799 2200 833 2234
rect -929 2092 -895 2126
rect -737 2092 -703 2126
rect -545 2092 -511 2126
rect -353 2092 -319 2126
rect -161 2092 -127 2126
rect 31 2092 65 2126
rect 223 2092 257 2126
rect 415 2092 449 2126
rect 607 2092 641 2126
rect 799 2092 833 2126
rect -833 1582 -799 1616
rect -641 1582 -607 1616
rect -449 1582 -415 1616
rect -257 1582 -223 1616
rect -65 1582 -31 1616
rect 127 1582 161 1616
rect 319 1582 353 1616
rect 511 1582 545 1616
rect 703 1582 737 1616
rect 895 1582 929 1616
rect -833 1474 -799 1508
rect -641 1474 -607 1508
rect -449 1474 -415 1508
rect -257 1474 -223 1508
rect -65 1474 -31 1508
rect 127 1474 161 1508
rect 319 1474 353 1508
rect 511 1474 545 1508
rect 703 1474 737 1508
rect 895 1474 929 1508
rect -929 964 -895 998
rect -737 964 -703 998
rect -545 964 -511 998
rect -353 964 -319 998
rect -161 964 -127 998
rect 31 964 65 998
rect 223 964 257 998
rect 415 964 449 998
rect 607 964 641 998
rect 799 964 833 998
rect -929 856 -895 890
rect -737 856 -703 890
rect -545 856 -511 890
rect -353 856 -319 890
rect -161 856 -127 890
rect 31 856 65 890
rect 223 856 257 890
rect 415 856 449 890
rect 607 856 641 890
rect 799 856 833 890
rect -833 346 -799 380
rect -641 346 -607 380
rect -449 346 -415 380
rect -257 346 -223 380
rect -65 346 -31 380
rect 127 346 161 380
rect 319 346 353 380
rect 511 346 545 380
rect 703 346 737 380
rect 895 346 929 380
rect -833 238 -799 272
rect -641 238 -607 272
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect 511 238 545 272
rect 703 238 737 272
rect 895 238 929 272
rect -929 -272 -895 -238
rect -737 -272 -703 -238
rect -545 -272 -511 -238
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
rect 607 -272 641 -238
rect 799 -272 833 -238
rect -929 -380 -895 -346
rect -737 -380 -703 -346
rect -545 -380 -511 -346
rect -353 -380 -319 -346
rect -161 -380 -127 -346
rect 31 -380 65 -346
rect 223 -380 257 -346
rect 415 -380 449 -346
rect 607 -380 641 -346
rect 799 -380 833 -346
rect -833 -890 -799 -856
rect -641 -890 -607 -856
rect -449 -890 -415 -856
rect -257 -890 -223 -856
rect -65 -890 -31 -856
rect 127 -890 161 -856
rect 319 -890 353 -856
rect 511 -890 545 -856
rect 703 -890 737 -856
rect 895 -890 929 -856
rect -833 -998 -799 -964
rect -641 -998 -607 -964
rect -449 -998 -415 -964
rect -257 -998 -223 -964
rect -65 -998 -31 -964
rect 127 -998 161 -964
rect 319 -998 353 -964
rect 511 -998 545 -964
rect 703 -998 737 -964
rect 895 -998 929 -964
rect -929 -1508 -895 -1474
rect -737 -1508 -703 -1474
rect -545 -1508 -511 -1474
rect -353 -1508 -319 -1474
rect -161 -1508 -127 -1474
rect 31 -1508 65 -1474
rect 223 -1508 257 -1474
rect 415 -1508 449 -1474
rect 607 -1508 641 -1474
rect 799 -1508 833 -1474
rect -929 -1616 -895 -1582
rect -737 -1616 -703 -1582
rect -545 -1616 -511 -1582
rect -353 -1616 -319 -1582
rect -161 -1616 -127 -1582
rect 31 -1616 65 -1582
rect 223 -1616 257 -1582
rect 415 -1616 449 -1582
rect 607 -1616 641 -1582
rect 799 -1616 833 -1582
rect -833 -2126 -799 -2092
rect -641 -2126 -607 -2092
rect -449 -2126 -415 -2092
rect -257 -2126 -223 -2092
rect -65 -2126 -31 -2092
rect 127 -2126 161 -2092
rect 319 -2126 353 -2092
rect 511 -2126 545 -2092
rect 703 -2126 737 -2092
rect 895 -2126 929 -2092
rect -833 -2234 -799 -2200
rect -641 -2234 -607 -2200
rect -449 -2234 -415 -2200
rect -257 -2234 -223 -2200
rect -65 -2234 -31 -2200
rect 127 -2234 161 -2200
rect 319 -2234 353 -2200
rect 511 -2234 545 -2200
rect 703 -2234 737 -2200
rect 895 -2234 929 -2200
rect -929 -2744 -895 -2710
rect -737 -2744 -703 -2710
rect -545 -2744 -511 -2710
rect -353 -2744 -319 -2710
rect -161 -2744 -127 -2710
rect 31 -2744 65 -2710
rect 223 -2744 257 -2710
rect 415 -2744 449 -2710
rect 607 -2744 641 -2710
rect 799 -2744 833 -2710
<< locali >>
rect -1091 2812 -995 2846
rect 995 2812 1091 2846
rect -1091 2750 -1057 2812
rect 1057 2750 1091 2812
rect -849 2710 -833 2744
rect -799 2710 -783 2744
rect -657 2710 -641 2744
rect -607 2710 -591 2744
rect -465 2710 -449 2744
rect -415 2710 -399 2744
rect -273 2710 -257 2744
rect -223 2710 -207 2744
rect -81 2710 -65 2744
rect -31 2710 -15 2744
rect 111 2710 127 2744
rect 161 2710 177 2744
rect 303 2710 319 2744
rect 353 2710 369 2744
rect 495 2710 511 2744
rect 545 2710 561 2744
rect 687 2710 703 2744
rect 737 2710 753 2744
rect 879 2710 895 2744
rect 929 2710 945 2744
rect -977 2660 -943 2676
rect -977 2268 -943 2284
rect -881 2660 -847 2676
rect -881 2268 -847 2284
rect -785 2660 -751 2676
rect -785 2268 -751 2284
rect -689 2660 -655 2676
rect -689 2268 -655 2284
rect -593 2660 -559 2676
rect -593 2268 -559 2284
rect -497 2660 -463 2676
rect -497 2268 -463 2284
rect -401 2660 -367 2676
rect -401 2268 -367 2284
rect -305 2660 -271 2676
rect -305 2268 -271 2284
rect -209 2660 -175 2676
rect -209 2268 -175 2284
rect -113 2660 -79 2676
rect -113 2268 -79 2284
rect -17 2660 17 2676
rect -17 2268 17 2284
rect 79 2660 113 2676
rect 79 2268 113 2284
rect 175 2660 209 2676
rect 175 2268 209 2284
rect 271 2660 305 2676
rect 271 2268 305 2284
rect 367 2660 401 2676
rect 367 2268 401 2284
rect 463 2660 497 2676
rect 463 2268 497 2284
rect 559 2660 593 2676
rect 559 2268 593 2284
rect 655 2660 689 2676
rect 655 2268 689 2284
rect 751 2660 785 2676
rect 751 2268 785 2284
rect 847 2660 881 2676
rect 847 2268 881 2284
rect 943 2660 977 2676
rect 943 2268 977 2284
rect -945 2200 -929 2234
rect -895 2200 -879 2234
rect -753 2200 -737 2234
rect -703 2200 -687 2234
rect -561 2200 -545 2234
rect -511 2200 -495 2234
rect -369 2200 -353 2234
rect -319 2200 -303 2234
rect -177 2200 -161 2234
rect -127 2200 -111 2234
rect 15 2200 31 2234
rect 65 2200 81 2234
rect 207 2200 223 2234
rect 257 2200 273 2234
rect 399 2200 415 2234
rect 449 2200 465 2234
rect 591 2200 607 2234
rect 641 2200 657 2234
rect 783 2200 799 2234
rect 833 2200 849 2234
rect -945 2092 -929 2126
rect -895 2092 -879 2126
rect -753 2092 -737 2126
rect -703 2092 -687 2126
rect -561 2092 -545 2126
rect -511 2092 -495 2126
rect -369 2092 -353 2126
rect -319 2092 -303 2126
rect -177 2092 -161 2126
rect -127 2092 -111 2126
rect 15 2092 31 2126
rect 65 2092 81 2126
rect 207 2092 223 2126
rect 257 2092 273 2126
rect 399 2092 415 2126
rect 449 2092 465 2126
rect 591 2092 607 2126
rect 641 2092 657 2126
rect 783 2092 799 2126
rect 833 2092 849 2126
rect -977 2042 -943 2058
rect -977 1650 -943 1666
rect -881 2042 -847 2058
rect -881 1650 -847 1666
rect -785 2042 -751 2058
rect -785 1650 -751 1666
rect -689 2042 -655 2058
rect -689 1650 -655 1666
rect -593 2042 -559 2058
rect -593 1650 -559 1666
rect -497 2042 -463 2058
rect -497 1650 -463 1666
rect -401 2042 -367 2058
rect -401 1650 -367 1666
rect -305 2042 -271 2058
rect -305 1650 -271 1666
rect -209 2042 -175 2058
rect -209 1650 -175 1666
rect -113 2042 -79 2058
rect -113 1650 -79 1666
rect -17 2042 17 2058
rect -17 1650 17 1666
rect 79 2042 113 2058
rect 79 1650 113 1666
rect 175 2042 209 2058
rect 175 1650 209 1666
rect 271 2042 305 2058
rect 271 1650 305 1666
rect 367 2042 401 2058
rect 367 1650 401 1666
rect 463 2042 497 2058
rect 463 1650 497 1666
rect 559 2042 593 2058
rect 559 1650 593 1666
rect 655 2042 689 2058
rect 655 1650 689 1666
rect 751 2042 785 2058
rect 751 1650 785 1666
rect 847 2042 881 2058
rect 847 1650 881 1666
rect 943 2042 977 2058
rect 943 1650 977 1666
rect -849 1582 -833 1616
rect -799 1582 -783 1616
rect -657 1582 -641 1616
rect -607 1582 -591 1616
rect -465 1582 -449 1616
rect -415 1582 -399 1616
rect -273 1582 -257 1616
rect -223 1582 -207 1616
rect -81 1582 -65 1616
rect -31 1582 -15 1616
rect 111 1582 127 1616
rect 161 1582 177 1616
rect 303 1582 319 1616
rect 353 1582 369 1616
rect 495 1582 511 1616
rect 545 1582 561 1616
rect 687 1582 703 1616
rect 737 1582 753 1616
rect 879 1582 895 1616
rect 929 1582 945 1616
rect -849 1474 -833 1508
rect -799 1474 -783 1508
rect -657 1474 -641 1508
rect -607 1474 -591 1508
rect -465 1474 -449 1508
rect -415 1474 -399 1508
rect -273 1474 -257 1508
rect -223 1474 -207 1508
rect -81 1474 -65 1508
rect -31 1474 -15 1508
rect 111 1474 127 1508
rect 161 1474 177 1508
rect 303 1474 319 1508
rect 353 1474 369 1508
rect 495 1474 511 1508
rect 545 1474 561 1508
rect 687 1474 703 1508
rect 737 1474 753 1508
rect 879 1474 895 1508
rect 929 1474 945 1508
rect -977 1424 -943 1440
rect -977 1032 -943 1048
rect -881 1424 -847 1440
rect -881 1032 -847 1048
rect -785 1424 -751 1440
rect -785 1032 -751 1048
rect -689 1424 -655 1440
rect -689 1032 -655 1048
rect -593 1424 -559 1440
rect -593 1032 -559 1048
rect -497 1424 -463 1440
rect -497 1032 -463 1048
rect -401 1424 -367 1440
rect -401 1032 -367 1048
rect -305 1424 -271 1440
rect -305 1032 -271 1048
rect -209 1424 -175 1440
rect -209 1032 -175 1048
rect -113 1424 -79 1440
rect -113 1032 -79 1048
rect -17 1424 17 1440
rect -17 1032 17 1048
rect 79 1424 113 1440
rect 79 1032 113 1048
rect 175 1424 209 1440
rect 175 1032 209 1048
rect 271 1424 305 1440
rect 271 1032 305 1048
rect 367 1424 401 1440
rect 367 1032 401 1048
rect 463 1424 497 1440
rect 463 1032 497 1048
rect 559 1424 593 1440
rect 559 1032 593 1048
rect 655 1424 689 1440
rect 655 1032 689 1048
rect 751 1424 785 1440
rect 751 1032 785 1048
rect 847 1424 881 1440
rect 847 1032 881 1048
rect 943 1424 977 1440
rect 943 1032 977 1048
rect -945 964 -929 998
rect -895 964 -879 998
rect -753 964 -737 998
rect -703 964 -687 998
rect -561 964 -545 998
rect -511 964 -495 998
rect -369 964 -353 998
rect -319 964 -303 998
rect -177 964 -161 998
rect -127 964 -111 998
rect 15 964 31 998
rect 65 964 81 998
rect 207 964 223 998
rect 257 964 273 998
rect 399 964 415 998
rect 449 964 465 998
rect 591 964 607 998
rect 641 964 657 998
rect 783 964 799 998
rect 833 964 849 998
rect -945 856 -929 890
rect -895 856 -879 890
rect -753 856 -737 890
rect -703 856 -687 890
rect -561 856 -545 890
rect -511 856 -495 890
rect -369 856 -353 890
rect -319 856 -303 890
rect -177 856 -161 890
rect -127 856 -111 890
rect 15 856 31 890
rect 65 856 81 890
rect 207 856 223 890
rect 257 856 273 890
rect 399 856 415 890
rect 449 856 465 890
rect 591 856 607 890
rect 641 856 657 890
rect 783 856 799 890
rect 833 856 849 890
rect -977 806 -943 822
rect -977 414 -943 430
rect -881 806 -847 822
rect -881 414 -847 430
rect -785 806 -751 822
rect -785 414 -751 430
rect -689 806 -655 822
rect -689 414 -655 430
rect -593 806 -559 822
rect -593 414 -559 430
rect -497 806 -463 822
rect -497 414 -463 430
rect -401 806 -367 822
rect -401 414 -367 430
rect -305 806 -271 822
rect -305 414 -271 430
rect -209 806 -175 822
rect -209 414 -175 430
rect -113 806 -79 822
rect -113 414 -79 430
rect -17 806 17 822
rect -17 414 17 430
rect 79 806 113 822
rect 79 414 113 430
rect 175 806 209 822
rect 175 414 209 430
rect 271 806 305 822
rect 271 414 305 430
rect 367 806 401 822
rect 367 414 401 430
rect 463 806 497 822
rect 463 414 497 430
rect 559 806 593 822
rect 559 414 593 430
rect 655 806 689 822
rect 655 414 689 430
rect 751 806 785 822
rect 751 414 785 430
rect 847 806 881 822
rect 847 414 881 430
rect 943 806 977 822
rect 943 414 977 430
rect -849 346 -833 380
rect -799 346 -783 380
rect -657 346 -641 380
rect -607 346 -591 380
rect -465 346 -449 380
rect -415 346 -399 380
rect -273 346 -257 380
rect -223 346 -207 380
rect -81 346 -65 380
rect -31 346 -15 380
rect 111 346 127 380
rect 161 346 177 380
rect 303 346 319 380
rect 353 346 369 380
rect 495 346 511 380
rect 545 346 561 380
rect 687 346 703 380
rect 737 346 753 380
rect 879 346 895 380
rect 929 346 945 380
rect -849 238 -833 272
rect -799 238 -783 272
rect -657 238 -641 272
rect -607 238 -591 272
rect -465 238 -449 272
rect -415 238 -399 272
rect -273 238 -257 272
rect -223 238 -207 272
rect -81 238 -65 272
rect -31 238 -15 272
rect 111 238 127 272
rect 161 238 177 272
rect 303 238 319 272
rect 353 238 369 272
rect 495 238 511 272
rect 545 238 561 272
rect 687 238 703 272
rect 737 238 753 272
rect 879 238 895 272
rect 929 238 945 272
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect -945 -272 -929 -238
rect -895 -272 -879 -238
rect -753 -272 -737 -238
rect -703 -272 -687 -238
rect -561 -272 -545 -238
rect -511 -272 -495 -238
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 399 -272 415 -238
rect 449 -272 465 -238
rect 591 -272 607 -238
rect 641 -272 657 -238
rect 783 -272 799 -238
rect 833 -272 849 -238
rect -945 -380 -929 -346
rect -895 -380 -879 -346
rect -753 -380 -737 -346
rect -703 -380 -687 -346
rect -561 -380 -545 -346
rect -511 -380 -495 -346
rect -369 -380 -353 -346
rect -319 -380 -303 -346
rect -177 -380 -161 -346
rect -127 -380 -111 -346
rect 15 -380 31 -346
rect 65 -380 81 -346
rect 207 -380 223 -346
rect 257 -380 273 -346
rect 399 -380 415 -346
rect 449 -380 465 -346
rect 591 -380 607 -346
rect 641 -380 657 -346
rect 783 -380 799 -346
rect 833 -380 849 -346
rect -977 -430 -943 -414
rect -977 -822 -943 -806
rect -881 -430 -847 -414
rect -881 -822 -847 -806
rect -785 -430 -751 -414
rect -785 -822 -751 -806
rect -689 -430 -655 -414
rect -689 -822 -655 -806
rect -593 -430 -559 -414
rect -593 -822 -559 -806
rect -497 -430 -463 -414
rect -497 -822 -463 -806
rect -401 -430 -367 -414
rect -401 -822 -367 -806
rect -305 -430 -271 -414
rect -305 -822 -271 -806
rect -209 -430 -175 -414
rect -209 -822 -175 -806
rect -113 -430 -79 -414
rect -113 -822 -79 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 79 -430 113 -414
rect 79 -822 113 -806
rect 175 -430 209 -414
rect 175 -822 209 -806
rect 271 -430 305 -414
rect 271 -822 305 -806
rect 367 -430 401 -414
rect 367 -822 401 -806
rect 463 -430 497 -414
rect 463 -822 497 -806
rect 559 -430 593 -414
rect 559 -822 593 -806
rect 655 -430 689 -414
rect 655 -822 689 -806
rect 751 -430 785 -414
rect 751 -822 785 -806
rect 847 -430 881 -414
rect 847 -822 881 -806
rect 943 -430 977 -414
rect 943 -822 977 -806
rect -849 -890 -833 -856
rect -799 -890 -783 -856
rect -657 -890 -641 -856
rect -607 -890 -591 -856
rect -465 -890 -449 -856
rect -415 -890 -399 -856
rect -273 -890 -257 -856
rect -223 -890 -207 -856
rect -81 -890 -65 -856
rect -31 -890 -15 -856
rect 111 -890 127 -856
rect 161 -890 177 -856
rect 303 -890 319 -856
rect 353 -890 369 -856
rect 495 -890 511 -856
rect 545 -890 561 -856
rect 687 -890 703 -856
rect 737 -890 753 -856
rect 879 -890 895 -856
rect 929 -890 945 -856
rect -849 -998 -833 -964
rect -799 -998 -783 -964
rect -657 -998 -641 -964
rect -607 -998 -591 -964
rect -465 -998 -449 -964
rect -415 -998 -399 -964
rect -273 -998 -257 -964
rect -223 -998 -207 -964
rect -81 -998 -65 -964
rect -31 -998 -15 -964
rect 111 -998 127 -964
rect 161 -998 177 -964
rect 303 -998 319 -964
rect 353 -998 369 -964
rect 495 -998 511 -964
rect 545 -998 561 -964
rect 687 -998 703 -964
rect 737 -998 753 -964
rect 879 -998 895 -964
rect 929 -998 945 -964
rect -977 -1048 -943 -1032
rect -977 -1440 -943 -1424
rect -881 -1048 -847 -1032
rect -881 -1440 -847 -1424
rect -785 -1048 -751 -1032
rect -785 -1440 -751 -1424
rect -689 -1048 -655 -1032
rect -689 -1440 -655 -1424
rect -593 -1048 -559 -1032
rect -593 -1440 -559 -1424
rect -497 -1048 -463 -1032
rect -497 -1440 -463 -1424
rect -401 -1048 -367 -1032
rect -401 -1440 -367 -1424
rect -305 -1048 -271 -1032
rect -305 -1440 -271 -1424
rect -209 -1048 -175 -1032
rect -209 -1440 -175 -1424
rect -113 -1048 -79 -1032
rect -113 -1440 -79 -1424
rect -17 -1048 17 -1032
rect -17 -1440 17 -1424
rect 79 -1048 113 -1032
rect 79 -1440 113 -1424
rect 175 -1048 209 -1032
rect 175 -1440 209 -1424
rect 271 -1048 305 -1032
rect 271 -1440 305 -1424
rect 367 -1048 401 -1032
rect 367 -1440 401 -1424
rect 463 -1048 497 -1032
rect 463 -1440 497 -1424
rect 559 -1048 593 -1032
rect 559 -1440 593 -1424
rect 655 -1048 689 -1032
rect 655 -1440 689 -1424
rect 751 -1048 785 -1032
rect 751 -1440 785 -1424
rect 847 -1048 881 -1032
rect 847 -1440 881 -1424
rect 943 -1048 977 -1032
rect 943 -1440 977 -1424
rect -945 -1508 -929 -1474
rect -895 -1508 -879 -1474
rect -753 -1508 -737 -1474
rect -703 -1508 -687 -1474
rect -561 -1508 -545 -1474
rect -511 -1508 -495 -1474
rect -369 -1508 -353 -1474
rect -319 -1508 -303 -1474
rect -177 -1508 -161 -1474
rect -127 -1508 -111 -1474
rect 15 -1508 31 -1474
rect 65 -1508 81 -1474
rect 207 -1508 223 -1474
rect 257 -1508 273 -1474
rect 399 -1508 415 -1474
rect 449 -1508 465 -1474
rect 591 -1508 607 -1474
rect 641 -1508 657 -1474
rect 783 -1508 799 -1474
rect 833 -1508 849 -1474
rect -945 -1616 -929 -1582
rect -895 -1616 -879 -1582
rect -753 -1616 -737 -1582
rect -703 -1616 -687 -1582
rect -561 -1616 -545 -1582
rect -511 -1616 -495 -1582
rect -369 -1616 -353 -1582
rect -319 -1616 -303 -1582
rect -177 -1616 -161 -1582
rect -127 -1616 -111 -1582
rect 15 -1616 31 -1582
rect 65 -1616 81 -1582
rect 207 -1616 223 -1582
rect 257 -1616 273 -1582
rect 399 -1616 415 -1582
rect 449 -1616 465 -1582
rect 591 -1616 607 -1582
rect 641 -1616 657 -1582
rect 783 -1616 799 -1582
rect 833 -1616 849 -1582
rect -977 -1666 -943 -1650
rect -977 -2058 -943 -2042
rect -881 -1666 -847 -1650
rect -881 -2058 -847 -2042
rect -785 -1666 -751 -1650
rect -785 -2058 -751 -2042
rect -689 -1666 -655 -1650
rect -689 -2058 -655 -2042
rect -593 -1666 -559 -1650
rect -593 -2058 -559 -2042
rect -497 -1666 -463 -1650
rect -497 -2058 -463 -2042
rect -401 -1666 -367 -1650
rect -401 -2058 -367 -2042
rect -305 -1666 -271 -1650
rect -305 -2058 -271 -2042
rect -209 -1666 -175 -1650
rect -209 -2058 -175 -2042
rect -113 -1666 -79 -1650
rect -113 -2058 -79 -2042
rect -17 -1666 17 -1650
rect -17 -2058 17 -2042
rect 79 -1666 113 -1650
rect 79 -2058 113 -2042
rect 175 -1666 209 -1650
rect 175 -2058 209 -2042
rect 271 -1666 305 -1650
rect 271 -2058 305 -2042
rect 367 -1666 401 -1650
rect 367 -2058 401 -2042
rect 463 -1666 497 -1650
rect 463 -2058 497 -2042
rect 559 -1666 593 -1650
rect 559 -2058 593 -2042
rect 655 -1666 689 -1650
rect 655 -2058 689 -2042
rect 751 -1666 785 -1650
rect 751 -2058 785 -2042
rect 847 -1666 881 -1650
rect 847 -2058 881 -2042
rect 943 -1666 977 -1650
rect 943 -2058 977 -2042
rect -849 -2126 -833 -2092
rect -799 -2126 -783 -2092
rect -657 -2126 -641 -2092
rect -607 -2126 -591 -2092
rect -465 -2126 -449 -2092
rect -415 -2126 -399 -2092
rect -273 -2126 -257 -2092
rect -223 -2126 -207 -2092
rect -81 -2126 -65 -2092
rect -31 -2126 -15 -2092
rect 111 -2126 127 -2092
rect 161 -2126 177 -2092
rect 303 -2126 319 -2092
rect 353 -2126 369 -2092
rect 495 -2126 511 -2092
rect 545 -2126 561 -2092
rect 687 -2126 703 -2092
rect 737 -2126 753 -2092
rect 879 -2126 895 -2092
rect 929 -2126 945 -2092
rect -849 -2234 -833 -2200
rect -799 -2234 -783 -2200
rect -657 -2234 -641 -2200
rect -607 -2234 -591 -2200
rect -465 -2234 -449 -2200
rect -415 -2234 -399 -2200
rect -273 -2234 -257 -2200
rect -223 -2234 -207 -2200
rect -81 -2234 -65 -2200
rect -31 -2234 -15 -2200
rect 111 -2234 127 -2200
rect 161 -2234 177 -2200
rect 303 -2234 319 -2200
rect 353 -2234 369 -2200
rect 495 -2234 511 -2200
rect 545 -2234 561 -2200
rect 687 -2234 703 -2200
rect 737 -2234 753 -2200
rect 879 -2234 895 -2200
rect 929 -2234 945 -2200
rect -977 -2284 -943 -2268
rect -977 -2676 -943 -2660
rect -881 -2284 -847 -2268
rect -881 -2676 -847 -2660
rect -785 -2284 -751 -2268
rect -785 -2676 -751 -2660
rect -689 -2284 -655 -2268
rect -689 -2676 -655 -2660
rect -593 -2284 -559 -2268
rect -593 -2676 -559 -2660
rect -497 -2284 -463 -2268
rect -497 -2676 -463 -2660
rect -401 -2284 -367 -2268
rect -401 -2676 -367 -2660
rect -305 -2284 -271 -2268
rect -305 -2676 -271 -2660
rect -209 -2284 -175 -2268
rect -209 -2676 -175 -2660
rect -113 -2284 -79 -2268
rect -113 -2676 -79 -2660
rect -17 -2284 17 -2268
rect -17 -2676 17 -2660
rect 79 -2284 113 -2268
rect 79 -2676 113 -2660
rect 175 -2284 209 -2268
rect 175 -2676 209 -2660
rect 271 -2284 305 -2268
rect 271 -2676 305 -2660
rect 367 -2284 401 -2268
rect 367 -2676 401 -2660
rect 463 -2284 497 -2268
rect 463 -2676 497 -2660
rect 559 -2284 593 -2268
rect 559 -2676 593 -2660
rect 655 -2284 689 -2268
rect 655 -2676 689 -2660
rect 751 -2284 785 -2268
rect 751 -2676 785 -2660
rect 847 -2284 881 -2268
rect 847 -2676 881 -2660
rect 943 -2284 977 -2268
rect 943 -2676 977 -2660
rect -945 -2744 -929 -2710
rect -895 -2744 -879 -2710
rect -753 -2744 -737 -2710
rect -703 -2744 -687 -2710
rect -561 -2744 -545 -2710
rect -511 -2744 -495 -2710
rect -369 -2744 -353 -2710
rect -319 -2744 -303 -2710
rect -177 -2744 -161 -2710
rect -127 -2744 -111 -2710
rect 15 -2744 31 -2710
rect 65 -2744 81 -2710
rect 207 -2744 223 -2710
rect 257 -2744 273 -2710
rect 399 -2744 415 -2710
rect 449 -2744 465 -2710
rect 591 -2744 607 -2710
rect 641 -2744 657 -2710
rect 783 -2744 799 -2710
rect 833 -2744 849 -2710
rect -1091 -2812 -1057 -2750
rect 1057 -2812 1091 -2750
rect -1091 -2846 -995 -2812
rect 995 -2846 1091 -2812
<< viali >>
rect -833 2710 -799 2744
rect -641 2710 -607 2744
rect -449 2710 -415 2744
rect -257 2710 -223 2744
rect -65 2710 -31 2744
rect 127 2710 161 2744
rect 319 2710 353 2744
rect 511 2710 545 2744
rect 703 2710 737 2744
rect 895 2710 929 2744
rect -977 2284 -943 2660
rect -881 2284 -847 2660
rect -785 2284 -751 2660
rect -689 2284 -655 2660
rect -593 2284 -559 2660
rect -497 2284 -463 2660
rect -401 2284 -367 2660
rect -305 2284 -271 2660
rect -209 2284 -175 2660
rect -113 2284 -79 2660
rect -17 2284 17 2660
rect 79 2284 113 2660
rect 175 2284 209 2660
rect 271 2284 305 2660
rect 367 2284 401 2660
rect 463 2284 497 2660
rect 559 2284 593 2660
rect 655 2284 689 2660
rect 751 2284 785 2660
rect 847 2284 881 2660
rect 943 2284 977 2660
rect -929 2200 -895 2234
rect -737 2200 -703 2234
rect -545 2200 -511 2234
rect -353 2200 -319 2234
rect -161 2200 -127 2234
rect 31 2200 65 2234
rect 223 2200 257 2234
rect 415 2200 449 2234
rect 607 2200 641 2234
rect 799 2200 833 2234
rect -929 2092 -895 2126
rect -737 2092 -703 2126
rect -545 2092 -511 2126
rect -353 2092 -319 2126
rect -161 2092 -127 2126
rect 31 2092 65 2126
rect 223 2092 257 2126
rect 415 2092 449 2126
rect 607 2092 641 2126
rect 799 2092 833 2126
rect -977 1666 -943 2042
rect -881 1666 -847 2042
rect -785 1666 -751 2042
rect -689 1666 -655 2042
rect -593 1666 -559 2042
rect -497 1666 -463 2042
rect -401 1666 -367 2042
rect -305 1666 -271 2042
rect -209 1666 -175 2042
rect -113 1666 -79 2042
rect -17 1666 17 2042
rect 79 1666 113 2042
rect 175 1666 209 2042
rect 271 1666 305 2042
rect 367 1666 401 2042
rect 463 1666 497 2042
rect 559 1666 593 2042
rect 655 1666 689 2042
rect 751 1666 785 2042
rect 847 1666 881 2042
rect 943 1666 977 2042
rect -833 1582 -799 1616
rect -641 1582 -607 1616
rect -449 1582 -415 1616
rect -257 1582 -223 1616
rect -65 1582 -31 1616
rect 127 1582 161 1616
rect 319 1582 353 1616
rect 511 1582 545 1616
rect 703 1582 737 1616
rect 895 1582 929 1616
rect -833 1474 -799 1508
rect -641 1474 -607 1508
rect -449 1474 -415 1508
rect -257 1474 -223 1508
rect -65 1474 -31 1508
rect 127 1474 161 1508
rect 319 1474 353 1508
rect 511 1474 545 1508
rect 703 1474 737 1508
rect 895 1474 929 1508
rect -977 1048 -943 1424
rect -881 1048 -847 1424
rect -785 1048 -751 1424
rect -689 1048 -655 1424
rect -593 1048 -559 1424
rect -497 1048 -463 1424
rect -401 1048 -367 1424
rect -305 1048 -271 1424
rect -209 1048 -175 1424
rect -113 1048 -79 1424
rect -17 1048 17 1424
rect 79 1048 113 1424
rect 175 1048 209 1424
rect 271 1048 305 1424
rect 367 1048 401 1424
rect 463 1048 497 1424
rect 559 1048 593 1424
rect 655 1048 689 1424
rect 751 1048 785 1424
rect 847 1048 881 1424
rect 943 1048 977 1424
rect -929 964 -895 998
rect -737 964 -703 998
rect -545 964 -511 998
rect -353 964 -319 998
rect -161 964 -127 998
rect 31 964 65 998
rect 223 964 257 998
rect 415 964 449 998
rect 607 964 641 998
rect 799 964 833 998
rect -929 856 -895 890
rect -737 856 -703 890
rect -545 856 -511 890
rect -353 856 -319 890
rect -161 856 -127 890
rect 31 856 65 890
rect 223 856 257 890
rect 415 856 449 890
rect 607 856 641 890
rect 799 856 833 890
rect -977 430 -943 806
rect -881 430 -847 806
rect -785 430 -751 806
rect -689 430 -655 806
rect -593 430 -559 806
rect -497 430 -463 806
rect -401 430 -367 806
rect -305 430 -271 806
rect -209 430 -175 806
rect -113 430 -79 806
rect -17 430 17 806
rect 79 430 113 806
rect 175 430 209 806
rect 271 430 305 806
rect 367 430 401 806
rect 463 430 497 806
rect 559 430 593 806
rect 655 430 689 806
rect 751 430 785 806
rect 847 430 881 806
rect 943 430 977 806
rect -833 346 -799 380
rect -641 346 -607 380
rect -449 346 -415 380
rect -257 346 -223 380
rect -65 346 -31 380
rect 127 346 161 380
rect 319 346 353 380
rect 511 346 545 380
rect 703 346 737 380
rect 895 346 929 380
rect -833 238 -799 272
rect -641 238 -607 272
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect 511 238 545 272
rect 703 238 737 272
rect 895 238 929 272
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect -929 -272 -895 -238
rect -737 -272 -703 -238
rect -545 -272 -511 -238
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
rect 607 -272 641 -238
rect 799 -272 833 -238
rect -929 -380 -895 -346
rect -737 -380 -703 -346
rect -545 -380 -511 -346
rect -353 -380 -319 -346
rect -161 -380 -127 -346
rect 31 -380 65 -346
rect 223 -380 257 -346
rect 415 -380 449 -346
rect 607 -380 641 -346
rect 799 -380 833 -346
rect -977 -806 -943 -430
rect -881 -806 -847 -430
rect -785 -806 -751 -430
rect -689 -806 -655 -430
rect -593 -806 -559 -430
rect -497 -806 -463 -430
rect -401 -806 -367 -430
rect -305 -806 -271 -430
rect -209 -806 -175 -430
rect -113 -806 -79 -430
rect -17 -806 17 -430
rect 79 -806 113 -430
rect 175 -806 209 -430
rect 271 -806 305 -430
rect 367 -806 401 -430
rect 463 -806 497 -430
rect 559 -806 593 -430
rect 655 -806 689 -430
rect 751 -806 785 -430
rect 847 -806 881 -430
rect 943 -806 977 -430
rect -833 -890 -799 -856
rect -641 -890 -607 -856
rect -449 -890 -415 -856
rect -257 -890 -223 -856
rect -65 -890 -31 -856
rect 127 -890 161 -856
rect 319 -890 353 -856
rect 511 -890 545 -856
rect 703 -890 737 -856
rect 895 -890 929 -856
rect -833 -998 -799 -964
rect -641 -998 -607 -964
rect -449 -998 -415 -964
rect -257 -998 -223 -964
rect -65 -998 -31 -964
rect 127 -998 161 -964
rect 319 -998 353 -964
rect 511 -998 545 -964
rect 703 -998 737 -964
rect 895 -998 929 -964
rect -977 -1424 -943 -1048
rect -881 -1424 -847 -1048
rect -785 -1424 -751 -1048
rect -689 -1424 -655 -1048
rect -593 -1424 -559 -1048
rect -497 -1424 -463 -1048
rect -401 -1424 -367 -1048
rect -305 -1424 -271 -1048
rect -209 -1424 -175 -1048
rect -113 -1424 -79 -1048
rect -17 -1424 17 -1048
rect 79 -1424 113 -1048
rect 175 -1424 209 -1048
rect 271 -1424 305 -1048
rect 367 -1424 401 -1048
rect 463 -1424 497 -1048
rect 559 -1424 593 -1048
rect 655 -1424 689 -1048
rect 751 -1424 785 -1048
rect 847 -1424 881 -1048
rect 943 -1424 977 -1048
rect -929 -1508 -895 -1474
rect -737 -1508 -703 -1474
rect -545 -1508 -511 -1474
rect -353 -1508 -319 -1474
rect -161 -1508 -127 -1474
rect 31 -1508 65 -1474
rect 223 -1508 257 -1474
rect 415 -1508 449 -1474
rect 607 -1508 641 -1474
rect 799 -1508 833 -1474
rect -929 -1616 -895 -1582
rect -737 -1616 -703 -1582
rect -545 -1616 -511 -1582
rect -353 -1616 -319 -1582
rect -161 -1616 -127 -1582
rect 31 -1616 65 -1582
rect 223 -1616 257 -1582
rect 415 -1616 449 -1582
rect 607 -1616 641 -1582
rect 799 -1616 833 -1582
rect -977 -2042 -943 -1666
rect -881 -2042 -847 -1666
rect -785 -2042 -751 -1666
rect -689 -2042 -655 -1666
rect -593 -2042 -559 -1666
rect -497 -2042 -463 -1666
rect -401 -2042 -367 -1666
rect -305 -2042 -271 -1666
rect -209 -2042 -175 -1666
rect -113 -2042 -79 -1666
rect -17 -2042 17 -1666
rect 79 -2042 113 -1666
rect 175 -2042 209 -1666
rect 271 -2042 305 -1666
rect 367 -2042 401 -1666
rect 463 -2042 497 -1666
rect 559 -2042 593 -1666
rect 655 -2042 689 -1666
rect 751 -2042 785 -1666
rect 847 -2042 881 -1666
rect 943 -2042 977 -1666
rect -833 -2126 -799 -2092
rect -641 -2126 -607 -2092
rect -449 -2126 -415 -2092
rect -257 -2126 -223 -2092
rect -65 -2126 -31 -2092
rect 127 -2126 161 -2092
rect 319 -2126 353 -2092
rect 511 -2126 545 -2092
rect 703 -2126 737 -2092
rect 895 -2126 929 -2092
rect -833 -2234 -799 -2200
rect -641 -2234 -607 -2200
rect -449 -2234 -415 -2200
rect -257 -2234 -223 -2200
rect -65 -2234 -31 -2200
rect 127 -2234 161 -2200
rect 319 -2234 353 -2200
rect 511 -2234 545 -2200
rect 703 -2234 737 -2200
rect 895 -2234 929 -2200
rect -977 -2660 -943 -2284
rect -881 -2660 -847 -2284
rect -785 -2660 -751 -2284
rect -689 -2660 -655 -2284
rect -593 -2660 -559 -2284
rect -497 -2660 -463 -2284
rect -401 -2660 -367 -2284
rect -305 -2660 -271 -2284
rect -209 -2660 -175 -2284
rect -113 -2660 -79 -2284
rect -17 -2660 17 -2284
rect 79 -2660 113 -2284
rect 175 -2660 209 -2284
rect 271 -2660 305 -2284
rect 367 -2660 401 -2284
rect 463 -2660 497 -2284
rect 559 -2660 593 -2284
rect 655 -2660 689 -2284
rect 751 -2660 785 -2284
rect 847 -2660 881 -2284
rect 943 -2660 977 -2284
rect -929 -2744 -895 -2710
rect -737 -2744 -703 -2710
rect -545 -2744 -511 -2710
rect -353 -2744 -319 -2710
rect -161 -2744 -127 -2710
rect 31 -2744 65 -2710
rect 223 -2744 257 -2710
rect 415 -2744 449 -2710
rect 607 -2744 641 -2710
rect 799 -2744 833 -2710
<< metal1 >>
rect -845 2744 -787 2750
rect -845 2710 -833 2744
rect -799 2710 -787 2744
rect -845 2704 -787 2710
rect -653 2744 -595 2750
rect -653 2710 -641 2744
rect -607 2710 -595 2744
rect -653 2704 -595 2710
rect -461 2744 -403 2750
rect -461 2710 -449 2744
rect -415 2710 -403 2744
rect -461 2704 -403 2710
rect -269 2744 -211 2750
rect -269 2710 -257 2744
rect -223 2710 -211 2744
rect -269 2704 -211 2710
rect -77 2744 -19 2750
rect -77 2710 -65 2744
rect -31 2710 -19 2744
rect -77 2704 -19 2710
rect 115 2744 173 2750
rect 115 2710 127 2744
rect 161 2710 173 2744
rect 115 2704 173 2710
rect 307 2744 365 2750
rect 307 2710 319 2744
rect 353 2710 365 2744
rect 307 2704 365 2710
rect 499 2744 557 2750
rect 499 2710 511 2744
rect 545 2710 557 2744
rect 499 2704 557 2710
rect 691 2744 749 2750
rect 691 2710 703 2744
rect 737 2710 749 2744
rect 691 2704 749 2710
rect 883 2744 941 2750
rect 883 2710 895 2744
rect 929 2710 941 2744
rect 883 2704 941 2710
rect -983 2660 -937 2672
rect -983 2284 -977 2660
rect -943 2284 -937 2660
rect -983 2272 -937 2284
rect -887 2660 -841 2672
rect -887 2284 -881 2660
rect -847 2284 -841 2660
rect -887 2272 -841 2284
rect -791 2660 -745 2672
rect -791 2284 -785 2660
rect -751 2284 -745 2660
rect -791 2272 -745 2284
rect -695 2660 -649 2672
rect -695 2284 -689 2660
rect -655 2284 -649 2660
rect -695 2272 -649 2284
rect -599 2660 -553 2672
rect -599 2284 -593 2660
rect -559 2284 -553 2660
rect -599 2272 -553 2284
rect -503 2660 -457 2672
rect -503 2284 -497 2660
rect -463 2284 -457 2660
rect -503 2272 -457 2284
rect -407 2660 -361 2672
rect -407 2284 -401 2660
rect -367 2284 -361 2660
rect -407 2272 -361 2284
rect -311 2660 -265 2672
rect -311 2284 -305 2660
rect -271 2284 -265 2660
rect -311 2272 -265 2284
rect -215 2660 -169 2672
rect -215 2284 -209 2660
rect -175 2284 -169 2660
rect -215 2272 -169 2284
rect -119 2660 -73 2672
rect -119 2284 -113 2660
rect -79 2284 -73 2660
rect -119 2272 -73 2284
rect -23 2660 23 2672
rect -23 2284 -17 2660
rect 17 2284 23 2660
rect -23 2272 23 2284
rect 73 2660 119 2672
rect 73 2284 79 2660
rect 113 2284 119 2660
rect 73 2272 119 2284
rect 169 2660 215 2672
rect 169 2284 175 2660
rect 209 2284 215 2660
rect 169 2272 215 2284
rect 265 2660 311 2672
rect 265 2284 271 2660
rect 305 2284 311 2660
rect 265 2272 311 2284
rect 361 2660 407 2672
rect 361 2284 367 2660
rect 401 2284 407 2660
rect 361 2272 407 2284
rect 457 2660 503 2672
rect 457 2284 463 2660
rect 497 2284 503 2660
rect 457 2272 503 2284
rect 553 2660 599 2672
rect 553 2284 559 2660
rect 593 2284 599 2660
rect 553 2272 599 2284
rect 649 2660 695 2672
rect 649 2284 655 2660
rect 689 2284 695 2660
rect 649 2272 695 2284
rect 745 2660 791 2672
rect 745 2284 751 2660
rect 785 2284 791 2660
rect 745 2272 791 2284
rect 841 2660 887 2672
rect 841 2284 847 2660
rect 881 2284 887 2660
rect 841 2272 887 2284
rect 937 2660 983 2672
rect 937 2284 943 2660
rect 977 2284 983 2660
rect 937 2272 983 2284
rect -941 2234 -883 2240
rect -941 2200 -929 2234
rect -895 2200 -883 2234
rect -941 2194 -883 2200
rect -749 2234 -691 2240
rect -749 2200 -737 2234
rect -703 2200 -691 2234
rect -749 2194 -691 2200
rect -557 2234 -499 2240
rect -557 2200 -545 2234
rect -511 2200 -499 2234
rect -557 2194 -499 2200
rect -365 2234 -307 2240
rect -365 2200 -353 2234
rect -319 2200 -307 2234
rect -365 2194 -307 2200
rect -173 2234 -115 2240
rect -173 2200 -161 2234
rect -127 2200 -115 2234
rect -173 2194 -115 2200
rect 19 2234 77 2240
rect 19 2200 31 2234
rect 65 2200 77 2234
rect 19 2194 77 2200
rect 211 2234 269 2240
rect 211 2200 223 2234
rect 257 2200 269 2234
rect 211 2194 269 2200
rect 403 2234 461 2240
rect 403 2200 415 2234
rect 449 2200 461 2234
rect 403 2194 461 2200
rect 595 2234 653 2240
rect 595 2200 607 2234
rect 641 2200 653 2234
rect 595 2194 653 2200
rect 787 2234 845 2240
rect 787 2200 799 2234
rect 833 2200 845 2234
rect 787 2194 845 2200
rect -941 2126 -883 2132
rect -941 2092 -929 2126
rect -895 2092 -883 2126
rect -941 2086 -883 2092
rect -749 2126 -691 2132
rect -749 2092 -737 2126
rect -703 2092 -691 2126
rect -749 2086 -691 2092
rect -557 2126 -499 2132
rect -557 2092 -545 2126
rect -511 2092 -499 2126
rect -557 2086 -499 2092
rect -365 2126 -307 2132
rect -365 2092 -353 2126
rect -319 2092 -307 2126
rect -365 2086 -307 2092
rect -173 2126 -115 2132
rect -173 2092 -161 2126
rect -127 2092 -115 2126
rect -173 2086 -115 2092
rect 19 2126 77 2132
rect 19 2092 31 2126
rect 65 2092 77 2126
rect 19 2086 77 2092
rect 211 2126 269 2132
rect 211 2092 223 2126
rect 257 2092 269 2126
rect 211 2086 269 2092
rect 403 2126 461 2132
rect 403 2092 415 2126
rect 449 2092 461 2126
rect 403 2086 461 2092
rect 595 2126 653 2132
rect 595 2092 607 2126
rect 641 2092 653 2126
rect 595 2086 653 2092
rect 787 2126 845 2132
rect 787 2092 799 2126
rect 833 2092 845 2126
rect 787 2086 845 2092
rect -983 2042 -937 2054
rect -983 1666 -977 2042
rect -943 1666 -937 2042
rect -983 1654 -937 1666
rect -887 2042 -841 2054
rect -887 1666 -881 2042
rect -847 1666 -841 2042
rect -887 1654 -841 1666
rect -791 2042 -745 2054
rect -791 1666 -785 2042
rect -751 1666 -745 2042
rect -791 1654 -745 1666
rect -695 2042 -649 2054
rect -695 1666 -689 2042
rect -655 1666 -649 2042
rect -695 1654 -649 1666
rect -599 2042 -553 2054
rect -599 1666 -593 2042
rect -559 1666 -553 2042
rect -599 1654 -553 1666
rect -503 2042 -457 2054
rect -503 1666 -497 2042
rect -463 1666 -457 2042
rect -503 1654 -457 1666
rect -407 2042 -361 2054
rect -407 1666 -401 2042
rect -367 1666 -361 2042
rect -407 1654 -361 1666
rect -311 2042 -265 2054
rect -311 1666 -305 2042
rect -271 1666 -265 2042
rect -311 1654 -265 1666
rect -215 2042 -169 2054
rect -215 1666 -209 2042
rect -175 1666 -169 2042
rect -215 1654 -169 1666
rect -119 2042 -73 2054
rect -119 1666 -113 2042
rect -79 1666 -73 2042
rect -119 1654 -73 1666
rect -23 2042 23 2054
rect -23 1666 -17 2042
rect 17 1666 23 2042
rect -23 1654 23 1666
rect 73 2042 119 2054
rect 73 1666 79 2042
rect 113 1666 119 2042
rect 73 1654 119 1666
rect 169 2042 215 2054
rect 169 1666 175 2042
rect 209 1666 215 2042
rect 169 1654 215 1666
rect 265 2042 311 2054
rect 265 1666 271 2042
rect 305 1666 311 2042
rect 265 1654 311 1666
rect 361 2042 407 2054
rect 361 1666 367 2042
rect 401 1666 407 2042
rect 361 1654 407 1666
rect 457 2042 503 2054
rect 457 1666 463 2042
rect 497 1666 503 2042
rect 457 1654 503 1666
rect 553 2042 599 2054
rect 553 1666 559 2042
rect 593 1666 599 2042
rect 553 1654 599 1666
rect 649 2042 695 2054
rect 649 1666 655 2042
rect 689 1666 695 2042
rect 649 1654 695 1666
rect 745 2042 791 2054
rect 745 1666 751 2042
rect 785 1666 791 2042
rect 745 1654 791 1666
rect 841 2042 887 2054
rect 841 1666 847 2042
rect 881 1666 887 2042
rect 841 1654 887 1666
rect 937 2042 983 2054
rect 937 1666 943 2042
rect 977 1666 983 2042
rect 937 1654 983 1666
rect -845 1616 -787 1622
rect -845 1582 -833 1616
rect -799 1582 -787 1616
rect -845 1576 -787 1582
rect -653 1616 -595 1622
rect -653 1582 -641 1616
rect -607 1582 -595 1616
rect -653 1576 -595 1582
rect -461 1616 -403 1622
rect -461 1582 -449 1616
rect -415 1582 -403 1616
rect -461 1576 -403 1582
rect -269 1616 -211 1622
rect -269 1582 -257 1616
rect -223 1582 -211 1616
rect -269 1576 -211 1582
rect -77 1616 -19 1622
rect -77 1582 -65 1616
rect -31 1582 -19 1616
rect -77 1576 -19 1582
rect 115 1616 173 1622
rect 115 1582 127 1616
rect 161 1582 173 1616
rect 115 1576 173 1582
rect 307 1616 365 1622
rect 307 1582 319 1616
rect 353 1582 365 1616
rect 307 1576 365 1582
rect 499 1616 557 1622
rect 499 1582 511 1616
rect 545 1582 557 1616
rect 499 1576 557 1582
rect 691 1616 749 1622
rect 691 1582 703 1616
rect 737 1582 749 1616
rect 691 1576 749 1582
rect 883 1616 941 1622
rect 883 1582 895 1616
rect 929 1582 941 1616
rect 883 1576 941 1582
rect -845 1508 -787 1514
rect -845 1474 -833 1508
rect -799 1474 -787 1508
rect -845 1468 -787 1474
rect -653 1508 -595 1514
rect -653 1474 -641 1508
rect -607 1474 -595 1508
rect -653 1468 -595 1474
rect -461 1508 -403 1514
rect -461 1474 -449 1508
rect -415 1474 -403 1508
rect -461 1468 -403 1474
rect -269 1508 -211 1514
rect -269 1474 -257 1508
rect -223 1474 -211 1508
rect -269 1468 -211 1474
rect -77 1508 -19 1514
rect -77 1474 -65 1508
rect -31 1474 -19 1508
rect -77 1468 -19 1474
rect 115 1508 173 1514
rect 115 1474 127 1508
rect 161 1474 173 1508
rect 115 1468 173 1474
rect 307 1508 365 1514
rect 307 1474 319 1508
rect 353 1474 365 1508
rect 307 1468 365 1474
rect 499 1508 557 1514
rect 499 1474 511 1508
rect 545 1474 557 1508
rect 499 1468 557 1474
rect 691 1508 749 1514
rect 691 1474 703 1508
rect 737 1474 749 1508
rect 691 1468 749 1474
rect 883 1508 941 1514
rect 883 1474 895 1508
rect 929 1474 941 1508
rect 883 1468 941 1474
rect -983 1424 -937 1436
rect -983 1048 -977 1424
rect -943 1048 -937 1424
rect -983 1036 -937 1048
rect -887 1424 -841 1436
rect -887 1048 -881 1424
rect -847 1048 -841 1424
rect -887 1036 -841 1048
rect -791 1424 -745 1436
rect -791 1048 -785 1424
rect -751 1048 -745 1424
rect -791 1036 -745 1048
rect -695 1424 -649 1436
rect -695 1048 -689 1424
rect -655 1048 -649 1424
rect -695 1036 -649 1048
rect -599 1424 -553 1436
rect -599 1048 -593 1424
rect -559 1048 -553 1424
rect -599 1036 -553 1048
rect -503 1424 -457 1436
rect -503 1048 -497 1424
rect -463 1048 -457 1424
rect -503 1036 -457 1048
rect -407 1424 -361 1436
rect -407 1048 -401 1424
rect -367 1048 -361 1424
rect -407 1036 -361 1048
rect -311 1424 -265 1436
rect -311 1048 -305 1424
rect -271 1048 -265 1424
rect -311 1036 -265 1048
rect -215 1424 -169 1436
rect -215 1048 -209 1424
rect -175 1048 -169 1424
rect -215 1036 -169 1048
rect -119 1424 -73 1436
rect -119 1048 -113 1424
rect -79 1048 -73 1424
rect -119 1036 -73 1048
rect -23 1424 23 1436
rect -23 1048 -17 1424
rect 17 1048 23 1424
rect -23 1036 23 1048
rect 73 1424 119 1436
rect 73 1048 79 1424
rect 113 1048 119 1424
rect 73 1036 119 1048
rect 169 1424 215 1436
rect 169 1048 175 1424
rect 209 1048 215 1424
rect 169 1036 215 1048
rect 265 1424 311 1436
rect 265 1048 271 1424
rect 305 1048 311 1424
rect 265 1036 311 1048
rect 361 1424 407 1436
rect 361 1048 367 1424
rect 401 1048 407 1424
rect 361 1036 407 1048
rect 457 1424 503 1436
rect 457 1048 463 1424
rect 497 1048 503 1424
rect 457 1036 503 1048
rect 553 1424 599 1436
rect 553 1048 559 1424
rect 593 1048 599 1424
rect 553 1036 599 1048
rect 649 1424 695 1436
rect 649 1048 655 1424
rect 689 1048 695 1424
rect 649 1036 695 1048
rect 745 1424 791 1436
rect 745 1048 751 1424
rect 785 1048 791 1424
rect 745 1036 791 1048
rect 841 1424 887 1436
rect 841 1048 847 1424
rect 881 1048 887 1424
rect 841 1036 887 1048
rect 937 1424 983 1436
rect 937 1048 943 1424
rect 977 1048 983 1424
rect 937 1036 983 1048
rect -941 998 -883 1004
rect -941 964 -929 998
rect -895 964 -883 998
rect -941 958 -883 964
rect -749 998 -691 1004
rect -749 964 -737 998
rect -703 964 -691 998
rect -749 958 -691 964
rect -557 998 -499 1004
rect -557 964 -545 998
rect -511 964 -499 998
rect -557 958 -499 964
rect -365 998 -307 1004
rect -365 964 -353 998
rect -319 964 -307 998
rect -365 958 -307 964
rect -173 998 -115 1004
rect -173 964 -161 998
rect -127 964 -115 998
rect -173 958 -115 964
rect 19 998 77 1004
rect 19 964 31 998
rect 65 964 77 998
rect 19 958 77 964
rect 211 998 269 1004
rect 211 964 223 998
rect 257 964 269 998
rect 211 958 269 964
rect 403 998 461 1004
rect 403 964 415 998
rect 449 964 461 998
rect 403 958 461 964
rect 595 998 653 1004
rect 595 964 607 998
rect 641 964 653 998
rect 595 958 653 964
rect 787 998 845 1004
rect 787 964 799 998
rect 833 964 845 998
rect 787 958 845 964
rect -941 890 -883 896
rect -941 856 -929 890
rect -895 856 -883 890
rect -941 850 -883 856
rect -749 890 -691 896
rect -749 856 -737 890
rect -703 856 -691 890
rect -749 850 -691 856
rect -557 890 -499 896
rect -557 856 -545 890
rect -511 856 -499 890
rect -557 850 -499 856
rect -365 890 -307 896
rect -365 856 -353 890
rect -319 856 -307 890
rect -365 850 -307 856
rect -173 890 -115 896
rect -173 856 -161 890
rect -127 856 -115 890
rect -173 850 -115 856
rect 19 890 77 896
rect 19 856 31 890
rect 65 856 77 890
rect 19 850 77 856
rect 211 890 269 896
rect 211 856 223 890
rect 257 856 269 890
rect 211 850 269 856
rect 403 890 461 896
rect 403 856 415 890
rect 449 856 461 890
rect 403 850 461 856
rect 595 890 653 896
rect 595 856 607 890
rect 641 856 653 890
rect 595 850 653 856
rect 787 890 845 896
rect 787 856 799 890
rect 833 856 845 890
rect 787 850 845 856
rect -983 806 -937 818
rect -983 430 -977 806
rect -943 430 -937 806
rect -983 418 -937 430
rect -887 806 -841 818
rect -887 430 -881 806
rect -847 430 -841 806
rect -887 418 -841 430
rect -791 806 -745 818
rect -791 430 -785 806
rect -751 430 -745 806
rect -791 418 -745 430
rect -695 806 -649 818
rect -695 430 -689 806
rect -655 430 -649 806
rect -695 418 -649 430
rect -599 806 -553 818
rect -599 430 -593 806
rect -559 430 -553 806
rect -599 418 -553 430
rect -503 806 -457 818
rect -503 430 -497 806
rect -463 430 -457 806
rect -503 418 -457 430
rect -407 806 -361 818
rect -407 430 -401 806
rect -367 430 -361 806
rect -407 418 -361 430
rect -311 806 -265 818
rect -311 430 -305 806
rect -271 430 -265 806
rect -311 418 -265 430
rect -215 806 -169 818
rect -215 430 -209 806
rect -175 430 -169 806
rect -215 418 -169 430
rect -119 806 -73 818
rect -119 430 -113 806
rect -79 430 -73 806
rect -119 418 -73 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 73 806 119 818
rect 73 430 79 806
rect 113 430 119 806
rect 73 418 119 430
rect 169 806 215 818
rect 169 430 175 806
rect 209 430 215 806
rect 169 418 215 430
rect 265 806 311 818
rect 265 430 271 806
rect 305 430 311 806
rect 265 418 311 430
rect 361 806 407 818
rect 361 430 367 806
rect 401 430 407 806
rect 361 418 407 430
rect 457 806 503 818
rect 457 430 463 806
rect 497 430 503 806
rect 457 418 503 430
rect 553 806 599 818
rect 553 430 559 806
rect 593 430 599 806
rect 553 418 599 430
rect 649 806 695 818
rect 649 430 655 806
rect 689 430 695 806
rect 649 418 695 430
rect 745 806 791 818
rect 745 430 751 806
rect 785 430 791 806
rect 745 418 791 430
rect 841 806 887 818
rect 841 430 847 806
rect 881 430 887 806
rect 841 418 887 430
rect 937 806 983 818
rect 937 430 943 806
rect 977 430 983 806
rect 937 418 983 430
rect -845 380 -787 386
rect -845 346 -833 380
rect -799 346 -787 380
rect -845 340 -787 346
rect -653 380 -595 386
rect -653 346 -641 380
rect -607 346 -595 380
rect -653 340 -595 346
rect -461 380 -403 386
rect -461 346 -449 380
rect -415 346 -403 380
rect -461 340 -403 346
rect -269 380 -211 386
rect -269 346 -257 380
rect -223 346 -211 380
rect -269 340 -211 346
rect -77 380 -19 386
rect -77 346 -65 380
rect -31 346 -19 380
rect -77 340 -19 346
rect 115 380 173 386
rect 115 346 127 380
rect 161 346 173 380
rect 115 340 173 346
rect 307 380 365 386
rect 307 346 319 380
rect 353 346 365 380
rect 307 340 365 346
rect 499 380 557 386
rect 499 346 511 380
rect 545 346 557 380
rect 499 340 557 346
rect 691 380 749 386
rect 691 346 703 380
rect 737 346 749 380
rect 691 340 749 346
rect 883 380 941 386
rect 883 346 895 380
rect 929 346 941 380
rect 883 340 941 346
rect -845 272 -787 278
rect -845 238 -833 272
rect -799 238 -787 272
rect -845 232 -787 238
rect -653 272 -595 278
rect -653 238 -641 272
rect -607 238 -595 272
rect -653 232 -595 238
rect -461 272 -403 278
rect -461 238 -449 272
rect -415 238 -403 272
rect -461 232 -403 238
rect -269 272 -211 278
rect -269 238 -257 272
rect -223 238 -211 272
rect -269 232 -211 238
rect -77 272 -19 278
rect -77 238 -65 272
rect -31 238 -19 272
rect -77 232 -19 238
rect 115 272 173 278
rect 115 238 127 272
rect 161 238 173 272
rect 115 232 173 238
rect 307 272 365 278
rect 307 238 319 272
rect 353 238 365 272
rect 307 232 365 238
rect 499 272 557 278
rect 499 238 511 272
rect 545 238 557 272
rect 499 232 557 238
rect 691 272 749 278
rect 691 238 703 272
rect 737 238 749 272
rect 691 232 749 238
rect 883 272 941 278
rect 883 238 895 272
rect 929 238 941 272
rect 883 232 941 238
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect -941 -238 -883 -232
rect -941 -272 -929 -238
rect -895 -272 -883 -238
rect -941 -278 -883 -272
rect -749 -238 -691 -232
rect -749 -272 -737 -238
rect -703 -272 -691 -238
rect -749 -278 -691 -272
rect -557 -238 -499 -232
rect -557 -272 -545 -238
rect -511 -272 -499 -238
rect -557 -278 -499 -272
rect -365 -238 -307 -232
rect -365 -272 -353 -238
rect -319 -272 -307 -238
rect -365 -278 -307 -272
rect -173 -238 -115 -232
rect -173 -272 -161 -238
rect -127 -272 -115 -238
rect -173 -278 -115 -272
rect 19 -238 77 -232
rect 19 -272 31 -238
rect 65 -272 77 -238
rect 19 -278 77 -272
rect 211 -238 269 -232
rect 211 -272 223 -238
rect 257 -272 269 -238
rect 211 -278 269 -272
rect 403 -238 461 -232
rect 403 -272 415 -238
rect 449 -272 461 -238
rect 403 -278 461 -272
rect 595 -238 653 -232
rect 595 -272 607 -238
rect 641 -272 653 -238
rect 595 -278 653 -272
rect 787 -238 845 -232
rect 787 -272 799 -238
rect 833 -272 845 -238
rect 787 -278 845 -272
rect -941 -346 -883 -340
rect -941 -380 -929 -346
rect -895 -380 -883 -346
rect -941 -386 -883 -380
rect -749 -346 -691 -340
rect -749 -380 -737 -346
rect -703 -380 -691 -346
rect -749 -386 -691 -380
rect -557 -346 -499 -340
rect -557 -380 -545 -346
rect -511 -380 -499 -346
rect -557 -386 -499 -380
rect -365 -346 -307 -340
rect -365 -380 -353 -346
rect -319 -380 -307 -346
rect -365 -386 -307 -380
rect -173 -346 -115 -340
rect -173 -380 -161 -346
rect -127 -380 -115 -346
rect -173 -386 -115 -380
rect 19 -346 77 -340
rect 19 -380 31 -346
rect 65 -380 77 -346
rect 19 -386 77 -380
rect 211 -346 269 -340
rect 211 -380 223 -346
rect 257 -380 269 -346
rect 211 -386 269 -380
rect 403 -346 461 -340
rect 403 -380 415 -346
rect 449 -380 461 -346
rect 403 -386 461 -380
rect 595 -346 653 -340
rect 595 -380 607 -346
rect 641 -380 653 -346
rect 595 -386 653 -380
rect 787 -346 845 -340
rect 787 -380 799 -346
rect 833 -380 845 -346
rect 787 -386 845 -380
rect -983 -430 -937 -418
rect -983 -806 -977 -430
rect -943 -806 -937 -430
rect -983 -818 -937 -806
rect -887 -430 -841 -418
rect -887 -806 -881 -430
rect -847 -806 -841 -430
rect -887 -818 -841 -806
rect -791 -430 -745 -418
rect -791 -806 -785 -430
rect -751 -806 -745 -430
rect -791 -818 -745 -806
rect -695 -430 -649 -418
rect -695 -806 -689 -430
rect -655 -806 -649 -430
rect -695 -818 -649 -806
rect -599 -430 -553 -418
rect -599 -806 -593 -430
rect -559 -806 -553 -430
rect -599 -818 -553 -806
rect -503 -430 -457 -418
rect -503 -806 -497 -430
rect -463 -806 -457 -430
rect -503 -818 -457 -806
rect -407 -430 -361 -418
rect -407 -806 -401 -430
rect -367 -806 -361 -430
rect -407 -818 -361 -806
rect -311 -430 -265 -418
rect -311 -806 -305 -430
rect -271 -806 -265 -430
rect -311 -818 -265 -806
rect -215 -430 -169 -418
rect -215 -806 -209 -430
rect -175 -806 -169 -430
rect -215 -818 -169 -806
rect -119 -430 -73 -418
rect -119 -806 -113 -430
rect -79 -806 -73 -430
rect -119 -818 -73 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 73 -430 119 -418
rect 73 -806 79 -430
rect 113 -806 119 -430
rect 73 -818 119 -806
rect 169 -430 215 -418
rect 169 -806 175 -430
rect 209 -806 215 -430
rect 169 -818 215 -806
rect 265 -430 311 -418
rect 265 -806 271 -430
rect 305 -806 311 -430
rect 265 -818 311 -806
rect 361 -430 407 -418
rect 361 -806 367 -430
rect 401 -806 407 -430
rect 361 -818 407 -806
rect 457 -430 503 -418
rect 457 -806 463 -430
rect 497 -806 503 -430
rect 457 -818 503 -806
rect 553 -430 599 -418
rect 553 -806 559 -430
rect 593 -806 599 -430
rect 553 -818 599 -806
rect 649 -430 695 -418
rect 649 -806 655 -430
rect 689 -806 695 -430
rect 649 -818 695 -806
rect 745 -430 791 -418
rect 745 -806 751 -430
rect 785 -806 791 -430
rect 745 -818 791 -806
rect 841 -430 887 -418
rect 841 -806 847 -430
rect 881 -806 887 -430
rect 841 -818 887 -806
rect 937 -430 983 -418
rect 937 -806 943 -430
rect 977 -806 983 -430
rect 937 -818 983 -806
rect -845 -856 -787 -850
rect -845 -890 -833 -856
rect -799 -890 -787 -856
rect -845 -896 -787 -890
rect -653 -856 -595 -850
rect -653 -890 -641 -856
rect -607 -890 -595 -856
rect -653 -896 -595 -890
rect -461 -856 -403 -850
rect -461 -890 -449 -856
rect -415 -890 -403 -856
rect -461 -896 -403 -890
rect -269 -856 -211 -850
rect -269 -890 -257 -856
rect -223 -890 -211 -856
rect -269 -896 -211 -890
rect -77 -856 -19 -850
rect -77 -890 -65 -856
rect -31 -890 -19 -856
rect -77 -896 -19 -890
rect 115 -856 173 -850
rect 115 -890 127 -856
rect 161 -890 173 -856
rect 115 -896 173 -890
rect 307 -856 365 -850
rect 307 -890 319 -856
rect 353 -890 365 -856
rect 307 -896 365 -890
rect 499 -856 557 -850
rect 499 -890 511 -856
rect 545 -890 557 -856
rect 499 -896 557 -890
rect 691 -856 749 -850
rect 691 -890 703 -856
rect 737 -890 749 -856
rect 691 -896 749 -890
rect 883 -856 941 -850
rect 883 -890 895 -856
rect 929 -890 941 -856
rect 883 -896 941 -890
rect -845 -964 -787 -958
rect -845 -998 -833 -964
rect -799 -998 -787 -964
rect -845 -1004 -787 -998
rect -653 -964 -595 -958
rect -653 -998 -641 -964
rect -607 -998 -595 -964
rect -653 -1004 -595 -998
rect -461 -964 -403 -958
rect -461 -998 -449 -964
rect -415 -998 -403 -964
rect -461 -1004 -403 -998
rect -269 -964 -211 -958
rect -269 -998 -257 -964
rect -223 -998 -211 -964
rect -269 -1004 -211 -998
rect -77 -964 -19 -958
rect -77 -998 -65 -964
rect -31 -998 -19 -964
rect -77 -1004 -19 -998
rect 115 -964 173 -958
rect 115 -998 127 -964
rect 161 -998 173 -964
rect 115 -1004 173 -998
rect 307 -964 365 -958
rect 307 -998 319 -964
rect 353 -998 365 -964
rect 307 -1004 365 -998
rect 499 -964 557 -958
rect 499 -998 511 -964
rect 545 -998 557 -964
rect 499 -1004 557 -998
rect 691 -964 749 -958
rect 691 -998 703 -964
rect 737 -998 749 -964
rect 691 -1004 749 -998
rect 883 -964 941 -958
rect 883 -998 895 -964
rect 929 -998 941 -964
rect 883 -1004 941 -998
rect -983 -1048 -937 -1036
rect -983 -1424 -977 -1048
rect -943 -1424 -937 -1048
rect -983 -1436 -937 -1424
rect -887 -1048 -841 -1036
rect -887 -1424 -881 -1048
rect -847 -1424 -841 -1048
rect -887 -1436 -841 -1424
rect -791 -1048 -745 -1036
rect -791 -1424 -785 -1048
rect -751 -1424 -745 -1048
rect -791 -1436 -745 -1424
rect -695 -1048 -649 -1036
rect -695 -1424 -689 -1048
rect -655 -1424 -649 -1048
rect -695 -1436 -649 -1424
rect -599 -1048 -553 -1036
rect -599 -1424 -593 -1048
rect -559 -1424 -553 -1048
rect -599 -1436 -553 -1424
rect -503 -1048 -457 -1036
rect -503 -1424 -497 -1048
rect -463 -1424 -457 -1048
rect -503 -1436 -457 -1424
rect -407 -1048 -361 -1036
rect -407 -1424 -401 -1048
rect -367 -1424 -361 -1048
rect -407 -1436 -361 -1424
rect -311 -1048 -265 -1036
rect -311 -1424 -305 -1048
rect -271 -1424 -265 -1048
rect -311 -1436 -265 -1424
rect -215 -1048 -169 -1036
rect -215 -1424 -209 -1048
rect -175 -1424 -169 -1048
rect -215 -1436 -169 -1424
rect -119 -1048 -73 -1036
rect -119 -1424 -113 -1048
rect -79 -1424 -73 -1048
rect -119 -1436 -73 -1424
rect -23 -1048 23 -1036
rect -23 -1424 -17 -1048
rect 17 -1424 23 -1048
rect -23 -1436 23 -1424
rect 73 -1048 119 -1036
rect 73 -1424 79 -1048
rect 113 -1424 119 -1048
rect 73 -1436 119 -1424
rect 169 -1048 215 -1036
rect 169 -1424 175 -1048
rect 209 -1424 215 -1048
rect 169 -1436 215 -1424
rect 265 -1048 311 -1036
rect 265 -1424 271 -1048
rect 305 -1424 311 -1048
rect 265 -1436 311 -1424
rect 361 -1048 407 -1036
rect 361 -1424 367 -1048
rect 401 -1424 407 -1048
rect 361 -1436 407 -1424
rect 457 -1048 503 -1036
rect 457 -1424 463 -1048
rect 497 -1424 503 -1048
rect 457 -1436 503 -1424
rect 553 -1048 599 -1036
rect 553 -1424 559 -1048
rect 593 -1424 599 -1048
rect 553 -1436 599 -1424
rect 649 -1048 695 -1036
rect 649 -1424 655 -1048
rect 689 -1424 695 -1048
rect 649 -1436 695 -1424
rect 745 -1048 791 -1036
rect 745 -1424 751 -1048
rect 785 -1424 791 -1048
rect 745 -1436 791 -1424
rect 841 -1048 887 -1036
rect 841 -1424 847 -1048
rect 881 -1424 887 -1048
rect 841 -1436 887 -1424
rect 937 -1048 983 -1036
rect 937 -1424 943 -1048
rect 977 -1424 983 -1048
rect 937 -1436 983 -1424
rect -941 -1474 -883 -1468
rect -941 -1508 -929 -1474
rect -895 -1508 -883 -1474
rect -941 -1514 -883 -1508
rect -749 -1474 -691 -1468
rect -749 -1508 -737 -1474
rect -703 -1508 -691 -1474
rect -749 -1514 -691 -1508
rect -557 -1474 -499 -1468
rect -557 -1508 -545 -1474
rect -511 -1508 -499 -1474
rect -557 -1514 -499 -1508
rect -365 -1474 -307 -1468
rect -365 -1508 -353 -1474
rect -319 -1508 -307 -1474
rect -365 -1514 -307 -1508
rect -173 -1474 -115 -1468
rect -173 -1508 -161 -1474
rect -127 -1508 -115 -1474
rect -173 -1514 -115 -1508
rect 19 -1474 77 -1468
rect 19 -1508 31 -1474
rect 65 -1508 77 -1474
rect 19 -1514 77 -1508
rect 211 -1474 269 -1468
rect 211 -1508 223 -1474
rect 257 -1508 269 -1474
rect 211 -1514 269 -1508
rect 403 -1474 461 -1468
rect 403 -1508 415 -1474
rect 449 -1508 461 -1474
rect 403 -1514 461 -1508
rect 595 -1474 653 -1468
rect 595 -1508 607 -1474
rect 641 -1508 653 -1474
rect 595 -1514 653 -1508
rect 787 -1474 845 -1468
rect 787 -1508 799 -1474
rect 833 -1508 845 -1474
rect 787 -1514 845 -1508
rect -941 -1582 -883 -1576
rect -941 -1616 -929 -1582
rect -895 -1616 -883 -1582
rect -941 -1622 -883 -1616
rect -749 -1582 -691 -1576
rect -749 -1616 -737 -1582
rect -703 -1616 -691 -1582
rect -749 -1622 -691 -1616
rect -557 -1582 -499 -1576
rect -557 -1616 -545 -1582
rect -511 -1616 -499 -1582
rect -557 -1622 -499 -1616
rect -365 -1582 -307 -1576
rect -365 -1616 -353 -1582
rect -319 -1616 -307 -1582
rect -365 -1622 -307 -1616
rect -173 -1582 -115 -1576
rect -173 -1616 -161 -1582
rect -127 -1616 -115 -1582
rect -173 -1622 -115 -1616
rect 19 -1582 77 -1576
rect 19 -1616 31 -1582
rect 65 -1616 77 -1582
rect 19 -1622 77 -1616
rect 211 -1582 269 -1576
rect 211 -1616 223 -1582
rect 257 -1616 269 -1582
rect 211 -1622 269 -1616
rect 403 -1582 461 -1576
rect 403 -1616 415 -1582
rect 449 -1616 461 -1582
rect 403 -1622 461 -1616
rect 595 -1582 653 -1576
rect 595 -1616 607 -1582
rect 641 -1616 653 -1582
rect 595 -1622 653 -1616
rect 787 -1582 845 -1576
rect 787 -1616 799 -1582
rect 833 -1616 845 -1582
rect 787 -1622 845 -1616
rect -983 -1666 -937 -1654
rect -983 -2042 -977 -1666
rect -943 -2042 -937 -1666
rect -983 -2054 -937 -2042
rect -887 -1666 -841 -1654
rect -887 -2042 -881 -1666
rect -847 -2042 -841 -1666
rect -887 -2054 -841 -2042
rect -791 -1666 -745 -1654
rect -791 -2042 -785 -1666
rect -751 -2042 -745 -1666
rect -791 -2054 -745 -2042
rect -695 -1666 -649 -1654
rect -695 -2042 -689 -1666
rect -655 -2042 -649 -1666
rect -695 -2054 -649 -2042
rect -599 -1666 -553 -1654
rect -599 -2042 -593 -1666
rect -559 -2042 -553 -1666
rect -599 -2054 -553 -2042
rect -503 -1666 -457 -1654
rect -503 -2042 -497 -1666
rect -463 -2042 -457 -1666
rect -503 -2054 -457 -2042
rect -407 -1666 -361 -1654
rect -407 -2042 -401 -1666
rect -367 -2042 -361 -1666
rect -407 -2054 -361 -2042
rect -311 -1666 -265 -1654
rect -311 -2042 -305 -1666
rect -271 -2042 -265 -1666
rect -311 -2054 -265 -2042
rect -215 -1666 -169 -1654
rect -215 -2042 -209 -1666
rect -175 -2042 -169 -1666
rect -215 -2054 -169 -2042
rect -119 -1666 -73 -1654
rect -119 -2042 -113 -1666
rect -79 -2042 -73 -1666
rect -119 -2054 -73 -2042
rect -23 -1666 23 -1654
rect -23 -2042 -17 -1666
rect 17 -2042 23 -1666
rect -23 -2054 23 -2042
rect 73 -1666 119 -1654
rect 73 -2042 79 -1666
rect 113 -2042 119 -1666
rect 73 -2054 119 -2042
rect 169 -1666 215 -1654
rect 169 -2042 175 -1666
rect 209 -2042 215 -1666
rect 169 -2054 215 -2042
rect 265 -1666 311 -1654
rect 265 -2042 271 -1666
rect 305 -2042 311 -1666
rect 265 -2054 311 -2042
rect 361 -1666 407 -1654
rect 361 -2042 367 -1666
rect 401 -2042 407 -1666
rect 361 -2054 407 -2042
rect 457 -1666 503 -1654
rect 457 -2042 463 -1666
rect 497 -2042 503 -1666
rect 457 -2054 503 -2042
rect 553 -1666 599 -1654
rect 553 -2042 559 -1666
rect 593 -2042 599 -1666
rect 553 -2054 599 -2042
rect 649 -1666 695 -1654
rect 649 -2042 655 -1666
rect 689 -2042 695 -1666
rect 649 -2054 695 -2042
rect 745 -1666 791 -1654
rect 745 -2042 751 -1666
rect 785 -2042 791 -1666
rect 745 -2054 791 -2042
rect 841 -1666 887 -1654
rect 841 -2042 847 -1666
rect 881 -2042 887 -1666
rect 841 -2054 887 -2042
rect 937 -1666 983 -1654
rect 937 -2042 943 -1666
rect 977 -2042 983 -1666
rect 937 -2054 983 -2042
rect -845 -2092 -787 -2086
rect -845 -2126 -833 -2092
rect -799 -2126 -787 -2092
rect -845 -2132 -787 -2126
rect -653 -2092 -595 -2086
rect -653 -2126 -641 -2092
rect -607 -2126 -595 -2092
rect -653 -2132 -595 -2126
rect -461 -2092 -403 -2086
rect -461 -2126 -449 -2092
rect -415 -2126 -403 -2092
rect -461 -2132 -403 -2126
rect -269 -2092 -211 -2086
rect -269 -2126 -257 -2092
rect -223 -2126 -211 -2092
rect -269 -2132 -211 -2126
rect -77 -2092 -19 -2086
rect -77 -2126 -65 -2092
rect -31 -2126 -19 -2092
rect -77 -2132 -19 -2126
rect 115 -2092 173 -2086
rect 115 -2126 127 -2092
rect 161 -2126 173 -2092
rect 115 -2132 173 -2126
rect 307 -2092 365 -2086
rect 307 -2126 319 -2092
rect 353 -2126 365 -2092
rect 307 -2132 365 -2126
rect 499 -2092 557 -2086
rect 499 -2126 511 -2092
rect 545 -2126 557 -2092
rect 499 -2132 557 -2126
rect 691 -2092 749 -2086
rect 691 -2126 703 -2092
rect 737 -2126 749 -2092
rect 691 -2132 749 -2126
rect 883 -2092 941 -2086
rect 883 -2126 895 -2092
rect 929 -2126 941 -2092
rect 883 -2132 941 -2126
rect -845 -2200 -787 -2194
rect -845 -2234 -833 -2200
rect -799 -2234 -787 -2200
rect -845 -2240 -787 -2234
rect -653 -2200 -595 -2194
rect -653 -2234 -641 -2200
rect -607 -2234 -595 -2200
rect -653 -2240 -595 -2234
rect -461 -2200 -403 -2194
rect -461 -2234 -449 -2200
rect -415 -2234 -403 -2200
rect -461 -2240 -403 -2234
rect -269 -2200 -211 -2194
rect -269 -2234 -257 -2200
rect -223 -2234 -211 -2200
rect -269 -2240 -211 -2234
rect -77 -2200 -19 -2194
rect -77 -2234 -65 -2200
rect -31 -2234 -19 -2200
rect -77 -2240 -19 -2234
rect 115 -2200 173 -2194
rect 115 -2234 127 -2200
rect 161 -2234 173 -2200
rect 115 -2240 173 -2234
rect 307 -2200 365 -2194
rect 307 -2234 319 -2200
rect 353 -2234 365 -2200
rect 307 -2240 365 -2234
rect 499 -2200 557 -2194
rect 499 -2234 511 -2200
rect 545 -2234 557 -2200
rect 499 -2240 557 -2234
rect 691 -2200 749 -2194
rect 691 -2234 703 -2200
rect 737 -2234 749 -2200
rect 691 -2240 749 -2234
rect 883 -2200 941 -2194
rect 883 -2234 895 -2200
rect 929 -2234 941 -2200
rect 883 -2240 941 -2234
rect -983 -2284 -937 -2272
rect -983 -2660 -977 -2284
rect -943 -2660 -937 -2284
rect -983 -2672 -937 -2660
rect -887 -2284 -841 -2272
rect -887 -2660 -881 -2284
rect -847 -2660 -841 -2284
rect -887 -2672 -841 -2660
rect -791 -2284 -745 -2272
rect -791 -2660 -785 -2284
rect -751 -2660 -745 -2284
rect -791 -2672 -745 -2660
rect -695 -2284 -649 -2272
rect -695 -2660 -689 -2284
rect -655 -2660 -649 -2284
rect -695 -2672 -649 -2660
rect -599 -2284 -553 -2272
rect -599 -2660 -593 -2284
rect -559 -2660 -553 -2284
rect -599 -2672 -553 -2660
rect -503 -2284 -457 -2272
rect -503 -2660 -497 -2284
rect -463 -2660 -457 -2284
rect -503 -2672 -457 -2660
rect -407 -2284 -361 -2272
rect -407 -2660 -401 -2284
rect -367 -2660 -361 -2284
rect -407 -2672 -361 -2660
rect -311 -2284 -265 -2272
rect -311 -2660 -305 -2284
rect -271 -2660 -265 -2284
rect -311 -2672 -265 -2660
rect -215 -2284 -169 -2272
rect -215 -2660 -209 -2284
rect -175 -2660 -169 -2284
rect -215 -2672 -169 -2660
rect -119 -2284 -73 -2272
rect -119 -2660 -113 -2284
rect -79 -2660 -73 -2284
rect -119 -2672 -73 -2660
rect -23 -2284 23 -2272
rect -23 -2660 -17 -2284
rect 17 -2660 23 -2284
rect -23 -2672 23 -2660
rect 73 -2284 119 -2272
rect 73 -2660 79 -2284
rect 113 -2660 119 -2284
rect 73 -2672 119 -2660
rect 169 -2284 215 -2272
rect 169 -2660 175 -2284
rect 209 -2660 215 -2284
rect 169 -2672 215 -2660
rect 265 -2284 311 -2272
rect 265 -2660 271 -2284
rect 305 -2660 311 -2284
rect 265 -2672 311 -2660
rect 361 -2284 407 -2272
rect 361 -2660 367 -2284
rect 401 -2660 407 -2284
rect 361 -2672 407 -2660
rect 457 -2284 503 -2272
rect 457 -2660 463 -2284
rect 497 -2660 503 -2284
rect 457 -2672 503 -2660
rect 553 -2284 599 -2272
rect 553 -2660 559 -2284
rect 593 -2660 599 -2284
rect 553 -2672 599 -2660
rect 649 -2284 695 -2272
rect 649 -2660 655 -2284
rect 689 -2660 695 -2284
rect 649 -2672 695 -2660
rect 745 -2284 791 -2272
rect 745 -2660 751 -2284
rect 785 -2660 791 -2284
rect 745 -2672 791 -2660
rect 841 -2284 887 -2272
rect 841 -2660 847 -2284
rect 881 -2660 887 -2284
rect 841 -2672 887 -2660
rect 937 -2284 983 -2272
rect 937 -2660 943 -2284
rect 977 -2660 983 -2284
rect 937 -2672 983 -2660
rect -941 -2710 -883 -2704
rect -941 -2744 -929 -2710
rect -895 -2744 -883 -2710
rect -941 -2750 -883 -2744
rect -749 -2710 -691 -2704
rect -749 -2744 -737 -2710
rect -703 -2744 -691 -2710
rect -749 -2750 -691 -2744
rect -557 -2710 -499 -2704
rect -557 -2744 -545 -2710
rect -511 -2744 -499 -2710
rect -557 -2750 -499 -2744
rect -365 -2710 -307 -2704
rect -365 -2744 -353 -2710
rect -319 -2744 -307 -2710
rect -365 -2750 -307 -2744
rect -173 -2710 -115 -2704
rect -173 -2744 -161 -2710
rect -127 -2744 -115 -2710
rect -173 -2750 -115 -2744
rect 19 -2710 77 -2704
rect 19 -2744 31 -2710
rect 65 -2744 77 -2710
rect 19 -2750 77 -2744
rect 211 -2710 269 -2704
rect 211 -2744 223 -2710
rect 257 -2744 269 -2710
rect 211 -2750 269 -2744
rect 403 -2710 461 -2704
rect 403 -2744 415 -2710
rect 449 -2744 461 -2710
rect 403 -2750 461 -2744
rect 595 -2710 653 -2704
rect 595 -2744 607 -2710
rect 641 -2744 653 -2710
rect 595 -2750 653 -2744
rect 787 -2710 845 -2704
rect 787 -2744 799 -2710
rect 833 -2744 845 -2710
rect 787 -2750 845 -2744
<< properties >>
string FIXED_BBOX -1074 -2829 1074 2829
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 9 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
