magic
tech sky130A
magscale 1 2
timestamp 1685031707
<< metal3 >>
rect -386 1012 386 1040
rect -386 -1012 302 1012
rect 366 -1012 386 1012
rect -386 -1040 386 -1012
<< via3 >>
rect 302 -1012 366 1012
<< mimcap >>
rect -346 960 54 1000
rect -346 -960 -306 960
rect 14 -960 54 960
rect -346 -1000 54 -960
<< mimcapcontact >>
rect -306 -960 14 960
<< metal4 >>
rect 286 1012 382 1028
rect -307 960 15 961
rect -307 -960 -306 960
rect 14 -960 15 960
rect -307 -961 15 -960
rect 286 -1012 302 1012
rect 366 -1012 382 1012
rect 286 -1028 382 -1012
<< properties >>
string FIXED_BBOX -386 -1040 94 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 10 val 44.56 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
