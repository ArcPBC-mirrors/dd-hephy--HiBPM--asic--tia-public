magic
tech sky130A
magscale 1 2
timestamp 1683130998
<< pwell >>
rect -812 -1955 812 1955
<< nmoslvt >>
rect -616 1345 -416 1745
rect -358 1345 -158 1745
rect -100 1345 100 1745
rect 158 1345 358 1745
rect 416 1345 616 1745
rect -616 727 -416 1127
rect -358 727 -158 1127
rect -100 727 100 1127
rect 158 727 358 1127
rect 416 727 616 1127
rect -616 109 -416 509
rect -358 109 -158 509
rect -100 109 100 509
rect 158 109 358 509
rect 416 109 616 509
rect -616 -509 -416 -109
rect -358 -509 -158 -109
rect -100 -509 100 -109
rect 158 -509 358 -109
rect 416 -509 616 -109
rect -616 -1127 -416 -727
rect -358 -1127 -158 -727
rect -100 -1127 100 -727
rect 158 -1127 358 -727
rect 416 -1127 616 -727
rect -616 -1745 -416 -1345
rect -358 -1745 -158 -1345
rect -100 -1745 100 -1345
rect 158 -1745 358 -1345
rect 416 -1745 616 -1345
<< ndiff >>
rect -674 1733 -616 1745
rect -674 1357 -662 1733
rect -628 1357 -616 1733
rect -674 1345 -616 1357
rect -416 1733 -358 1745
rect -416 1357 -404 1733
rect -370 1357 -358 1733
rect -416 1345 -358 1357
rect -158 1733 -100 1745
rect -158 1357 -146 1733
rect -112 1357 -100 1733
rect -158 1345 -100 1357
rect 100 1733 158 1745
rect 100 1357 112 1733
rect 146 1357 158 1733
rect 100 1345 158 1357
rect 358 1733 416 1745
rect 358 1357 370 1733
rect 404 1357 416 1733
rect 358 1345 416 1357
rect 616 1733 674 1745
rect 616 1357 628 1733
rect 662 1357 674 1733
rect 616 1345 674 1357
rect -674 1115 -616 1127
rect -674 739 -662 1115
rect -628 739 -616 1115
rect -674 727 -616 739
rect -416 1115 -358 1127
rect -416 739 -404 1115
rect -370 739 -358 1115
rect -416 727 -358 739
rect -158 1115 -100 1127
rect -158 739 -146 1115
rect -112 739 -100 1115
rect -158 727 -100 739
rect 100 1115 158 1127
rect 100 739 112 1115
rect 146 739 158 1115
rect 100 727 158 739
rect 358 1115 416 1127
rect 358 739 370 1115
rect 404 739 416 1115
rect 358 727 416 739
rect 616 1115 674 1127
rect 616 739 628 1115
rect 662 739 674 1115
rect 616 727 674 739
rect -674 497 -616 509
rect -674 121 -662 497
rect -628 121 -616 497
rect -674 109 -616 121
rect -416 497 -358 509
rect -416 121 -404 497
rect -370 121 -358 497
rect -416 109 -358 121
rect -158 497 -100 509
rect -158 121 -146 497
rect -112 121 -100 497
rect -158 109 -100 121
rect 100 497 158 509
rect 100 121 112 497
rect 146 121 158 497
rect 100 109 158 121
rect 358 497 416 509
rect 358 121 370 497
rect 404 121 416 497
rect 358 109 416 121
rect 616 497 674 509
rect 616 121 628 497
rect 662 121 674 497
rect 616 109 674 121
rect -674 -121 -616 -109
rect -674 -497 -662 -121
rect -628 -497 -616 -121
rect -674 -509 -616 -497
rect -416 -121 -358 -109
rect -416 -497 -404 -121
rect -370 -497 -358 -121
rect -416 -509 -358 -497
rect -158 -121 -100 -109
rect -158 -497 -146 -121
rect -112 -497 -100 -121
rect -158 -509 -100 -497
rect 100 -121 158 -109
rect 100 -497 112 -121
rect 146 -497 158 -121
rect 100 -509 158 -497
rect 358 -121 416 -109
rect 358 -497 370 -121
rect 404 -497 416 -121
rect 358 -509 416 -497
rect 616 -121 674 -109
rect 616 -497 628 -121
rect 662 -497 674 -121
rect 616 -509 674 -497
rect -674 -739 -616 -727
rect -674 -1115 -662 -739
rect -628 -1115 -616 -739
rect -674 -1127 -616 -1115
rect -416 -739 -358 -727
rect -416 -1115 -404 -739
rect -370 -1115 -358 -739
rect -416 -1127 -358 -1115
rect -158 -739 -100 -727
rect -158 -1115 -146 -739
rect -112 -1115 -100 -739
rect -158 -1127 -100 -1115
rect 100 -739 158 -727
rect 100 -1115 112 -739
rect 146 -1115 158 -739
rect 100 -1127 158 -1115
rect 358 -739 416 -727
rect 358 -1115 370 -739
rect 404 -1115 416 -739
rect 358 -1127 416 -1115
rect 616 -739 674 -727
rect 616 -1115 628 -739
rect 662 -1115 674 -739
rect 616 -1127 674 -1115
rect -674 -1357 -616 -1345
rect -674 -1733 -662 -1357
rect -628 -1733 -616 -1357
rect -674 -1745 -616 -1733
rect -416 -1357 -358 -1345
rect -416 -1733 -404 -1357
rect -370 -1733 -358 -1357
rect -416 -1745 -358 -1733
rect -158 -1357 -100 -1345
rect -158 -1733 -146 -1357
rect -112 -1733 -100 -1357
rect -158 -1745 -100 -1733
rect 100 -1357 158 -1345
rect 100 -1733 112 -1357
rect 146 -1733 158 -1357
rect 100 -1745 158 -1733
rect 358 -1357 416 -1345
rect 358 -1733 370 -1357
rect 404 -1733 416 -1357
rect 358 -1745 416 -1733
rect 616 -1357 674 -1345
rect 616 -1733 628 -1357
rect 662 -1733 674 -1357
rect 616 -1745 674 -1733
<< ndiffc >>
rect -662 1357 -628 1733
rect -404 1357 -370 1733
rect -146 1357 -112 1733
rect 112 1357 146 1733
rect 370 1357 404 1733
rect 628 1357 662 1733
rect -662 739 -628 1115
rect -404 739 -370 1115
rect -146 739 -112 1115
rect 112 739 146 1115
rect 370 739 404 1115
rect 628 739 662 1115
rect -662 121 -628 497
rect -404 121 -370 497
rect -146 121 -112 497
rect 112 121 146 497
rect 370 121 404 497
rect 628 121 662 497
rect -662 -497 -628 -121
rect -404 -497 -370 -121
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect 370 -497 404 -121
rect 628 -497 662 -121
rect -662 -1115 -628 -739
rect -404 -1115 -370 -739
rect -146 -1115 -112 -739
rect 112 -1115 146 -739
rect 370 -1115 404 -739
rect 628 -1115 662 -739
rect -662 -1733 -628 -1357
rect -404 -1733 -370 -1357
rect -146 -1733 -112 -1357
rect 112 -1733 146 -1357
rect 370 -1733 404 -1357
rect 628 -1733 662 -1357
<< psubdiff >>
rect -776 1885 -680 1919
rect 680 1885 776 1919
rect -776 1823 -742 1885
rect 742 1823 776 1885
rect -776 -1885 -742 -1823
rect 742 -1885 776 -1823
rect -776 -1919 -680 -1885
rect 680 -1919 776 -1885
<< psubdiffcont >>
rect -680 1885 680 1919
rect -776 -1823 -742 1823
rect 742 -1823 776 1823
rect -680 -1919 680 -1885
<< poly >>
rect -616 1817 -416 1833
rect -616 1783 -600 1817
rect -432 1783 -416 1817
rect -616 1745 -416 1783
rect -358 1817 -158 1833
rect -358 1783 -342 1817
rect -174 1783 -158 1817
rect -358 1745 -158 1783
rect -100 1817 100 1833
rect -100 1783 -84 1817
rect 84 1783 100 1817
rect -100 1745 100 1783
rect 158 1817 358 1833
rect 158 1783 174 1817
rect 342 1783 358 1817
rect 158 1745 358 1783
rect 416 1817 616 1833
rect 416 1783 432 1817
rect 600 1783 616 1817
rect 416 1745 616 1783
rect -616 1307 -416 1345
rect -616 1273 -600 1307
rect -432 1273 -416 1307
rect -616 1257 -416 1273
rect -358 1307 -158 1345
rect -358 1273 -342 1307
rect -174 1273 -158 1307
rect -358 1257 -158 1273
rect -100 1307 100 1345
rect -100 1273 -84 1307
rect 84 1273 100 1307
rect -100 1257 100 1273
rect 158 1307 358 1345
rect 158 1273 174 1307
rect 342 1273 358 1307
rect 158 1257 358 1273
rect 416 1307 616 1345
rect 416 1273 432 1307
rect 600 1273 616 1307
rect 416 1257 616 1273
rect -616 1199 -416 1215
rect -616 1165 -600 1199
rect -432 1165 -416 1199
rect -616 1127 -416 1165
rect -358 1199 -158 1215
rect -358 1165 -342 1199
rect -174 1165 -158 1199
rect -358 1127 -158 1165
rect -100 1199 100 1215
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -100 1127 100 1165
rect 158 1199 358 1215
rect 158 1165 174 1199
rect 342 1165 358 1199
rect 158 1127 358 1165
rect 416 1199 616 1215
rect 416 1165 432 1199
rect 600 1165 616 1199
rect 416 1127 616 1165
rect -616 689 -416 727
rect -616 655 -600 689
rect -432 655 -416 689
rect -616 639 -416 655
rect -358 689 -158 727
rect -358 655 -342 689
rect -174 655 -158 689
rect -358 639 -158 655
rect -100 689 100 727
rect -100 655 -84 689
rect 84 655 100 689
rect -100 639 100 655
rect 158 689 358 727
rect 158 655 174 689
rect 342 655 358 689
rect 158 639 358 655
rect 416 689 616 727
rect 416 655 432 689
rect 600 655 616 689
rect 416 639 616 655
rect -616 581 -416 597
rect -616 547 -600 581
rect -432 547 -416 581
rect -616 509 -416 547
rect -358 581 -158 597
rect -358 547 -342 581
rect -174 547 -158 581
rect -358 509 -158 547
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 509 100 547
rect 158 581 358 597
rect 158 547 174 581
rect 342 547 358 581
rect 158 509 358 547
rect 416 581 616 597
rect 416 547 432 581
rect 600 547 616 581
rect 416 509 616 547
rect -616 71 -416 109
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 109
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 109
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 109
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect -616 -37 -416 -21
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -616 -109 -416 -71
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -109 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -109 358 -71
rect 416 -37 616 -21
rect 416 -71 432 -37
rect 600 -71 616 -37
rect 416 -109 616 -71
rect -616 -547 -416 -509
rect -616 -581 -600 -547
rect -432 -581 -416 -547
rect -616 -597 -416 -581
rect -358 -547 -158 -509
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -358 -597 -158 -581
rect -100 -547 100 -509
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
rect 158 -547 358 -509
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 158 -597 358 -581
rect 416 -547 616 -509
rect 416 -581 432 -547
rect 600 -581 616 -547
rect 416 -597 616 -581
rect -616 -655 -416 -639
rect -616 -689 -600 -655
rect -432 -689 -416 -655
rect -616 -727 -416 -689
rect -358 -655 -158 -639
rect -358 -689 -342 -655
rect -174 -689 -158 -655
rect -358 -727 -158 -689
rect -100 -655 100 -639
rect -100 -689 -84 -655
rect 84 -689 100 -655
rect -100 -727 100 -689
rect 158 -655 358 -639
rect 158 -689 174 -655
rect 342 -689 358 -655
rect 158 -727 358 -689
rect 416 -655 616 -639
rect 416 -689 432 -655
rect 600 -689 616 -655
rect 416 -727 616 -689
rect -616 -1165 -416 -1127
rect -616 -1199 -600 -1165
rect -432 -1199 -416 -1165
rect -616 -1215 -416 -1199
rect -358 -1165 -158 -1127
rect -358 -1199 -342 -1165
rect -174 -1199 -158 -1165
rect -358 -1215 -158 -1199
rect -100 -1165 100 -1127
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1215 100 -1199
rect 158 -1165 358 -1127
rect 158 -1199 174 -1165
rect 342 -1199 358 -1165
rect 158 -1215 358 -1199
rect 416 -1165 616 -1127
rect 416 -1199 432 -1165
rect 600 -1199 616 -1165
rect 416 -1215 616 -1199
rect -616 -1273 -416 -1257
rect -616 -1307 -600 -1273
rect -432 -1307 -416 -1273
rect -616 -1345 -416 -1307
rect -358 -1273 -158 -1257
rect -358 -1307 -342 -1273
rect -174 -1307 -158 -1273
rect -358 -1345 -158 -1307
rect -100 -1273 100 -1257
rect -100 -1307 -84 -1273
rect 84 -1307 100 -1273
rect -100 -1345 100 -1307
rect 158 -1273 358 -1257
rect 158 -1307 174 -1273
rect 342 -1307 358 -1273
rect 158 -1345 358 -1307
rect 416 -1273 616 -1257
rect 416 -1307 432 -1273
rect 600 -1307 616 -1273
rect 416 -1345 616 -1307
rect -616 -1783 -416 -1745
rect -616 -1817 -600 -1783
rect -432 -1817 -416 -1783
rect -616 -1833 -416 -1817
rect -358 -1783 -158 -1745
rect -358 -1817 -342 -1783
rect -174 -1817 -158 -1783
rect -358 -1833 -158 -1817
rect -100 -1783 100 -1745
rect -100 -1817 -84 -1783
rect 84 -1817 100 -1783
rect -100 -1833 100 -1817
rect 158 -1783 358 -1745
rect 158 -1817 174 -1783
rect 342 -1817 358 -1783
rect 158 -1833 358 -1817
rect 416 -1783 616 -1745
rect 416 -1817 432 -1783
rect 600 -1817 616 -1783
rect 416 -1833 616 -1817
<< polycont >>
rect -600 1783 -432 1817
rect -342 1783 -174 1817
rect -84 1783 84 1817
rect 174 1783 342 1817
rect 432 1783 600 1817
rect -600 1273 -432 1307
rect -342 1273 -174 1307
rect -84 1273 84 1307
rect 174 1273 342 1307
rect 432 1273 600 1307
rect -600 1165 -432 1199
rect -342 1165 -174 1199
rect -84 1165 84 1199
rect 174 1165 342 1199
rect 432 1165 600 1199
rect -600 655 -432 689
rect -342 655 -174 689
rect -84 655 84 689
rect 174 655 342 689
rect 432 655 600 689
rect -600 547 -432 581
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect 432 547 600 581
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -600 -581 -432 -547
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
rect 432 -581 600 -547
rect -600 -689 -432 -655
rect -342 -689 -174 -655
rect -84 -689 84 -655
rect 174 -689 342 -655
rect 432 -689 600 -655
rect -600 -1199 -432 -1165
rect -342 -1199 -174 -1165
rect -84 -1199 84 -1165
rect 174 -1199 342 -1165
rect 432 -1199 600 -1165
rect -600 -1307 -432 -1273
rect -342 -1307 -174 -1273
rect -84 -1307 84 -1273
rect 174 -1307 342 -1273
rect 432 -1307 600 -1273
rect -600 -1817 -432 -1783
rect -342 -1817 -174 -1783
rect -84 -1817 84 -1783
rect 174 -1817 342 -1783
rect 432 -1817 600 -1783
<< locali >>
rect -776 1885 -680 1919
rect 680 1885 776 1919
rect -776 1823 -742 1885
rect 742 1823 776 1885
rect -616 1783 -600 1817
rect -432 1783 -416 1817
rect -358 1783 -342 1817
rect -174 1783 -158 1817
rect -100 1783 -84 1817
rect 84 1783 100 1817
rect 158 1783 174 1817
rect 342 1783 358 1817
rect 416 1783 432 1817
rect 600 1783 616 1817
rect -662 1733 -628 1749
rect -662 1341 -628 1357
rect -404 1733 -370 1749
rect -404 1341 -370 1357
rect -146 1733 -112 1749
rect -146 1341 -112 1357
rect 112 1733 146 1749
rect 112 1341 146 1357
rect 370 1733 404 1749
rect 370 1341 404 1357
rect 628 1733 662 1749
rect 628 1341 662 1357
rect -616 1273 -600 1307
rect -432 1273 -416 1307
rect -358 1273 -342 1307
rect -174 1273 -158 1307
rect -100 1273 -84 1307
rect 84 1273 100 1307
rect 158 1273 174 1307
rect 342 1273 358 1307
rect 416 1273 432 1307
rect 600 1273 616 1307
rect -616 1165 -600 1199
rect -432 1165 -416 1199
rect -358 1165 -342 1199
rect -174 1165 -158 1199
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect 158 1165 174 1199
rect 342 1165 358 1199
rect 416 1165 432 1199
rect 600 1165 616 1199
rect -662 1115 -628 1131
rect -662 723 -628 739
rect -404 1115 -370 1131
rect -404 723 -370 739
rect -146 1115 -112 1131
rect -146 723 -112 739
rect 112 1115 146 1131
rect 112 723 146 739
rect 370 1115 404 1131
rect 370 723 404 739
rect 628 1115 662 1131
rect 628 723 662 739
rect -616 655 -600 689
rect -432 655 -416 689
rect -358 655 -342 689
rect -174 655 -158 689
rect -100 655 -84 689
rect 84 655 100 689
rect 158 655 174 689
rect 342 655 358 689
rect 416 655 432 689
rect 600 655 616 689
rect -616 547 -600 581
rect -432 547 -416 581
rect -358 547 -342 581
rect -174 547 -158 581
rect -100 547 -84 581
rect 84 547 100 581
rect 158 547 174 581
rect 342 547 358 581
rect 416 547 432 581
rect 600 547 616 581
rect -662 497 -628 513
rect -662 105 -628 121
rect -404 497 -370 513
rect -404 105 -370 121
rect -146 497 -112 513
rect -146 105 -112 121
rect 112 497 146 513
rect 112 105 146 121
rect 370 497 404 513
rect 370 105 404 121
rect 628 497 662 513
rect 628 105 662 121
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 416 -71 432 -37
rect 600 -71 616 -37
rect -662 -121 -628 -105
rect -662 -513 -628 -497
rect -404 -121 -370 -105
rect -404 -513 -370 -497
rect -146 -121 -112 -105
rect -146 -513 -112 -497
rect 112 -121 146 -105
rect 112 -513 146 -497
rect 370 -121 404 -105
rect 370 -513 404 -497
rect 628 -121 662 -105
rect 628 -513 662 -497
rect -616 -581 -600 -547
rect -432 -581 -416 -547
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 416 -581 432 -547
rect 600 -581 616 -547
rect -616 -689 -600 -655
rect -432 -689 -416 -655
rect -358 -689 -342 -655
rect -174 -689 -158 -655
rect -100 -689 -84 -655
rect 84 -689 100 -655
rect 158 -689 174 -655
rect 342 -689 358 -655
rect 416 -689 432 -655
rect 600 -689 616 -655
rect -662 -739 -628 -723
rect -662 -1131 -628 -1115
rect -404 -739 -370 -723
rect -404 -1131 -370 -1115
rect -146 -739 -112 -723
rect -146 -1131 -112 -1115
rect 112 -739 146 -723
rect 112 -1131 146 -1115
rect 370 -739 404 -723
rect 370 -1131 404 -1115
rect 628 -739 662 -723
rect 628 -1131 662 -1115
rect -616 -1199 -600 -1165
rect -432 -1199 -416 -1165
rect -358 -1199 -342 -1165
rect -174 -1199 -158 -1165
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect 158 -1199 174 -1165
rect 342 -1199 358 -1165
rect 416 -1199 432 -1165
rect 600 -1199 616 -1165
rect -616 -1307 -600 -1273
rect -432 -1307 -416 -1273
rect -358 -1307 -342 -1273
rect -174 -1307 -158 -1273
rect -100 -1307 -84 -1273
rect 84 -1307 100 -1273
rect 158 -1307 174 -1273
rect 342 -1307 358 -1273
rect 416 -1307 432 -1273
rect 600 -1307 616 -1273
rect -662 -1357 -628 -1341
rect -662 -1749 -628 -1733
rect -404 -1357 -370 -1341
rect -404 -1749 -370 -1733
rect -146 -1357 -112 -1341
rect -146 -1749 -112 -1733
rect 112 -1357 146 -1341
rect 112 -1749 146 -1733
rect 370 -1357 404 -1341
rect 370 -1749 404 -1733
rect 628 -1357 662 -1341
rect 628 -1749 662 -1733
rect -616 -1817 -600 -1783
rect -432 -1817 -416 -1783
rect -358 -1817 -342 -1783
rect -174 -1817 -158 -1783
rect -100 -1817 -84 -1783
rect 84 -1817 100 -1783
rect 158 -1817 174 -1783
rect 342 -1817 358 -1783
rect 416 -1817 432 -1783
rect 600 -1817 616 -1783
rect -776 -1885 -742 -1823
rect 742 -1885 776 -1823
rect -776 -1919 -680 -1885
rect 680 -1919 776 -1885
<< viali >>
rect -600 1783 -432 1817
rect -342 1783 -174 1817
rect -84 1783 84 1817
rect 174 1783 342 1817
rect 432 1783 600 1817
rect -662 1357 -628 1733
rect -404 1357 -370 1733
rect -146 1357 -112 1733
rect 112 1357 146 1733
rect 370 1357 404 1733
rect 628 1357 662 1733
rect -600 1273 -432 1307
rect -342 1273 -174 1307
rect -84 1273 84 1307
rect 174 1273 342 1307
rect 432 1273 600 1307
rect -600 1165 -432 1199
rect -342 1165 -174 1199
rect -84 1165 84 1199
rect 174 1165 342 1199
rect 432 1165 600 1199
rect -662 739 -628 1115
rect -404 739 -370 1115
rect -146 739 -112 1115
rect 112 739 146 1115
rect 370 739 404 1115
rect 628 739 662 1115
rect -600 655 -432 689
rect -342 655 -174 689
rect -84 655 84 689
rect 174 655 342 689
rect 432 655 600 689
rect -600 547 -432 581
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect 432 547 600 581
rect -662 121 -628 497
rect -404 121 -370 497
rect -146 121 -112 497
rect 112 121 146 497
rect 370 121 404 497
rect 628 121 662 497
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -662 -497 -628 -121
rect -404 -497 -370 -121
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect 370 -497 404 -121
rect 628 -497 662 -121
rect -600 -581 -432 -547
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
rect 432 -581 600 -547
rect -600 -689 -432 -655
rect -342 -689 -174 -655
rect -84 -689 84 -655
rect 174 -689 342 -655
rect 432 -689 600 -655
rect -662 -1115 -628 -739
rect -404 -1115 -370 -739
rect -146 -1115 -112 -739
rect 112 -1115 146 -739
rect 370 -1115 404 -739
rect 628 -1115 662 -739
rect -600 -1199 -432 -1165
rect -342 -1199 -174 -1165
rect -84 -1199 84 -1165
rect 174 -1199 342 -1165
rect 432 -1199 600 -1165
rect -600 -1307 -432 -1273
rect -342 -1307 -174 -1273
rect -84 -1307 84 -1273
rect 174 -1307 342 -1273
rect 432 -1307 600 -1273
rect -662 -1733 -628 -1357
rect -404 -1733 -370 -1357
rect -146 -1733 -112 -1357
rect 112 -1733 146 -1357
rect 370 -1733 404 -1357
rect 628 -1733 662 -1357
rect -600 -1817 -432 -1783
rect -342 -1817 -174 -1783
rect -84 -1817 84 -1783
rect 174 -1817 342 -1783
rect 432 -1817 600 -1783
<< metal1 >>
rect -612 1817 -420 1823
rect -612 1783 -600 1817
rect -432 1783 -420 1817
rect -612 1777 -420 1783
rect -354 1817 -162 1823
rect -354 1783 -342 1817
rect -174 1783 -162 1817
rect -354 1777 -162 1783
rect -96 1817 96 1823
rect -96 1783 -84 1817
rect 84 1783 96 1817
rect -96 1777 96 1783
rect 162 1817 354 1823
rect 162 1783 174 1817
rect 342 1783 354 1817
rect 162 1777 354 1783
rect 420 1817 612 1823
rect 420 1783 432 1817
rect 600 1783 612 1817
rect 420 1777 612 1783
rect -668 1733 -622 1745
rect -668 1357 -662 1733
rect -628 1357 -622 1733
rect -668 1345 -622 1357
rect -410 1733 -364 1745
rect -410 1357 -404 1733
rect -370 1357 -364 1733
rect -410 1345 -364 1357
rect -152 1733 -106 1745
rect -152 1357 -146 1733
rect -112 1357 -106 1733
rect -152 1345 -106 1357
rect 106 1733 152 1745
rect 106 1357 112 1733
rect 146 1357 152 1733
rect 106 1345 152 1357
rect 364 1733 410 1745
rect 364 1357 370 1733
rect 404 1357 410 1733
rect 364 1345 410 1357
rect 622 1733 668 1745
rect 622 1357 628 1733
rect 662 1357 668 1733
rect 622 1345 668 1357
rect -612 1307 -420 1313
rect -612 1273 -600 1307
rect -432 1273 -420 1307
rect -612 1267 -420 1273
rect -354 1307 -162 1313
rect -354 1273 -342 1307
rect -174 1273 -162 1307
rect -354 1267 -162 1273
rect -96 1307 96 1313
rect -96 1273 -84 1307
rect 84 1273 96 1307
rect -96 1267 96 1273
rect 162 1307 354 1313
rect 162 1273 174 1307
rect 342 1273 354 1307
rect 162 1267 354 1273
rect 420 1307 612 1313
rect 420 1273 432 1307
rect 600 1273 612 1307
rect 420 1267 612 1273
rect -612 1199 -420 1205
rect -612 1165 -600 1199
rect -432 1165 -420 1199
rect -612 1159 -420 1165
rect -354 1199 -162 1205
rect -354 1165 -342 1199
rect -174 1165 -162 1199
rect -354 1159 -162 1165
rect -96 1199 96 1205
rect -96 1165 -84 1199
rect 84 1165 96 1199
rect -96 1159 96 1165
rect 162 1199 354 1205
rect 162 1165 174 1199
rect 342 1165 354 1199
rect 162 1159 354 1165
rect 420 1199 612 1205
rect 420 1165 432 1199
rect 600 1165 612 1199
rect 420 1159 612 1165
rect -668 1115 -622 1127
rect -668 739 -662 1115
rect -628 739 -622 1115
rect -668 727 -622 739
rect -410 1115 -364 1127
rect -410 739 -404 1115
rect -370 739 -364 1115
rect -410 727 -364 739
rect -152 1115 -106 1127
rect -152 739 -146 1115
rect -112 739 -106 1115
rect -152 727 -106 739
rect 106 1115 152 1127
rect 106 739 112 1115
rect 146 739 152 1115
rect 106 727 152 739
rect 364 1115 410 1127
rect 364 739 370 1115
rect 404 739 410 1115
rect 364 727 410 739
rect 622 1115 668 1127
rect 622 739 628 1115
rect 662 739 668 1115
rect 622 727 668 739
rect -612 689 -420 695
rect -612 655 -600 689
rect -432 655 -420 689
rect -612 649 -420 655
rect -354 689 -162 695
rect -354 655 -342 689
rect -174 655 -162 689
rect -354 649 -162 655
rect -96 689 96 695
rect -96 655 -84 689
rect 84 655 96 689
rect -96 649 96 655
rect 162 689 354 695
rect 162 655 174 689
rect 342 655 354 689
rect 162 649 354 655
rect 420 689 612 695
rect 420 655 432 689
rect 600 655 612 689
rect 420 649 612 655
rect -612 581 -420 587
rect -612 547 -600 581
rect -432 547 -420 581
rect -612 541 -420 547
rect -354 581 -162 587
rect -354 547 -342 581
rect -174 547 -162 581
rect -354 541 -162 547
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect 162 581 354 587
rect 162 547 174 581
rect 342 547 354 581
rect 162 541 354 547
rect 420 581 612 587
rect 420 547 432 581
rect 600 547 612 581
rect 420 541 612 547
rect -668 497 -622 509
rect -668 121 -662 497
rect -628 121 -622 497
rect -668 109 -622 121
rect -410 497 -364 509
rect -410 121 -404 497
rect -370 121 -364 497
rect -410 109 -364 121
rect -152 497 -106 509
rect -152 121 -146 497
rect -112 121 -106 497
rect -152 109 -106 121
rect 106 497 152 509
rect 106 121 112 497
rect 146 121 152 497
rect 106 109 152 121
rect 364 497 410 509
rect 364 121 370 497
rect 404 121 410 497
rect 364 109 410 121
rect 622 497 668 509
rect 622 121 628 497
rect 662 121 668 497
rect 622 109 668 121
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect -612 -37 -420 -31
rect -612 -71 -600 -37
rect -432 -71 -420 -37
rect -612 -77 -420 -71
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect 420 -37 612 -31
rect 420 -71 432 -37
rect 600 -71 612 -37
rect 420 -77 612 -71
rect -668 -121 -622 -109
rect -668 -497 -662 -121
rect -628 -497 -622 -121
rect -668 -509 -622 -497
rect -410 -121 -364 -109
rect -410 -497 -404 -121
rect -370 -497 -364 -121
rect -410 -509 -364 -497
rect -152 -121 -106 -109
rect -152 -497 -146 -121
rect -112 -497 -106 -121
rect -152 -509 -106 -497
rect 106 -121 152 -109
rect 106 -497 112 -121
rect 146 -497 152 -121
rect 106 -509 152 -497
rect 364 -121 410 -109
rect 364 -497 370 -121
rect 404 -497 410 -121
rect 364 -509 410 -497
rect 622 -121 668 -109
rect 622 -497 628 -121
rect 662 -497 668 -121
rect 622 -509 668 -497
rect -612 -547 -420 -541
rect -612 -581 -600 -547
rect -432 -581 -420 -547
rect -612 -587 -420 -581
rect -354 -547 -162 -541
rect -354 -581 -342 -547
rect -174 -581 -162 -547
rect -354 -587 -162 -581
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
rect 162 -547 354 -541
rect 162 -581 174 -547
rect 342 -581 354 -547
rect 162 -587 354 -581
rect 420 -547 612 -541
rect 420 -581 432 -547
rect 600 -581 612 -547
rect 420 -587 612 -581
rect -612 -655 -420 -649
rect -612 -689 -600 -655
rect -432 -689 -420 -655
rect -612 -695 -420 -689
rect -354 -655 -162 -649
rect -354 -689 -342 -655
rect -174 -689 -162 -655
rect -354 -695 -162 -689
rect -96 -655 96 -649
rect -96 -689 -84 -655
rect 84 -689 96 -655
rect -96 -695 96 -689
rect 162 -655 354 -649
rect 162 -689 174 -655
rect 342 -689 354 -655
rect 162 -695 354 -689
rect 420 -655 612 -649
rect 420 -689 432 -655
rect 600 -689 612 -655
rect 420 -695 612 -689
rect -668 -739 -622 -727
rect -668 -1115 -662 -739
rect -628 -1115 -622 -739
rect -668 -1127 -622 -1115
rect -410 -739 -364 -727
rect -410 -1115 -404 -739
rect -370 -1115 -364 -739
rect -410 -1127 -364 -1115
rect -152 -739 -106 -727
rect -152 -1115 -146 -739
rect -112 -1115 -106 -739
rect -152 -1127 -106 -1115
rect 106 -739 152 -727
rect 106 -1115 112 -739
rect 146 -1115 152 -739
rect 106 -1127 152 -1115
rect 364 -739 410 -727
rect 364 -1115 370 -739
rect 404 -1115 410 -739
rect 364 -1127 410 -1115
rect 622 -739 668 -727
rect 622 -1115 628 -739
rect 662 -1115 668 -739
rect 622 -1127 668 -1115
rect -612 -1165 -420 -1159
rect -612 -1199 -600 -1165
rect -432 -1199 -420 -1165
rect -612 -1205 -420 -1199
rect -354 -1165 -162 -1159
rect -354 -1199 -342 -1165
rect -174 -1199 -162 -1165
rect -354 -1205 -162 -1199
rect -96 -1165 96 -1159
rect -96 -1199 -84 -1165
rect 84 -1199 96 -1165
rect -96 -1205 96 -1199
rect 162 -1165 354 -1159
rect 162 -1199 174 -1165
rect 342 -1199 354 -1165
rect 162 -1205 354 -1199
rect 420 -1165 612 -1159
rect 420 -1199 432 -1165
rect 600 -1199 612 -1165
rect 420 -1205 612 -1199
rect -612 -1273 -420 -1267
rect -612 -1307 -600 -1273
rect -432 -1307 -420 -1273
rect -612 -1313 -420 -1307
rect -354 -1273 -162 -1267
rect -354 -1307 -342 -1273
rect -174 -1307 -162 -1273
rect -354 -1313 -162 -1307
rect -96 -1273 96 -1267
rect -96 -1307 -84 -1273
rect 84 -1307 96 -1273
rect -96 -1313 96 -1307
rect 162 -1273 354 -1267
rect 162 -1307 174 -1273
rect 342 -1307 354 -1273
rect 162 -1313 354 -1307
rect 420 -1273 612 -1267
rect 420 -1307 432 -1273
rect 600 -1307 612 -1273
rect 420 -1313 612 -1307
rect -668 -1357 -622 -1345
rect -668 -1733 -662 -1357
rect -628 -1733 -622 -1357
rect -668 -1745 -622 -1733
rect -410 -1357 -364 -1345
rect -410 -1733 -404 -1357
rect -370 -1733 -364 -1357
rect -410 -1745 -364 -1733
rect -152 -1357 -106 -1345
rect -152 -1733 -146 -1357
rect -112 -1733 -106 -1357
rect -152 -1745 -106 -1733
rect 106 -1357 152 -1345
rect 106 -1733 112 -1357
rect 146 -1733 152 -1357
rect 106 -1745 152 -1733
rect 364 -1357 410 -1345
rect 364 -1733 370 -1357
rect 404 -1733 410 -1357
rect 364 -1745 410 -1733
rect 622 -1357 668 -1345
rect 622 -1733 628 -1357
rect 662 -1733 668 -1357
rect 622 -1745 668 -1733
rect -612 -1783 -420 -1777
rect -612 -1817 -600 -1783
rect -432 -1817 -420 -1783
rect -612 -1823 -420 -1817
rect -354 -1783 -162 -1777
rect -354 -1817 -342 -1783
rect -174 -1817 -162 -1783
rect -354 -1823 -162 -1817
rect -96 -1783 96 -1777
rect -96 -1817 -84 -1783
rect 84 -1817 96 -1783
rect -96 -1823 96 -1817
rect 162 -1783 354 -1777
rect 162 -1817 174 -1783
rect 342 -1817 354 -1783
rect 162 -1823 354 -1817
rect 420 -1783 612 -1777
rect 420 -1817 432 -1783
rect 600 -1817 612 -1783
rect 420 -1823 612 -1817
<< properties >>
string FIXED_BBOX -759 -1902 759 1902
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 1 m 6 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
