magic
tech sky130A
magscale 1 2
timestamp 1684931108
<< pwell >>
rect -3709 -798 3709 798
<< psubdiff >>
rect -3673 728 -3577 762
rect 3577 728 3673 762
rect -3673 666 -3639 728
rect 3639 666 3673 728
rect -3673 -728 -3639 -666
rect 3639 -728 3673 -666
rect -3673 -762 -3577 -728
rect 3577 -762 3673 -728
<< psubdiffcont >>
rect -3577 728 3577 762
rect -3673 -666 -3639 666
rect 3639 -666 3673 666
rect -3577 -762 3577 -728
<< xpolycontact >>
rect -3543 200 -3261 632
rect -3543 -632 -3261 -200
rect -3165 200 -2883 632
rect -3165 -632 -2883 -200
rect -2787 200 -2505 632
rect -2787 -632 -2505 -200
rect -2409 200 -2127 632
rect -2409 -632 -2127 -200
rect -2031 200 -1749 632
rect -2031 -632 -1749 -200
rect -1653 200 -1371 632
rect -1653 -632 -1371 -200
rect -1275 200 -993 632
rect -1275 -632 -993 -200
rect -897 200 -615 632
rect -897 -632 -615 -200
rect -519 200 -237 632
rect -519 -632 -237 -200
rect -141 200 141 632
rect -141 -632 141 -200
rect 237 200 519 632
rect 237 -632 519 -200
rect 615 200 897 632
rect 615 -632 897 -200
rect 993 200 1275 632
rect 993 -632 1275 -200
rect 1371 200 1653 632
rect 1371 -632 1653 -200
rect 1749 200 2031 632
rect 1749 -632 2031 -200
rect 2127 200 2409 632
rect 2127 -632 2409 -200
rect 2505 200 2787 632
rect 2505 -632 2787 -200
rect 2883 200 3165 632
rect 2883 -632 3165 -200
rect 3261 200 3543 632
rect 3261 -632 3543 -200
<< ppolyres >>
rect -3543 -200 -3261 200
rect -3165 -200 -2883 200
rect -2787 -200 -2505 200
rect -2409 -200 -2127 200
rect -2031 -200 -1749 200
rect -1653 -200 -1371 200
rect -1275 -200 -993 200
rect -897 -200 -615 200
rect -519 -200 -237 200
rect -141 -200 141 200
rect 237 -200 519 200
rect 615 -200 897 200
rect 993 -200 1275 200
rect 1371 -200 1653 200
rect 1749 -200 2031 200
rect 2127 -200 2409 200
rect 2505 -200 2787 200
rect 2883 -200 3165 200
rect 3261 -200 3543 200
<< locali >>
rect -3673 728 -3577 762
rect 3577 728 3673 762
rect -3673 666 -3639 728
rect 3639 666 3673 728
rect -3673 -728 -3639 -666
rect 3639 -728 3673 -666
rect -3673 -762 -3577 -728
rect 3577 -762 3673 -728
<< viali >>
rect -3527 217 -3277 614
rect -3149 217 -2899 614
rect -2771 217 -2521 614
rect -2393 217 -2143 614
rect -2015 217 -1765 614
rect -1637 217 -1387 614
rect -1259 217 -1009 614
rect -881 217 -631 614
rect -503 217 -253 614
rect -125 217 125 614
rect 253 217 503 614
rect 631 217 881 614
rect 1009 217 1259 614
rect 1387 217 1637 614
rect 1765 217 2015 614
rect 2143 217 2393 614
rect 2521 217 2771 614
rect 2899 217 3149 614
rect 3277 217 3527 614
rect -3527 -614 -3277 -217
rect -3149 -614 -2899 -217
rect -2771 -614 -2521 -217
rect -2393 -614 -2143 -217
rect -2015 -614 -1765 -217
rect -1637 -614 -1387 -217
rect -1259 -614 -1009 -217
rect -881 -614 -631 -217
rect -503 -614 -253 -217
rect -125 -614 125 -217
rect 253 -614 503 -217
rect 631 -614 881 -217
rect 1009 -614 1259 -217
rect 1387 -614 1637 -217
rect 1765 -614 2015 -217
rect 2143 -614 2393 -217
rect 2521 -614 2771 -217
rect 2899 -614 3149 -217
rect 3277 -614 3527 -217
<< metal1 >>
rect -3533 614 -3271 626
rect -3533 217 -3527 614
rect -3277 217 -3271 614
rect -3533 205 -3271 217
rect -3155 614 -2893 626
rect -3155 217 -3149 614
rect -2899 217 -2893 614
rect -3155 205 -2893 217
rect -2777 614 -2515 626
rect -2777 217 -2771 614
rect -2521 217 -2515 614
rect -2777 205 -2515 217
rect -2399 614 -2137 626
rect -2399 217 -2393 614
rect -2143 217 -2137 614
rect -2399 205 -2137 217
rect -2021 614 -1759 626
rect -2021 217 -2015 614
rect -1765 217 -1759 614
rect -2021 205 -1759 217
rect -1643 614 -1381 626
rect -1643 217 -1637 614
rect -1387 217 -1381 614
rect -1643 205 -1381 217
rect -1265 614 -1003 626
rect -1265 217 -1259 614
rect -1009 217 -1003 614
rect -1265 205 -1003 217
rect -887 614 -625 626
rect -887 217 -881 614
rect -631 217 -625 614
rect -887 205 -625 217
rect -509 614 -247 626
rect -509 217 -503 614
rect -253 217 -247 614
rect -509 205 -247 217
rect -131 614 131 626
rect -131 217 -125 614
rect 125 217 131 614
rect -131 205 131 217
rect 247 614 509 626
rect 247 217 253 614
rect 503 217 509 614
rect 247 205 509 217
rect 625 614 887 626
rect 625 217 631 614
rect 881 217 887 614
rect 625 205 887 217
rect 1003 614 1265 626
rect 1003 217 1009 614
rect 1259 217 1265 614
rect 1003 205 1265 217
rect 1381 614 1643 626
rect 1381 217 1387 614
rect 1637 217 1643 614
rect 1381 205 1643 217
rect 1759 614 2021 626
rect 1759 217 1765 614
rect 2015 217 2021 614
rect 1759 205 2021 217
rect 2137 614 2399 626
rect 2137 217 2143 614
rect 2393 217 2399 614
rect 2137 205 2399 217
rect 2515 614 2777 626
rect 2515 217 2521 614
rect 2771 217 2777 614
rect 2515 205 2777 217
rect 2893 614 3155 626
rect 2893 217 2899 614
rect 3149 217 3155 614
rect 2893 205 3155 217
rect 3271 614 3533 626
rect 3271 217 3277 614
rect 3527 217 3533 614
rect 3271 205 3533 217
rect -3533 -217 -3271 -205
rect -3533 -614 -3527 -217
rect -3277 -614 -3271 -217
rect -3533 -626 -3271 -614
rect -3155 -217 -2893 -205
rect -3155 -614 -3149 -217
rect -2899 -614 -2893 -217
rect -3155 -626 -2893 -614
rect -2777 -217 -2515 -205
rect -2777 -614 -2771 -217
rect -2521 -614 -2515 -217
rect -2777 -626 -2515 -614
rect -2399 -217 -2137 -205
rect -2399 -614 -2393 -217
rect -2143 -614 -2137 -217
rect -2399 -626 -2137 -614
rect -2021 -217 -1759 -205
rect -2021 -614 -2015 -217
rect -1765 -614 -1759 -217
rect -2021 -626 -1759 -614
rect -1643 -217 -1381 -205
rect -1643 -614 -1637 -217
rect -1387 -614 -1381 -217
rect -1643 -626 -1381 -614
rect -1265 -217 -1003 -205
rect -1265 -614 -1259 -217
rect -1009 -614 -1003 -217
rect -1265 -626 -1003 -614
rect -887 -217 -625 -205
rect -887 -614 -881 -217
rect -631 -614 -625 -217
rect -887 -626 -625 -614
rect -509 -217 -247 -205
rect -509 -614 -503 -217
rect -253 -614 -247 -217
rect -509 -626 -247 -614
rect -131 -217 131 -205
rect -131 -614 -125 -217
rect 125 -614 131 -217
rect -131 -626 131 -614
rect 247 -217 509 -205
rect 247 -614 253 -217
rect 503 -614 509 -217
rect 247 -626 509 -614
rect 625 -217 887 -205
rect 625 -614 631 -217
rect 881 -614 887 -217
rect 625 -626 887 -614
rect 1003 -217 1265 -205
rect 1003 -614 1009 -217
rect 1259 -614 1265 -217
rect 1003 -626 1265 -614
rect 1381 -217 1643 -205
rect 1381 -614 1387 -217
rect 1637 -614 1643 -217
rect 1381 -626 1643 -614
rect 1759 -217 2021 -205
rect 1759 -614 1765 -217
rect 2015 -614 2021 -217
rect 1759 -626 2021 -614
rect 2137 -217 2399 -205
rect 2137 -614 2143 -217
rect 2393 -614 2399 -217
rect 2137 -626 2399 -614
rect 2515 -217 2777 -205
rect 2515 -614 2521 -217
rect 2771 -614 2777 -217
rect 2515 -626 2777 -614
rect 2893 -217 3155 -205
rect 2893 -614 2899 -217
rect 3149 -614 3155 -217
rect 2893 -626 3155 -614
rect 3271 -217 3533 -205
rect 3271 -614 3277 -217
rect 3527 -614 3533 -217
rect 3271 -626 3533 -614
<< res1p41 >>
rect -3545 -202 -3259 202
rect -3167 -202 -2881 202
rect -2789 -202 -2503 202
rect -2411 -202 -2125 202
rect -2033 -202 -1747 202
rect -1655 -202 -1369 202
rect -1277 -202 -991 202
rect -899 -202 -613 202
rect -521 -202 -235 202
rect -143 -202 143 202
rect 235 -202 521 202
rect 613 -202 899 202
rect 991 -202 1277 202
rect 1369 -202 1655 202
rect 1747 -202 2033 202
rect 2125 -202 2411 202
rect 2503 -202 2789 202
rect 2881 -202 3167 202
rect 3259 -202 3545 202
<< properties >>
string FIXED_BBOX -3656 -745 3656 745
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 2.0 m 1 nx 19 wmin 1.410 lmin 0.50 rho 319.8 val 729.957 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
