magic
tech sky130A
magscale 1 2
timestamp 1684167095
<< metal1 >>
rect 236 2408 1408 2516
rect 430 2188 440 2368
rect 492 2188 502 2368
rect 946 2188 956 2368
rect 1008 2188 1018 2368
rect 170 1964 180 2144
rect 232 1964 242 2144
rect 686 1964 696 2144
rect 748 1964 758 2144
rect 1202 1964 1212 2144
rect 1264 1964 1274 2144
rect 1316 1928 1408 2408
rect 236 1768 1408 1928
rect 430 1552 440 1732
rect 492 1552 502 1732
rect 946 1552 956 1732
rect 1008 1552 1018 1732
rect 170 1328 180 1508
rect 232 1328 242 1508
rect 686 1328 696 1508
rect 748 1328 758 1508
rect 1202 1328 1212 1508
rect 1264 1328 1274 1508
rect 1316 1292 1408 1768
rect 236 1132 1408 1292
rect 430 916 440 1096
rect 492 916 502 1096
rect 946 916 956 1096
rect 1008 916 1018 1096
rect 170 692 180 872
rect 232 692 242 872
rect 686 692 696 872
rect 748 692 758 872
rect 1202 692 1212 872
rect 1264 692 1274 872
rect 1316 656 1408 1132
rect 232 496 1408 656
rect 430 280 440 460
rect 492 280 502 460
rect 946 280 956 460
rect 1008 280 1018 460
rect 170 56 180 236
rect 232 56 242 236
rect 686 56 696 236
rect 748 56 758 236
rect 1202 56 1212 236
rect 1264 56 1274 236
rect 1316 20 1408 496
rect 236 -88 1408 20
rect 1056 -220 1152 -88
rect 1316 -100 1408 -88
rect 220 -324 1152 -220
rect 266 -544 276 -364
rect 328 -544 338 -364
rect 458 -544 468 -364
rect 520 -544 530 -364
rect 650 -544 660 -364
rect 712 -544 722 -364
rect 842 -544 852 -364
rect 904 -544 914 -364
rect 170 -768 180 -588
rect 232 -768 242 -588
rect 362 -768 372 -588
rect 424 -768 434 -588
rect 554 -768 564 -588
rect 616 -768 626 -588
rect 746 -768 756 -588
rect 808 -768 818 -588
rect 938 -768 948 -588
rect 1000 -768 1010 -588
rect 1056 -804 1152 -324
rect 316 -960 1152 -804
rect 266 -1180 276 -1000
rect 328 -1180 338 -1000
rect 458 -1180 468 -1000
rect 520 -1180 530 -1000
rect 650 -1180 660 -1000
rect 712 -1180 722 -1000
rect 842 -1180 852 -1000
rect 904 -1180 914 -1000
rect 170 -1404 180 -1224
rect 232 -1404 242 -1224
rect 362 -1404 372 -1224
rect 424 -1404 434 -1224
rect 554 -1404 564 -1224
rect 616 -1404 626 -1224
rect 746 -1404 756 -1224
rect 808 -1404 818 -1224
rect 938 -1404 948 -1224
rect 1000 -1404 1010 -1224
rect 1056 -1440 1152 -960
rect 216 -1552 1152 -1440
<< via1 >>
rect 440 2188 492 2368
rect 956 2188 1008 2368
rect 180 1964 232 2144
rect 696 1964 748 2144
rect 1212 1964 1264 2144
rect 440 1552 492 1732
rect 956 1552 1008 1732
rect 180 1328 232 1508
rect 696 1328 748 1508
rect 1212 1328 1264 1508
rect 440 916 492 1096
rect 956 916 1008 1096
rect 180 692 232 872
rect 696 692 748 872
rect 1212 692 1264 872
rect 440 280 492 460
rect 956 280 1008 460
rect 180 56 232 236
rect 696 56 748 236
rect 1212 56 1264 236
rect 276 -544 328 -364
rect 468 -544 520 -364
rect 660 -544 712 -364
rect 852 -544 904 -364
rect 180 -768 232 -588
rect 372 -768 424 -588
rect 564 -768 616 -588
rect 756 -768 808 -588
rect 948 -768 1000 -588
rect 276 -1180 328 -1000
rect 468 -1180 520 -1000
rect 660 -1180 712 -1000
rect 852 -1180 904 -1000
rect 180 -1404 232 -1224
rect 372 -1404 424 -1224
rect 564 -1404 616 -1224
rect 756 -1404 808 -1224
rect 948 -1404 1000 -1224
<< metal2 >>
rect 100 2456 1004 2540
rect 100 2208 124 2456
rect 676 2378 1004 2456
rect 676 2368 1008 2378
rect 676 2208 956 2368
rect 100 2188 440 2208
rect 492 2188 956 2208
rect 440 2178 492 2188
rect 956 2178 1008 2188
rect 180 2144 232 2154
rect 696 2144 748 2154
rect 1212 2144 1264 2154
rect 232 1964 696 2144
rect 748 2132 1212 2144
rect 1264 2132 1344 2144
rect 748 1964 772 2132
rect 180 1880 772 1964
rect 1332 1880 1344 2132
rect 180 1860 1344 1880
rect 180 1826 1008 1832
rect 124 1816 1008 1826
rect 676 1732 1008 1816
rect 676 1568 956 1732
rect 124 1558 440 1568
rect 180 1552 440 1558
rect 492 1552 956 1568
rect 440 1542 492 1552
rect 956 1542 1008 1552
rect 180 1508 232 1518
rect 696 1508 748 1518
rect 1212 1508 1264 1518
rect 232 1328 696 1508
rect 748 1496 1212 1508
rect 1264 1496 1344 1508
rect 748 1328 772 1496
rect 180 1244 772 1328
rect 1332 1244 1344 1496
rect 180 1224 1344 1244
rect 180 1186 1008 1196
rect 124 1176 1008 1186
rect 676 1096 1008 1176
rect 676 928 956 1096
rect 124 918 440 928
rect 180 916 440 918
rect 492 916 956 928
rect 440 906 492 916
rect 956 906 1008 916
rect 180 872 232 882
rect 696 872 748 882
rect 1212 872 1264 882
rect 232 692 696 872
rect 748 856 1212 872
rect 1264 856 1344 872
rect 748 692 772 856
rect 180 604 772 692
rect 1332 604 1344 856
rect 180 588 1344 604
rect 184 554 1012 560
rect 124 544 1012 554
rect 676 460 1012 544
rect 676 296 956 460
rect 124 286 440 296
rect 184 280 440 286
rect 492 280 956 296
rect 1008 280 1012 460
rect 440 270 492 280
rect 956 270 1008 280
rect 180 236 232 246
rect 696 236 748 246
rect 1212 236 1264 246
rect 232 56 696 236
rect 748 220 1212 236
rect 1264 220 1348 236
rect 748 56 772 220
rect 180 -84 772 56
rect 1332 -84 1348 220
rect 180 -100 1348 -84
rect 276 -292 1348 -276
rect 276 -364 772 -292
rect 328 -544 468 -364
rect 520 -544 660 -364
rect 712 -528 772 -364
rect 1332 -528 1348 -292
rect 712 -544 852 -528
rect 904 -544 1348 -528
rect 276 -554 328 -544
rect 468 -554 520 -544
rect 660 -554 712 -544
rect 852 -554 904 -544
rect 180 -588 232 -578
rect 372 -588 424 -578
rect 564 -588 616 -578
rect 756 -588 808 -578
rect 948 -588 1000 -578
rect 64 -612 180 -588
rect 232 -612 372 -588
rect 424 -612 564 -588
rect 64 -860 80 -612
rect 616 -768 756 -588
rect 808 -768 948 -588
rect 600 -860 1000 -768
rect 64 -876 1000 -860
rect 276 -928 1348 -912
rect 276 -1000 772 -928
rect 328 -1180 468 -1000
rect 520 -1180 660 -1000
rect 712 -1164 772 -1000
rect 1332 -1164 1348 -928
rect 712 -1180 852 -1164
rect 904 -1180 1348 -1164
rect 276 -1190 328 -1180
rect 468 -1190 520 -1180
rect 660 -1190 712 -1180
rect 852 -1190 904 -1180
rect 180 -1224 232 -1214
rect 372 -1224 424 -1214
rect 564 -1224 616 -1214
rect 756 -1224 808 -1214
rect 948 -1224 1000 -1214
rect 76 -1248 180 -1224
rect 232 -1248 372 -1224
rect 424 -1248 564 -1224
rect 76 -1496 88 -1248
rect 616 -1404 756 -1224
rect 808 -1404 948 -1224
rect 1000 -1404 1012 -1224
rect 608 -1496 1012 -1404
rect 76 -1512 1012 -1496
<< via2 >>
rect 124 2368 676 2456
rect 124 2208 440 2368
rect 440 2208 492 2368
rect 492 2208 676 2368
rect 772 1964 1212 2132
rect 1212 1964 1264 2132
rect 1264 1964 1332 2132
rect 772 1880 1332 1964
rect 124 1732 676 1816
rect 124 1568 440 1732
rect 440 1568 492 1732
rect 492 1568 676 1732
rect 772 1328 1212 1496
rect 1212 1328 1264 1496
rect 1264 1328 1332 1496
rect 772 1244 1332 1328
rect 124 1096 676 1176
rect 124 928 440 1096
rect 440 928 492 1096
rect 492 928 676 1096
rect 772 692 1212 856
rect 1212 692 1264 856
rect 1264 692 1332 856
rect 772 604 1332 692
rect 124 460 676 544
rect 124 296 440 460
rect 440 296 492 460
rect 492 296 676 460
rect 772 56 1212 220
rect 1212 56 1264 220
rect 1264 56 1332 220
rect 772 -84 1332 56
rect 772 -364 1332 -292
rect 772 -528 852 -364
rect 852 -528 904 -364
rect 904 -528 1332 -364
rect 80 -768 180 -612
rect 180 -768 232 -612
rect 232 -768 372 -612
rect 372 -768 424 -612
rect 424 -768 564 -612
rect 564 -768 600 -612
rect 80 -860 600 -768
rect 772 -1000 1332 -928
rect 772 -1164 852 -1000
rect 852 -1164 904 -1000
rect 904 -1164 1332 -1000
rect 88 -1404 180 -1248
rect 180 -1404 232 -1248
rect 232 -1404 372 -1248
rect 372 -1404 424 -1248
rect 424 -1404 564 -1248
rect 564 -1404 608 -1248
rect 88 -1496 608 -1404
<< metal3 >>
rect 100 2456 692 2476
rect 100 2208 124 2456
rect 676 2208 692 2456
rect 100 1816 692 2208
rect 100 1568 124 1816
rect 676 1568 692 1816
rect 100 1176 692 1568
rect 100 928 124 1176
rect 676 928 692 1176
rect 100 544 692 928
rect 100 296 124 544
rect 676 296 692 544
rect 100 280 692 296
rect 756 2132 1348 2144
rect 756 1880 772 2132
rect 1332 1880 1348 2132
rect 756 1496 1348 1880
rect 756 1244 772 1496
rect 1332 1244 1348 1496
rect 756 856 1348 1244
rect 756 604 772 856
rect 1332 604 1348 856
rect 756 220 1348 604
rect 756 -84 772 220
rect 1332 -84 1348 220
rect 756 -292 1348 -84
rect 756 -528 772 -292
rect 1332 -528 1348 -292
rect 72 -607 628 -588
rect 70 -612 628 -607
rect 70 -860 80 -612
rect 600 -860 628 -612
rect 70 -865 628 -860
rect 72 -1248 628 -865
rect 756 -928 1348 -528
rect 756 -1164 772 -928
rect 1332 -1164 1348 -928
rect 756 -1180 1348 -1164
rect 72 -1496 88 -1248
rect 608 -1496 628 -1248
rect 72 -1620 628 -1496
use sky130_fd_pr__pfet_01v8_LXX5YL  sky130_fd_pr__pfet_01v8_LXX5YL_1
timestamp 1684167095
transform 1 0 723 0 1 1213
box -683 -1373 683 1373
use sky130_fd_pr__pfet_01v8_U4PLGH  sky130_fd_pr__pfet_01v8_U4PLGH_0
timestamp 1684167095
transform 1 0 591 0 1 -883
box -551 -737 551 737
<< end >>
