magic
tech sky130A
magscale 1 2
timestamp 1689672086
<< metal1 >>
rect 74 3208 84 3636
rect 1500 3208 1510 3636
rect 74 2376 84 2808
rect 1504 2376 1514 2808
rect 78 1840 88 2268
rect 1504 1840 1514 2268
rect 74 1004 84 1440
rect 1504 1004 1514 1440
rect 336 660 964 776
rect 286 448 296 628
rect 348 448 358 628
rect 478 448 488 628
rect 540 448 550 628
rect 670 448 680 628
rect 732 448 742 628
rect 862 448 872 628
rect 924 448 934 628
rect 382 232 392 412
rect 444 232 454 412
rect 574 232 584 412
rect 636 232 646 412
rect 766 232 776 412
rect 828 232 838 412
rect 308 84 916 200
<< via1 >>
rect 84 3208 1500 3636
rect 84 2376 1504 2808
rect 88 1840 1504 2268
rect 84 1004 1504 1440
rect 296 448 348 628
rect 488 448 540 628
rect 680 448 732 628
rect 872 448 924 628
rect 392 232 444 412
rect 584 232 636 412
rect 776 232 828 412
<< metal2 >>
rect 80 3644 1508 3654
rect 80 3198 1508 3208
rect 84 2808 1504 2818
rect 84 2368 464 2376
rect 1128 2368 1504 2376
rect 84 2366 1504 2368
rect 464 2358 1128 2366
rect 84 2278 368 2286
rect 1220 2278 1504 2286
rect 84 2276 1504 2278
rect 368 2268 1220 2276
rect 84 1830 1504 1840
rect 84 1440 1504 1450
rect 84 996 88 1004
rect 1500 996 1504 1004
rect 84 994 1504 996
rect 88 986 1500 994
rect 256 820 1308 986
rect 256 628 964 820
rect 256 464 296 628
rect 348 520 488 628
rect 348 464 388 520
rect 452 464 488 520
rect 296 438 348 448
rect 540 520 680 628
rect 540 464 580 520
rect 644 464 680 520
rect 488 438 540 448
rect 732 520 872 628
rect 732 464 772 520
rect 836 464 872 520
rect 680 438 732 448
rect 924 464 964 628
rect 872 438 924 448
rect 392 412 444 422
rect 356 340 392 396
rect 308 232 392 340
rect 584 412 636 422
rect 444 340 484 396
rect 548 340 584 396
rect 444 232 584 340
rect 776 412 828 422
rect 636 340 672 396
rect 736 340 776 396
rect 636 232 776 340
rect 828 340 868 396
rect 828 232 916 340
rect 308 60 916 232
<< via2 >>
rect 80 3636 1508 3644
rect 80 3208 84 3636
rect 84 3208 1500 3636
rect 1500 3208 1508 3636
rect 464 2376 1128 2808
rect 464 2368 1128 2376
rect 84 2268 368 2276
rect 1220 2268 1504 2276
rect 84 1840 88 2268
rect 88 1840 368 2268
rect 1220 1840 1504 2268
rect 88 1004 1500 1440
rect 88 996 1500 1004
<< metal3 >>
rect 70 3644 1518 3649
rect 70 3208 80 3644
rect 1508 3208 1518 3644
rect 70 3203 1518 3208
rect 84 2281 368 3203
rect 454 2808 1138 2813
rect 454 2368 464 2808
rect 1128 2368 1138 2808
rect 454 2363 1138 2368
rect 74 2276 378 2281
rect 74 1840 84 2276
rect 368 1840 378 2276
rect 74 1835 378 1840
rect 464 1445 748 2363
rect 840 1445 1124 2363
rect 1220 2281 1504 3203
rect 1210 2276 1514 2281
rect 1210 1840 1220 2276
rect 1504 1840 1514 2276
rect 1210 1835 1514 1840
rect 78 1440 1510 1445
rect 78 996 88 1440
rect 1500 996 1510 1440
rect 78 991 1510 996
use sky130_fd_pr__nfet_01v8_lvt_V6SMGN  sky130_fd_pr__nfet_01v8_lvt_V6SMGN_0
timestamp 1687116177
transform 1 0 611 0 1 430
box -455 -410 455 410
use sky130_fd_pr__res_xhigh_po_1p41_FUYU7G  sky130_fd_pr__res_xhigh_po_1p41_FUYU7G_0
timestamp 1689672086
transform 1 0 794 0 1 2322
box -874 -1482 874 1482
<< end >>
