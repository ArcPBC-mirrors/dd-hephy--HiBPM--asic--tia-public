magic
tech sky130A
timestamp 1689607358
<< via4 >>
rect -3600 -2850 -3450 -850
rect -2850 -2850 -2700 -850
<< metal5 >>
rect -3612 -850 -3438 -838
rect -2862 -850 -2688 -838
rect -3612 -2850 -3600 -850
rect -3450 -2850 -3400 -850
rect -2900 -2850 -2850 -850
rect -2700 -2850 -2688 -850
rect -3612 -2862 -3438 -2850
rect -2862 -2862 -2688 -2850
<< rm5 >>
rect -3400 -2850 -2900 -850
<< end >>
