magic
tech sky130A
magscale 1 2
timestamp 1683627527
<< error_p >>
rect -221 272 -163 278
rect -29 272 29 278
rect 163 272 221 278
rect -221 238 -209 272
rect -29 238 -17 272
rect 163 238 175 272
rect -221 232 -163 238
rect -29 232 29 238
rect 163 232 221 238
rect -317 -238 -259 -232
rect -125 -238 -67 -232
rect 67 -238 125 -232
rect 259 -238 317 -232
rect -317 -272 -305 -238
rect -125 -272 -113 -238
rect 67 -272 79 -238
rect 259 -272 271 -238
rect -317 -278 -259 -272
rect -125 -278 -67 -272
rect 67 -278 125 -272
rect 259 -278 317 -272
<< pwell >>
rect -503 -410 503 410
<< nmoslvt >>
rect -303 -200 -273 200
rect -207 -200 -177 200
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
rect 177 -200 207 200
rect 273 -200 303 200
<< ndiff >>
rect -365 188 -303 200
rect -365 -188 -353 188
rect -319 -188 -303 188
rect -365 -200 -303 -188
rect -273 188 -207 200
rect -273 -188 -257 188
rect -223 -188 -207 188
rect -273 -200 -207 -188
rect -177 188 -111 200
rect -177 -188 -161 188
rect -127 -188 -111 188
rect -177 -200 -111 -188
rect -81 188 -15 200
rect -81 -188 -65 188
rect -31 -188 -15 188
rect -81 -200 -15 -188
rect 15 188 81 200
rect 15 -188 31 188
rect 65 -188 81 188
rect 15 -200 81 -188
rect 111 188 177 200
rect 111 -188 127 188
rect 161 -188 177 188
rect 111 -200 177 -188
rect 207 188 273 200
rect 207 -188 223 188
rect 257 -188 273 188
rect 207 -200 273 -188
rect 303 188 365 200
rect 303 -188 319 188
rect 353 -188 365 188
rect 303 -200 365 -188
<< ndiffc >>
rect -353 -188 -319 188
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect 319 -188 353 188
<< psubdiff >>
rect -467 340 -371 374
rect 371 340 467 374
rect -467 278 -433 340
rect 433 278 467 340
rect -467 -340 -433 -278
rect 433 -340 467 -278
rect -467 -374 -371 -340
rect 371 -374 467 -340
<< psubdiffcont >>
rect -371 340 371 374
rect -467 -278 -433 278
rect 433 -278 467 278
rect -371 -374 371 -340
<< poly >>
rect -225 272 -159 288
rect -225 238 -209 272
rect -175 238 -159 272
rect -303 200 -273 226
rect -225 222 -159 238
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -207 200 -177 222
rect -111 200 -81 226
rect -33 222 33 238
rect 159 272 225 288
rect 159 238 175 272
rect 209 238 225 272
rect -15 200 15 222
rect 81 200 111 226
rect 159 222 225 238
rect 177 200 207 222
rect 273 200 303 226
rect -303 -222 -273 -200
rect -321 -238 -255 -222
rect -207 -226 -177 -200
rect -111 -222 -81 -200
rect -321 -272 -305 -238
rect -271 -272 -255 -238
rect -321 -288 -255 -272
rect -129 -238 -63 -222
rect -15 -226 15 -200
rect 81 -222 111 -200
rect -129 -272 -113 -238
rect -79 -272 -63 -238
rect -129 -288 -63 -272
rect 63 -238 129 -222
rect 177 -226 207 -200
rect 273 -222 303 -200
rect 63 -272 79 -238
rect 113 -272 129 -238
rect 63 -288 129 -272
rect 255 -238 321 -222
rect 255 -272 271 -238
rect 305 -272 321 -238
rect 255 -288 321 -272
<< polycont >>
rect -209 238 -175 272
rect -17 238 17 272
rect 175 238 209 272
rect -305 -272 -271 -238
rect -113 -272 -79 -238
rect 79 -272 113 -238
rect 271 -272 305 -238
<< locali >>
rect -467 340 -371 374
rect 371 340 467 374
rect -467 278 -433 340
rect 433 278 467 340
rect -225 238 -209 272
rect -175 238 -159 272
rect -33 238 -17 272
rect 17 238 33 272
rect 159 238 175 272
rect 209 238 225 272
rect -353 188 -319 204
rect -353 -204 -319 -188
rect -257 188 -223 204
rect -257 -204 -223 -188
rect -161 188 -127 204
rect -161 -204 -127 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 127 188 161 204
rect 127 -204 161 -188
rect 223 188 257 204
rect 223 -204 257 -188
rect 319 188 353 204
rect 319 -204 353 -188
rect -321 -272 -305 -238
rect -271 -272 -255 -238
rect -129 -272 -113 -238
rect -79 -272 -63 -238
rect 63 -272 79 -238
rect 113 -272 129 -238
rect 255 -272 271 -238
rect 305 -272 321 -238
rect -467 -340 -433 -278
rect 433 -340 467 -278
rect -467 -374 -371 -340
rect 371 -374 467 -340
<< viali >>
rect -209 238 -175 272
rect -17 238 17 272
rect 175 238 209 272
rect -353 -188 -319 188
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect 319 -188 353 188
rect -305 -272 -271 -238
rect -113 -272 -79 -238
rect 79 -272 113 -238
rect 271 -272 305 -238
<< metal1 >>
rect -221 272 -163 278
rect -221 238 -209 272
rect -175 238 -163 272
rect -221 232 -163 238
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect 163 272 221 278
rect 163 238 175 272
rect 209 238 221 272
rect 163 232 221 238
rect -359 188 -313 200
rect -359 -188 -353 188
rect -319 -188 -313 188
rect -359 -200 -313 -188
rect -263 188 -217 200
rect -263 -188 -257 188
rect -223 -188 -217 188
rect -263 -200 -217 -188
rect -167 188 -121 200
rect -167 -188 -161 188
rect -127 -188 -121 188
rect -167 -200 -121 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 121 188 167 200
rect 121 -188 127 188
rect 161 -188 167 188
rect 121 -200 167 -188
rect 217 188 263 200
rect 217 -188 223 188
rect 257 -188 263 188
rect 217 -200 263 -188
rect 313 188 359 200
rect 313 -188 319 188
rect 353 -188 359 188
rect 313 -200 359 -188
rect -317 -238 -259 -232
rect -317 -272 -305 -238
rect -271 -272 -259 -238
rect -317 -278 -259 -272
rect -125 -238 -67 -232
rect -125 -272 -113 -238
rect -79 -272 -67 -238
rect -125 -278 -67 -272
rect 67 -238 125 -232
rect 67 -272 79 -238
rect 113 -272 125 -238
rect 67 -278 125 -272
rect 259 -238 317 -232
rect 259 -272 271 -238
rect 305 -272 317 -238
rect 259 -278 317 -272
<< properties >>
string FIXED_BBOX -450 -357 450 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
