magic
tech sky130A
magscale 1 2
timestamp 1683628480
<< error_p >>
rect 19418 310256 19434 310260
rect 129578 310256 129594 310260
rect 19198 310253 19418 310256
rect 129358 310253 129578 310256
rect 6675 309987 6691 310215
rect 116835 309996 116842 310220
rect 6691 309984 6702 309987
rect 116842 309984 116862 309996
rect 19138 308004 19158 308016
rect 129298 308013 129309 308016
rect 19158 307780 19165 308004
rect 129309 307785 129325 308013
rect 6422 307744 6642 307747
rect 116582 307744 116802 307747
rect 6406 307740 6422 307744
rect 116566 307740 116582 307744
rect 6086 307260 6102 307280
rect 12941 307260 13841 307280
rect 19802 307260 19808 307280
rect 12941 307120 13841 307140
rect 19802 307137 19808 307140
rect 5766 307040 5782 307060
rect 12941 307040 13841 307060
rect 19892 307050 20112 307053
rect 20112 307040 20128 307050
rect 20112 306940 20128 306960
rect 20112 306817 20128 306820
rect 19418 295256 19434 295260
rect 19198 295253 19418 295256
rect 6675 294987 6691 295215
rect 6691 294984 6702 294987
rect 19138 293004 19158 293016
rect 19158 292780 19165 293004
rect 6422 292744 6642 292747
rect 6406 292740 6422 292744
rect 19418 280256 19434 280260
rect 19198 280253 19418 280256
rect 6675 279987 6691 280215
rect 6691 279984 6702 279987
rect 19138 278004 19158 278016
rect 19158 277780 19165 278004
rect 6422 277744 6642 277747
rect 6406 277740 6422 277744
rect 19418 265256 19434 265260
rect 19198 265253 19418 265256
rect 6675 264987 6691 265215
rect 6691 264984 6702 264987
rect 19138 263004 19158 263016
rect 19158 262780 19165 263004
rect 6422 262744 6642 262747
rect 6406 262740 6422 262744
rect 19418 250256 19434 250260
rect 19198 250253 19418 250256
rect 6675 249987 6691 250215
rect 6691 249984 6702 249987
rect 19138 248004 19158 248016
rect 19158 247780 19165 248004
rect 6422 247744 6642 247747
rect 6406 247740 6422 247744
rect 19418 200256 19434 200260
rect 129578 200256 129594 200260
rect 19198 200253 19418 200256
rect 129358 200253 129578 200256
rect 6675 199987 6691 200215
rect 116835 199996 116842 200220
rect 6691 199984 6702 199987
rect 116842 199984 116862 199996
rect 19138 198004 19158 198016
rect 129298 198013 129309 198016
rect 19158 197780 19165 198004
rect 129309 197785 129325 198013
rect 6422 197744 6642 197747
rect 116582 197744 116802 197747
rect 6406 197740 6422 197744
rect 116566 197740 116582 197744
rect 6086 197260 6102 197280
rect 12941 197260 13841 197280
rect 19802 197260 19808 197280
rect 12941 197120 13841 197140
rect 19802 197137 19808 197140
rect 5766 197040 5782 197060
rect 12941 197040 13841 197060
rect 19892 197050 20112 197053
rect 20112 197040 20128 197050
rect 20112 196940 20128 196960
rect 20112 196817 20128 196820
rect 19418 185256 19434 185260
rect 19198 185253 19418 185256
rect 6675 184987 6691 185215
rect 6691 184984 6702 184987
rect 19138 183004 19158 183016
rect 19158 182780 19165 183004
rect 6422 182744 6642 182747
rect 6406 182740 6422 182744
rect 19418 170256 19434 170260
rect 19198 170253 19418 170256
rect 6675 169987 6691 170215
rect 6691 169984 6702 169987
rect 19138 168004 19158 168016
rect 19158 167780 19165 168004
rect 6422 167744 6642 167747
rect 6406 167740 6422 167744
rect 19418 155256 19434 155260
rect 19198 155253 19418 155256
rect 6675 154987 6691 155215
rect 6691 154984 6702 154987
rect 19138 153004 19158 153016
rect 19158 152780 19165 153004
rect 6422 152744 6642 152747
rect 6406 152740 6422 152744
rect 19418 140256 19434 140260
rect 19198 140253 19418 140256
rect 6675 139987 6691 140215
rect 6691 139984 6702 139987
rect 19138 138004 19158 138016
rect 19158 137780 19165 138004
rect 6422 137744 6642 137747
rect 6406 137740 6422 137744
rect 19418 88256 19434 88260
rect 129578 88256 129594 88260
rect 19198 88253 19418 88256
rect 129358 88253 129578 88256
rect 6675 87987 6691 88215
rect 116835 87996 116842 88220
rect 6691 87984 6702 87987
rect 116842 87984 116862 87996
rect 19138 86004 19158 86016
rect 129298 86013 129309 86016
rect 19158 85780 19165 86004
rect 129309 85785 129325 86013
rect 6422 85744 6642 85747
rect 116582 85744 116802 85747
rect 6406 85740 6422 85744
rect 116566 85740 116582 85744
rect 6086 85260 6102 85280
rect 12941 85260 13841 85280
rect 19802 85260 19808 85280
rect 12941 85120 13841 85140
rect 19802 85137 19808 85140
rect 5766 85040 5782 85060
rect 12941 85040 13841 85060
rect 19892 85050 20112 85053
rect 20112 85040 20128 85050
rect 20112 84940 20128 84960
rect 20112 84817 20128 84820
rect 19418 73256 19434 73260
rect 19198 73253 19418 73256
rect 6675 72987 6691 73215
rect 6691 72984 6702 72987
rect 19138 71004 19158 71016
rect 19158 70780 19165 71004
rect 6422 70744 6642 70747
rect 6406 70740 6422 70744
rect 19418 58256 19434 58260
rect 19198 58253 19418 58256
rect 6675 57987 6691 58215
rect 6691 57984 6702 57987
rect 19138 56004 19158 56016
rect 19158 55780 19165 56004
rect 6422 55744 6642 55747
rect 6406 55740 6422 55744
rect 19418 43256 19434 43260
rect 19198 43253 19418 43256
rect 6675 42987 6691 43215
rect 6691 42984 6702 42987
rect 19138 41004 19158 41016
rect 19158 40780 19165 41004
rect 6422 40744 6642 40747
rect 6406 40740 6422 40744
rect 19418 28256 19434 28260
rect 19198 28253 19418 28256
rect 6675 27987 6691 28215
rect 6691 27984 6702 27987
rect 19138 26004 19158 26016
rect 19158 25780 19165 26004
rect 6422 25744 6642 25747
rect 6406 25740 6422 25744
use top  top_0
timestamp 1683628480
transform 1 0 6000 0 1 260000
box -6000 -26000 130000 64000
use top  top_1
timestamp 1683628480
transform 1 0 6000 0 1 38000
box -6000 -26000 130000 64000
use top  top_2
timestamp 1683628480
transform 1 0 6000 0 1 150000
box -6000 -26000 130000 64000
<< end >>
