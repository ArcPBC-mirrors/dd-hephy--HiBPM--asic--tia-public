magic
tech sky130A
magscale 1 2
timestamp 1688995864
<< pwell >>
rect -1457 -1028 1457 1028
<< nmos >>
rect -1261 418 -1061 818
rect -1003 418 -803 818
rect -745 418 -545 818
rect -487 418 -287 818
rect -229 418 -29 818
rect 29 418 229 818
rect 287 418 487 818
rect 545 418 745 818
rect 803 418 1003 818
rect 1061 418 1261 818
rect -1261 -200 -1061 200
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
rect 1061 -200 1261 200
rect -1261 -818 -1061 -418
rect -1003 -818 -803 -418
rect -745 -818 -545 -418
rect -487 -818 -287 -418
rect -229 -818 -29 -418
rect 29 -818 229 -418
rect 287 -818 487 -418
rect 545 -818 745 -418
rect 803 -818 1003 -418
rect 1061 -818 1261 -418
<< ndiff >>
rect -1319 806 -1261 818
rect -1319 430 -1307 806
rect -1273 430 -1261 806
rect -1319 418 -1261 430
rect -1061 806 -1003 818
rect -1061 430 -1049 806
rect -1015 430 -1003 806
rect -1061 418 -1003 430
rect -803 806 -745 818
rect -803 430 -791 806
rect -757 430 -745 806
rect -803 418 -745 430
rect -545 806 -487 818
rect -545 430 -533 806
rect -499 430 -487 806
rect -545 418 -487 430
rect -287 806 -229 818
rect -287 430 -275 806
rect -241 430 -229 806
rect -287 418 -229 430
rect -29 806 29 818
rect -29 430 -17 806
rect 17 430 29 806
rect -29 418 29 430
rect 229 806 287 818
rect 229 430 241 806
rect 275 430 287 806
rect 229 418 287 430
rect 487 806 545 818
rect 487 430 499 806
rect 533 430 545 806
rect 487 418 545 430
rect 745 806 803 818
rect 745 430 757 806
rect 791 430 803 806
rect 745 418 803 430
rect 1003 806 1061 818
rect 1003 430 1015 806
rect 1049 430 1061 806
rect 1003 418 1061 430
rect 1261 806 1319 818
rect 1261 430 1273 806
rect 1307 430 1319 806
rect 1261 418 1319 430
rect -1319 188 -1261 200
rect -1319 -188 -1307 188
rect -1273 -188 -1261 188
rect -1319 -200 -1261 -188
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
rect 1261 188 1319 200
rect 1261 -188 1273 188
rect 1307 -188 1319 188
rect 1261 -200 1319 -188
rect -1319 -430 -1261 -418
rect -1319 -806 -1307 -430
rect -1273 -806 -1261 -430
rect -1319 -818 -1261 -806
rect -1061 -430 -1003 -418
rect -1061 -806 -1049 -430
rect -1015 -806 -1003 -430
rect -1061 -818 -1003 -806
rect -803 -430 -745 -418
rect -803 -806 -791 -430
rect -757 -806 -745 -430
rect -803 -818 -745 -806
rect -545 -430 -487 -418
rect -545 -806 -533 -430
rect -499 -806 -487 -430
rect -545 -818 -487 -806
rect -287 -430 -229 -418
rect -287 -806 -275 -430
rect -241 -806 -229 -430
rect -287 -818 -229 -806
rect -29 -430 29 -418
rect -29 -806 -17 -430
rect 17 -806 29 -430
rect -29 -818 29 -806
rect 229 -430 287 -418
rect 229 -806 241 -430
rect 275 -806 287 -430
rect 229 -818 287 -806
rect 487 -430 545 -418
rect 487 -806 499 -430
rect 533 -806 545 -430
rect 487 -818 545 -806
rect 745 -430 803 -418
rect 745 -806 757 -430
rect 791 -806 803 -430
rect 745 -818 803 -806
rect 1003 -430 1061 -418
rect 1003 -806 1015 -430
rect 1049 -806 1061 -430
rect 1003 -818 1061 -806
rect 1261 -430 1319 -418
rect 1261 -806 1273 -430
rect 1307 -806 1319 -430
rect 1261 -818 1319 -806
<< ndiffc >>
rect -1307 430 -1273 806
rect -1049 430 -1015 806
rect -791 430 -757 806
rect -533 430 -499 806
rect -275 430 -241 806
rect -17 430 17 806
rect 241 430 275 806
rect 499 430 533 806
rect 757 430 791 806
rect 1015 430 1049 806
rect 1273 430 1307 806
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect -1307 -806 -1273 -430
rect -1049 -806 -1015 -430
rect -791 -806 -757 -430
rect -533 -806 -499 -430
rect -275 -806 -241 -430
rect -17 -806 17 -430
rect 241 -806 275 -430
rect 499 -806 533 -430
rect 757 -806 791 -430
rect 1015 -806 1049 -430
rect 1273 -806 1307 -430
<< psubdiff >>
rect -1421 958 -1325 992
rect 1325 958 1421 992
rect -1421 896 -1387 958
rect 1387 896 1421 958
rect -1421 -958 -1387 -896
rect 1387 -958 1421 -896
rect -1421 -992 -1325 -958
rect 1325 -992 1421 -958
<< psubdiffcont >>
rect -1325 958 1325 992
rect -1421 -896 -1387 896
rect 1387 -896 1421 896
rect -1325 -992 1325 -958
<< poly >>
rect -1261 890 -1061 906
rect -1261 856 -1245 890
rect -1077 856 -1061 890
rect -1261 818 -1061 856
rect -1003 890 -803 906
rect -1003 856 -987 890
rect -819 856 -803 890
rect -1003 818 -803 856
rect -745 890 -545 906
rect -745 856 -729 890
rect -561 856 -545 890
rect -745 818 -545 856
rect -487 890 -287 906
rect -487 856 -471 890
rect -303 856 -287 890
rect -487 818 -287 856
rect -229 890 -29 906
rect -229 856 -213 890
rect -45 856 -29 890
rect -229 818 -29 856
rect 29 890 229 906
rect 29 856 45 890
rect 213 856 229 890
rect 29 818 229 856
rect 287 890 487 906
rect 287 856 303 890
rect 471 856 487 890
rect 287 818 487 856
rect 545 890 745 906
rect 545 856 561 890
rect 729 856 745 890
rect 545 818 745 856
rect 803 890 1003 906
rect 803 856 819 890
rect 987 856 1003 890
rect 803 818 1003 856
rect 1061 890 1261 906
rect 1061 856 1077 890
rect 1245 856 1261 890
rect 1061 818 1261 856
rect -1261 380 -1061 418
rect -1261 346 -1245 380
rect -1077 346 -1061 380
rect -1261 330 -1061 346
rect -1003 380 -803 418
rect -1003 346 -987 380
rect -819 346 -803 380
rect -1003 330 -803 346
rect -745 380 -545 418
rect -745 346 -729 380
rect -561 346 -545 380
rect -745 330 -545 346
rect -487 380 -287 418
rect -487 346 -471 380
rect -303 346 -287 380
rect -487 330 -287 346
rect -229 380 -29 418
rect -229 346 -213 380
rect -45 346 -29 380
rect -229 330 -29 346
rect 29 380 229 418
rect 29 346 45 380
rect 213 346 229 380
rect 29 330 229 346
rect 287 380 487 418
rect 287 346 303 380
rect 471 346 487 380
rect 287 330 487 346
rect 545 380 745 418
rect 545 346 561 380
rect 729 346 745 380
rect 545 330 745 346
rect 803 380 1003 418
rect 803 346 819 380
rect 987 346 1003 380
rect 803 330 1003 346
rect 1061 380 1261 418
rect 1061 346 1077 380
rect 1245 346 1261 380
rect 1061 330 1261 346
rect -1261 272 -1061 288
rect -1261 238 -1245 272
rect -1077 238 -1061 272
rect -1261 200 -1061 238
rect -1003 272 -803 288
rect -1003 238 -987 272
rect -819 238 -803 272
rect -1003 200 -803 238
rect -745 272 -545 288
rect -745 238 -729 272
rect -561 238 -545 272
rect -745 200 -545 238
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect 545 272 745 288
rect 545 238 561 272
rect 729 238 745 272
rect 545 200 745 238
rect 803 272 1003 288
rect 803 238 819 272
rect 987 238 1003 272
rect 803 200 1003 238
rect 1061 272 1261 288
rect 1061 238 1077 272
rect 1245 238 1261 272
rect 1061 200 1261 238
rect -1261 -238 -1061 -200
rect -1261 -272 -1245 -238
rect -1077 -272 -1061 -238
rect -1261 -288 -1061 -272
rect -1003 -238 -803 -200
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -1003 -288 -803 -272
rect -745 -238 -545 -200
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -745 -288 -545 -272
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
rect 545 -238 745 -200
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 545 -288 745 -272
rect 803 -238 1003 -200
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect 803 -288 1003 -272
rect 1061 -238 1261 -200
rect 1061 -272 1077 -238
rect 1245 -272 1261 -238
rect 1061 -288 1261 -272
rect -1261 -346 -1061 -330
rect -1261 -380 -1245 -346
rect -1077 -380 -1061 -346
rect -1261 -418 -1061 -380
rect -1003 -346 -803 -330
rect -1003 -380 -987 -346
rect -819 -380 -803 -346
rect -1003 -418 -803 -380
rect -745 -346 -545 -330
rect -745 -380 -729 -346
rect -561 -380 -545 -346
rect -745 -418 -545 -380
rect -487 -346 -287 -330
rect -487 -380 -471 -346
rect -303 -380 -287 -346
rect -487 -418 -287 -380
rect -229 -346 -29 -330
rect -229 -380 -213 -346
rect -45 -380 -29 -346
rect -229 -418 -29 -380
rect 29 -346 229 -330
rect 29 -380 45 -346
rect 213 -380 229 -346
rect 29 -418 229 -380
rect 287 -346 487 -330
rect 287 -380 303 -346
rect 471 -380 487 -346
rect 287 -418 487 -380
rect 545 -346 745 -330
rect 545 -380 561 -346
rect 729 -380 745 -346
rect 545 -418 745 -380
rect 803 -346 1003 -330
rect 803 -380 819 -346
rect 987 -380 1003 -346
rect 803 -418 1003 -380
rect 1061 -346 1261 -330
rect 1061 -380 1077 -346
rect 1245 -380 1261 -346
rect 1061 -418 1261 -380
rect -1261 -856 -1061 -818
rect -1261 -890 -1245 -856
rect -1077 -890 -1061 -856
rect -1261 -906 -1061 -890
rect -1003 -856 -803 -818
rect -1003 -890 -987 -856
rect -819 -890 -803 -856
rect -1003 -906 -803 -890
rect -745 -856 -545 -818
rect -745 -890 -729 -856
rect -561 -890 -545 -856
rect -745 -906 -545 -890
rect -487 -856 -287 -818
rect -487 -890 -471 -856
rect -303 -890 -287 -856
rect -487 -906 -287 -890
rect -229 -856 -29 -818
rect -229 -890 -213 -856
rect -45 -890 -29 -856
rect -229 -906 -29 -890
rect 29 -856 229 -818
rect 29 -890 45 -856
rect 213 -890 229 -856
rect 29 -906 229 -890
rect 287 -856 487 -818
rect 287 -890 303 -856
rect 471 -890 487 -856
rect 287 -906 487 -890
rect 545 -856 745 -818
rect 545 -890 561 -856
rect 729 -890 745 -856
rect 545 -906 745 -890
rect 803 -856 1003 -818
rect 803 -890 819 -856
rect 987 -890 1003 -856
rect 803 -906 1003 -890
rect 1061 -856 1261 -818
rect 1061 -890 1077 -856
rect 1245 -890 1261 -856
rect 1061 -906 1261 -890
<< polycont >>
rect -1245 856 -1077 890
rect -987 856 -819 890
rect -729 856 -561 890
rect -471 856 -303 890
rect -213 856 -45 890
rect 45 856 213 890
rect 303 856 471 890
rect 561 856 729 890
rect 819 856 987 890
rect 1077 856 1245 890
rect -1245 346 -1077 380
rect -987 346 -819 380
rect -729 346 -561 380
rect -471 346 -303 380
rect -213 346 -45 380
rect 45 346 213 380
rect 303 346 471 380
rect 561 346 729 380
rect 819 346 987 380
rect 1077 346 1245 380
rect -1245 238 -1077 272
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect 1077 238 1245 272
rect -1245 -272 -1077 -238
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
rect 1077 -272 1245 -238
rect -1245 -380 -1077 -346
rect -987 -380 -819 -346
rect -729 -380 -561 -346
rect -471 -380 -303 -346
rect -213 -380 -45 -346
rect 45 -380 213 -346
rect 303 -380 471 -346
rect 561 -380 729 -346
rect 819 -380 987 -346
rect 1077 -380 1245 -346
rect -1245 -890 -1077 -856
rect -987 -890 -819 -856
rect -729 -890 -561 -856
rect -471 -890 -303 -856
rect -213 -890 -45 -856
rect 45 -890 213 -856
rect 303 -890 471 -856
rect 561 -890 729 -856
rect 819 -890 987 -856
rect 1077 -890 1245 -856
<< locali >>
rect -1421 958 -1325 992
rect 1325 958 1421 992
rect -1421 896 -1387 958
rect 1387 896 1421 958
rect -1261 856 -1245 890
rect -1077 856 -1061 890
rect -1003 856 -987 890
rect -819 856 -803 890
rect -745 856 -729 890
rect -561 856 -545 890
rect -487 856 -471 890
rect -303 856 -287 890
rect -229 856 -213 890
rect -45 856 -29 890
rect 29 856 45 890
rect 213 856 229 890
rect 287 856 303 890
rect 471 856 487 890
rect 545 856 561 890
rect 729 856 745 890
rect 803 856 819 890
rect 987 856 1003 890
rect 1061 856 1077 890
rect 1245 856 1261 890
rect -1307 806 -1273 822
rect -1307 414 -1273 430
rect -1049 806 -1015 822
rect -1049 414 -1015 430
rect -791 806 -757 822
rect -791 414 -757 430
rect -533 806 -499 822
rect -533 414 -499 430
rect -275 806 -241 822
rect -275 414 -241 430
rect -17 806 17 822
rect -17 414 17 430
rect 241 806 275 822
rect 241 414 275 430
rect 499 806 533 822
rect 499 414 533 430
rect 757 806 791 822
rect 757 414 791 430
rect 1015 806 1049 822
rect 1015 414 1049 430
rect 1273 806 1307 822
rect 1273 414 1307 430
rect -1261 346 -1245 380
rect -1077 346 -1061 380
rect -1003 346 -987 380
rect -819 346 -803 380
rect -745 346 -729 380
rect -561 346 -545 380
rect -487 346 -471 380
rect -303 346 -287 380
rect -229 346 -213 380
rect -45 346 -29 380
rect 29 346 45 380
rect 213 346 229 380
rect 287 346 303 380
rect 471 346 487 380
rect 545 346 561 380
rect 729 346 745 380
rect 803 346 819 380
rect 987 346 1003 380
rect 1061 346 1077 380
rect 1245 346 1261 380
rect -1261 238 -1245 272
rect -1077 238 -1061 272
rect -1003 238 -987 272
rect -819 238 -803 272
rect -745 238 -729 272
rect -561 238 -545 272
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect 545 238 561 272
rect 729 238 745 272
rect 803 238 819 272
rect 987 238 1003 272
rect 1061 238 1077 272
rect 1245 238 1261 272
rect -1307 188 -1273 204
rect -1307 -204 -1273 -188
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect 1273 188 1307 204
rect 1273 -204 1307 -188
rect -1261 -272 -1245 -238
rect -1077 -272 -1061 -238
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect 1061 -272 1077 -238
rect 1245 -272 1261 -238
rect -1261 -380 -1245 -346
rect -1077 -380 -1061 -346
rect -1003 -380 -987 -346
rect -819 -380 -803 -346
rect -745 -380 -729 -346
rect -561 -380 -545 -346
rect -487 -380 -471 -346
rect -303 -380 -287 -346
rect -229 -380 -213 -346
rect -45 -380 -29 -346
rect 29 -380 45 -346
rect 213 -380 229 -346
rect 287 -380 303 -346
rect 471 -380 487 -346
rect 545 -380 561 -346
rect 729 -380 745 -346
rect 803 -380 819 -346
rect 987 -380 1003 -346
rect 1061 -380 1077 -346
rect 1245 -380 1261 -346
rect -1307 -430 -1273 -414
rect -1307 -822 -1273 -806
rect -1049 -430 -1015 -414
rect -1049 -822 -1015 -806
rect -791 -430 -757 -414
rect -791 -822 -757 -806
rect -533 -430 -499 -414
rect -533 -822 -499 -806
rect -275 -430 -241 -414
rect -275 -822 -241 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 241 -430 275 -414
rect 241 -822 275 -806
rect 499 -430 533 -414
rect 499 -822 533 -806
rect 757 -430 791 -414
rect 757 -822 791 -806
rect 1015 -430 1049 -414
rect 1015 -822 1049 -806
rect 1273 -430 1307 -414
rect 1273 -822 1307 -806
rect -1261 -890 -1245 -856
rect -1077 -890 -1061 -856
rect -1003 -890 -987 -856
rect -819 -890 -803 -856
rect -745 -890 -729 -856
rect -561 -890 -545 -856
rect -487 -890 -471 -856
rect -303 -890 -287 -856
rect -229 -890 -213 -856
rect -45 -890 -29 -856
rect 29 -890 45 -856
rect 213 -890 229 -856
rect 287 -890 303 -856
rect 471 -890 487 -856
rect 545 -890 561 -856
rect 729 -890 745 -856
rect 803 -890 819 -856
rect 987 -890 1003 -856
rect 1061 -890 1077 -856
rect 1245 -890 1261 -856
rect -1421 -958 -1387 -896
rect 1387 -958 1421 -896
rect -1421 -992 -1325 -958
rect 1325 -992 1421 -958
<< viali >>
rect -1245 856 -1077 890
rect -987 856 -819 890
rect -729 856 -561 890
rect -471 856 -303 890
rect -213 856 -45 890
rect 45 856 213 890
rect 303 856 471 890
rect 561 856 729 890
rect 819 856 987 890
rect 1077 856 1245 890
rect -1307 430 -1273 806
rect -1049 430 -1015 806
rect -791 430 -757 806
rect -533 430 -499 806
rect -275 430 -241 806
rect -17 430 17 806
rect 241 430 275 806
rect 499 430 533 806
rect 757 430 791 806
rect 1015 430 1049 806
rect 1273 430 1307 806
rect -1245 346 -1077 380
rect -987 346 -819 380
rect -729 346 -561 380
rect -471 346 -303 380
rect -213 346 -45 380
rect 45 346 213 380
rect 303 346 471 380
rect 561 346 729 380
rect 819 346 987 380
rect 1077 346 1245 380
rect -1245 238 -1077 272
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect 1077 238 1245 272
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect -1245 -272 -1077 -238
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
rect 1077 -272 1245 -238
rect -1245 -380 -1077 -346
rect -987 -380 -819 -346
rect -729 -380 -561 -346
rect -471 -380 -303 -346
rect -213 -380 -45 -346
rect 45 -380 213 -346
rect 303 -380 471 -346
rect 561 -380 729 -346
rect 819 -380 987 -346
rect 1077 -380 1245 -346
rect -1307 -806 -1273 -430
rect -1049 -806 -1015 -430
rect -791 -806 -757 -430
rect -533 -806 -499 -430
rect -275 -806 -241 -430
rect -17 -806 17 -430
rect 241 -806 275 -430
rect 499 -806 533 -430
rect 757 -806 791 -430
rect 1015 -806 1049 -430
rect 1273 -806 1307 -430
rect -1245 -890 -1077 -856
rect -987 -890 -819 -856
rect -729 -890 -561 -856
rect -471 -890 -303 -856
rect -213 -890 -45 -856
rect 45 -890 213 -856
rect 303 -890 471 -856
rect 561 -890 729 -856
rect 819 -890 987 -856
rect 1077 -890 1245 -856
<< metal1 >>
rect -1257 890 -1065 896
rect -1257 856 -1245 890
rect -1077 856 -1065 890
rect -1257 850 -1065 856
rect -999 890 -807 896
rect -999 856 -987 890
rect -819 856 -807 890
rect -999 850 -807 856
rect -741 890 -549 896
rect -741 856 -729 890
rect -561 856 -549 890
rect -741 850 -549 856
rect -483 890 -291 896
rect -483 856 -471 890
rect -303 856 -291 890
rect -483 850 -291 856
rect -225 890 -33 896
rect -225 856 -213 890
rect -45 856 -33 890
rect -225 850 -33 856
rect 33 890 225 896
rect 33 856 45 890
rect 213 856 225 890
rect 33 850 225 856
rect 291 890 483 896
rect 291 856 303 890
rect 471 856 483 890
rect 291 850 483 856
rect 549 890 741 896
rect 549 856 561 890
rect 729 856 741 890
rect 549 850 741 856
rect 807 890 999 896
rect 807 856 819 890
rect 987 856 999 890
rect 807 850 999 856
rect 1065 890 1257 896
rect 1065 856 1077 890
rect 1245 856 1257 890
rect 1065 850 1257 856
rect -1313 806 -1267 818
rect -1313 430 -1307 806
rect -1273 430 -1267 806
rect -1313 418 -1267 430
rect -1055 806 -1009 818
rect -1055 430 -1049 806
rect -1015 430 -1009 806
rect -1055 418 -1009 430
rect -797 806 -751 818
rect -797 430 -791 806
rect -757 430 -751 806
rect -797 418 -751 430
rect -539 806 -493 818
rect -539 430 -533 806
rect -499 430 -493 806
rect -539 418 -493 430
rect -281 806 -235 818
rect -281 430 -275 806
rect -241 430 -235 806
rect -281 418 -235 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 235 806 281 818
rect 235 430 241 806
rect 275 430 281 806
rect 235 418 281 430
rect 493 806 539 818
rect 493 430 499 806
rect 533 430 539 806
rect 493 418 539 430
rect 751 806 797 818
rect 751 430 757 806
rect 791 430 797 806
rect 751 418 797 430
rect 1009 806 1055 818
rect 1009 430 1015 806
rect 1049 430 1055 806
rect 1009 418 1055 430
rect 1267 806 1313 818
rect 1267 430 1273 806
rect 1307 430 1313 806
rect 1267 418 1313 430
rect -1257 380 -1065 386
rect -1257 346 -1245 380
rect -1077 346 -1065 380
rect -1257 340 -1065 346
rect -999 380 -807 386
rect -999 346 -987 380
rect -819 346 -807 380
rect -999 340 -807 346
rect -741 380 -549 386
rect -741 346 -729 380
rect -561 346 -549 380
rect -741 340 -549 346
rect -483 380 -291 386
rect -483 346 -471 380
rect -303 346 -291 380
rect -483 340 -291 346
rect -225 380 -33 386
rect -225 346 -213 380
rect -45 346 -33 380
rect -225 340 -33 346
rect 33 380 225 386
rect 33 346 45 380
rect 213 346 225 380
rect 33 340 225 346
rect 291 380 483 386
rect 291 346 303 380
rect 471 346 483 380
rect 291 340 483 346
rect 549 380 741 386
rect 549 346 561 380
rect 729 346 741 380
rect 549 340 741 346
rect 807 380 999 386
rect 807 346 819 380
rect 987 346 999 380
rect 807 340 999 346
rect 1065 380 1257 386
rect 1065 346 1077 380
rect 1245 346 1257 380
rect 1065 340 1257 346
rect -1257 272 -1065 278
rect -1257 238 -1245 272
rect -1077 238 -1065 272
rect -1257 232 -1065 238
rect -999 272 -807 278
rect -999 238 -987 272
rect -819 238 -807 272
rect -999 232 -807 238
rect -741 272 -549 278
rect -741 238 -729 272
rect -561 238 -549 272
rect -741 232 -549 238
rect -483 272 -291 278
rect -483 238 -471 272
rect -303 238 -291 272
rect -483 232 -291 238
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect 291 272 483 278
rect 291 238 303 272
rect 471 238 483 272
rect 291 232 483 238
rect 549 272 741 278
rect 549 238 561 272
rect 729 238 741 272
rect 549 232 741 238
rect 807 272 999 278
rect 807 238 819 272
rect 987 238 999 272
rect 807 232 999 238
rect 1065 272 1257 278
rect 1065 238 1077 272
rect 1245 238 1257 272
rect 1065 232 1257 238
rect -1313 188 -1267 200
rect -1313 -188 -1307 188
rect -1273 -188 -1267 188
rect -1313 -200 -1267 -188
rect -1055 188 -1009 200
rect -1055 -188 -1049 188
rect -1015 -188 -1009 188
rect -1055 -200 -1009 -188
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect 1009 188 1055 200
rect 1009 -188 1015 188
rect 1049 -188 1055 188
rect 1009 -200 1055 -188
rect 1267 188 1313 200
rect 1267 -188 1273 188
rect 1307 -188 1313 188
rect 1267 -200 1313 -188
rect -1257 -238 -1065 -232
rect -1257 -272 -1245 -238
rect -1077 -272 -1065 -238
rect -1257 -278 -1065 -272
rect -999 -238 -807 -232
rect -999 -272 -987 -238
rect -819 -272 -807 -238
rect -999 -278 -807 -272
rect -741 -238 -549 -232
rect -741 -272 -729 -238
rect -561 -272 -549 -238
rect -741 -278 -549 -272
rect -483 -238 -291 -232
rect -483 -272 -471 -238
rect -303 -272 -291 -238
rect -483 -278 -291 -272
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
rect 291 -238 483 -232
rect 291 -272 303 -238
rect 471 -272 483 -238
rect 291 -278 483 -272
rect 549 -238 741 -232
rect 549 -272 561 -238
rect 729 -272 741 -238
rect 549 -278 741 -272
rect 807 -238 999 -232
rect 807 -272 819 -238
rect 987 -272 999 -238
rect 807 -278 999 -272
rect 1065 -238 1257 -232
rect 1065 -272 1077 -238
rect 1245 -272 1257 -238
rect 1065 -278 1257 -272
rect -1257 -346 -1065 -340
rect -1257 -380 -1245 -346
rect -1077 -380 -1065 -346
rect -1257 -386 -1065 -380
rect -999 -346 -807 -340
rect -999 -380 -987 -346
rect -819 -380 -807 -346
rect -999 -386 -807 -380
rect -741 -346 -549 -340
rect -741 -380 -729 -346
rect -561 -380 -549 -346
rect -741 -386 -549 -380
rect -483 -346 -291 -340
rect -483 -380 -471 -346
rect -303 -380 -291 -346
rect -483 -386 -291 -380
rect -225 -346 -33 -340
rect -225 -380 -213 -346
rect -45 -380 -33 -346
rect -225 -386 -33 -380
rect 33 -346 225 -340
rect 33 -380 45 -346
rect 213 -380 225 -346
rect 33 -386 225 -380
rect 291 -346 483 -340
rect 291 -380 303 -346
rect 471 -380 483 -346
rect 291 -386 483 -380
rect 549 -346 741 -340
rect 549 -380 561 -346
rect 729 -380 741 -346
rect 549 -386 741 -380
rect 807 -346 999 -340
rect 807 -380 819 -346
rect 987 -380 999 -346
rect 807 -386 999 -380
rect 1065 -346 1257 -340
rect 1065 -380 1077 -346
rect 1245 -380 1257 -346
rect 1065 -386 1257 -380
rect -1313 -430 -1267 -418
rect -1313 -806 -1307 -430
rect -1273 -806 -1267 -430
rect -1313 -818 -1267 -806
rect -1055 -430 -1009 -418
rect -1055 -806 -1049 -430
rect -1015 -806 -1009 -430
rect -1055 -818 -1009 -806
rect -797 -430 -751 -418
rect -797 -806 -791 -430
rect -757 -806 -751 -430
rect -797 -818 -751 -806
rect -539 -430 -493 -418
rect -539 -806 -533 -430
rect -499 -806 -493 -430
rect -539 -818 -493 -806
rect -281 -430 -235 -418
rect -281 -806 -275 -430
rect -241 -806 -235 -430
rect -281 -818 -235 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 235 -430 281 -418
rect 235 -806 241 -430
rect 275 -806 281 -430
rect 235 -818 281 -806
rect 493 -430 539 -418
rect 493 -806 499 -430
rect 533 -806 539 -430
rect 493 -818 539 -806
rect 751 -430 797 -418
rect 751 -806 757 -430
rect 791 -806 797 -430
rect 751 -818 797 -806
rect 1009 -430 1055 -418
rect 1009 -806 1015 -430
rect 1049 -806 1055 -430
rect 1009 -818 1055 -806
rect 1267 -430 1313 -418
rect 1267 -806 1273 -430
rect 1307 -806 1313 -430
rect 1267 -818 1313 -806
rect -1257 -856 -1065 -850
rect -1257 -890 -1245 -856
rect -1077 -890 -1065 -856
rect -1257 -896 -1065 -890
rect -999 -856 -807 -850
rect -999 -890 -987 -856
rect -819 -890 -807 -856
rect -999 -896 -807 -890
rect -741 -856 -549 -850
rect -741 -890 -729 -856
rect -561 -890 -549 -856
rect -741 -896 -549 -890
rect -483 -856 -291 -850
rect -483 -890 -471 -856
rect -303 -890 -291 -856
rect -483 -896 -291 -890
rect -225 -856 -33 -850
rect -225 -890 -213 -856
rect -45 -890 -33 -856
rect -225 -896 -33 -890
rect 33 -856 225 -850
rect 33 -890 45 -856
rect 213 -890 225 -856
rect 33 -896 225 -890
rect 291 -856 483 -850
rect 291 -890 303 -856
rect 471 -890 483 -856
rect 291 -896 483 -890
rect 549 -856 741 -850
rect 549 -890 561 -856
rect 729 -890 741 -856
rect 549 -896 741 -890
rect 807 -856 999 -850
rect 807 -890 819 -856
rect 987 -890 999 -856
rect 807 -896 999 -890
rect 1065 -856 1257 -850
rect 1065 -890 1077 -856
rect 1245 -890 1257 -856
rect 1065 -896 1257 -890
<< properties >>
string FIXED_BBOX -1404 -975 1404 975
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 3 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
