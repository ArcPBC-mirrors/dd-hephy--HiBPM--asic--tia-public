magic
tech sky130A
magscale 1 2
timestamp 1685113734
<< locali >>
rect -4 1692 836 1768
rect -4 1688 776 1692
<< metal1 >>
rect 136 2980 848 3064
rect 90 2768 100 2948
rect 152 2768 162 2948
rect 282 2768 292 2948
rect 344 2768 354 2948
rect 474 2768 484 2948
rect 536 2768 546 2948
rect 666 2768 676 2948
rect 728 2768 738 2948
rect 186 2548 196 2728
rect 248 2548 258 2728
rect 378 2548 388 2728
rect 440 2548 450 2728
rect 570 2548 580 2728
rect 632 2548 642 2728
rect 768 2516 848 2980
rect 196 2360 848 2516
rect 186 2152 196 2332
rect 248 2152 258 2332
rect 378 2152 388 2332
rect 440 2152 450 2332
rect 570 2152 580 2332
rect 632 2152 642 2332
rect 90 1932 100 2112
rect 152 1932 162 2112
rect 282 1932 292 2112
rect 344 1932 354 2112
rect 474 1932 484 2112
rect 536 1932 546 2112
rect 666 1932 676 2112
rect 728 1932 738 2112
rect 768 1896 848 2360
rect 140 1800 848 1896
rect 712 1624 796 1800
rect 148 1556 964 1624
rect 210 1348 220 1528
rect 272 1348 282 1528
rect 446 1348 456 1528
rect 508 1348 518 1528
rect 682 1348 692 1528
rect 744 1348 754 1528
rect 90 1124 100 1304
rect 152 1124 162 1304
rect 326 1124 336 1304
rect 388 1124 398 1304
rect 562 1124 572 1304
rect 624 1124 634 1304
rect 798 1124 808 1304
rect 860 1124 870 1304
rect 900 1096 964 1556
rect 152 1028 964 1096
<< via1 >>
rect 100 2768 152 2948
rect 292 2768 344 2948
rect 484 2768 536 2948
rect 676 2768 728 2948
rect 196 2548 248 2728
rect 388 2548 440 2728
rect 580 2548 632 2728
rect 196 2152 248 2332
rect 388 2152 440 2332
rect 580 2152 632 2332
rect 100 1932 152 2112
rect 292 1932 344 2112
rect 484 1932 536 2112
rect 676 1932 728 2112
rect 220 1348 272 1528
rect 456 1348 508 1528
rect 692 1348 744 1528
rect 100 1124 152 1304
rect 336 1124 388 1304
rect 572 1124 624 1304
rect 808 1124 860 1304
<< metal2 >>
rect -40 2948 860 3000
rect -40 2768 100 2948
rect 152 2776 292 2948
rect -40 2758 152 2768
rect 344 2776 484 2948
rect 292 2758 344 2768
rect 536 2776 676 2948
rect 484 2758 536 2768
rect 668 2768 676 2776
rect 728 2768 860 2948
rect -40 2120 140 2758
rect 668 2748 860 2768
rect 196 2728 248 2738
rect 388 2728 440 2738
rect 248 2548 388 2720
rect 580 2728 632 2738
rect 440 2548 580 2720
rect 196 2332 632 2548
rect 248 2160 388 2332
rect 196 2142 248 2152
rect 440 2160 580 2332
rect 388 2142 440 2152
rect 680 2160 860 2748
rect 580 2142 632 2152
rect -40 2112 152 2120
rect -40 1932 100 2112
rect 292 2112 344 2122
rect 152 1932 292 2104
rect 484 2112 536 2122
rect 344 1932 484 2104
rect 668 2112 860 2160
rect 668 2104 676 2112
rect 536 1932 676 2104
rect 728 1932 860 2112
rect -40 1820 860 1932
rect 220 1528 760 1820
rect 272 1360 456 1528
rect 220 1338 272 1348
rect 508 1360 692 1528
rect 456 1338 508 1348
rect 744 1360 760 1528
rect 692 1338 744 1348
rect 100 1304 152 1314
rect 336 1304 388 1314
rect 152 1124 336 1296
rect 572 1304 624 1314
rect 388 1124 572 1296
rect 808 1304 860 1314
rect 624 1124 808 1296
rect 100 1024 860 1124
use sky130_fd_pr__nfet_01v8_lvt_2CP4KV#0  sky130_fd_pr__nfet_01v8_lvt_2CP4KV_0
timestamp 1683888831
transform 1 0 415 0 1 2439
box -455 -719 455 719
use sky130_fd_pr__nfet_01v8_lvt_E7L2KW#0  sky130_fd_pr__nfet_01v8_lvt_E7L2KW_0
timestamp 1683887376
transform 1 0 481 0 1 1326
box -521 -410 521 410
<< end >>
