magic
tech sky130A
magscale 1 2
timestamp 1687207134
<< locali >>
rect 10800 2620 12160 2740
rect 10920 1920 11020 2620
rect 11960 1920 12060 2620
rect 6840 1820 16000 1920
rect 7780 -320 7880 1820
rect 8840 -320 8940 1820
rect 9880 -320 9980 1820
rect 10920 -320 11020 1820
rect 11960 -320 12060 1820
rect 13000 -320 13100 1820
rect 14040 -320 14140 1820
rect 15080 -320 15180 1820
rect 6840 -420 16000 -320
rect 7780 -2560 7880 -420
rect 8840 -2560 8940 -420
rect 9880 -2560 9980 -420
rect 10920 -2560 11020 -420
rect 11960 -2560 12060 -420
rect 13000 -2560 13100 -420
rect 14040 -2560 14140 -420
rect 15080 -2560 15180 -420
rect 6840 -2660 16000 -2560
rect 7780 -4820 7880 -2660
rect 8840 -4820 8940 -2660
rect 9880 -4820 9980 -2660
rect 10920 -4820 11020 -2660
rect 11960 -4820 12060 -2660
rect 13000 -4820 13100 -2660
rect 14040 -4820 14140 -2660
rect 7780 -4920 14960 -4820
rect 7780 -7060 7880 -4920
rect 8840 -6980 8940 -4920
rect 9880 -6980 9980 -4920
rect 10920 -6980 11020 -4920
rect 8840 -7060 8920 -6980
rect 9880 -7060 9960 -6980
rect 10920 -7060 11000 -6980
rect 11960 -7060 12060 -4920
rect 13000 -6980 13100 -4920
rect 14040 -6980 14140 -4920
rect 13000 -7060 13080 -6980
rect 14040 -7060 14120 -6980
rect 15080 -7060 15180 -2660
<< viali >>
rect 8920 -7080 9020 -6980
rect 9960 -7080 10060 -6980
rect 11000 -7080 11100 -6980
rect 13080 -7080 13180 -6980
rect 14120 -7080 14220 -6980
<< metal1 >>
rect 11030 5860 11040 6300
rect 11320 5860 11330 6300
rect 11630 5840 11640 6280
rect 11920 5840 11930 6280
rect 11030 4620 11040 5060
rect 11320 4620 11330 5060
rect 11630 4620 11640 5060
rect 11920 4620 11930 5060
rect 11030 4080 11040 4520
rect 11320 4080 11330 4520
rect 11630 4080 11640 4520
rect 11920 4080 11930 4520
rect 11030 2840 11040 3280
rect 11320 2840 11330 3280
rect 11630 2840 11640 3280
rect 11920 2840 11930 3280
rect 6820 -500 16040 -240
rect 6800 -2740 16020 -2480
rect 6800 -4980 16020 -4720
rect 7750 -7080 7760 -6940
rect 7900 -7080 7910 -6940
rect 8908 -6980 9032 -6974
rect 8908 -7080 8920 -6980
rect 9020 -7080 9032 -6980
rect 8908 -7086 9032 -7080
rect 9948 -6980 10072 -6974
rect 9948 -7080 9960 -6980
rect 10060 -7080 10072 -6980
rect 9948 -7086 10072 -7080
rect 10988 -6980 11112 -6974
rect 10988 -7080 11000 -6980
rect 11100 -7080 11112 -6980
rect 10988 -7086 11112 -7080
rect 13068 -6980 13192 -6974
rect 13068 -7080 13080 -6980
rect 13180 -7080 13192 -6980
rect 13068 -7086 13192 -7080
rect 14108 -6980 14232 -6974
rect 14108 -7080 14120 -6980
rect 14220 -7080 14232 -6980
rect 14108 -7086 14232 -7080
<< via1 >>
rect 11040 5860 11320 6300
rect 11640 5840 11920 6280
rect 11040 4620 11320 5060
rect 11640 4620 11920 5060
rect 11040 4080 11320 4520
rect 11640 4080 11920 4520
rect 11040 2840 11320 3280
rect 11640 2840 11920 3280
rect 7760 -7080 7900 -6940
rect 8920 -7080 9020 -6980
rect 9960 -7080 10060 -6980
rect 11000 -7080 11100 -6980
rect 13080 -7080 13180 -6980
rect 14120 -7080 14220 -6980
<< metal2 >>
rect 11040 6300 11320 6310
rect 10060 5860 11040 6300
rect 10060 5720 11320 5860
rect 11640 6280 11920 6290
rect 11920 5840 12900 6280
rect 11640 5700 12900 5840
rect 10060 5060 11320 5180
rect 10060 4620 11040 5060
rect 10060 4600 11320 4620
rect 11640 5060 12900 5200
rect 11920 4620 12900 5060
rect 11640 4610 11920 4620
rect 11040 4520 11320 4530
rect 10060 4080 11040 4520
rect 10060 3940 11320 4080
rect 11640 4520 11920 4530
rect 11920 4080 12900 4520
rect 11640 3940 12900 4080
rect 10080 3280 11340 3420
rect 10080 2840 11040 3280
rect 11320 2840 11340 3280
rect 11640 3280 12900 3420
rect 11920 2840 12900 3280
rect 11040 2830 11320 2840
rect 11640 2830 11920 2840
rect 6900 2160 16140 2170
rect 6900 1810 16140 1820
rect 6800 1560 15960 1680
rect 7060 1400 7460 1410
rect 7060 910 7460 920
rect 8100 1400 8500 1410
rect 8100 910 8500 920
rect 9140 1400 9540 1410
rect 9140 910 9540 920
rect 10180 1400 10580 1410
rect 10180 910 10580 920
rect 11220 1400 11620 1410
rect 11220 910 11620 920
rect 12260 1400 12660 1410
rect 12260 910 12660 920
rect 13300 1400 13700 1410
rect 13300 910 13700 920
rect 14340 1400 14740 1410
rect 14340 910 14740 920
rect 15400 1400 15800 1410
rect 15400 910 15800 920
rect 6740 -580 6840 720
rect 6920 -40 16040 -20
rect 6920 -300 7560 -40
rect 7980 -300 8600 -40
rect 9020 -300 9640 -40
rect 10060 -300 10680 -40
rect 11100 -300 11720 -40
rect 12140 -300 12780 -40
rect 13200 -300 13800 -40
rect 14220 -300 14860 -40
rect 15280 -300 16040 -40
rect 7560 -310 7980 -300
rect 8600 -310 9020 -300
rect 9640 -310 10060 -300
rect 10680 -310 11100 -300
rect 11720 -310 12140 -300
rect 12780 -310 13200 -300
rect 13800 -310 14220 -300
rect 14860 -310 15280 -300
rect 6740 -700 15900 -580
rect 6740 -2820 6840 -700
rect 7060 -860 7460 -850
rect 7060 -1350 7460 -1340
rect 8100 -860 8500 -850
rect 8100 -1350 8500 -1340
rect 9140 -860 9540 -850
rect 9140 -1350 9540 -1340
rect 10180 -860 10580 -850
rect 10180 -1350 10580 -1340
rect 11220 -860 11620 -850
rect 11220 -1350 11620 -1340
rect 12260 -860 12660 -850
rect 12260 -1350 12660 -1340
rect 13300 -860 13700 -850
rect 13300 -1350 13700 -1340
rect 14340 -860 14740 -850
rect 14340 -1350 14740 -1340
rect 15400 -860 15800 -850
rect 15400 -1350 15800 -1340
rect 6920 -2280 16040 -2240
rect 6920 -2520 7560 -2280
rect 7980 -2520 8600 -2280
rect 7560 -2550 7980 -2540
rect 9020 -2520 9640 -2280
rect 8600 -2550 9020 -2540
rect 10060 -2520 10680 -2280
rect 9640 -2550 10060 -2540
rect 11100 -2520 11720 -2280
rect 10680 -2550 11100 -2540
rect 12140 -2520 12780 -2280
rect 11720 -2550 12140 -2540
rect 13200 -2520 13800 -2280
rect 12780 -2550 13200 -2540
rect 14220 -2520 14860 -2280
rect 13800 -2550 14220 -2540
rect 15280 -2520 16040 -2280
rect 14860 -2550 15280 -2540
rect 6740 -2940 15900 -2820
rect 6740 -5060 6840 -2940
rect 7060 -3080 7460 -3070
rect 7060 -3570 7460 -3560
rect 8100 -3080 8500 -3070
rect 8100 -3570 8500 -3560
rect 9140 -3080 9540 -3070
rect 9140 -3570 9540 -3560
rect 10180 -3080 10580 -3070
rect 10180 -3570 10580 -3560
rect 11220 -3080 11620 -3070
rect 11220 -3570 11620 -3560
rect 12260 -3080 12660 -3070
rect 12260 -3570 12660 -3560
rect 13300 -3080 13700 -3070
rect 13300 -3570 13700 -3560
rect 14340 -3080 14740 -3070
rect 14340 -3570 14740 -3560
rect 15400 -3080 15800 -3070
rect 15400 -3570 15800 -3560
rect 6920 -4520 16040 -4500
rect 6920 -4780 7560 -4520
rect 7980 -4780 8600 -4520
rect 9020 -4780 9640 -4520
rect 10060 -4780 10680 -4520
rect 11100 -4780 11720 -4520
rect 12140 -4780 12780 -4520
rect 13200 -4780 13800 -4520
rect 14220 -4780 14860 -4520
rect 15280 -4780 16040 -4520
rect 7560 -4790 7980 -4780
rect 8600 -4790 9020 -4780
rect 9640 -4790 10060 -4780
rect 10680 -4790 11100 -4780
rect 11720 -4790 12140 -4780
rect 12780 -4790 13200 -4780
rect 13800 -4790 14220 -4780
rect 14860 -4790 15280 -4780
rect 6740 -5180 14880 -5060
rect 8100 -5340 8500 -5330
rect 8100 -5830 8500 -5820
rect 9140 -5340 9540 -5330
rect 9140 -5830 9540 -5820
rect 10180 -5340 10580 -5330
rect 10180 -5830 10580 -5820
rect 11220 -5340 11620 -5330
rect 11220 -5830 11620 -5820
rect 12260 -5340 12660 -5330
rect 12260 -5830 12660 -5820
rect 13300 -5340 13700 -5330
rect 13300 -5830 13700 -5820
rect 14340 -5340 14740 -5330
rect 14340 -5830 14740 -5820
rect 7540 -6800 15300 -6760
rect 7540 -7060 7560 -6800
rect 7540 -7080 7760 -7060
rect 7980 -7060 8600 -6800
rect 7900 -7080 8920 -7060
rect 9020 -7060 9640 -6800
rect 9020 -7080 9960 -7060
rect 10060 -7060 10680 -6800
rect 10060 -7080 11000 -7060
rect 11100 -7060 11720 -6800
rect 12140 -7060 12780 -6800
rect 11100 -7080 13080 -7060
rect 13200 -7060 13800 -6800
rect 13180 -7080 14120 -7060
rect 14220 -7060 14860 -6800
rect 15280 -7060 15300 -6800
rect 14220 -7080 15300 -7060
rect 7760 -7090 7900 -7080
rect 8920 -7090 9020 -7080
rect 9960 -7090 10060 -7080
rect 11000 -7090 11100 -7080
rect 13080 -7090 13180 -7080
rect 14120 -7090 14220 -7080
<< via2 >>
rect 6900 1820 16140 2160
rect 7060 920 7460 1400
rect 8100 920 8500 1400
rect 9140 920 9540 1400
rect 10180 920 10580 1400
rect 11220 920 11620 1400
rect 12260 920 12660 1400
rect 13300 920 13700 1400
rect 14340 920 14740 1400
rect 15400 920 15800 1400
rect 7560 -300 7980 -40
rect 8600 -300 9020 -40
rect 9640 -300 10060 -40
rect 10680 -300 11100 -40
rect 11720 -300 12140 -40
rect 12780 -300 13200 -40
rect 13800 -300 14220 -40
rect 14860 -300 15280 -40
rect 7060 -1340 7460 -860
rect 8100 -1340 8500 -860
rect 9140 -1340 9540 -860
rect 10180 -1340 10580 -860
rect 11220 -1340 11620 -860
rect 12260 -1340 12660 -860
rect 13300 -1340 13700 -860
rect 14340 -1340 14740 -860
rect 15400 -1340 15800 -860
rect 7560 -2540 7980 -2280
rect 8600 -2540 9020 -2280
rect 9640 -2540 10060 -2280
rect 10680 -2540 11100 -2280
rect 11720 -2540 12140 -2280
rect 12780 -2540 13200 -2280
rect 13800 -2540 14220 -2280
rect 14860 -2540 15280 -2280
rect 7060 -3560 7460 -3080
rect 8100 -3560 8500 -3080
rect 9140 -3560 9540 -3080
rect 10180 -3560 10580 -3080
rect 11220 -3560 11620 -3080
rect 12260 -3560 12660 -3080
rect 13300 -3560 13700 -3080
rect 14340 -3560 14740 -3080
rect 15400 -3560 15800 -3080
rect 7560 -4780 7980 -4520
rect 8600 -4780 9020 -4520
rect 9640 -4780 10060 -4520
rect 10680 -4780 11100 -4520
rect 11720 -4780 12140 -4520
rect 12780 -4780 13200 -4520
rect 13800 -4780 14220 -4520
rect 14860 -4780 15280 -4520
rect 8100 -5820 8500 -5340
rect 9140 -5820 9540 -5340
rect 10180 -5820 10580 -5340
rect 11220 -5820 11620 -5340
rect 12260 -5820 12660 -5340
rect 13300 -5820 13700 -5340
rect 14340 -5820 14740 -5340
rect 7560 -6940 7980 -6800
rect 7560 -7060 7760 -6940
rect 7760 -7080 7900 -6940
rect 7900 -7060 7980 -6940
rect 8600 -6980 9020 -6800
rect 8600 -7060 8920 -6980
rect 8920 -7080 9020 -6980
rect 9640 -6980 10060 -6800
rect 9640 -7060 9960 -6980
rect 9960 -7080 10060 -6980
rect 10680 -6980 11100 -6800
rect 10680 -7060 11000 -6980
rect 11000 -7080 11100 -6980
rect 11720 -7060 12140 -6800
rect 12780 -6980 13200 -6800
rect 12780 -7060 13080 -6980
rect 13080 -7080 13180 -6980
rect 13180 -7060 13200 -6980
rect 13800 -6980 14220 -6800
rect 13800 -7060 14120 -6980
rect 14120 -7080 14220 -6980
rect 14860 -7060 15280 -6800
<< metal3 >>
rect 6880 6400 16100 6720
rect 6890 2160 16150 2165
rect 6890 1820 6900 2160
rect 16140 1820 16150 2160
rect 6890 1815 16150 1820
rect 7060 1405 7460 1815
rect 8100 1405 8500 1815
rect 9140 1405 9540 1815
rect 10180 1405 10580 1815
rect 11220 1405 11620 1815
rect 12260 1405 12660 1815
rect 13300 1405 13700 1815
rect 14340 1405 14740 1815
rect 15420 1405 15820 1815
rect 7050 1400 7470 1405
rect 7050 920 7060 1400
rect 7460 920 7470 1400
rect 7050 915 7470 920
rect 8090 1400 8510 1405
rect 8090 920 8100 1400
rect 8500 920 8510 1400
rect 8090 915 8510 920
rect 9130 1400 9550 1405
rect 9130 920 9140 1400
rect 9540 920 9550 1400
rect 9130 915 9550 920
rect 10170 1400 10590 1405
rect 10170 920 10180 1400
rect 10580 920 10590 1400
rect 10170 915 10590 920
rect 11210 1400 11630 1405
rect 11210 920 11220 1400
rect 11620 920 11630 1400
rect 11210 915 11630 920
rect 12250 1400 12670 1405
rect 12250 920 12260 1400
rect 12660 920 12670 1400
rect 12250 915 12670 920
rect 13290 1400 13710 1405
rect 13290 920 13300 1400
rect 13700 920 13710 1400
rect 13290 915 13710 920
rect 14330 1400 14750 1405
rect 14330 920 14340 1400
rect 14740 920 14750 1400
rect 14330 915 14750 920
rect 15390 1400 15820 1405
rect 15390 920 15400 1400
rect 15800 920 15820 1400
rect 15390 915 15820 920
rect 7060 -855 7460 915
rect 7540 -40 8000 0
rect 7540 -300 7560 -40
rect 7980 -300 8000 -40
rect 7050 -860 7470 -855
rect 7050 -1340 7060 -860
rect 7460 -1340 7470 -860
rect 7050 -1345 7470 -1340
rect 7060 -3075 7460 -1345
rect 7540 -2280 8000 -300
rect 8100 -855 8500 915
rect 8580 -40 9040 0
rect 8580 -300 8600 -40
rect 9020 -300 9040 -40
rect 8090 -860 8510 -855
rect 8090 -1340 8100 -860
rect 8500 -1340 8510 -860
rect 8090 -1345 8510 -1340
rect 7540 -2540 7560 -2280
rect 7980 -2540 8000 -2280
rect 7050 -3080 7470 -3075
rect 7050 -3560 7060 -3080
rect 7460 -3560 7470 -3080
rect 7050 -3565 7470 -3560
rect 7060 -3580 7460 -3565
rect 7540 -4520 8000 -2540
rect 8100 -3075 8500 -1345
rect 8580 -2280 9040 -300
rect 9140 -855 9540 915
rect 9620 -40 10080 0
rect 9620 -300 9640 -40
rect 10060 -300 10080 -40
rect 9130 -860 9550 -855
rect 9130 -1340 9140 -860
rect 9540 -1340 9550 -860
rect 9130 -1345 9550 -1340
rect 8580 -2540 8600 -2280
rect 9020 -2540 9040 -2280
rect 8090 -3080 8510 -3075
rect 8090 -3560 8100 -3080
rect 8500 -3560 8510 -3080
rect 8090 -3565 8510 -3560
rect 7540 -4780 7560 -4520
rect 7980 -4780 8000 -4520
rect 7540 -6800 8000 -4780
rect 8100 -5335 8500 -3565
rect 8580 -4520 9040 -2540
rect 9140 -3075 9540 -1345
rect 9620 -2280 10080 -300
rect 10180 -855 10580 915
rect 10660 -40 11120 0
rect 10660 -300 10680 -40
rect 11100 -300 11120 -40
rect 10170 -860 10590 -855
rect 10170 -1340 10180 -860
rect 10580 -1340 10590 -860
rect 10170 -1345 10590 -1340
rect 9620 -2540 9640 -2280
rect 10060 -2540 10080 -2280
rect 9130 -3080 9550 -3075
rect 9130 -3560 9140 -3080
rect 9540 -3560 9550 -3080
rect 9130 -3565 9550 -3560
rect 8580 -4780 8600 -4520
rect 9020 -4780 9040 -4520
rect 8090 -5340 8510 -5335
rect 8090 -5820 8100 -5340
rect 8500 -5820 8510 -5340
rect 8090 -5825 8510 -5820
rect 8580 -6800 9040 -4780
rect 9140 -5335 9540 -3565
rect 9620 -4520 10080 -2540
rect 10180 -3075 10580 -1345
rect 10660 -2280 11120 -300
rect 11220 -855 11620 915
rect 11700 -40 12160 0
rect 11700 -300 11720 -40
rect 12140 -300 12160 -40
rect 11210 -860 11630 -855
rect 11210 -1340 11220 -860
rect 11620 -1340 11630 -860
rect 11210 -1345 11630 -1340
rect 10660 -2540 10680 -2280
rect 11100 -2540 11120 -2280
rect 10170 -3080 10590 -3075
rect 10170 -3560 10180 -3080
rect 10580 -3560 10590 -3080
rect 10170 -3565 10590 -3560
rect 9620 -4780 9640 -4520
rect 10060 -4780 10080 -4520
rect 9130 -5340 9550 -5335
rect 9130 -5820 9140 -5340
rect 9540 -5820 9550 -5340
rect 9130 -5825 9550 -5820
rect 9620 -6800 10080 -4780
rect 10180 -5335 10580 -3565
rect 10660 -4520 11120 -2540
rect 11220 -3075 11620 -1345
rect 11700 -2280 12160 -300
rect 12260 -855 12660 915
rect 12760 -40 13220 0
rect 12760 -300 12780 -40
rect 13200 -300 13220 -40
rect 12250 -860 12670 -855
rect 12250 -1340 12260 -860
rect 12660 -1340 12670 -860
rect 12250 -1345 12670 -1340
rect 11700 -2540 11720 -2280
rect 12140 -2540 12160 -2280
rect 11210 -3080 11630 -3075
rect 11210 -3560 11220 -3080
rect 11620 -3560 11630 -3080
rect 11210 -3565 11630 -3560
rect 10660 -4780 10680 -4520
rect 11100 -4780 11120 -4520
rect 10170 -5340 10590 -5335
rect 10170 -5820 10180 -5340
rect 10580 -5820 10590 -5340
rect 10170 -5825 10590 -5820
rect 10660 -6800 11120 -4780
rect 11220 -5335 11620 -3565
rect 11700 -4520 12160 -2540
rect 12260 -3075 12660 -1345
rect 12760 -2280 13220 -300
rect 13300 -855 13700 915
rect 13780 -40 14240 0
rect 13780 -300 13800 -40
rect 14220 -300 14240 -40
rect 13290 -860 13710 -855
rect 13290 -1340 13300 -860
rect 13700 -1340 13710 -860
rect 13290 -1345 13710 -1340
rect 12760 -2540 12780 -2280
rect 13200 -2540 13220 -2280
rect 12250 -3080 12670 -3075
rect 12250 -3560 12260 -3080
rect 12660 -3560 12670 -3080
rect 12250 -3565 12670 -3560
rect 11700 -4780 11720 -4520
rect 12140 -4780 12160 -4520
rect 11210 -5340 11630 -5335
rect 11210 -5820 11220 -5340
rect 11620 -5820 11630 -5340
rect 11210 -5825 11630 -5820
rect 11700 -6800 12160 -4780
rect 12260 -5335 12660 -3565
rect 12760 -4520 13220 -2540
rect 13300 -3075 13700 -1345
rect 13780 -2280 14240 -300
rect 14340 -855 14740 915
rect 14840 -40 15300 0
rect 14840 -300 14860 -40
rect 15280 -300 15300 -40
rect 14330 -860 14750 -855
rect 14330 -1340 14340 -860
rect 14740 -1340 14750 -860
rect 14330 -1345 14750 -1340
rect 13780 -2540 13800 -2280
rect 14220 -2540 14240 -2280
rect 13290 -3080 13710 -3075
rect 13290 -3560 13300 -3080
rect 13700 -3560 13710 -3080
rect 13290 -3565 13710 -3560
rect 12760 -4780 12780 -4520
rect 13200 -4780 13220 -4520
rect 12250 -5340 12670 -5335
rect 12250 -5820 12260 -5340
rect 12660 -5820 12670 -5340
rect 12250 -5825 12670 -5820
rect 12760 -6800 13220 -4780
rect 13300 -5335 13700 -3565
rect 13780 -4520 14240 -2540
rect 14340 -3075 14740 -1345
rect 14840 -2280 15300 -300
rect 15420 -855 15820 915
rect 15390 -860 15820 -855
rect 15390 -1340 15400 -860
rect 15800 -1340 15820 -860
rect 15390 -1345 15820 -1340
rect 14840 -2540 14860 -2280
rect 15280 -2540 15300 -2280
rect 14330 -3080 14750 -3075
rect 14330 -3560 14340 -3080
rect 14740 -3560 14750 -3080
rect 14330 -3565 14750 -3560
rect 13780 -4780 13800 -4520
rect 14220 -4780 14240 -4520
rect 13290 -5340 13710 -5335
rect 13290 -5820 13300 -5340
rect 13700 -5820 13710 -5340
rect 13290 -5825 13710 -5820
rect 13780 -6800 14240 -4780
rect 14340 -5335 14740 -3565
rect 14840 -4520 15300 -2540
rect 15420 -3075 15820 -1345
rect 15390 -3080 15820 -3075
rect 15390 -3560 15400 -3080
rect 15800 -3560 15820 -3080
rect 15390 -3565 15820 -3560
rect 15420 -3580 15820 -3565
rect 14840 -4780 14860 -4520
rect 15280 -4780 15300 -4520
rect 14330 -5340 14750 -5335
rect 14330 -5820 14340 -5340
rect 14740 -5820 14750 -5340
rect 14330 -5825 14750 -5820
rect 14840 -6800 15300 -4780
rect 7540 -7060 7560 -6800
rect 7980 -7060 8600 -6800
rect 9020 -7060 9640 -6800
rect 10060 -7060 10680 -6800
rect 11100 -7060 11720 -6800
rect 12140 -7060 12780 -6800
rect 13200 -7060 13800 -6800
rect 14220 -7060 14860 -6800
rect 15280 -7060 15300 -6800
rect 7540 -7080 7760 -7060
rect 7900 -7080 8920 -7060
rect 9020 -7080 9960 -7060
rect 10060 -7080 11000 -7060
rect 11100 -7080 13080 -7060
rect 13180 -7080 14120 -7060
rect 14220 -7080 15300 -7060
rect 7540 -7100 15300 -7080
use outd_curm  outd_curm_25
timestamp 1683888831
transform 1 0 9966 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_26
timestamp 1683888831
transform 1 0 8924 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_27
timestamp 1683888831
transform 1 0 6840 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_28
timestamp 1683888831
transform 1 0 7882 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_29
timestamp 1683888831
transform 1 0 14134 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_30
timestamp 1683888831
transform 1 0 13092 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_31
timestamp 1683888831
transform 1 0 12050 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_32
timestamp 1683888831
transform 1 0 11008 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_33
timestamp 1683888831
transform 1 0 15176 0 1 -5774
box -40 916 1002 3158
use outd_curm  outd_curm_34
timestamp 1683888831
transform 1 0 6840 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_35
timestamp 1683888831
transform 1 0 7882 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_36
timestamp 1683888831
transform 1 0 8924 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_37
timestamp 1683888831
transform 1 0 9966 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_38
timestamp 1683888831
transform 1 0 11008 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_39
timestamp 1683888831
transform 1 0 12050 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_40
timestamp 1683888831
transform 1 0 13092 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_41
timestamp 1683888831
transform 1 0 14134 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_42
timestamp 1683888831
transform 1 0 9966 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_43
timestamp 1683888831
transform 1 0 9966 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_44
timestamp 1683888831
transform 1 0 8924 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_46
timestamp 1683888831
transform 1 0 7882 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_47
timestamp 1683888831
transform 1 0 14134 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_48
timestamp 1683888831
transform 1 0 13092 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_49
timestamp 1683888831
transform 1 0 12050 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_50
timestamp 1683888831
transform 1 0 11008 0 1 -8016
box -40 916 1002 3158
use outd_curm  outd_curm_52
timestamp 1683888831
transform 1 0 8924 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_53
timestamp 1683888831
transform 1 0 6840 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_54
timestamp 1683888831
transform 1 0 7882 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_55
timestamp 1683888831
transform 1 0 14134 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_56
timestamp 1683888831
transform 1 0 13092 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_57
timestamp 1683888831
transform 1 0 12050 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_58
timestamp 1683888831
transform 1 0 11008 0 1 -1294
box -40 916 1002 3158
use outd_curm  outd_curm_59
timestamp 1683888831
transform 1 0 15176 0 1 -3536
box -40 916 1002 3158
use outd_curm  outd_curm_60
timestamp 1683888831
transform 1 0 15176 0 1 -1294
box -40 916 1002 3158
use outd_diffamp_50ohm  outd_diffamp_50ohm_0
timestamp 1687116508
transform 1 0 12000 0 1 2680
box 0 -820 4174 4040
use outd_diffamp_50ohm  outd_diffamp_50ohm_1
timestamp 1687116508
transform 1 0 6800 0 1 2680
box 0 -820 4174 4040
use sky130_fd_pr__res_high_po_1p41_3FC2Y3  sky130_fd_pr__res_high_po_1p41_3FC2Y3_0
timestamp 1685111951
transform 1 0 11187 0 1 4562
box -307 -1882 307 1882
use sky130_fd_pr__res_high_po_1p41_3FC2Y3  sky130_fd_pr__res_high_po_1p41_3FC2Y3_1
timestamp 1685111951
transform 1 0 11787 0 1 4562
box -307 -1882 307 1882
<< end >>
