magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< nwell >>
rect -996 -319 996 319
<< pmos >>
rect -800 -100 800 100
<< pdiff >>
rect -858 88 -800 100
rect -858 -88 -846 88
rect -812 -88 -800 88
rect -858 -100 -800 -88
rect 800 88 858 100
rect 800 -88 812 88
rect 846 -88 858 88
rect 800 -100 858 -88
<< pdiffc >>
rect -846 -88 -812 88
rect 812 -88 846 88
<< nsubdiff >>
rect -960 249 -864 283
rect 864 249 960 283
rect -960 187 -926 249
rect 926 187 960 249
rect -960 -249 -926 -187
rect 926 -249 960 -187
rect -960 -283 -864 -249
rect 864 -283 960 -249
<< nsubdiffcont >>
rect -864 249 864 283
rect -960 -187 -926 187
rect 926 -187 960 187
rect -864 -283 864 -249
<< poly >>
rect -800 181 800 197
rect -800 147 -784 181
rect 784 147 800 181
rect -800 100 800 147
rect -800 -147 800 -100
rect -800 -181 -784 -147
rect 784 -181 800 -147
rect -800 -197 800 -181
<< polycont >>
rect -784 147 784 181
rect -784 -181 784 -147
<< locali >>
rect -960 249 -864 283
rect 864 249 960 283
rect -960 187 -926 249
rect 926 187 960 249
rect -800 147 -784 181
rect 784 147 800 181
rect -846 88 -812 104
rect -846 -104 -812 -88
rect 812 88 846 104
rect 812 -104 846 -88
rect -800 -181 -784 -147
rect 784 -181 800 -147
rect -960 -249 -926 -187
rect 926 -249 960 -187
rect -960 -283 -864 -249
rect 864 -283 960 -249
<< viali >>
rect -784 147 784 181
rect -846 -88 -812 88
rect 812 -88 846 88
rect -784 -181 784 -147
<< metal1 >>
rect -796 181 796 187
rect -796 147 -784 181
rect 784 147 796 181
rect -796 141 796 147
rect -852 88 -806 100
rect -852 -88 -846 88
rect -812 -88 -806 88
rect -852 -100 -806 -88
rect 806 88 852 100
rect 806 -88 812 88
rect 846 -88 852 88
rect 806 -100 852 -88
rect -796 -147 796 -141
rect -796 -181 -784 -147
rect 784 -181 796 -147
rect -796 -187 796 -181
<< properties >>
string FIXED_BBOX -943 -266 943 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
