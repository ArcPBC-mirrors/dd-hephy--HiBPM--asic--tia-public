magic
tech sky130A
magscale 1 2
timestamp 1683801646
<< error_p >>
rect -173 1235 -115 1241
rect 19 1235 77 1241
rect -173 1201 -161 1235
rect 19 1201 31 1235
rect -173 1195 -115 1201
rect 19 1195 77 1201
rect -77 707 -19 713
rect 115 707 173 713
rect -77 673 -65 707
rect 115 673 127 707
rect -77 667 -19 673
rect 115 667 173 673
rect -77 599 -19 605
rect 115 599 173 605
rect -77 565 -65 599
rect 115 565 127 599
rect -77 559 -19 565
rect 115 559 173 565
rect -173 71 -115 77
rect 19 71 77 77
rect -173 37 -161 71
rect 19 37 31 71
rect -173 31 -115 37
rect 19 31 77 37
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect -77 -565 -19 -559
rect 115 -565 173 -559
rect -77 -599 -65 -565
rect 115 -599 127 -565
rect -77 -605 -19 -599
rect 115 -605 173 -599
rect -77 -673 -19 -667
rect 115 -673 173 -667
rect -77 -707 -65 -673
rect 115 -707 127 -673
rect -77 -713 -19 -707
rect 115 -713 173 -707
rect -173 -1201 -115 -1195
rect 19 -1201 77 -1195
rect -173 -1235 -161 -1201
rect 19 -1235 31 -1201
rect -173 -1241 -115 -1235
rect 19 -1241 77 -1235
<< nwell >>
rect -359 -1373 359 1373
<< pmos >>
rect -159 754 -129 1154
rect -63 754 -33 1154
rect 33 754 63 1154
rect 129 754 159 1154
rect -159 118 -129 518
rect -63 118 -33 518
rect 33 118 63 518
rect 129 118 159 518
rect -159 -518 -129 -118
rect -63 -518 -33 -118
rect 33 -518 63 -118
rect 129 -518 159 -118
rect -159 -1154 -129 -754
rect -63 -1154 -33 -754
rect 33 -1154 63 -754
rect 129 -1154 159 -754
<< pdiff >>
rect -221 1142 -159 1154
rect -221 766 -209 1142
rect -175 766 -159 1142
rect -221 754 -159 766
rect -129 1142 -63 1154
rect -129 766 -113 1142
rect -79 766 -63 1142
rect -129 754 -63 766
rect -33 1142 33 1154
rect -33 766 -17 1142
rect 17 766 33 1142
rect -33 754 33 766
rect 63 1142 129 1154
rect 63 766 79 1142
rect 113 766 129 1142
rect 63 754 129 766
rect 159 1142 221 1154
rect 159 766 175 1142
rect 209 766 221 1142
rect 159 754 221 766
rect -221 506 -159 518
rect -221 130 -209 506
rect -175 130 -159 506
rect -221 118 -159 130
rect -129 506 -63 518
rect -129 130 -113 506
rect -79 130 -63 506
rect -129 118 -63 130
rect -33 506 33 518
rect -33 130 -17 506
rect 17 130 33 506
rect -33 118 33 130
rect 63 506 129 518
rect 63 130 79 506
rect 113 130 129 506
rect 63 118 129 130
rect 159 506 221 518
rect 159 130 175 506
rect 209 130 221 506
rect 159 118 221 130
rect -221 -130 -159 -118
rect -221 -506 -209 -130
rect -175 -506 -159 -130
rect -221 -518 -159 -506
rect -129 -130 -63 -118
rect -129 -506 -113 -130
rect -79 -506 -63 -130
rect -129 -518 -63 -506
rect -33 -130 33 -118
rect -33 -506 -17 -130
rect 17 -506 33 -130
rect -33 -518 33 -506
rect 63 -130 129 -118
rect 63 -506 79 -130
rect 113 -506 129 -130
rect 63 -518 129 -506
rect 159 -130 221 -118
rect 159 -506 175 -130
rect 209 -506 221 -130
rect 159 -518 221 -506
rect -221 -766 -159 -754
rect -221 -1142 -209 -766
rect -175 -1142 -159 -766
rect -221 -1154 -159 -1142
rect -129 -766 -63 -754
rect -129 -1142 -113 -766
rect -79 -1142 -63 -766
rect -129 -1154 -63 -1142
rect -33 -766 33 -754
rect -33 -1142 -17 -766
rect 17 -1142 33 -766
rect -33 -1154 33 -1142
rect 63 -766 129 -754
rect 63 -1142 79 -766
rect 113 -1142 129 -766
rect 63 -1154 129 -1142
rect 159 -766 221 -754
rect 159 -1142 175 -766
rect 209 -1142 221 -766
rect 159 -1154 221 -1142
<< pdiffc >>
rect -209 766 -175 1142
rect -113 766 -79 1142
rect -17 766 17 1142
rect 79 766 113 1142
rect 175 766 209 1142
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect -209 -1142 -175 -766
rect -113 -1142 -79 -766
rect -17 -1142 17 -766
rect 79 -1142 113 -766
rect 175 -1142 209 -766
<< nsubdiff >>
rect -323 1303 -227 1337
rect 227 1303 323 1337
rect -323 1241 -289 1303
rect 289 1241 323 1303
rect -323 -1303 -289 -1241
rect 289 -1303 323 -1241
rect -323 -1337 -227 -1303
rect 227 -1337 323 -1303
<< nsubdiffcont >>
rect -227 1303 227 1337
rect -323 -1241 -289 1241
rect 289 -1241 323 1241
rect -227 -1337 227 -1303
<< poly >>
rect -177 1235 -111 1251
rect -177 1201 -161 1235
rect -127 1201 -111 1235
rect -177 1185 -111 1201
rect 15 1235 81 1251
rect 15 1201 31 1235
rect 65 1201 81 1235
rect 15 1185 81 1201
rect -159 1154 -129 1185
rect -63 1154 -33 1180
rect 33 1154 63 1185
rect 129 1154 159 1180
rect -159 728 -129 754
rect -63 723 -33 754
rect 33 728 63 754
rect 129 723 159 754
rect -81 707 -15 723
rect -81 673 -65 707
rect -31 673 -15 707
rect -81 657 -15 673
rect 111 707 177 723
rect 111 673 127 707
rect 161 673 177 707
rect 111 657 177 673
rect -81 599 -15 615
rect -81 565 -65 599
rect -31 565 -15 599
rect -81 549 -15 565
rect 111 599 177 615
rect 111 565 127 599
rect 161 565 177 599
rect 111 549 177 565
rect -159 518 -129 544
rect -63 518 -33 549
rect 33 518 63 544
rect 129 518 159 549
rect -159 87 -129 118
rect -63 92 -33 118
rect 33 87 63 118
rect 129 92 159 118
rect -177 71 -111 87
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect -159 -118 -129 -87
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect 129 -118 159 -92
rect -159 -544 -129 -518
rect -63 -549 -33 -518
rect 33 -544 63 -518
rect 129 -549 159 -518
rect -81 -565 -15 -549
rect -81 -599 -65 -565
rect -31 -599 -15 -565
rect -81 -615 -15 -599
rect 111 -565 177 -549
rect 111 -599 127 -565
rect 161 -599 177 -565
rect 111 -615 177 -599
rect -81 -673 -15 -657
rect -81 -707 -65 -673
rect -31 -707 -15 -673
rect -81 -723 -15 -707
rect 111 -673 177 -657
rect 111 -707 127 -673
rect 161 -707 177 -673
rect 111 -723 177 -707
rect -159 -754 -129 -728
rect -63 -754 -33 -723
rect 33 -754 63 -728
rect 129 -754 159 -723
rect -159 -1185 -129 -1154
rect -63 -1180 -33 -1154
rect 33 -1185 63 -1154
rect 129 -1180 159 -1154
rect -177 -1201 -111 -1185
rect -177 -1235 -161 -1201
rect -127 -1235 -111 -1201
rect -177 -1251 -111 -1235
rect 15 -1201 81 -1185
rect 15 -1235 31 -1201
rect 65 -1235 81 -1201
rect 15 -1251 81 -1235
<< polycont >>
rect -161 1201 -127 1235
rect 31 1201 65 1235
rect -65 673 -31 707
rect 127 673 161 707
rect -65 565 -31 599
rect 127 565 161 599
rect -161 37 -127 71
rect 31 37 65 71
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect -65 -599 -31 -565
rect 127 -599 161 -565
rect -65 -707 -31 -673
rect 127 -707 161 -673
rect -161 -1235 -127 -1201
rect 31 -1235 65 -1201
<< locali >>
rect -323 1303 -227 1337
rect 227 1303 323 1337
rect -323 1241 -289 1303
rect 289 1241 323 1303
rect -177 1201 -161 1235
rect -127 1201 -111 1235
rect 15 1201 31 1235
rect 65 1201 81 1235
rect -209 1142 -175 1158
rect -209 750 -175 766
rect -113 1142 -79 1158
rect -113 750 -79 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 79 1142 113 1158
rect 79 750 113 766
rect 175 1142 209 1158
rect 175 750 209 766
rect -81 673 -65 707
rect -31 673 -15 707
rect 111 673 127 707
rect 161 673 177 707
rect -81 565 -65 599
rect -31 565 -15 599
rect 111 565 127 599
rect 161 565 177 599
rect -209 506 -175 522
rect -209 114 -175 130
rect -113 506 -79 522
rect -113 114 -79 130
rect -17 506 17 522
rect -17 114 17 130
rect 79 506 113 522
rect 79 114 113 130
rect 175 506 209 522
rect 175 114 209 130
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -209 -130 -175 -114
rect -209 -522 -175 -506
rect -113 -130 -79 -114
rect -113 -522 -79 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 79 -130 113 -114
rect 79 -522 113 -506
rect 175 -130 209 -114
rect 175 -522 209 -506
rect -81 -599 -65 -565
rect -31 -599 -15 -565
rect 111 -599 127 -565
rect 161 -599 177 -565
rect -81 -707 -65 -673
rect -31 -707 -15 -673
rect 111 -707 127 -673
rect 161 -707 177 -673
rect -209 -766 -175 -750
rect -209 -1158 -175 -1142
rect -113 -766 -79 -750
rect -113 -1158 -79 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 79 -766 113 -750
rect 79 -1158 113 -1142
rect 175 -766 209 -750
rect 175 -1158 209 -1142
rect -177 -1235 -161 -1201
rect -127 -1235 -111 -1201
rect 15 -1235 31 -1201
rect 65 -1235 81 -1201
rect -323 -1303 -289 -1241
rect 289 -1303 323 -1241
rect -323 -1337 -227 -1303
rect 227 -1337 323 -1303
<< viali >>
rect -161 1201 -127 1235
rect 31 1201 65 1235
rect -209 766 -175 1142
rect -113 766 -79 1142
rect -17 766 17 1142
rect 79 766 113 1142
rect 175 766 209 1142
rect -65 673 -31 707
rect 127 673 161 707
rect -65 565 -31 599
rect 127 565 161 599
rect -209 130 -175 506
rect -113 130 -79 506
rect -17 130 17 506
rect 79 130 113 506
rect 175 130 209 506
rect -161 37 -127 71
rect 31 37 65 71
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect -209 -506 -175 -130
rect -113 -506 -79 -130
rect -17 -506 17 -130
rect 79 -506 113 -130
rect 175 -506 209 -130
rect -65 -599 -31 -565
rect 127 -599 161 -565
rect -65 -707 -31 -673
rect 127 -707 161 -673
rect -209 -1142 -175 -766
rect -113 -1142 -79 -766
rect -17 -1142 17 -766
rect 79 -1142 113 -766
rect 175 -1142 209 -766
rect -161 -1235 -127 -1201
rect 31 -1235 65 -1201
<< metal1 >>
rect -173 1235 -115 1241
rect -173 1201 -161 1235
rect -127 1201 -115 1235
rect -173 1195 -115 1201
rect 19 1235 77 1241
rect 19 1201 31 1235
rect 65 1201 77 1235
rect 19 1195 77 1201
rect -215 1142 -169 1154
rect -215 766 -209 1142
rect -175 766 -169 1142
rect -215 754 -169 766
rect -119 1142 -73 1154
rect -119 766 -113 1142
rect -79 766 -73 1142
rect -119 754 -73 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 73 1142 119 1154
rect 73 766 79 1142
rect 113 766 119 1142
rect 73 754 119 766
rect 169 1142 215 1154
rect 169 766 175 1142
rect 209 766 215 1142
rect 169 754 215 766
rect -77 707 -19 713
rect -77 673 -65 707
rect -31 673 -19 707
rect -77 667 -19 673
rect 115 707 173 713
rect 115 673 127 707
rect 161 673 173 707
rect 115 667 173 673
rect -77 599 -19 605
rect -77 565 -65 599
rect -31 565 -19 599
rect -77 559 -19 565
rect 115 599 173 605
rect 115 565 127 599
rect 161 565 173 599
rect 115 559 173 565
rect -215 506 -169 518
rect -215 130 -209 506
rect -175 130 -169 506
rect -215 118 -169 130
rect -119 506 -73 518
rect -119 130 -113 506
rect -79 130 -73 506
rect -119 118 -73 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 73 506 119 518
rect 73 130 79 506
rect 113 130 119 506
rect 73 118 119 130
rect 169 506 215 518
rect 169 130 175 506
rect 209 130 215 506
rect 169 118 215 130
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect -215 -130 -169 -118
rect -215 -506 -209 -130
rect -175 -506 -169 -130
rect -215 -518 -169 -506
rect -119 -130 -73 -118
rect -119 -506 -113 -130
rect -79 -506 -73 -130
rect -119 -518 -73 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 73 -130 119 -118
rect 73 -506 79 -130
rect 113 -506 119 -130
rect 73 -518 119 -506
rect 169 -130 215 -118
rect 169 -506 175 -130
rect 209 -506 215 -130
rect 169 -518 215 -506
rect -77 -565 -19 -559
rect -77 -599 -65 -565
rect -31 -599 -19 -565
rect -77 -605 -19 -599
rect 115 -565 173 -559
rect 115 -599 127 -565
rect 161 -599 173 -565
rect 115 -605 173 -599
rect -77 -673 -19 -667
rect -77 -707 -65 -673
rect -31 -707 -19 -673
rect -77 -713 -19 -707
rect 115 -673 173 -667
rect 115 -707 127 -673
rect 161 -707 173 -673
rect 115 -713 173 -707
rect -215 -766 -169 -754
rect -215 -1142 -209 -766
rect -175 -1142 -169 -766
rect -215 -1154 -169 -1142
rect -119 -766 -73 -754
rect -119 -1142 -113 -766
rect -79 -1142 -73 -766
rect -119 -1154 -73 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 73 -766 119 -754
rect 73 -1142 79 -766
rect 113 -1142 119 -766
rect 73 -1154 119 -1142
rect 169 -766 215 -754
rect 169 -1142 175 -766
rect 209 -1142 215 -766
rect 169 -1154 215 -1142
rect -173 -1201 -115 -1195
rect -173 -1235 -161 -1201
rect -127 -1235 -115 -1201
rect -173 -1241 -115 -1235
rect 19 -1201 77 -1195
rect 19 -1235 31 -1201
rect 65 -1235 77 -1201
rect 19 -1241 77 -1235
<< properties >>
string FIXED_BBOX -306 -1320 306 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
