magic
tech sky130A
magscale 1 2
timestamp 1683737876
<< error_p >>
rect -1133 3053 -1075 3059
rect -941 3053 -883 3059
rect -749 3053 -691 3059
rect -557 3053 -499 3059
rect -365 3053 -307 3059
rect -173 3053 -115 3059
rect 19 3053 77 3059
rect 211 3053 269 3059
rect 403 3053 461 3059
rect 595 3053 653 3059
rect 787 3053 845 3059
rect 979 3053 1037 3059
rect -1133 3019 -1121 3053
rect -941 3019 -929 3053
rect -749 3019 -737 3053
rect -557 3019 -545 3053
rect -365 3019 -353 3053
rect -173 3019 -161 3053
rect 19 3019 31 3053
rect 211 3019 223 3053
rect 403 3019 415 3053
rect 595 3019 607 3053
rect 787 3019 799 3053
rect 979 3019 991 3053
rect -1133 3013 -1075 3019
rect -941 3013 -883 3019
rect -749 3013 -691 3019
rect -557 3013 -499 3019
rect -365 3013 -307 3019
rect -173 3013 -115 3019
rect 19 3013 77 3019
rect 211 3013 269 3019
rect 403 3013 461 3019
rect 595 3013 653 3019
rect 787 3013 845 3019
rect 979 3013 1037 3019
rect -1037 2543 -979 2549
rect -845 2543 -787 2549
rect -653 2543 -595 2549
rect -461 2543 -403 2549
rect -269 2543 -211 2549
rect -77 2543 -19 2549
rect 115 2543 173 2549
rect 307 2543 365 2549
rect 499 2543 557 2549
rect 691 2543 749 2549
rect 883 2543 941 2549
rect 1075 2543 1133 2549
rect -1037 2509 -1025 2543
rect -845 2509 -833 2543
rect -653 2509 -641 2543
rect -461 2509 -449 2543
rect -269 2509 -257 2543
rect -77 2509 -65 2543
rect 115 2509 127 2543
rect 307 2509 319 2543
rect 499 2509 511 2543
rect 691 2509 703 2543
rect 883 2509 895 2543
rect 1075 2509 1087 2543
rect -1037 2503 -979 2509
rect -845 2503 -787 2509
rect -653 2503 -595 2509
rect -461 2503 -403 2509
rect -269 2503 -211 2509
rect -77 2503 -19 2509
rect 115 2503 173 2509
rect 307 2503 365 2509
rect 499 2503 557 2509
rect 691 2503 749 2509
rect 883 2503 941 2509
rect 1075 2503 1133 2509
rect -1037 2435 -979 2441
rect -845 2435 -787 2441
rect -653 2435 -595 2441
rect -461 2435 -403 2441
rect -269 2435 -211 2441
rect -77 2435 -19 2441
rect 115 2435 173 2441
rect 307 2435 365 2441
rect 499 2435 557 2441
rect 691 2435 749 2441
rect 883 2435 941 2441
rect 1075 2435 1133 2441
rect -1037 2401 -1025 2435
rect -845 2401 -833 2435
rect -653 2401 -641 2435
rect -461 2401 -449 2435
rect -269 2401 -257 2435
rect -77 2401 -65 2435
rect 115 2401 127 2435
rect 307 2401 319 2435
rect 499 2401 511 2435
rect 691 2401 703 2435
rect 883 2401 895 2435
rect 1075 2401 1087 2435
rect -1037 2395 -979 2401
rect -845 2395 -787 2401
rect -653 2395 -595 2401
rect -461 2395 -403 2401
rect -269 2395 -211 2401
rect -77 2395 -19 2401
rect 115 2395 173 2401
rect 307 2395 365 2401
rect 499 2395 557 2401
rect 691 2395 749 2401
rect 883 2395 941 2401
rect 1075 2395 1133 2401
rect -1133 1925 -1075 1931
rect -941 1925 -883 1931
rect -749 1925 -691 1931
rect -557 1925 -499 1931
rect -365 1925 -307 1931
rect -173 1925 -115 1931
rect 19 1925 77 1931
rect 211 1925 269 1931
rect 403 1925 461 1931
rect 595 1925 653 1931
rect 787 1925 845 1931
rect 979 1925 1037 1931
rect -1133 1891 -1121 1925
rect -941 1891 -929 1925
rect -749 1891 -737 1925
rect -557 1891 -545 1925
rect -365 1891 -353 1925
rect -173 1891 -161 1925
rect 19 1891 31 1925
rect 211 1891 223 1925
rect 403 1891 415 1925
rect 595 1891 607 1925
rect 787 1891 799 1925
rect 979 1891 991 1925
rect -1133 1885 -1075 1891
rect -941 1885 -883 1891
rect -749 1885 -691 1891
rect -557 1885 -499 1891
rect -365 1885 -307 1891
rect -173 1885 -115 1891
rect 19 1885 77 1891
rect 211 1885 269 1891
rect 403 1885 461 1891
rect 595 1885 653 1891
rect 787 1885 845 1891
rect 979 1885 1037 1891
rect -1133 1817 -1075 1823
rect -941 1817 -883 1823
rect -749 1817 -691 1823
rect -557 1817 -499 1823
rect -365 1817 -307 1823
rect -173 1817 -115 1823
rect 19 1817 77 1823
rect 211 1817 269 1823
rect 403 1817 461 1823
rect 595 1817 653 1823
rect 787 1817 845 1823
rect 979 1817 1037 1823
rect -1133 1783 -1121 1817
rect -941 1783 -929 1817
rect -749 1783 -737 1817
rect -557 1783 -545 1817
rect -365 1783 -353 1817
rect -173 1783 -161 1817
rect 19 1783 31 1817
rect 211 1783 223 1817
rect 403 1783 415 1817
rect 595 1783 607 1817
rect 787 1783 799 1817
rect 979 1783 991 1817
rect -1133 1777 -1075 1783
rect -941 1777 -883 1783
rect -749 1777 -691 1783
rect -557 1777 -499 1783
rect -365 1777 -307 1783
rect -173 1777 -115 1783
rect 19 1777 77 1783
rect 211 1777 269 1783
rect 403 1777 461 1783
rect 595 1777 653 1783
rect 787 1777 845 1783
rect 979 1777 1037 1783
rect -1037 1307 -979 1313
rect -845 1307 -787 1313
rect -653 1307 -595 1313
rect -461 1307 -403 1313
rect -269 1307 -211 1313
rect -77 1307 -19 1313
rect 115 1307 173 1313
rect 307 1307 365 1313
rect 499 1307 557 1313
rect 691 1307 749 1313
rect 883 1307 941 1313
rect 1075 1307 1133 1313
rect -1037 1273 -1025 1307
rect -845 1273 -833 1307
rect -653 1273 -641 1307
rect -461 1273 -449 1307
rect -269 1273 -257 1307
rect -77 1273 -65 1307
rect 115 1273 127 1307
rect 307 1273 319 1307
rect 499 1273 511 1307
rect 691 1273 703 1307
rect 883 1273 895 1307
rect 1075 1273 1087 1307
rect -1037 1267 -979 1273
rect -845 1267 -787 1273
rect -653 1267 -595 1273
rect -461 1267 -403 1273
rect -269 1267 -211 1273
rect -77 1267 -19 1273
rect 115 1267 173 1273
rect 307 1267 365 1273
rect 499 1267 557 1273
rect 691 1267 749 1273
rect 883 1267 941 1273
rect 1075 1267 1133 1273
rect -1037 1199 -979 1205
rect -845 1199 -787 1205
rect -653 1199 -595 1205
rect -461 1199 -403 1205
rect -269 1199 -211 1205
rect -77 1199 -19 1205
rect 115 1199 173 1205
rect 307 1199 365 1205
rect 499 1199 557 1205
rect 691 1199 749 1205
rect 883 1199 941 1205
rect 1075 1199 1133 1205
rect -1037 1165 -1025 1199
rect -845 1165 -833 1199
rect -653 1165 -641 1199
rect -461 1165 -449 1199
rect -269 1165 -257 1199
rect -77 1165 -65 1199
rect 115 1165 127 1199
rect 307 1165 319 1199
rect 499 1165 511 1199
rect 691 1165 703 1199
rect 883 1165 895 1199
rect 1075 1165 1087 1199
rect -1037 1159 -979 1165
rect -845 1159 -787 1165
rect -653 1159 -595 1165
rect -461 1159 -403 1165
rect -269 1159 -211 1165
rect -77 1159 -19 1165
rect 115 1159 173 1165
rect 307 1159 365 1165
rect 499 1159 557 1165
rect 691 1159 749 1165
rect 883 1159 941 1165
rect 1075 1159 1133 1165
rect -1133 689 -1075 695
rect -941 689 -883 695
rect -749 689 -691 695
rect -557 689 -499 695
rect -365 689 -307 695
rect -173 689 -115 695
rect 19 689 77 695
rect 211 689 269 695
rect 403 689 461 695
rect 595 689 653 695
rect 787 689 845 695
rect 979 689 1037 695
rect -1133 655 -1121 689
rect -941 655 -929 689
rect -749 655 -737 689
rect -557 655 -545 689
rect -365 655 -353 689
rect -173 655 -161 689
rect 19 655 31 689
rect 211 655 223 689
rect 403 655 415 689
rect 595 655 607 689
rect 787 655 799 689
rect 979 655 991 689
rect -1133 649 -1075 655
rect -941 649 -883 655
rect -749 649 -691 655
rect -557 649 -499 655
rect -365 649 -307 655
rect -173 649 -115 655
rect 19 649 77 655
rect 211 649 269 655
rect 403 649 461 655
rect 595 649 653 655
rect 787 649 845 655
rect 979 649 1037 655
rect -1133 581 -1075 587
rect -941 581 -883 587
rect -749 581 -691 587
rect -557 581 -499 587
rect -365 581 -307 587
rect -173 581 -115 587
rect 19 581 77 587
rect 211 581 269 587
rect 403 581 461 587
rect 595 581 653 587
rect 787 581 845 587
rect 979 581 1037 587
rect -1133 547 -1121 581
rect -941 547 -929 581
rect -749 547 -737 581
rect -557 547 -545 581
rect -365 547 -353 581
rect -173 547 -161 581
rect 19 547 31 581
rect 211 547 223 581
rect 403 547 415 581
rect 595 547 607 581
rect 787 547 799 581
rect 979 547 991 581
rect -1133 541 -1075 547
rect -941 541 -883 547
rect -749 541 -691 547
rect -557 541 -499 547
rect -365 541 -307 547
rect -173 541 -115 547
rect 19 541 77 547
rect 211 541 269 547
rect 403 541 461 547
rect 595 541 653 547
rect 787 541 845 547
rect 979 541 1037 547
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect -1133 -547 -1075 -541
rect -941 -547 -883 -541
rect -749 -547 -691 -541
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect 595 -547 653 -541
rect 787 -547 845 -541
rect 979 -547 1037 -541
rect -1133 -581 -1121 -547
rect -941 -581 -929 -547
rect -749 -581 -737 -547
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect 595 -581 607 -547
rect 787 -581 799 -547
rect 979 -581 991 -547
rect -1133 -587 -1075 -581
rect -941 -587 -883 -581
rect -749 -587 -691 -581
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
rect 595 -587 653 -581
rect 787 -587 845 -581
rect 979 -587 1037 -581
rect -1133 -655 -1075 -649
rect -941 -655 -883 -649
rect -749 -655 -691 -649
rect -557 -655 -499 -649
rect -365 -655 -307 -649
rect -173 -655 -115 -649
rect 19 -655 77 -649
rect 211 -655 269 -649
rect 403 -655 461 -649
rect 595 -655 653 -649
rect 787 -655 845 -649
rect 979 -655 1037 -649
rect -1133 -689 -1121 -655
rect -941 -689 -929 -655
rect -749 -689 -737 -655
rect -557 -689 -545 -655
rect -365 -689 -353 -655
rect -173 -689 -161 -655
rect 19 -689 31 -655
rect 211 -689 223 -655
rect 403 -689 415 -655
rect 595 -689 607 -655
rect 787 -689 799 -655
rect 979 -689 991 -655
rect -1133 -695 -1075 -689
rect -941 -695 -883 -689
rect -749 -695 -691 -689
rect -557 -695 -499 -689
rect -365 -695 -307 -689
rect -173 -695 -115 -689
rect 19 -695 77 -689
rect 211 -695 269 -689
rect 403 -695 461 -689
rect 595 -695 653 -689
rect 787 -695 845 -689
rect 979 -695 1037 -689
rect -1037 -1165 -979 -1159
rect -845 -1165 -787 -1159
rect -653 -1165 -595 -1159
rect -461 -1165 -403 -1159
rect -269 -1165 -211 -1159
rect -77 -1165 -19 -1159
rect 115 -1165 173 -1159
rect 307 -1165 365 -1159
rect 499 -1165 557 -1159
rect 691 -1165 749 -1159
rect 883 -1165 941 -1159
rect 1075 -1165 1133 -1159
rect -1037 -1199 -1025 -1165
rect -845 -1199 -833 -1165
rect -653 -1199 -641 -1165
rect -461 -1199 -449 -1165
rect -269 -1199 -257 -1165
rect -77 -1199 -65 -1165
rect 115 -1199 127 -1165
rect 307 -1199 319 -1165
rect 499 -1199 511 -1165
rect 691 -1199 703 -1165
rect 883 -1199 895 -1165
rect 1075 -1199 1087 -1165
rect -1037 -1205 -979 -1199
rect -845 -1205 -787 -1199
rect -653 -1205 -595 -1199
rect -461 -1205 -403 -1199
rect -269 -1205 -211 -1199
rect -77 -1205 -19 -1199
rect 115 -1205 173 -1199
rect 307 -1205 365 -1199
rect 499 -1205 557 -1199
rect 691 -1205 749 -1199
rect 883 -1205 941 -1199
rect 1075 -1205 1133 -1199
rect -1037 -1273 -979 -1267
rect -845 -1273 -787 -1267
rect -653 -1273 -595 -1267
rect -461 -1273 -403 -1267
rect -269 -1273 -211 -1267
rect -77 -1273 -19 -1267
rect 115 -1273 173 -1267
rect 307 -1273 365 -1267
rect 499 -1273 557 -1267
rect 691 -1273 749 -1267
rect 883 -1273 941 -1267
rect 1075 -1273 1133 -1267
rect -1037 -1307 -1025 -1273
rect -845 -1307 -833 -1273
rect -653 -1307 -641 -1273
rect -461 -1307 -449 -1273
rect -269 -1307 -257 -1273
rect -77 -1307 -65 -1273
rect 115 -1307 127 -1273
rect 307 -1307 319 -1273
rect 499 -1307 511 -1273
rect 691 -1307 703 -1273
rect 883 -1307 895 -1273
rect 1075 -1307 1087 -1273
rect -1037 -1313 -979 -1307
rect -845 -1313 -787 -1307
rect -653 -1313 -595 -1307
rect -461 -1313 -403 -1307
rect -269 -1313 -211 -1307
rect -77 -1313 -19 -1307
rect 115 -1313 173 -1307
rect 307 -1313 365 -1307
rect 499 -1313 557 -1307
rect 691 -1313 749 -1307
rect 883 -1313 941 -1307
rect 1075 -1313 1133 -1307
rect -1133 -1783 -1075 -1777
rect -941 -1783 -883 -1777
rect -749 -1783 -691 -1777
rect -557 -1783 -499 -1777
rect -365 -1783 -307 -1777
rect -173 -1783 -115 -1777
rect 19 -1783 77 -1777
rect 211 -1783 269 -1777
rect 403 -1783 461 -1777
rect 595 -1783 653 -1777
rect 787 -1783 845 -1777
rect 979 -1783 1037 -1777
rect -1133 -1817 -1121 -1783
rect -941 -1817 -929 -1783
rect -749 -1817 -737 -1783
rect -557 -1817 -545 -1783
rect -365 -1817 -353 -1783
rect -173 -1817 -161 -1783
rect 19 -1817 31 -1783
rect 211 -1817 223 -1783
rect 403 -1817 415 -1783
rect 595 -1817 607 -1783
rect 787 -1817 799 -1783
rect 979 -1817 991 -1783
rect -1133 -1823 -1075 -1817
rect -941 -1823 -883 -1817
rect -749 -1823 -691 -1817
rect -557 -1823 -499 -1817
rect -365 -1823 -307 -1817
rect -173 -1823 -115 -1817
rect 19 -1823 77 -1817
rect 211 -1823 269 -1817
rect 403 -1823 461 -1817
rect 595 -1823 653 -1817
rect 787 -1823 845 -1817
rect 979 -1823 1037 -1817
rect -1133 -1891 -1075 -1885
rect -941 -1891 -883 -1885
rect -749 -1891 -691 -1885
rect -557 -1891 -499 -1885
rect -365 -1891 -307 -1885
rect -173 -1891 -115 -1885
rect 19 -1891 77 -1885
rect 211 -1891 269 -1885
rect 403 -1891 461 -1885
rect 595 -1891 653 -1885
rect 787 -1891 845 -1885
rect 979 -1891 1037 -1885
rect -1133 -1925 -1121 -1891
rect -941 -1925 -929 -1891
rect -749 -1925 -737 -1891
rect -557 -1925 -545 -1891
rect -365 -1925 -353 -1891
rect -173 -1925 -161 -1891
rect 19 -1925 31 -1891
rect 211 -1925 223 -1891
rect 403 -1925 415 -1891
rect 595 -1925 607 -1891
rect 787 -1925 799 -1891
rect 979 -1925 991 -1891
rect -1133 -1931 -1075 -1925
rect -941 -1931 -883 -1925
rect -749 -1931 -691 -1925
rect -557 -1931 -499 -1925
rect -365 -1931 -307 -1925
rect -173 -1931 -115 -1925
rect 19 -1931 77 -1925
rect 211 -1931 269 -1925
rect 403 -1931 461 -1925
rect 595 -1931 653 -1925
rect 787 -1931 845 -1925
rect 979 -1931 1037 -1925
rect -1037 -2401 -979 -2395
rect -845 -2401 -787 -2395
rect -653 -2401 -595 -2395
rect -461 -2401 -403 -2395
rect -269 -2401 -211 -2395
rect -77 -2401 -19 -2395
rect 115 -2401 173 -2395
rect 307 -2401 365 -2395
rect 499 -2401 557 -2395
rect 691 -2401 749 -2395
rect 883 -2401 941 -2395
rect 1075 -2401 1133 -2395
rect -1037 -2435 -1025 -2401
rect -845 -2435 -833 -2401
rect -653 -2435 -641 -2401
rect -461 -2435 -449 -2401
rect -269 -2435 -257 -2401
rect -77 -2435 -65 -2401
rect 115 -2435 127 -2401
rect 307 -2435 319 -2401
rect 499 -2435 511 -2401
rect 691 -2435 703 -2401
rect 883 -2435 895 -2401
rect 1075 -2435 1087 -2401
rect -1037 -2441 -979 -2435
rect -845 -2441 -787 -2435
rect -653 -2441 -595 -2435
rect -461 -2441 -403 -2435
rect -269 -2441 -211 -2435
rect -77 -2441 -19 -2435
rect 115 -2441 173 -2435
rect 307 -2441 365 -2435
rect 499 -2441 557 -2435
rect 691 -2441 749 -2435
rect 883 -2441 941 -2435
rect 1075 -2441 1133 -2435
rect -1037 -2509 -979 -2503
rect -845 -2509 -787 -2503
rect -653 -2509 -595 -2503
rect -461 -2509 -403 -2503
rect -269 -2509 -211 -2503
rect -77 -2509 -19 -2503
rect 115 -2509 173 -2503
rect 307 -2509 365 -2503
rect 499 -2509 557 -2503
rect 691 -2509 749 -2503
rect 883 -2509 941 -2503
rect 1075 -2509 1133 -2503
rect -1037 -2543 -1025 -2509
rect -845 -2543 -833 -2509
rect -653 -2543 -641 -2509
rect -461 -2543 -449 -2509
rect -269 -2543 -257 -2509
rect -77 -2543 -65 -2509
rect 115 -2543 127 -2509
rect 307 -2543 319 -2509
rect 499 -2543 511 -2509
rect 691 -2543 703 -2509
rect 883 -2543 895 -2509
rect 1075 -2543 1087 -2509
rect -1037 -2549 -979 -2543
rect -845 -2549 -787 -2543
rect -653 -2549 -595 -2543
rect -461 -2549 -403 -2543
rect -269 -2549 -211 -2543
rect -77 -2549 -19 -2543
rect 115 -2549 173 -2543
rect 307 -2549 365 -2543
rect 499 -2549 557 -2543
rect 691 -2549 749 -2543
rect 883 -2549 941 -2543
rect 1075 -2549 1133 -2543
rect -1133 -3019 -1075 -3013
rect -941 -3019 -883 -3013
rect -749 -3019 -691 -3013
rect -557 -3019 -499 -3013
rect -365 -3019 -307 -3013
rect -173 -3019 -115 -3013
rect 19 -3019 77 -3013
rect 211 -3019 269 -3013
rect 403 -3019 461 -3013
rect 595 -3019 653 -3013
rect 787 -3019 845 -3013
rect 979 -3019 1037 -3013
rect -1133 -3053 -1121 -3019
rect -941 -3053 -929 -3019
rect -749 -3053 -737 -3019
rect -557 -3053 -545 -3019
rect -365 -3053 -353 -3019
rect -173 -3053 -161 -3019
rect 19 -3053 31 -3019
rect 211 -3053 223 -3019
rect 403 -3053 415 -3019
rect 595 -3053 607 -3019
rect 787 -3053 799 -3019
rect 979 -3053 991 -3019
rect -1133 -3059 -1075 -3053
rect -941 -3059 -883 -3053
rect -749 -3059 -691 -3053
rect -557 -3059 -499 -3053
rect -365 -3059 -307 -3053
rect -173 -3059 -115 -3053
rect 19 -3059 77 -3053
rect 211 -3059 269 -3053
rect 403 -3059 461 -3053
rect 595 -3059 653 -3053
rect 787 -3059 845 -3053
rect 979 -3059 1037 -3053
<< pwell >>
rect -1319 -3191 1319 3191
<< nmoslvt >>
rect -1119 2581 -1089 2981
rect -1023 2581 -993 2981
rect -927 2581 -897 2981
rect -831 2581 -801 2981
rect -735 2581 -705 2981
rect -639 2581 -609 2981
rect -543 2581 -513 2981
rect -447 2581 -417 2981
rect -351 2581 -321 2981
rect -255 2581 -225 2981
rect -159 2581 -129 2981
rect -63 2581 -33 2981
rect 33 2581 63 2981
rect 129 2581 159 2981
rect 225 2581 255 2981
rect 321 2581 351 2981
rect 417 2581 447 2981
rect 513 2581 543 2981
rect 609 2581 639 2981
rect 705 2581 735 2981
rect 801 2581 831 2981
rect 897 2581 927 2981
rect 993 2581 1023 2981
rect 1089 2581 1119 2981
rect -1119 1963 -1089 2363
rect -1023 1963 -993 2363
rect -927 1963 -897 2363
rect -831 1963 -801 2363
rect -735 1963 -705 2363
rect -639 1963 -609 2363
rect -543 1963 -513 2363
rect -447 1963 -417 2363
rect -351 1963 -321 2363
rect -255 1963 -225 2363
rect -159 1963 -129 2363
rect -63 1963 -33 2363
rect 33 1963 63 2363
rect 129 1963 159 2363
rect 225 1963 255 2363
rect 321 1963 351 2363
rect 417 1963 447 2363
rect 513 1963 543 2363
rect 609 1963 639 2363
rect 705 1963 735 2363
rect 801 1963 831 2363
rect 897 1963 927 2363
rect 993 1963 1023 2363
rect 1089 1963 1119 2363
rect -1119 1345 -1089 1745
rect -1023 1345 -993 1745
rect -927 1345 -897 1745
rect -831 1345 -801 1745
rect -735 1345 -705 1745
rect -639 1345 -609 1745
rect -543 1345 -513 1745
rect -447 1345 -417 1745
rect -351 1345 -321 1745
rect -255 1345 -225 1745
rect -159 1345 -129 1745
rect -63 1345 -33 1745
rect 33 1345 63 1745
rect 129 1345 159 1745
rect 225 1345 255 1745
rect 321 1345 351 1745
rect 417 1345 447 1745
rect 513 1345 543 1745
rect 609 1345 639 1745
rect 705 1345 735 1745
rect 801 1345 831 1745
rect 897 1345 927 1745
rect 993 1345 1023 1745
rect 1089 1345 1119 1745
rect -1119 727 -1089 1127
rect -1023 727 -993 1127
rect -927 727 -897 1127
rect -831 727 -801 1127
rect -735 727 -705 1127
rect -639 727 -609 1127
rect -543 727 -513 1127
rect -447 727 -417 1127
rect -351 727 -321 1127
rect -255 727 -225 1127
rect -159 727 -129 1127
rect -63 727 -33 1127
rect 33 727 63 1127
rect 129 727 159 1127
rect 225 727 255 1127
rect 321 727 351 1127
rect 417 727 447 1127
rect 513 727 543 1127
rect 609 727 639 1127
rect 705 727 735 1127
rect 801 727 831 1127
rect 897 727 927 1127
rect 993 727 1023 1127
rect 1089 727 1119 1127
rect -1119 109 -1089 509
rect -1023 109 -993 509
rect -927 109 -897 509
rect -831 109 -801 509
rect -735 109 -705 509
rect -639 109 -609 509
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect 609 109 639 509
rect 705 109 735 509
rect 801 109 831 509
rect 897 109 927 509
rect 993 109 1023 509
rect 1089 109 1119 509
rect -1119 -509 -1089 -109
rect -1023 -509 -993 -109
rect -927 -509 -897 -109
rect -831 -509 -801 -109
rect -735 -509 -705 -109
rect -639 -509 -609 -109
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect 609 -509 639 -109
rect 705 -509 735 -109
rect 801 -509 831 -109
rect 897 -509 927 -109
rect 993 -509 1023 -109
rect 1089 -509 1119 -109
rect -1119 -1127 -1089 -727
rect -1023 -1127 -993 -727
rect -927 -1127 -897 -727
rect -831 -1127 -801 -727
rect -735 -1127 -705 -727
rect -639 -1127 -609 -727
rect -543 -1127 -513 -727
rect -447 -1127 -417 -727
rect -351 -1127 -321 -727
rect -255 -1127 -225 -727
rect -159 -1127 -129 -727
rect -63 -1127 -33 -727
rect 33 -1127 63 -727
rect 129 -1127 159 -727
rect 225 -1127 255 -727
rect 321 -1127 351 -727
rect 417 -1127 447 -727
rect 513 -1127 543 -727
rect 609 -1127 639 -727
rect 705 -1127 735 -727
rect 801 -1127 831 -727
rect 897 -1127 927 -727
rect 993 -1127 1023 -727
rect 1089 -1127 1119 -727
rect -1119 -1745 -1089 -1345
rect -1023 -1745 -993 -1345
rect -927 -1745 -897 -1345
rect -831 -1745 -801 -1345
rect -735 -1745 -705 -1345
rect -639 -1745 -609 -1345
rect -543 -1745 -513 -1345
rect -447 -1745 -417 -1345
rect -351 -1745 -321 -1345
rect -255 -1745 -225 -1345
rect -159 -1745 -129 -1345
rect -63 -1745 -33 -1345
rect 33 -1745 63 -1345
rect 129 -1745 159 -1345
rect 225 -1745 255 -1345
rect 321 -1745 351 -1345
rect 417 -1745 447 -1345
rect 513 -1745 543 -1345
rect 609 -1745 639 -1345
rect 705 -1745 735 -1345
rect 801 -1745 831 -1345
rect 897 -1745 927 -1345
rect 993 -1745 1023 -1345
rect 1089 -1745 1119 -1345
rect -1119 -2363 -1089 -1963
rect -1023 -2363 -993 -1963
rect -927 -2363 -897 -1963
rect -831 -2363 -801 -1963
rect -735 -2363 -705 -1963
rect -639 -2363 -609 -1963
rect -543 -2363 -513 -1963
rect -447 -2363 -417 -1963
rect -351 -2363 -321 -1963
rect -255 -2363 -225 -1963
rect -159 -2363 -129 -1963
rect -63 -2363 -33 -1963
rect 33 -2363 63 -1963
rect 129 -2363 159 -1963
rect 225 -2363 255 -1963
rect 321 -2363 351 -1963
rect 417 -2363 447 -1963
rect 513 -2363 543 -1963
rect 609 -2363 639 -1963
rect 705 -2363 735 -1963
rect 801 -2363 831 -1963
rect 897 -2363 927 -1963
rect 993 -2363 1023 -1963
rect 1089 -2363 1119 -1963
rect -1119 -2981 -1089 -2581
rect -1023 -2981 -993 -2581
rect -927 -2981 -897 -2581
rect -831 -2981 -801 -2581
rect -735 -2981 -705 -2581
rect -639 -2981 -609 -2581
rect -543 -2981 -513 -2581
rect -447 -2981 -417 -2581
rect -351 -2981 -321 -2581
rect -255 -2981 -225 -2581
rect -159 -2981 -129 -2581
rect -63 -2981 -33 -2581
rect 33 -2981 63 -2581
rect 129 -2981 159 -2581
rect 225 -2981 255 -2581
rect 321 -2981 351 -2581
rect 417 -2981 447 -2581
rect 513 -2981 543 -2581
rect 609 -2981 639 -2581
rect 705 -2981 735 -2581
rect 801 -2981 831 -2581
rect 897 -2981 927 -2581
rect 993 -2981 1023 -2581
rect 1089 -2981 1119 -2581
<< ndiff >>
rect -1181 2969 -1119 2981
rect -1181 2593 -1169 2969
rect -1135 2593 -1119 2969
rect -1181 2581 -1119 2593
rect -1089 2969 -1023 2981
rect -1089 2593 -1073 2969
rect -1039 2593 -1023 2969
rect -1089 2581 -1023 2593
rect -993 2969 -927 2981
rect -993 2593 -977 2969
rect -943 2593 -927 2969
rect -993 2581 -927 2593
rect -897 2969 -831 2981
rect -897 2593 -881 2969
rect -847 2593 -831 2969
rect -897 2581 -831 2593
rect -801 2969 -735 2981
rect -801 2593 -785 2969
rect -751 2593 -735 2969
rect -801 2581 -735 2593
rect -705 2969 -639 2981
rect -705 2593 -689 2969
rect -655 2593 -639 2969
rect -705 2581 -639 2593
rect -609 2969 -543 2981
rect -609 2593 -593 2969
rect -559 2593 -543 2969
rect -609 2581 -543 2593
rect -513 2969 -447 2981
rect -513 2593 -497 2969
rect -463 2593 -447 2969
rect -513 2581 -447 2593
rect -417 2969 -351 2981
rect -417 2593 -401 2969
rect -367 2593 -351 2969
rect -417 2581 -351 2593
rect -321 2969 -255 2981
rect -321 2593 -305 2969
rect -271 2593 -255 2969
rect -321 2581 -255 2593
rect -225 2969 -159 2981
rect -225 2593 -209 2969
rect -175 2593 -159 2969
rect -225 2581 -159 2593
rect -129 2969 -63 2981
rect -129 2593 -113 2969
rect -79 2593 -63 2969
rect -129 2581 -63 2593
rect -33 2969 33 2981
rect -33 2593 -17 2969
rect 17 2593 33 2969
rect -33 2581 33 2593
rect 63 2969 129 2981
rect 63 2593 79 2969
rect 113 2593 129 2969
rect 63 2581 129 2593
rect 159 2969 225 2981
rect 159 2593 175 2969
rect 209 2593 225 2969
rect 159 2581 225 2593
rect 255 2969 321 2981
rect 255 2593 271 2969
rect 305 2593 321 2969
rect 255 2581 321 2593
rect 351 2969 417 2981
rect 351 2593 367 2969
rect 401 2593 417 2969
rect 351 2581 417 2593
rect 447 2969 513 2981
rect 447 2593 463 2969
rect 497 2593 513 2969
rect 447 2581 513 2593
rect 543 2969 609 2981
rect 543 2593 559 2969
rect 593 2593 609 2969
rect 543 2581 609 2593
rect 639 2969 705 2981
rect 639 2593 655 2969
rect 689 2593 705 2969
rect 639 2581 705 2593
rect 735 2969 801 2981
rect 735 2593 751 2969
rect 785 2593 801 2969
rect 735 2581 801 2593
rect 831 2969 897 2981
rect 831 2593 847 2969
rect 881 2593 897 2969
rect 831 2581 897 2593
rect 927 2969 993 2981
rect 927 2593 943 2969
rect 977 2593 993 2969
rect 927 2581 993 2593
rect 1023 2969 1089 2981
rect 1023 2593 1039 2969
rect 1073 2593 1089 2969
rect 1023 2581 1089 2593
rect 1119 2969 1181 2981
rect 1119 2593 1135 2969
rect 1169 2593 1181 2969
rect 1119 2581 1181 2593
rect -1181 2351 -1119 2363
rect -1181 1975 -1169 2351
rect -1135 1975 -1119 2351
rect -1181 1963 -1119 1975
rect -1089 2351 -1023 2363
rect -1089 1975 -1073 2351
rect -1039 1975 -1023 2351
rect -1089 1963 -1023 1975
rect -993 2351 -927 2363
rect -993 1975 -977 2351
rect -943 1975 -927 2351
rect -993 1963 -927 1975
rect -897 2351 -831 2363
rect -897 1975 -881 2351
rect -847 1975 -831 2351
rect -897 1963 -831 1975
rect -801 2351 -735 2363
rect -801 1975 -785 2351
rect -751 1975 -735 2351
rect -801 1963 -735 1975
rect -705 2351 -639 2363
rect -705 1975 -689 2351
rect -655 1975 -639 2351
rect -705 1963 -639 1975
rect -609 2351 -543 2363
rect -609 1975 -593 2351
rect -559 1975 -543 2351
rect -609 1963 -543 1975
rect -513 2351 -447 2363
rect -513 1975 -497 2351
rect -463 1975 -447 2351
rect -513 1963 -447 1975
rect -417 2351 -351 2363
rect -417 1975 -401 2351
rect -367 1975 -351 2351
rect -417 1963 -351 1975
rect -321 2351 -255 2363
rect -321 1975 -305 2351
rect -271 1975 -255 2351
rect -321 1963 -255 1975
rect -225 2351 -159 2363
rect -225 1975 -209 2351
rect -175 1975 -159 2351
rect -225 1963 -159 1975
rect -129 2351 -63 2363
rect -129 1975 -113 2351
rect -79 1975 -63 2351
rect -129 1963 -63 1975
rect -33 2351 33 2363
rect -33 1975 -17 2351
rect 17 1975 33 2351
rect -33 1963 33 1975
rect 63 2351 129 2363
rect 63 1975 79 2351
rect 113 1975 129 2351
rect 63 1963 129 1975
rect 159 2351 225 2363
rect 159 1975 175 2351
rect 209 1975 225 2351
rect 159 1963 225 1975
rect 255 2351 321 2363
rect 255 1975 271 2351
rect 305 1975 321 2351
rect 255 1963 321 1975
rect 351 2351 417 2363
rect 351 1975 367 2351
rect 401 1975 417 2351
rect 351 1963 417 1975
rect 447 2351 513 2363
rect 447 1975 463 2351
rect 497 1975 513 2351
rect 447 1963 513 1975
rect 543 2351 609 2363
rect 543 1975 559 2351
rect 593 1975 609 2351
rect 543 1963 609 1975
rect 639 2351 705 2363
rect 639 1975 655 2351
rect 689 1975 705 2351
rect 639 1963 705 1975
rect 735 2351 801 2363
rect 735 1975 751 2351
rect 785 1975 801 2351
rect 735 1963 801 1975
rect 831 2351 897 2363
rect 831 1975 847 2351
rect 881 1975 897 2351
rect 831 1963 897 1975
rect 927 2351 993 2363
rect 927 1975 943 2351
rect 977 1975 993 2351
rect 927 1963 993 1975
rect 1023 2351 1089 2363
rect 1023 1975 1039 2351
rect 1073 1975 1089 2351
rect 1023 1963 1089 1975
rect 1119 2351 1181 2363
rect 1119 1975 1135 2351
rect 1169 1975 1181 2351
rect 1119 1963 1181 1975
rect -1181 1733 -1119 1745
rect -1181 1357 -1169 1733
rect -1135 1357 -1119 1733
rect -1181 1345 -1119 1357
rect -1089 1733 -1023 1745
rect -1089 1357 -1073 1733
rect -1039 1357 -1023 1733
rect -1089 1345 -1023 1357
rect -993 1733 -927 1745
rect -993 1357 -977 1733
rect -943 1357 -927 1733
rect -993 1345 -927 1357
rect -897 1733 -831 1745
rect -897 1357 -881 1733
rect -847 1357 -831 1733
rect -897 1345 -831 1357
rect -801 1733 -735 1745
rect -801 1357 -785 1733
rect -751 1357 -735 1733
rect -801 1345 -735 1357
rect -705 1733 -639 1745
rect -705 1357 -689 1733
rect -655 1357 -639 1733
rect -705 1345 -639 1357
rect -609 1733 -543 1745
rect -609 1357 -593 1733
rect -559 1357 -543 1733
rect -609 1345 -543 1357
rect -513 1733 -447 1745
rect -513 1357 -497 1733
rect -463 1357 -447 1733
rect -513 1345 -447 1357
rect -417 1733 -351 1745
rect -417 1357 -401 1733
rect -367 1357 -351 1733
rect -417 1345 -351 1357
rect -321 1733 -255 1745
rect -321 1357 -305 1733
rect -271 1357 -255 1733
rect -321 1345 -255 1357
rect -225 1733 -159 1745
rect -225 1357 -209 1733
rect -175 1357 -159 1733
rect -225 1345 -159 1357
rect -129 1733 -63 1745
rect -129 1357 -113 1733
rect -79 1357 -63 1733
rect -129 1345 -63 1357
rect -33 1733 33 1745
rect -33 1357 -17 1733
rect 17 1357 33 1733
rect -33 1345 33 1357
rect 63 1733 129 1745
rect 63 1357 79 1733
rect 113 1357 129 1733
rect 63 1345 129 1357
rect 159 1733 225 1745
rect 159 1357 175 1733
rect 209 1357 225 1733
rect 159 1345 225 1357
rect 255 1733 321 1745
rect 255 1357 271 1733
rect 305 1357 321 1733
rect 255 1345 321 1357
rect 351 1733 417 1745
rect 351 1357 367 1733
rect 401 1357 417 1733
rect 351 1345 417 1357
rect 447 1733 513 1745
rect 447 1357 463 1733
rect 497 1357 513 1733
rect 447 1345 513 1357
rect 543 1733 609 1745
rect 543 1357 559 1733
rect 593 1357 609 1733
rect 543 1345 609 1357
rect 639 1733 705 1745
rect 639 1357 655 1733
rect 689 1357 705 1733
rect 639 1345 705 1357
rect 735 1733 801 1745
rect 735 1357 751 1733
rect 785 1357 801 1733
rect 735 1345 801 1357
rect 831 1733 897 1745
rect 831 1357 847 1733
rect 881 1357 897 1733
rect 831 1345 897 1357
rect 927 1733 993 1745
rect 927 1357 943 1733
rect 977 1357 993 1733
rect 927 1345 993 1357
rect 1023 1733 1089 1745
rect 1023 1357 1039 1733
rect 1073 1357 1089 1733
rect 1023 1345 1089 1357
rect 1119 1733 1181 1745
rect 1119 1357 1135 1733
rect 1169 1357 1181 1733
rect 1119 1345 1181 1357
rect -1181 1115 -1119 1127
rect -1181 739 -1169 1115
rect -1135 739 -1119 1115
rect -1181 727 -1119 739
rect -1089 1115 -1023 1127
rect -1089 739 -1073 1115
rect -1039 739 -1023 1115
rect -1089 727 -1023 739
rect -993 1115 -927 1127
rect -993 739 -977 1115
rect -943 739 -927 1115
rect -993 727 -927 739
rect -897 1115 -831 1127
rect -897 739 -881 1115
rect -847 739 -831 1115
rect -897 727 -831 739
rect -801 1115 -735 1127
rect -801 739 -785 1115
rect -751 739 -735 1115
rect -801 727 -735 739
rect -705 1115 -639 1127
rect -705 739 -689 1115
rect -655 739 -639 1115
rect -705 727 -639 739
rect -609 1115 -543 1127
rect -609 739 -593 1115
rect -559 739 -543 1115
rect -609 727 -543 739
rect -513 1115 -447 1127
rect -513 739 -497 1115
rect -463 739 -447 1115
rect -513 727 -447 739
rect -417 1115 -351 1127
rect -417 739 -401 1115
rect -367 739 -351 1115
rect -417 727 -351 739
rect -321 1115 -255 1127
rect -321 739 -305 1115
rect -271 739 -255 1115
rect -321 727 -255 739
rect -225 1115 -159 1127
rect -225 739 -209 1115
rect -175 739 -159 1115
rect -225 727 -159 739
rect -129 1115 -63 1127
rect -129 739 -113 1115
rect -79 739 -63 1115
rect -129 727 -63 739
rect -33 1115 33 1127
rect -33 739 -17 1115
rect 17 739 33 1115
rect -33 727 33 739
rect 63 1115 129 1127
rect 63 739 79 1115
rect 113 739 129 1115
rect 63 727 129 739
rect 159 1115 225 1127
rect 159 739 175 1115
rect 209 739 225 1115
rect 159 727 225 739
rect 255 1115 321 1127
rect 255 739 271 1115
rect 305 739 321 1115
rect 255 727 321 739
rect 351 1115 417 1127
rect 351 739 367 1115
rect 401 739 417 1115
rect 351 727 417 739
rect 447 1115 513 1127
rect 447 739 463 1115
rect 497 739 513 1115
rect 447 727 513 739
rect 543 1115 609 1127
rect 543 739 559 1115
rect 593 739 609 1115
rect 543 727 609 739
rect 639 1115 705 1127
rect 639 739 655 1115
rect 689 739 705 1115
rect 639 727 705 739
rect 735 1115 801 1127
rect 735 739 751 1115
rect 785 739 801 1115
rect 735 727 801 739
rect 831 1115 897 1127
rect 831 739 847 1115
rect 881 739 897 1115
rect 831 727 897 739
rect 927 1115 993 1127
rect 927 739 943 1115
rect 977 739 993 1115
rect 927 727 993 739
rect 1023 1115 1089 1127
rect 1023 739 1039 1115
rect 1073 739 1089 1115
rect 1023 727 1089 739
rect 1119 1115 1181 1127
rect 1119 739 1135 1115
rect 1169 739 1181 1115
rect 1119 727 1181 739
rect -1181 497 -1119 509
rect -1181 121 -1169 497
rect -1135 121 -1119 497
rect -1181 109 -1119 121
rect -1089 497 -1023 509
rect -1089 121 -1073 497
rect -1039 121 -1023 497
rect -1089 109 -1023 121
rect -993 497 -927 509
rect -993 121 -977 497
rect -943 121 -927 497
rect -993 109 -927 121
rect -897 497 -831 509
rect -897 121 -881 497
rect -847 121 -831 497
rect -897 109 -831 121
rect -801 497 -735 509
rect -801 121 -785 497
rect -751 121 -735 497
rect -801 109 -735 121
rect -705 497 -639 509
rect -705 121 -689 497
rect -655 121 -639 497
rect -705 109 -639 121
rect -609 497 -543 509
rect -609 121 -593 497
rect -559 121 -543 497
rect -609 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 609 509
rect 543 121 559 497
rect 593 121 609 497
rect 543 109 609 121
rect 639 497 705 509
rect 639 121 655 497
rect 689 121 705 497
rect 639 109 705 121
rect 735 497 801 509
rect 735 121 751 497
rect 785 121 801 497
rect 735 109 801 121
rect 831 497 897 509
rect 831 121 847 497
rect 881 121 897 497
rect 831 109 897 121
rect 927 497 993 509
rect 927 121 943 497
rect 977 121 993 497
rect 927 109 993 121
rect 1023 497 1089 509
rect 1023 121 1039 497
rect 1073 121 1089 497
rect 1023 109 1089 121
rect 1119 497 1181 509
rect 1119 121 1135 497
rect 1169 121 1181 497
rect 1119 109 1181 121
rect -1181 -121 -1119 -109
rect -1181 -497 -1169 -121
rect -1135 -497 -1119 -121
rect -1181 -509 -1119 -497
rect -1089 -121 -1023 -109
rect -1089 -497 -1073 -121
rect -1039 -497 -1023 -121
rect -1089 -509 -1023 -497
rect -993 -121 -927 -109
rect -993 -497 -977 -121
rect -943 -497 -927 -121
rect -993 -509 -927 -497
rect -897 -121 -831 -109
rect -897 -497 -881 -121
rect -847 -497 -831 -121
rect -897 -509 -831 -497
rect -801 -121 -735 -109
rect -801 -497 -785 -121
rect -751 -497 -735 -121
rect -801 -509 -735 -497
rect -705 -121 -639 -109
rect -705 -497 -689 -121
rect -655 -497 -639 -121
rect -705 -509 -639 -497
rect -609 -121 -543 -109
rect -609 -497 -593 -121
rect -559 -497 -543 -121
rect -609 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 609 -109
rect 543 -497 559 -121
rect 593 -497 609 -121
rect 543 -509 609 -497
rect 639 -121 705 -109
rect 639 -497 655 -121
rect 689 -497 705 -121
rect 639 -509 705 -497
rect 735 -121 801 -109
rect 735 -497 751 -121
rect 785 -497 801 -121
rect 735 -509 801 -497
rect 831 -121 897 -109
rect 831 -497 847 -121
rect 881 -497 897 -121
rect 831 -509 897 -497
rect 927 -121 993 -109
rect 927 -497 943 -121
rect 977 -497 993 -121
rect 927 -509 993 -497
rect 1023 -121 1089 -109
rect 1023 -497 1039 -121
rect 1073 -497 1089 -121
rect 1023 -509 1089 -497
rect 1119 -121 1181 -109
rect 1119 -497 1135 -121
rect 1169 -497 1181 -121
rect 1119 -509 1181 -497
rect -1181 -739 -1119 -727
rect -1181 -1115 -1169 -739
rect -1135 -1115 -1119 -739
rect -1181 -1127 -1119 -1115
rect -1089 -739 -1023 -727
rect -1089 -1115 -1073 -739
rect -1039 -1115 -1023 -739
rect -1089 -1127 -1023 -1115
rect -993 -739 -927 -727
rect -993 -1115 -977 -739
rect -943 -1115 -927 -739
rect -993 -1127 -927 -1115
rect -897 -739 -831 -727
rect -897 -1115 -881 -739
rect -847 -1115 -831 -739
rect -897 -1127 -831 -1115
rect -801 -739 -735 -727
rect -801 -1115 -785 -739
rect -751 -1115 -735 -739
rect -801 -1127 -735 -1115
rect -705 -739 -639 -727
rect -705 -1115 -689 -739
rect -655 -1115 -639 -739
rect -705 -1127 -639 -1115
rect -609 -739 -543 -727
rect -609 -1115 -593 -739
rect -559 -1115 -543 -739
rect -609 -1127 -543 -1115
rect -513 -739 -447 -727
rect -513 -1115 -497 -739
rect -463 -1115 -447 -739
rect -513 -1127 -447 -1115
rect -417 -739 -351 -727
rect -417 -1115 -401 -739
rect -367 -1115 -351 -739
rect -417 -1127 -351 -1115
rect -321 -739 -255 -727
rect -321 -1115 -305 -739
rect -271 -1115 -255 -739
rect -321 -1127 -255 -1115
rect -225 -739 -159 -727
rect -225 -1115 -209 -739
rect -175 -1115 -159 -739
rect -225 -1127 -159 -1115
rect -129 -739 -63 -727
rect -129 -1115 -113 -739
rect -79 -1115 -63 -739
rect -129 -1127 -63 -1115
rect -33 -739 33 -727
rect -33 -1115 -17 -739
rect 17 -1115 33 -739
rect -33 -1127 33 -1115
rect 63 -739 129 -727
rect 63 -1115 79 -739
rect 113 -1115 129 -739
rect 63 -1127 129 -1115
rect 159 -739 225 -727
rect 159 -1115 175 -739
rect 209 -1115 225 -739
rect 159 -1127 225 -1115
rect 255 -739 321 -727
rect 255 -1115 271 -739
rect 305 -1115 321 -739
rect 255 -1127 321 -1115
rect 351 -739 417 -727
rect 351 -1115 367 -739
rect 401 -1115 417 -739
rect 351 -1127 417 -1115
rect 447 -739 513 -727
rect 447 -1115 463 -739
rect 497 -1115 513 -739
rect 447 -1127 513 -1115
rect 543 -739 609 -727
rect 543 -1115 559 -739
rect 593 -1115 609 -739
rect 543 -1127 609 -1115
rect 639 -739 705 -727
rect 639 -1115 655 -739
rect 689 -1115 705 -739
rect 639 -1127 705 -1115
rect 735 -739 801 -727
rect 735 -1115 751 -739
rect 785 -1115 801 -739
rect 735 -1127 801 -1115
rect 831 -739 897 -727
rect 831 -1115 847 -739
rect 881 -1115 897 -739
rect 831 -1127 897 -1115
rect 927 -739 993 -727
rect 927 -1115 943 -739
rect 977 -1115 993 -739
rect 927 -1127 993 -1115
rect 1023 -739 1089 -727
rect 1023 -1115 1039 -739
rect 1073 -1115 1089 -739
rect 1023 -1127 1089 -1115
rect 1119 -739 1181 -727
rect 1119 -1115 1135 -739
rect 1169 -1115 1181 -739
rect 1119 -1127 1181 -1115
rect -1181 -1357 -1119 -1345
rect -1181 -1733 -1169 -1357
rect -1135 -1733 -1119 -1357
rect -1181 -1745 -1119 -1733
rect -1089 -1357 -1023 -1345
rect -1089 -1733 -1073 -1357
rect -1039 -1733 -1023 -1357
rect -1089 -1745 -1023 -1733
rect -993 -1357 -927 -1345
rect -993 -1733 -977 -1357
rect -943 -1733 -927 -1357
rect -993 -1745 -927 -1733
rect -897 -1357 -831 -1345
rect -897 -1733 -881 -1357
rect -847 -1733 -831 -1357
rect -897 -1745 -831 -1733
rect -801 -1357 -735 -1345
rect -801 -1733 -785 -1357
rect -751 -1733 -735 -1357
rect -801 -1745 -735 -1733
rect -705 -1357 -639 -1345
rect -705 -1733 -689 -1357
rect -655 -1733 -639 -1357
rect -705 -1745 -639 -1733
rect -609 -1357 -543 -1345
rect -609 -1733 -593 -1357
rect -559 -1733 -543 -1357
rect -609 -1745 -543 -1733
rect -513 -1357 -447 -1345
rect -513 -1733 -497 -1357
rect -463 -1733 -447 -1357
rect -513 -1745 -447 -1733
rect -417 -1357 -351 -1345
rect -417 -1733 -401 -1357
rect -367 -1733 -351 -1357
rect -417 -1745 -351 -1733
rect -321 -1357 -255 -1345
rect -321 -1733 -305 -1357
rect -271 -1733 -255 -1357
rect -321 -1745 -255 -1733
rect -225 -1357 -159 -1345
rect -225 -1733 -209 -1357
rect -175 -1733 -159 -1357
rect -225 -1745 -159 -1733
rect -129 -1357 -63 -1345
rect -129 -1733 -113 -1357
rect -79 -1733 -63 -1357
rect -129 -1745 -63 -1733
rect -33 -1357 33 -1345
rect -33 -1733 -17 -1357
rect 17 -1733 33 -1357
rect -33 -1745 33 -1733
rect 63 -1357 129 -1345
rect 63 -1733 79 -1357
rect 113 -1733 129 -1357
rect 63 -1745 129 -1733
rect 159 -1357 225 -1345
rect 159 -1733 175 -1357
rect 209 -1733 225 -1357
rect 159 -1745 225 -1733
rect 255 -1357 321 -1345
rect 255 -1733 271 -1357
rect 305 -1733 321 -1357
rect 255 -1745 321 -1733
rect 351 -1357 417 -1345
rect 351 -1733 367 -1357
rect 401 -1733 417 -1357
rect 351 -1745 417 -1733
rect 447 -1357 513 -1345
rect 447 -1733 463 -1357
rect 497 -1733 513 -1357
rect 447 -1745 513 -1733
rect 543 -1357 609 -1345
rect 543 -1733 559 -1357
rect 593 -1733 609 -1357
rect 543 -1745 609 -1733
rect 639 -1357 705 -1345
rect 639 -1733 655 -1357
rect 689 -1733 705 -1357
rect 639 -1745 705 -1733
rect 735 -1357 801 -1345
rect 735 -1733 751 -1357
rect 785 -1733 801 -1357
rect 735 -1745 801 -1733
rect 831 -1357 897 -1345
rect 831 -1733 847 -1357
rect 881 -1733 897 -1357
rect 831 -1745 897 -1733
rect 927 -1357 993 -1345
rect 927 -1733 943 -1357
rect 977 -1733 993 -1357
rect 927 -1745 993 -1733
rect 1023 -1357 1089 -1345
rect 1023 -1733 1039 -1357
rect 1073 -1733 1089 -1357
rect 1023 -1745 1089 -1733
rect 1119 -1357 1181 -1345
rect 1119 -1733 1135 -1357
rect 1169 -1733 1181 -1357
rect 1119 -1745 1181 -1733
rect -1181 -1975 -1119 -1963
rect -1181 -2351 -1169 -1975
rect -1135 -2351 -1119 -1975
rect -1181 -2363 -1119 -2351
rect -1089 -1975 -1023 -1963
rect -1089 -2351 -1073 -1975
rect -1039 -2351 -1023 -1975
rect -1089 -2363 -1023 -2351
rect -993 -1975 -927 -1963
rect -993 -2351 -977 -1975
rect -943 -2351 -927 -1975
rect -993 -2363 -927 -2351
rect -897 -1975 -831 -1963
rect -897 -2351 -881 -1975
rect -847 -2351 -831 -1975
rect -897 -2363 -831 -2351
rect -801 -1975 -735 -1963
rect -801 -2351 -785 -1975
rect -751 -2351 -735 -1975
rect -801 -2363 -735 -2351
rect -705 -1975 -639 -1963
rect -705 -2351 -689 -1975
rect -655 -2351 -639 -1975
rect -705 -2363 -639 -2351
rect -609 -1975 -543 -1963
rect -609 -2351 -593 -1975
rect -559 -2351 -543 -1975
rect -609 -2363 -543 -2351
rect -513 -1975 -447 -1963
rect -513 -2351 -497 -1975
rect -463 -2351 -447 -1975
rect -513 -2363 -447 -2351
rect -417 -1975 -351 -1963
rect -417 -2351 -401 -1975
rect -367 -2351 -351 -1975
rect -417 -2363 -351 -2351
rect -321 -1975 -255 -1963
rect -321 -2351 -305 -1975
rect -271 -2351 -255 -1975
rect -321 -2363 -255 -2351
rect -225 -1975 -159 -1963
rect -225 -2351 -209 -1975
rect -175 -2351 -159 -1975
rect -225 -2363 -159 -2351
rect -129 -1975 -63 -1963
rect -129 -2351 -113 -1975
rect -79 -2351 -63 -1975
rect -129 -2363 -63 -2351
rect -33 -1975 33 -1963
rect -33 -2351 -17 -1975
rect 17 -2351 33 -1975
rect -33 -2363 33 -2351
rect 63 -1975 129 -1963
rect 63 -2351 79 -1975
rect 113 -2351 129 -1975
rect 63 -2363 129 -2351
rect 159 -1975 225 -1963
rect 159 -2351 175 -1975
rect 209 -2351 225 -1975
rect 159 -2363 225 -2351
rect 255 -1975 321 -1963
rect 255 -2351 271 -1975
rect 305 -2351 321 -1975
rect 255 -2363 321 -2351
rect 351 -1975 417 -1963
rect 351 -2351 367 -1975
rect 401 -2351 417 -1975
rect 351 -2363 417 -2351
rect 447 -1975 513 -1963
rect 447 -2351 463 -1975
rect 497 -2351 513 -1975
rect 447 -2363 513 -2351
rect 543 -1975 609 -1963
rect 543 -2351 559 -1975
rect 593 -2351 609 -1975
rect 543 -2363 609 -2351
rect 639 -1975 705 -1963
rect 639 -2351 655 -1975
rect 689 -2351 705 -1975
rect 639 -2363 705 -2351
rect 735 -1975 801 -1963
rect 735 -2351 751 -1975
rect 785 -2351 801 -1975
rect 735 -2363 801 -2351
rect 831 -1975 897 -1963
rect 831 -2351 847 -1975
rect 881 -2351 897 -1975
rect 831 -2363 897 -2351
rect 927 -1975 993 -1963
rect 927 -2351 943 -1975
rect 977 -2351 993 -1975
rect 927 -2363 993 -2351
rect 1023 -1975 1089 -1963
rect 1023 -2351 1039 -1975
rect 1073 -2351 1089 -1975
rect 1023 -2363 1089 -2351
rect 1119 -1975 1181 -1963
rect 1119 -2351 1135 -1975
rect 1169 -2351 1181 -1975
rect 1119 -2363 1181 -2351
rect -1181 -2593 -1119 -2581
rect -1181 -2969 -1169 -2593
rect -1135 -2969 -1119 -2593
rect -1181 -2981 -1119 -2969
rect -1089 -2593 -1023 -2581
rect -1089 -2969 -1073 -2593
rect -1039 -2969 -1023 -2593
rect -1089 -2981 -1023 -2969
rect -993 -2593 -927 -2581
rect -993 -2969 -977 -2593
rect -943 -2969 -927 -2593
rect -993 -2981 -927 -2969
rect -897 -2593 -831 -2581
rect -897 -2969 -881 -2593
rect -847 -2969 -831 -2593
rect -897 -2981 -831 -2969
rect -801 -2593 -735 -2581
rect -801 -2969 -785 -2593
rect -751 -2969 -735 -2593
rect -801 -2981 -735 -2969
rect -705 -2593 -639 -2581
rect -705 -2969 -689 -2593
rect -655 -2969 -639 -2593
rect -705 -2981 -639 -2969
rect -609 -2593 -543 -2581
rect -609 -2969 -593 -2593
rect -559 -2969 -543 -2593
rect -609 -2981 -543 -2969
rect -513 -2593 -447 -2581
rect -513 -2969 -497 -2593
rect -463 -2969 -447 -2593
rect -513 -2981 -447 -2969
rect -417 -2593 -351 -2581
rect -417 -2969 -401 -2593
rect -367 -2969 -351 -2593
rect -417 -2981 -351 -2969
rect -321 -2593 -255 -2581
rect -321 -2969 -305 -2593
rect -271 -2969 -255 -2593
rect -321 -2981 -255 -2969
rect -225 -2593 -159 -2581
rect -225 -2969 -209 -2593
rect -175 -2969 -159 -2593
rect -225 -2981 -159 -2969
rect -129 -2593 -63 -2581
rect -129 -2969 -113 -2593
rect -79 -2969 -63 -2593
rect -129 -2981 -63 -2969
rect -33 -2593 33 -2581
rect -33 -2969 -17 -2593
rect 17 -2969 33 -2593
rect -33 -2981 33 -2969
rect 63 -2593 129 -2581
rect 63 -2969 79 -2593
rect 113 -2969 129 -2593
rect 63 -2981 129 -2969
rect 159 -2593 225 -2581
rect 159 -2969 175 -2593
rect 209 -2969 225 -2593
rect 159 -2981 225 -2969
rect 255 -2593 321 -2581
rect 255 -2969 271 -2593
rect 305 -2969 321 -2593
rect 255 -2981 321 -2969
rect 351 -2593 417 -2581
rect 351 -2969 367 -2593
rect 401 -2969 417 -2593
rect 351 -2981 417 -2969
rect 447 -2593 513 -2581
rect 447 -2969 463 -2593
rect 497 -2969 513 -2593
rect 447 -2981 513 -2969
rect 543 -2593 609 -2581
rect 543 -2969 559 -2593
rect 593 -2969 609 -2593
rect 543 -2981 609 -2969
rect 639 -2593 705 -2581
rect 639 -2969 655 -2593
rect 689 -2969 705 -2593
rect 639 -2981 705 -2969
rect 735 -2593 801 -2581
rect 735 -2969 751 -2593
rect 785 -2969 801 -2593
rect 735 -2981 801 -2969
rect 831 -2593 897 -2581
rect 831 -2969 847 -2593
rect 881 -2969 897 -2593
rect 831 -2981 897 -2969
rect 927 -2593 993 -2581
rect 927 -2969 943 -2593
rect 977 -2969 993 -2593
rect 927 -2981 993 -2969
rect 1023 -2593 1089 -2581
rect 1023 -2969 1039 -2593
rect 1073 -2969 1089 -2593
rect 1023 -2981 1089 -2969
rect 1119 -2593 1181 -2581
rect 1119 -2969 1135 -2593
rect 1169 -2969 1181 -2593
rect 1119 -2981 1181 -2969
<< ndiffc >>
rect -1169 2593 -1135 2969
rect -1073 2593 -1039 2969
rect -977 2593 -943 2969
rect -881 2593 -847 2969
rect -785 2593 -751 2969
rect -689 2593 -655 2969
rect -593 2593 -559 2969
rect -497 2593 -463 2969
rect -401 2593 -367 2969
rect -305 2593 -271 2969
rect -209 2593 -175 2969
rect -113 2593 -79 2969
rect -17 2593 17 2969
rect 79 2593 113 2969
rect 175 2593 209 2969
rect 271 2593 305 2969
rect 367 2593 401 2969
rect 463 2593 497 2969
rect 559 2593 593 2969
rect 655 2593 689 2969
rect 751 2593 785 2969
rect 847 2593 881 2969
rect 943 2593 977 2969
rect 1039 2593 1073 2969
rect 1135 2593 1169 2969
rect -1169 1975 -1135 2351
rect -1073 1975 -1039 2351
rect -977 1975 -943 2351
rect -881 1975 -847 2351
rect -785 1975 -751 2351
rect -689 1975 -655 2351
rect -593 1975 -559 2351
rect -497 1975 -463 2351
rect -401 1975 -367 2351
rect -305 1975 -271 2351
rect -209 1975 -175 2351
rect -113 1975 -79 2351
rect -17 1975 17 2351
rect 79 1975 113 2351
rect 175 1975 209 2351
rect 271 1975 305 2351
rect 367 1975 401 2351
rect 463 1975 497 2351
rect 559 1975 593 2351
rect 655 1975 689 2351
rect 751 1975 785 2351
rect 847 1975 881 2351
rect 943 1975 977 2351
rect 1039 1975 1073 2351
rect 1135 1975 1169 2351
rect -1169 1357 -1135 1733
rect -1073 1357 -1039 1733
rect -977 1357 -943 1733
rect -881 1357 -847 1733
rect -785 1357 -751 1733
rect -689 1357 -655 1733
rect -593 1357 -559 1733
rect -497 1357 -463 1733
rect -401 1357 -367 1733
rect -305 1357 -271 1733
rect -209 1357 -175 1733
rect -113 1357 -79 1733
rect -17 1357 17 1733
rect 79 1357 113 1733
rect 175 1357 209 1733
rect 271 1357 305 1733
rect 367 1357 401 1733
rect 463 1357 497 1733
rect 559 1357 593 1733
rect 655 1357 689 1733
rect 751 1357 785 1733
rect 847 1357 881 1733
rect 943 1357 977 1733
rect 1039 1357 1073 1733
rect 1135 1357 1169 1733
rect -1169 739 -1135 1115
rect -1073 739 -1039 1115
rect -977 739 -943 1115
rect -881 739 -847 1115
rect -785 739 -751 1115
rect -689 739 -655 1115
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect 655 739 689 1115
rect 751 739 785 1115
rect 847 739 881 1115
rect 943 739 977 1115
rect 1039 739 1073 1115
rect 1135 739 1169 1115
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect -1169 -1115 -1135 -739
rect -1073 -1115 -1039 -739
rect -977 -1115 -943 -739
rect -881 -1115 -847 -739
rect -785 -1115 -751 -739
rect -689 -1115 -655 -739
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect 655 -1115 689 -739
rect 751 -1115 785 -739
rect 847 -1115 881 -739
rect 943 -1115 977 -739
rect 1039 -1115 1073 -739
rect 1135 -1115 1169 -739
rect -1169 -1733 -1135 -1357
rect -1073 -1733 -1039 -1357
rect -977 -1733 -943 -1357
rect -881 -1733 -847 -1357
rect -785 -1733 -751 -1357
rect -689 -1733 -655 -1357
rect -593 -1733 -559 -1357
rect -497 -1733 -463 -1357
rect -401 -1733 -367 -1357
rect -305 -1733 -271 -1357
rect -209 -1733 -175 -1357
rect -113 -1733 -79 -1357
rect -17 -1733 17 -1357
rect 79 -1733 113 -1357
rect 175 -1733 209 -1357
rect 271 -1733 305 -1357
rect 367 -1733 401 -1357
rect 463 -1733 497 -1357
rect 559 -1733 593 -1357
rect 655 -1733 689 -1357
rect 751 -1733 785 -1357
rect 847 -1733 881 -1357
rect 943 -1733 977 -1357
rect 1039 -1733 1073 -1357
rect 1135 -1733 1169 -1357
rect -1169 -2351 -1135 -1975
rect -1073 -2351 -1039 -1975
rect -977 -2351 -943 -1975
rect -881 -2351 -847 -1975
rect -785 -2351 -751 -1975
rect -689 -2351 -655 -1975
rect -593 -2351 -559 -1975
rect -497 -2351 -463 -1975
rect -401 -2351 -367 -1975
rect -305 -2351 -271 -1975
rect -209 -2351 -175 -1975
rect -113 -2351 -79 -1975
rect -17 -2351 17 -1975
rect 79 -2351 113 -1975
rect 175 -2351 209 -1975
rect 271 -2351 305 -1975
rect 367 -2351 401 -1975
rect 463 -2351 497 -1975
rect 559 -2351 593 -1975
rect 655 -2351 689 -1975
rect 751 -2351 785 -1975
rect 847 -2351 881 -1975
rect 943 -2351 977 -1975
rect 1039 -2351 1073 -1975
rect 1135 -2351 1169 -1975
rect -1169 -2969 -1135 -2593
rect -1073 -2969 -1039 -2593
rect -977 -2969 -943 -2593
rect -881 -2969 -847 -2593
rect -785 -2969 -751 -2593
rect -689 -2969 -655 -2593
rect -593 -2969 -559 -2593
rect -497 -2969 -463 -2593
rect -401 -2969 -367 -2593
rect -305 -2969 -271 -2593
rect -209 -2969 -175 -2593
rect -113 -2969 -79 -2593
rect -17 -2969 17 -2593
rect 79 -2969 113 -2593
rect 175 -2969 209 -2593
rect 271 -2969 305 -2593
rect 367 -2969 401 -2593
rect 463 -2969 497 -2593
rect 559 -2969 593 -2593
rect 655 -2969 689 -2593
rect 751 -2969 785 -2593
rect 847 -2969 881 -2593
rect 943 -2969 977 -2593
rect 1039 -2969 1073 -2593
rect 1135 -2969 1169 -2593
<< psubdiff >>
rect -1283 3121 -1187 3155
rect 1187 3121 1283 3155
rect -1283 3059 -1249 3121
rect 1249 3059 1283 3121
rect -1283 -3121 -1249 -3059
rect 1249 -3121 1283 -3059
rect -1283 -3155 -1187 -3121
rect 1187 -3155 1283 -3121
<< psubdiffcont >>
rect -1187 3121 1187 3155
rect -1283 -3059 -1249 3059
rect 1249 -3059 1283 3059
rect -1187 -3155 1187 -3121
<< poly >>
rect -1137 3053 -1071 3069
rect -1137 3019 -1121 3053
rect -1087 3019 -1071 3053
rect -1137 3003 -1071 3019
rect -945 3053 -879 3069
rect -945 3019 -929 3053
rect -895 3019 -879 3053
rect -1119 2981 -1089 3003
rect -1023 2981 -993 3007
rect -945 3003 -879 3019
rect -753 3053 -687 3069
rect -753 3019 -737 3053
rect -703 3019 -687 3053
rect -927 2981 -897 3003
rect -831 2981 -801 3007
rect -753 3003 -687 3019
rect -561 3053 -495 3069
rect -561 3019 -545 3053
rect -511 3019 -495 3053
rect -735 2981 -705 3003
rect -639 2981 -609 3007
rect -561 3003 -495 3019
rect -369 3053 -303 3069
rect -369 3019 -353 3053
rect -319 3019 -303 3053
rect -543 2981 -513 3003
rect -447 2981 -417 3007
rect -369 3003 -303 3019
rect -177 3053 -111 3069
rect -177 3019 -161 3053
rect -127 3019 -111 3053
rect -351 2981 -321 3003
rect -255 2981 -225 3007
rect -177 3003 -111 3019
rect 15 3053 81 3069
rect 15 3019 31 3053
rect 65 3019 81 3053
rect -159 2981 -129 3003
rect -63 2981 -33 3007
rect 15 3003 81 3019
rect 207 3053 273 3069
rect 207 3019 223 3053
rect 257 3019 273 3053
rect 33 2981 63 3003
rect 129 2981 159 3007
rect 207 3003 273 3019
rect 399 3053 465 3069
rect 399 3019 415 3053
rect 449 3019 465 3053
rect 225 2981 255 3003
rect 321 2981 351 3007
rect 399 3003 465 3019
rect 591 3053 657 3069
rect 591 3019 607 3053
rect 641 3019 657 3053
rect 417 2981 447 3003
rect 513 2981 543 3007
rect 591 3003 657 3019
rect 783 3053 849 3069
rect 783 3019 799 3053
rect 833 3019 849 3053
rect 609 2981 639 3003
rect 705 2981 735 3007
rect 783 3003 849 3019
rect 975 3053 1041 3069
rect 975 3019 991 3053
rect 1025 3019 1041 3053
rect 801 2981 831 3003
rect 897 2981 927 3007
rect 975 3003 1041 3019
rect 993 2981 1023 3003
rect 1089 2981 1119 3007
rect -1119 2555 -1089 2581
rect -1023 2559 -993 2581
rect -1041 2543 -975 2559
rect -927 2555 -897 2581
rect -831 2559 -801 2581
rect -1041 2509 -1025 2543
rect -991 2509 -975 2543
rect -1041 2493 -975 2509
rect -849 2543 -783 2559
rect -735 2555 -705 2581
rect -639 2559 -609 2581
rect -849 2509 -833 2543
rect -799 2509 -783 2543
rect -849 2493 -783 2509
rect -657 2543 -591 2559
rect -543 2555 -513 2581
rect -447 2559 -417 2581
rect -657 2509 -641 2543
rect -607 2509 -591 2543
rect -657 2493 -591 2509
rect -465 2543 -399 2559
rect -351 2555 -321 2581
rect -255 2559 -225 2581
rect -465 2509 -449 2543
rect -415 2509 -399 2543
rect -465 2493 -399 2509
rect -273 2543 -207 2559
rect -159 2555 -129 2581
rect -63 2559 -33 2581
rect -273 2509 -257 2543
rect -223 2509 -207 2543
rect -273 2493 -207 2509
rect -81 2543 -15 2559
rect 33 2555 63 2581
rect 129 2559 159 2581
rect -81 2509 -65 2543
rect -31 2509 -15 2543
rect -81 2493 -15 2509
rect 111 2543 177 2559
rect 225 2555 255 2581
rect 321 2559 351 2581
rect 111 2509 127 2543
rect 161 2509 177 2543
rect 111 2493 177 2509
rect 303 2543 369 2559
rect 417 2555 447 2581
rect 513 2559 543 2581
rect 303 2509 319 2543
rect 353 2509 369 2543
rect 303 2493 369 2509
rect 495 2543 561 2559
rect 609 2555 639 2581
rect 705 2559 735 2581
rect 495 2509 511 2543
rect 545 2509 561 2543
rect 495 2493 561 2509
rect 687 2543 753 2559
rect 801 2555 831 2581
rect 897 2559 927 2581
rect 687 2509 703 2543
rect 737 2509 753 2543
rect 687 2493 753 2509
rect 879 2543 945 2559
rect 993 2555 1023 2581
rect 1089 2559 1119 2581
rect 879 2509 895 2543
rect 929 2509 945 2543
rect 879 2493 945 2509
rect 1071 2543 1137 2559
rect 1071 2509 1087 2543
rect 1121 2509 1137 2543
rect 1071 2493 1137 2509
rect -1041 2435 -975 2451
rect -1041 2401 -1025 2435
rect -991 2401 -975 2435
rect -1119 2363 -1089 2389
rect -1041 2385 -975 2401
rect -849 2435 -783 2451
rect -849 2401 -833 2435
rect -799 2401 -783 2435
rect -1023 2363 -993 2385
rect -927 2363 -897 2389
rect -849 2385 -783 2401
rect -657 2435 -591 2451
rect -657 2401 -641 2435
rect -607 2401 -591 2435
rect -831 2363 -801 2385
rect -735 2363 -705 2389
rect -657 2385 -591 2401
rect -465 2435 -399 2451
rect -465 2401 -449 2435
rect -415 2401 -399 2435
rect -639 2363 -609 2385
rect -543 2363 -513 2389
rect -465 2385 -399 2401
rect -273 2435 -207 2451
rect -273 2401 -257 2435
rect -223 2401 -207 2435
rect -447 2363 -417 2385
rect -351 2363 -321 2389
rect -273 2385 -207 2401
rect -81 2435 -15 2451
rect -81 2401 -65 2435
rect -31 2401 -15 2435
rect -255 2363 -225 2385
rect -159 2363 -129 2389
rect -81 2385 -15 2401
rect 111 2435 177 2451
rect 111 2401 127 2435
rect 161 2401 177 2435
rect -63 2363 -33 2385
rect 33 2363 63 2389
rect 111 2385 177 2401
rect 303 2435 369 2451
rect 303 2401 319 2435
rect 353 2401 369 2435
rect 129 2363 159 2385
rect 225 2363 255 2389
rect 303 2385 369 2401
rect 495 2435 561 2451
rect 495 2401 511 2435
rect 545 2401 561 2435
rect 321 2363 351 2385
rect 417 2363 447 2389
rect 495 2385 561 2401
rect 687 2435 753 2451
rect 687 2401 703 2435
rect 737 2401 753 2435
rect 513 2363 543 2385
rect 609 2363 639 2389
rect 687 2385 753 2401
rect 879 2435 945 2451
rect 879 2401 895 2435
rect 929 2401 945 2435
rect 705 2363 735 2385
rect 801 2363 831 2389
rect 879 2385 945 2401
rect 1071 2435 1137 2451
rect 1071 2401 1087 2435
rect 1121 2401 1137 2435
rect 897 2363 927 2385
rect 993 2363 1023 2389
rect 1071 2385 1137 2401
rect 1089 2363 1119 2385
rect -1119 1941 -1089 1963
rect -1137 1925 -1071 1941
rect -1023 1937 -993 1963
rect -927 1941 -897 1963
rect -1137 1891 -1121 1925
rect -1087 1891 -1071 1925
rect -1137 1875 -1071 1891
rect -945 1925 -879 1941
rect -831 1937 -801 1963
rect -735 1941 -705 1963
rect -945 1891 -929 1925
rect -895 1891 -879 1925
rect -945 1875 -879 1891
rect -753 1925 -687 1941
rect -639 1937 -609 1963
rect -543 1941 -513 1963
rect -753 1891 -737 1925
rect -703 1891 -687 1925
rect -753 1875 -687 1891
rect -561 1925 -495 1941
rect -447 1937 -417 1963
rect -351 1941 -321 1963
rect -561 1891 -545 1925
rect -511 1891 -495 1925
rect -561 1875 -495 1891
rect -369 1925 -303 1941
rect -255 1937 -225 1963
rect -159 1941 -129 1963
rect -369 1891 -353 1925
rect -319 1891 -303 1925
rect -369 1875 -303 1891
rect -177 1925 -111 1941
rect -63 1937 -33 1963
rect 33 1941 63 1963
rect -177 1891 -161 1925
rect -127 1891 -111 1925
rect -177 1875 -111 1891
rect 15 1925 81 1941
rect 129 1937 159 1963
rect 225 1941 255 1963
rect 15 1891 31 1925
rect 65 1891 81 1925
rect 15 1875 81 1891
rect 207 1925 273 1941
rect 321 1937 351 1963
rect 417 1941 447 1963
rect 207 1891 223 1925
rect 257 1891 273 1925
rect 207 1875 273 1891
rect 399 1925 465 1941
rect 513 1937 543 1963
rect 609 1941 639 1963
rect 399 1891 415 1925
rect 449 1891 465 1925
rect 399 1875 465 1891
rect 591 1925 657 1941
rect 705 1937 735 1963
rect 801 1941 831 1963
rect 591 1891 607 1925
rect 641 1891 657 1925
rect 591 1875 657 1891
rect 783 1925 849 1941
rect 897 1937 927 1963
rect 993 1941 1023 1963
rect 783 1891 799 1925
rect 833 1891 849 1925
rect 783 1875 849 1891
rect 975 1925 1041 1941
rect 1089 1937 1119 1963
rect 975 1891 991 1925
rect 1025 1891 1041 1925
rect 975 1875 1041 1891
rect -1137 1817 -1071 1833
rect -1137 1783 -1121 1817
rect -1087 1783 -1071 1817
rect -1137 1767 -1071 1783
rect -945 1817 -879 1833
rect -945 1783 -929 1817
rect -895 1783 -879 1817
rect -1119 1745 -1089 1767
rect -1023 1745 -993 1771
rect -945 1767 -879 1783
rect -753 1817 -687 1833
rect -753 1783 -737 1817
rect -703 1783 -687 1817
rect -927 1745 -897 1767
rect -831 1745 -801 1771
rect -753 1767 -687 1783
rect -561 1817 -495 1833
rect -561 1783 -545 1817
rect -511 1783 -495 1817
rect -735 1745 -705 1767
rect -639 1745 -609 1771
rect -561 1767 -495 1783
rect -369 1817 -303 1833
rect -369 1783 -353 1817
rect -319 1783 -303 1817
rect -543 1745 -513 1767
rect -447 1745 -417 1771
rect -369 1767 -303 1783
rect -177 1817 -111 1833
rect -177 1783 -161 1817
rect -127 1783 -111 1817
rect -351 1745 -321 1767
rect -255 1745 -225 1771
rect -177 1767 -111 1783
rect 15 1817 81 1833
rect 15 1783 31 1817
rect 65 1783 81 1817
rect -159 1745 -129 1767
rect -63 1745 -33 1771
rect 15 1767 81 1783
rect 207 1817 273 1833
rect 207 1783 223 1817
rect 257 1783 273 1817
rect 33 1745 63 1767
rect 129 1745 159 1771
rect 207 1767 273 1783
rect 399 1817 465 1833
rect 399 1783 415 1817
rect 449 1783 465 1817
rect 225 1745 255 1767
rect 321 1745 351 1771
rect 399 1767 465 1783
rect 591 1817 657 1833
rect 591 1783 607 1817
rect 641 1783 657 1817
rect 417 1745 447 1767
rect 513 1745 543 1771
rect 591 1767 657 1783
rect 783 1817 849 1833
rect 783 1783 799 1817
rect 833 1783 849 1817
rect 609 1745 639 1767
rect 705 1745 735 1771
rect 783 1767 849 1783
rect 975 1817 1041 1833
rect 975 1783 991 1817
rect 1025 1783 1041 1817
rect 801 1745 831 1767
rect 897 1745 927 1771
rect 975 1767 1041 1783
rect 993 1745 1023 1767
rect 1089 1745 1119 1771
rect -1119 1319 -1089 1345
rect -1023 1323 -993 1345
rect -1041 1307 -975 1323
rect -927 1319 -897 1345
rect -831 1323 -801 1345
rect -1041 1273 -1025 1307
rect -991 1273 -975 1307
rect -1041 1257 -975 1273
rect -849 1307 -783 1323
rect -735 1319 -705 1345
rect -639 1323 -609 1345
rect -849 1273 -833 1307
rect -799 1273 -783 1307
rect -849 1257 -783 1273
rect -657 1307 -591 1323
rect -543 1319 -513 1345
rect -447 1323 -417 1345
rect -657 1273 -641 1307
rect -607 1273 -591 1307
rect -657 1257 -591 1273
rect -465 1307 -399 1323
rect -351 1319 -321 1345
rect -255 1323 -225 1345
rect -465 1273 -449 1307
rect -415 1273 -399 1307
rect -465 1257 -399 1273
rect -273 1307 -207 1323
rect -159 1319 -129 1345
rect -63 1323 -33 1345
rect -273 1273 -257 1307
rect -223 1273 -207 1307
rect -273 1257 -207 1273
rect -81 1307 -15 1323
rect 33 1319 63 1345
rect 129 1323 159 1345
rect -81 1273 -65 1307
rect -31 1273 -15 1307
rect -81 1257 -15 1273
rect 111 1307 177 1323
rect 225 1319 255 1345
rect 321 1323 351 1345
rect 111 1273 127 1307
rect 161 1273 177 1307
rect 111 1257 177 1273
rect 303 1307 369 1323
rect 417 1319 447 1345
rect 513 1323 543 1345
rect 303 1273 319 1307
rect 353 1273 369 1307
rect 303 1257 369 1273
rect 495 1307 561 1323
rect 609 1319 639 1345
rect 705 1323 735 1345
rect 495 1273 511 1307
rect 545 1273 561 1307
rect 495 1257 561 1273
rect 687 1307 753 1323
rect 801 1319 831 1345
rect 897 1323 927 1345
rect 687 1273 703 1307
rect 737 1273 753 1307
rect 687 1257 753 1273
rect 879 1307 945 1323
rect 993 1319 1023 1345
rect 1089 1323 1119 1345
rect 879 1273 895 1307
rect 929 1273 945 1307
rect 879 1257 945 1273
rect 1071 1307 1137 1323
rect 1071 1273 1087 1307
rect 1121 1273 1137 1307
rect 1071 1257 1137 1273
rect -1041 1199 -975 1215
rect -1041 1165 -1025 1199
rect -991 1165 -975 1199
rect -1119 1127 -1089 1153
rect -1041 1149 -975 1165
rect -849 1199 -783 1215
rect -849 1165 -833 1199
rect -799 1165 -783 1199
rect -1023 1127 -993 1149
rect -927 1127 -897 1153
rect -849 1149 -783 1165
rect -657 1199 -591 1215
rect -657 1165 -641 1199
rect -607 1165 -591 1199
rect -831 1127 -801 1149
rect -735 1127 -705 1153
rect -657 1149 -591 1165
rect -465 1199 -399 1215
rect -465 1165 -449 1199
rect -415 1165 -399 1199
rect -639 1127 -609 1149
rect -543 1127 -513 1153
rect -465 1149 -399 1165
rect -273 1199 -207 1215
rect -273 1165 -257 1199
rect -223 1165 -207 1199
rect -447 1127 -417 1149
rect -351 1127 -321 1153
rect -273 1149 -207 1165
rect -81 1199 -15 1215
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect -255 1127 -225 1149
rect -159 1127 -129 1153
rect -81 1149 -15 1165
rect 111 1199 177 1215
rect 111 1165 127 1199
rect 161 1165 177 1199
rect -63 1127 -33 1149
rect 33 1127 63 1153
rect 111 1149 177 1165
rect 303 1199 369 1215
rect 303 1165 319 1199
rect 353 1165 369 1199
rect 129 1127 159 1149
rect 225 1127 255 1153
rect 303 1149 369 1165
rect 495 1199 561 1215
rect 495 1165 511 1199
rect 545 1165 561 1199
rect 321 1127 351 1149
rect 417 1127 447 1153
rect 495 1149 561 1165
rect 687 1199 753 1215
rect 687 1165 703 1199
rect 737 1165 753 1199
rect 513 1127 543 1149
rect 609 1127 639 1153
rect 687 1149 753 1165
rect 879 1199 945 1215
rect 879 1165 895 1199
rect 929 1165 945 1199
rect 705 1127 735 1149
rect 801 1127 831 1153
rect 879 1149 945 1165
rect 1071 1199 1137 1215
rect 1071 1165 1087 1199
rect 1121 1165 1137 1199
rect 897 1127 927 1149
rect 993 1127 1023 1153
rect 1071 1149 1137 1165
rect 1089 1127 1119 1149
rect -1119 705 -1089 727
rect -1137 689 -1071 705
rect -1023 701 -993 727
rect -927 705 -897 727
rect -1137 655 -1121 689
rect -1087 655 -1071 689
rect -1137 639 -1071 655
rect -945 689 -879 705
rect -831 701 -801 727
rect -735 705 -705 727
rect -945 655 -929 689
rect -895 655 -879 689
rect -945 639 -879 655
rect -753 689 -687 705
rect -639 701 -609 727
rect -543 705 -513 727
rect -753 655 -737 689
rect -703 655 -687 689
rect -753 639 -687 655
rect -561 689 -495 705
rect -447 701 -417 727
rect -351 705 -321 727
rect -561 655 -545 689
rect -511 655 -495 689
rect -561 639 -495 655
rect -369 689 -303 705
rect -255 701 -225 727
rect -159 705 -129 727
rect -369 655 -353 689
rect -319 655 -303 689
rect -369 639 -303 655
rect -177 689 -111 705
rect -63 701 -33 727
rect 33 705 63 727
rect -177 655 -161 689
rect -127 655 -111 689
rect -177 639 -111 655
rect 15 689 81 705
rect 129 701 159 727
rect 225 705 255 727
rect 15 655 31 689
rect 65 655 81 689
rect 15 639 81 655
rect 207 689 273 705
rect 321 701 351 727
rect 417 705 447 727
rect 207 655 223 689
rect 257 655 273 689
rect 207 639 273 655
rect 399 689 465 705
rect 513 701 543 727
rect 609 705 639 727
rect 399 655 415 689
rect 449 655 465 689
rect 399 639 465 655
rect 591 689 657 705
rect 705 701 735 727
rect 801 705 831 727
rect 591 655 607 689
rect 641 655 657 689
rect 591 639 657 655
rect 783 689 849 705
rect 897 701 927 727
rect 993 705 1023 727
rect 783 655 799 689
rect 833 655 849 689
rect 783 639 849 655
rect 975 689 1041 705
rect 1089 701 1119 727
rect 975 655 991 689
rect 1025 655 1041 689
rect 975 639 1041 655
rect -1137 581 -1071 597
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -1137 531 -1071 547
rect -945 581 -879 597
rect -945 547 -929 581
rect -895 547 -879 581
rect -1119 509 -1089 531
rect -1023 509 -993 535
rect -945 531 -879 547
rect -753 581 -687 597
rect -753 547 -737 581
rect -703 547 -687 581
rect -927 509 -897 531
rect -831 509 -801 535
rect -753 531 -687 547
rect -561 581 -495 597
rect -561 547 -545 581
rect -511 547 -495 581
rect -735 509 -705 531
rect -639 509 -609 535
rect -561 531 -495 547
rect -369 581 -303 597
rect -369 547 -353 581
rect -319 547 -303 581
rect -543 509 -513 531
rect -447 509 -417 535
rect -369 531 -303 547
rect -177 581 -111 597
rect -177 547 -161 581
rect -127 547 -111 581
rect -351 509 -321 531
rect -255 509 -225 535
rect -177 531 -111 547
rect 15 581 81 597
rect 15 547 31 581
rect 65 547 81 581
rect -159 509 -129 531
rect -63 509 -33 535
rect 15 531 81 547
rect 207 581 273 597
rect 207 547 223 581
rect 257 547 273 581
rect 33 509 63 531
rect 129 509 159 535
rect 207 531 273 547
rect 399 581 465 597
rect 399 547 415 581
rect 449 547 465 581
rect 225 509 255 531
rect 321 509 351 535
rect 399 531 465 547
rect 591 581 657 597
rect 591 547 607 581
rect 641 547 657 581
rect 417 509 447 531
rect 513 509 543 535
rect 591 531 657 547
rect 783 581 849 597
rect 783 547 799 581
rect 833 547 849 581
rect 609 509 639 531
rect 705 509 735 535
rect 783 531 849 547
rect 975 581 1041 597
rect 975 547 991 581
rect 1025 547 1041 581
rect 801 509 831 531
rect 897 509 927 535
rect 975 531 1041 547
rect 993 509 1023 531
rect 1089 509 1119 535
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1089 -109 1119 -87
rect -1119 -531 -1089 -509
rect -1137 -547 -1071 -531
rect -1023 -535 -993 -509
rect -927 -531 -897 -509
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -1137 -597 -1071 -581
rect -945 -547 -879 -531
rect -831 -535 -801 -509
rect -735 -531 -705 -509
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -945 -597 -879 -581
rect -753 -547 -687 -531
rect -639 -535 -609 -509
rect -543 -531 -513 -509
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -753 -597 -687 -581
rect -561 -547 -495 -531
rect -447 -535 -417 -509
rect -351 -531 -321 -509
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -255 -535 -225 -509
rect -159 -531 -129 -509
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -63 -535 -33 -509
rect 33 -531 63 -509
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 129 -535 159 -509
rect 225 -531 255 -509
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 321 -535 351 -509
rect 417 -531 447 -509
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 513 -535 543 -509
rect 609 -531 639 -509
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
rect 591 -547 657 -531
rect 705 -535 735 -509
rect 801 -531 831 -509
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 591 -597 657 -581
rect 783 -547 849 -531
rect 897 -535 927 -509
rect 993 -531 1023 -509
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 783 -597 849 -581
rect 975 -547 1041 -531
rect 1089 -535 1119 -509
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 975 -597 1041 -581
rect -1137 -655 -1071 -639
rect -1137 -689 -1121 -655
rect -1087 -689 -1071 -655
rect -1137 -705 -1071 -689
rect -945 -655 -879 -639
rect -945 -689 -929 -655
rect -895 -689 -879 -655
rect -1119 -727 -1089 -705
rect -1023 -727 -993 -701
rect -945 -705 -879 -689
rect -753 -655 -687 -639
rect -753 -689 -737 -655
rect -703 -689 -687 -655
rect -927 -727 -897 -705
rect -831 -727 -801 -701
rect -753 -705 -687 -689
rect -561 -655 -495 -639
rect -561 -689 -545 -655
rect -511 -689 -495 -655
rect -735 -727 -705 -705
rect -639 -727 -609 -701
rect -561 -705 -495 -689
rect -369 -655 -303 -639
rect -369 -689 -353 -655
rect -319 -689 -303 -655
rect -543 -727 -513 -705
rect -447 -727 -417 -701
rect -369 -705 -303 -689
rect -177 -655 -111 -639
rect -177 -689 -161 -655
rect -127 -689 -111 -655
rect -351 -727 -321 -705
rect -255 -727 -225 -701
rect -177 -705 -111 -689
rect 15 -655 81 -639
rect 15 -689 31 -655
rect 65 -689 81 -655
rect -159 -727 -129 -705
rect -63 -727 -33 -701
rect 15 -705 81 -689
rect 207 -655 273 -639
rect 207 -689 223 -655
rect 257 -689 273 -655
rect 33 -727 63 -705
rect 129 -727 159 -701
rect 207 -705 273 -689
rect 399 -655 465 -639
rect 399 -689 415 -655
rect 449 -689 465 -655
rect 225 -727 255 -705
rect 321 -727 351 -701
rect 399 -705 465 -689
rect 591 -655 657 -639
rect 591 -689 607 -655
rect 641 -689 657 -655
rect 417 -727 447 -705
rect 513 -727 543 -701
rect 591 -705 657 -689
rect 783 -655 849 -639
rect 783 -689 799 -655
rect 833 -689 849 -655
rect 609 -727 639 -705
rect 705 -727 735 -701
rect 783 -705 849 -689
rect 975 -655 1041 -639
rect 975 -689 991 -655
rect 1025 -689 1041 -655
rect 801 -727 831 -705
rect 897 -727 927 -701
rect 975 -705 1041 -689
rect 993 -727 1023 -705
rect 1089 -727 1119 -701
rect -1119 -1153 -1089 -1127
rect -1023 -1149 -993 -1127
rect -1041 -1165 -975 -1149
rect -927 -1153 -897 -1127
rect -831 -1149 -801 -1127
rect -1041 -1199 -1025 -1165
rect -991 -1199 -975 -1165
rect -1041 -1215 -975 -1199
rect -849 -1165 -783 -1149
rect -735 -1153 -705 -1127
rect -639 -1149 -609 -1127
rect -849 -1199 -833 -1165
rect -799 -1199 -783 -1165
rect -849 -1215 -783 -1199
rect -657 -1165 -591 -1149
rect -543 -1153 -513 -1127
rect -447 -1149 -417 -1127
rect -657 -1199 -641 -1165
rect -607 -1199 -591 -1165
rect -657 -1215 -591 -1199
rect -465 -1165 -399 -1149
rect -351 -1153 -321 -1127
rect -255 -1149 -225 -1127
rect -465 -1199 -449 -1165
rect -415 -1199 -399 -1165
rect -465 -1215 -399 -1199
rect -273 -1165 -207 -1149
rect -159 -1153 -129 -1127
rect -63 -1149 -33 -1127
rect -273 -1199 -257 -1165
rect -223 -1199 -207 -1165
rect -273 -1215 -207 -1199
rect -81 -1165 -15 -1149
rect 33 -1153 63 -1127
rect 129 -1149 159 -1127
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect -81 -1215 -15 -1199
rect 111 -1165 177 -1149
rect 225 -1153 255 -1127
rect 321 -1149 351 -1127
rect 111 -1199 127 -1165
rect 161 -1199 177 -1165
rect 111 -1215 177 -1199
rect 303 -1165 369 -1149
rect 417 -1153 447 -1127
rect 513 -1149 543 -1127
rect 303 -1199 319 -1165
rect 353 -1199 369 -1165
rect 303 -1215 369 -1199
rect 495 -1165 561 -1149
rect 609 -1153 639 -1127
rect 705 -1149 735 -1127
rect 495 -1199 511 -1165
rect 545 -1199 561 -1165
rect 495 -1215 561 -1199
rect 687 -1165 753 -1149
rect 801 -1153 831 -1127
rect 897 -1149 927 -1127
rect 687 -1199 703 -1165
rect 737 -1199 753 -1165
rect 687 -1215 753 -1199
rect 879 -1165 945 -1149
rect 993 -1153 1023 -1127
rect 1089 -1149 1119 -1127
rect 879 -1199 895 -1165
rect 929 -1199 945 -1165
rect 879 -1215 945 -1199
rect 1071 -1165 1137 -1149
rect 1071 -1199 1087 -1165
rect 1121 -1199 1137 -1165
rect 1071 -1215 1137 -1199
rect -1041 -1273 -975 -1257
rect -1041 -1307 -1025 -1273
rect -991 -1307 -975 -1273
rect -1119 -1345 -1089 -1319
rect -1041 -1323 -975 -1307
rect -849 -1273 -783 -1257
rect -849 -1307 -833 -1273
rect -799 -1307 -783 -1273
rect -1023 -1345 -993 -1323
rect -927 -1345 -897 -1319
rect -849 -1323 -783 -1307
rect -657 -1273 -591 -1257
rect -657 -1307 -641 -1273
rect -607 -1307 -591 -1273
rect -831 -1345 -801 -1323
rect -735 -1345 -705 -1319
rect -657 -1323 -591 -1307
rect -465 -1273 -399 -1257
rect -465 -1307 -449 -1273
rect -415 -1307 -399 -1273
rect -639 -1345 -609 -1323
rect -543 -1345 -513 -1319
rect -465 -1323 -399 -1307
rect -273 -1273 -207 -1257
rect -273 -1307 -257 -1273
rect -223 -1307 -207 -1273
rect -447 -1345 -417 -1323
rect -351 -1345 -321 -1319
rect -273 -1323 -207 -1307
rect -81 -1273 -15 -1257
rect -81 -1307 -65 -1273
rect -31 -1307 -15 -1273
rect -255 -1345 -225 -1323
rect -159 -1345 -129 -1319
rect -81 -1323 -15 -1307
rect 111 -1273 177 -1257
rect 111 -1307 127 -1273
rect 161 -1307 177 -1273
rect -63 -1345 -33 -1323
rect 33 -1345 63 -1319
rect 111 -1323 177 -1307
rect 303 -1273 369 -1257
rect 303 -1307 319 -1273
rect 353 -1307 369 -1273
rect 129 -1345 159 -1323
rect 225 -1345 255 -1319
rect 303 -1323 369 -1307
rect 495 -1273 561 -1257
rect 495 -1307 511 -1273
rect 545 -1307 561 -1273
rect 321 -1345 351 -1323
rect 417 -1345 447 -1319
rect 495 -1323 561 -1307
rect 687 -1273 753 -1257
rect 687 -1307 703 -1273
rect 737 -1307 753 -1273
rect 513 -1345 543 -1323
rect 609 -1345 639 -1319
rect 687 -1323 753 -1307
rect 879 -1273 945 -1257
rect 879 -1307 895 -1273
rect 929 -1307 945 -1273
rect 705 -1345 735 -1323
rect 801 -1345 831 -1319
rect 879 -1323 945 -1307
rect 1071 -1273 1137 -1257
rect 1071 -1307 1087 -1273
rect 1121 -1307 1137 -1273
rect 897 -1345 927 -1323
rect 993 -1345 1023 -1319
rect 1071 -1323 1137 -1307
rect 1089 -1345 1119 -1323
rect -1119 -1767 -1089 -1745
rect -1137 -1783 -1071 -1767
rect -1023 -1771 -993 -1745
rect -927 -1767 -897 -1745
rect -1137 -1817 -1121 -1783
rect -1087 -1817 -1071 -1783
rect -1137 -1833 -1071 -1817
rect -945 -1783 -879 -1767
rect -831 -1771 -801 -1745
rect -735 -1767 -705 -1745
rect -945 -1817 -929 -1783
rect -895 -1817 -879 -1783
rect -945 -1833 -879 -1817
rect -753 -1783 -687 -1767
rect -639 -1771 -609 -1745
rect -543 -1767 -513 -1745
rect -753 -1817 -737 -1783
rect -703 -1817 -687 -1783
rect -753 -1833 -687 -1817
rect -561 -1783 -495 -1767
rect -447 -1771 -417 -1745
rect -351 -1767 -321 -1745
rect -561 -1817 -545 -1783
rect -511 -1817 -495 -1783
rect -561 -1833 -495 -1817
rect -369 -1783 -303 -1767
rect -255 -1771 -225 -1745
rect -159 -1767 -129 -1745
rect -369 -1817 -353 -1783
rect -319 -1817 -303 -1783
rect -369 -1833 -303 -1817
rect -177 -1783 -111 -1767
rect -63 -1771 -33 -1745
rect 33 -1767 63 -1745
rect -177 -1817 -161 -1783
rect -127 -1817 -111 -1783
rect -177 -1833 -111 -1817
rect 15 -1783 81 -1767
rect 129 -1771 159 -1745
rect 225 -1767 255 -1745
rect 15 -1817 31 -1783
rect 65 -1817 81 -1783
rect 15 -1833 81 -1817
rect 207 -1783 273 -1767
rect 321 -1771 351 -1745
rect 417 -1767 447 -1745
rect 207 -1817 223 -1783
rect 257 -1817 273 -1783
rect 207 -1833 273 -1817
rect 399 -1783 465 -1767
rect 513 -1771 543 -1745
rect 609 -1767 639 -1745
rect 399 -1817 415 -1783
rect 449 -1817 465 -1783
rect 399 -1833 465 -1817
rect 591 -1783 657 -1767
rect 705 -1771 735 -1745
rect 801 -1767 831 -1745
rect 591 -1817 607 -1783
rect 641 -1817 657 -1783
rect 591 -1833 657 -1817
rect 783 -1783 849 -1767
rect 897 -1771 927 -1745
rect 993 -1767 1023 -1745
rect 783 -1817 799 -1783
rect 833 -1817 849 -1783
rect 783 -1833 849 -1817
rect 975 -1783 1041 -1767
rect 1089 -1771 1119 -1745
rect 975 -1817 991 -1783
rect 1025 -1817 1041 -1783
rect 975 -1833 1041 -1817
rect -1137 -1891 -1071 -1875
rect -1137 -1925 -1121 -1891
rect -1087 -1925 -1071 -1891
rect -1137 -1941 -1071 -1925
rect -945 -1891 -879 -1875
rect -945 -1925 -929 -1891
rect -895 -1925 -879 -1891
rect -1119 -1963 -1089 -1941
rect -1023 -1963 -993 -1937
rect -945 -1941 -879 -1925
rect -753 -1891 -687 -1875
rect -753 -1925 -737 -1891
rect -703 -1925 -687 -1891
rect -927 -1963 -897 -1941
rect -831 -1963 -801 -1937
rect -753 -1941 -687 -1925
rect -561 -1891 -495 -1875
rect -561 -1925 -545 -1891
rect -511 -1925 -495 -1891
rect -735 -1963 -705 -1941
rect -639 -1963 -609 -1937
rect -561 -1941 -495 -1925
rect -369 -1891 -303 -1875
rect -369 -1925 -353 -1891
rect -319 -1925 -303 -1891
rect -543 -1963 -513 -1941
rect -447 -1963 -417 -1937
rect -369 -1941 -303 -1925
rect -177 -1891 -111 -1875
rect -177 -1925 -161 -1891
rect -127 -1925 -111 -1891
rect -351 -1963 -321 -1941
rect -255 -1963 -225 -1937
rect -177 -1941 -111 -1925
rect 15 -1891 81 -1875
rect 15 -1925 31 -1891
rect 65 -1925 81 -1891
rect -159 -1963 -129 -1941
rect -63 -1963 -33 -1937
rect 15 -1941 81 -1925
rect 207 -1891 273 -1875
rect 207 -1925 223 -1891
rect 257 -1925 273 -1891
rect 33 -1963 63 -1941
rect 129 -1963 159 -1937
rect 207 -1941 273 -1925
rect 399 -1891 465 -1875
rect 399 -1925 415 -1891
rect 449 -1925 465 -1891
rect 225 -1963 255 -1941
rect 321 -1963 351 -1937
rect 399 -1941 465 -1925
rect 591 -1891 657 -1875
rect 591 -1925 607 -1891
rect 641 -1925 657 -1891
rect 417 -1963 447 -1941
rect 513 -1963 543 -1937
rect 591 -1941 657 -1925
rect 783 -1891 849 -1875
rect 783 -1925 799 -1891
rect 833 -1925 849 -1891
rect 609 -1963 639 -1941
rect 705 -1963 735 -1937
rect 783 -1941 849 -1925
rect 975 -1891 1041 -1875
rect 975 -1925 991 -1891
rect 1025 -1925 1041 -1891
rect 801 -1963 831 -1941
rect 897 -1963 927 -1937
rect 975 -1941 1041 -1925
rect 993 -1963 1023 -1941
rect 1089 -1963 1119 -1937
rect -1119 -2389 -1089 -2363
rect -1023 -2385 -993 -2363
rect -1041 -2401 -975 -2385
rect -927 -2389 -897 -2363
rect -831 -2385 -801 -2363
rect -1041 -2435 -1025 -2401
rect -991 -2435 -975 -2401
rect -1041 -2451 -975 -2435
rect -849 -2401 -783 -2385
rect -735 -2389 -705 -2363
rect -639 -2385 -609 -2363
rect -849 -2435 -833 -2401
rect -799 -2435 -783 -2401
rect -849 -2451 -783 -2435
rect -657 -2401 -591 -2385
rect -543 -2389 -513 -2363
rect -447 -2385 -417 -2363
rect -657 -2435 -641 -2401
rect -607 -2435 -591 -2401
rect -657 -2451 -591 -2435
rect -465 -2401 -399 -2385
rect -351 -2389 -321 -2363
rect -255 -2385 -225 -2363
rect -465 -2435 -449 -2401
rect -415 -2435 -399 -2401
rect -465 -2451 -399 -2435
rect -273 -2401 -207 -2385
rect -159 -2389 -129 -2363
rect -63 -2385 -33 -2363
rect -273 -2435 -257 -2401
rect -223 -2435 -207 -2401
rect -273 -2451 -207 -2435
rect -81 -2401 -15 -2385
rect 33 -2389 63 -2363
rect 129 -2385 159 -2363
rect -81 -2435 -65 -2401
rect -31 -2435 -15 -2401
rect -81 -2451 -15 -2435
rect 111 -2401 177 -2385
rect 225 -2389 255 -2363
rect 321 -2385 351 -2363
rect 111 -2435 127 -2401
rect 161 -2435 177 -2401
rect 111 -2451 177 -2435
rect 303 -2401 369 -2385
rect 417 -2389 447 -2363
rect 513 -2385 543 -2363
rect 303 -2435 319 -2401
rect 353 -2435 369 -2401
rect 303 -2451 369 -2435
rect 495 -2401 561 -2385
rect 609 -2389 639 -2363
rect 705 -2385 735 -2363
rect 495 -2435 511 -2401
rect 545 -2435 561 -2401
rect 495 -2451 561 -2435
rect 687 -2401 753 -2385
rect 801 -2389 831 -2363
rect 897 -2385 927 -2363
rect 687 -2435 703 -2401
rect 737 -2435 753 -2401
rect 687 -2451 753 -2435
rect 879 -2401 945 -2385
rect 993 -2389 1023 -2363
rect 1089 -2385 1119 -2363
rect 879 -2435 895 -2401
rect 929 -2435 945 -2401
rect 879 -2451 945 -2435
rect 1071 -2401 1137 -2385
rect 1071 -2435 1087 -2401
rect 1121 -2435 1137 -2401
rect 1071 -2451 1137 -2435
rect -1041 -2509 -975 -2493
rect -1041 -2543 -1025 -2509
rect -991 -2543 -975 -2509
rect -1119 -2581 -1089 -2555
rect -1041 -2559 -975 -2543
rect -849 -2509 -783 -2493
rect -849 -2543 -833 -2509
rect -799 -2543 -783 -2509
rect -1023 -2581 -993 -2559
rect -927 -2581 -897 -2555
rect -849 -2559 -783 -2543
rect -657 -2509 -591 -2493
rect -657 -2543 -641 -2509
rect -607 -2543 -591 -2509
rect -831 -2581 -801 -2559
rect -735 -2581 -705 -2555
rect -657 -2559 -591 -2543
rect -465 -2509 -399 -2493
rect -465 -2543 -449 -2509
rect -415 -2543 -399 -2509
rect -639 -2581 -609 -2559
rect -543 -2581 -513 -2555
rect -465 -2559 -399 -2543
rect -273 -2509 -207 -2493
rect -273 -2543 -257 -2509
rect -223 -2543 -207 -2509
rect -447 -2581 -417 -2559
rect -351 -2581 -321 -2555
rect -273 -2559 -207 -2543
rect -81 -2509 -15 -2493
rect -81 -2543 -65 -2509
rect -31 -2543 -15 -2509
rect -255 -2581 -225 -2559
rect -159 -2581 -129 -2555
rect -81 -2559 -15 -2543
rect 111 -2509 177 -2493
rect 111 -2543 127 -2509
rect 161 -2543 177 -2509
rect -63 -2581 -33 -2559
rect 33 -2581 63 -2555
rect 111 -2559 177 -2543
rect 303 -2509 369 -2493
rect 303 -2543 319 -2509
rect 353 -2543 369 -2509
rect 129 -2581 159 -2559
rect 225 -2581 255 -2555
rect 303 -2559 369 -2543
rect 495 -2509 561 -2493
rect 495 -2543 511 -2509
rect 545 -2543 561 -2509
rect 321 -2581 351 -2559
rect 417 -2581 447 -2555
rect 495 -2559 561 -2543
rect 687 -2509 753 -2493
rect 687 -2543 703 -2509
rect 737 -2543 753 -2509
rect 513 -2581 543 -2559
rect 609 -2581 639 -2555
rect 687 -2559 753 -2543
rect 879 -2509 945 -2493
rect 879 -2543 895 -2509
rect 929 -2543 945 -2509
rect 705 -2581 735 -2559
rect 801 -2581 831 -2555
rect 879 -2559 945 -2543
rect 1071 -2509 1137 -2493
rect 1071 -2543 1087 -2509
rect 1121 -2543 1137 -2509
rect 897 -2581 927 -2559
rect 993 -2581 1023 -2555
rect 1071 -2559 1137 -2543
rect 1089 -2581 1119 -2559
rect -1119 -3003 -1089 -2981
rect -1137 -3019 -1071 -3003
rect -1023 -3007 -993 -2981
rect -927 -3003 -897 -2981
rect -1137 -3053 -1121 -3019
rect -1087 -3053 -1071 -3019
rect -1137 -3069 -1071 -3053
rect -945 -3019 -879 -3003
rect -831 -3007 -801 -2981
rect -735 -3003 -705 -2981
rect -945 -3053 -929 -3019
rect -895 -3053 -879 -3019
rect -945 -3069 -879 -3053
rect -753 -3019 -687 -3003
rect -639 -3007 -609 -2981
rect -543 -3003 -513 -2981
rect -753 -3053 -737 -3019
rect -703 -3053 -687 -3019
rect -753 -3069 -687 -3053
rect -561 -3019 -495 -3003
rect -447 -3007 -417 -2981
rect -351 -3003 -321 -2981
rect -561 -3053 -545 -3019
rect -511 -3053 -495 -3019
rect -561 -3069 -495 -3053
rect -369 -3019 -303 -3003
rect -255 -3007 -225 -2981
rect -159 -3003 -129 -2981
rect -369 -3053 -353 -3019
rect -319 -3053 -303 -3019
rect -369 -3069 -303 -3053
rect -177 -3019 -111 -3003
rect -63 -3007 -33 -2981
rect 33 -3003 63 -2981
rect -177 -3053 -161 -3019
rect -127 -3053 -111 -3019
rect -177 -3069 -111 -3053
rect 15 -3019 81 -3003
rect 129 -3007 159 -2981
rect 225 -3003 255 -2981
rect 15 -3053 31 -3019
rect 65 -3053 81 -3019
rect 15 -3069 81 -3053
rect 207 -3019 273 -3003
rect 321 -3007 351 -2981
rect 417 -3003 447 -2981
rect 207 -3053 223 -3019
rect 257 -3053 273 -3019
rect 207 -3069 273 -3053
rect 399 -3019 465 -3003
rect 513 -3007 543 -2981
rect 609 -3003 639 -2981
rect 399 -3053 415 -3019
rect 449 -3053 465 -3019
rect 399 -3069 465 -3053
rect 591 -3019 657 -3003
rect 705 -3007 735 -2981
rect 801 -3003 831 -2981
rect 591 -3053 607 -3019
rect 641 -3053 657 -3019
rect 591 -3069 657 -3053
rect 783 -3019 849 -3003
rect 897 -3007 927 -2981
rect 993 -3003 1023 -2981
rect 783 -3053 799 -3019
rect 833 -3053 849 -3019
rect 783 -3069 849 -3053
rect 975 -3019 1041 -3003
rect 1089 -3007 1119 -2981
rect 975 -3053 991 -3019
rect 1025 -3053 1041 -3019
rect 975 -3069 1041 -3053
<< polycont >>
rect -1121 3019 -1087 3053
rect -929 3019 -895 3053
rect -737 3019 -703 3053
rect -545 3019 -511 3053
rect -353 3019 -319 3053
rect -161 3019 -127 3053
rect 31 3019 65 3053
rect 223 3019 257 3053
rect 415 3019 449 3053
rect 607 3019 641 3053
rect 799 3019 833 3053
rect 991 3019 1025 3053
rect -1025 2509 -991 2543
rect -833 2509 -799 2543
rect -641 2509 -607 2543
rect -449 2509 -415 2543
rect -257 2509 -223 2543
rect -65 2509 -31 2543
rect 127 2509 161 2543
rect 319 2509 353 2543
rect 511 2509 545 2543
rect 703 2509 737 2543
rect 895 2509 929 2543
rect 1087 2509 1121 2543
rect -1025 2401 -991 2435
rect -833 2401 -799 2435
rect -641 2401 -607 2435
rect -449 2401 -415 2435
rect -257 2401 -223 2435
rect -65 2401 -31 2435
rect 127 2401 161 2435
rect 319 2401 353 2435
rect 511 2401 545 2435
rect 703 2401 737 2435
rect 895 2401 929 2435
rect 1087 2401 1121 2435
rect -1121 1891 -1087 1925
rect -929 1891 -895 1925
rect -737 1891 -703 1925
rect -545 1891 -511 1925
rect -353 1891 -319 1925
rect -161 1891 -127 1925
rect 31 1891 65 1925
rect 223 1891 257 1925
rect 415 1891 449 1925
rect 607 1891 641 1925
rect 799 1891 833 1925
rect 991 1891 1025 1925
rect -1121 1783 -1087 1817
rect -929 1783 -895 1817
rect -737 1783 -703 1817
rect -545 1783 -511 1817
rect -353 1783 -319 1817
rect -161 1783 -127 1817
rect 31 1783 65 1817
rect 223 1783 257 1817
rect 415 1783 449 1817
rect 607 1783 641 1817
rect 799 1783 833 1817
rect 991 1783 1025 1817
rect -1025 1273 -991 1307
rect -833 1273 -799 1307
rect -641 1273 -607 1307
rect -449 1273 -415 1307
rect -257 1273 -223 1307
rect -65 1273 -31 1307
rect 127 1273 161 1307
rect 319 1273 353 1307
rect 511 1273 545 1307
rect 703 1273 737 1307
rect 895 1273 929 1307
rect 1087 1273 1121 1307
rect -1025 1165 -991 1199
rect -833 1165 -799 1199
rect -641 1165 -607 1199
rect -449 1165 -415 1199
rect -257 1165 -223 1199
rect -65 1165 -31 1199
rect 127 1165 161 1199
rect 319 1165 353 1199
rect 511 1165 545 1199
rect 703 1165 737 1199
rect 895 1165 929 1199
rect 1087 1165 1121 1199
rect -1121 655 -1087 689
rect -929 655 -895 689
rect -737 655 -703 689
rect -545 655 -511 689
rect -353 655 -319 689
rect -161 655 -127 689
rect 31 655 65 689
rect 223 655 257 689
rect 415 655 449 689
rect 607 655 641 689
rect 799 655 833 689
rect 991 655 1025 689
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect -1121 -689 -1087 -655
rect -929 -689 -895 -655
rect -737 -689 -703 -655
rect -545 -689 -511 -655
rect -353 -689 -319 -655
rect -161 -689 -127 -655
rect 31 -689 65 -655
rect 223 -689 257 -655
rect 415 -689 449 -655
rect 607 -689 641 -655
rect 799 -689 833 -655
rect 991 -689 1025 -655
rect -1025 -1199 -991 -1165
rect -833 -1199 -799 -1165
rect -641 -1199 -607 -1165
rect -449 -1199 -415 -1165
rect -257 -1199 -223 -1165
rect -65 -1199 -31 -1165
rect 127 -1199 161 -1165
rect 319 -1199 353 -1165
rect 511 -1199 545 -1165
rect 703 -1199 737 -1165
rect 895 -1199 929 -1165
rect 1087 -1199 1121 -1165
rect -1025 -1307 -991 -1273
rect -833 -1307 -799 -1273
rect -641 -1307 -607 -1273
rect -449 -1307 -415 -1273
rect -257 -1307 -223 -1273
rect -65 -1307 -31 -1273
rect 127 -1307 161 -1273
rect 319 -1307 353 -1273
rect 511 -1307 545 -1273
rect 703 -1307 737 -1273
rect 895 -1307 929 -1273
rect 1087 -1307 1121 -1273
rect -1121 -1817 -1087 -1783
rect -929 -1817 -895 -1783
rect -737 -1817 -703 -1783
rect -545 -1817 -511 -1783
rect -353 -1817 -319 -1783
rect -161 -1817 -127 -1783
rect 31 -1817 65 -1783
rect 223 -1817 257 -1783
rect 415 -1817 449 -1783
rect 607 -1817 641 -1783
rect 799 -1817 833 -1783
rect 991 -1817 1025 -1783
rect -1121 -1925 -1087 -1891
rect -929 -1925 -895 -1891
rect -737 -1925 -703 -1891
rect -545 -1925 -511 -1891
rect -353 -1925 -319 -1891
rect -161 -1925 -127 -1891
rect 31 -1925 65 -1891
rect 223 -1925 257 -1891
rect 415 -1925 449 -1891
rect 607 -1925 641 -1891
rect 799 -1925 833 -1891
rect 991 -1925 1025 -1891
rect -1025 -2435 -991 -2401
rect -833 -2435 -799 -2401
rect -641 -2435 -607 -2401
rect -449 -2435 -415 -2401
rect -257 -2435 -223 -2401
rect -65 -2435 -31 -2401
rect 127 -2435 161 -2401
rect 319 -2435 353 -2401
rect 511 -2435 545 -2401
rect 703 -2435 737 -2401
rect 895 -2435 929 -2401
rect 1087 -2435 1121 -2401
rect -1025 -2543 -991 -2509
rect -833 -2543 -799 -2509
rect -641 -2543 -607 -2509
rect -449 -2543 -415 -2509
rect -257 -2543 -223 -2509
rect -65 -2543 -31 -2509
rect 127 -2543 161 -2509
rect 319 -2543 353 -2509
rect 511 -2543 545 -2509
rect 703 -2543 737 -2509
rect 895 -2543 929 -2509
rect 1087 -2543 1121 -2509
rect -1121 -3053 -1087 -3019
rect -929 -3053 -895 -3019
rect -737 -3053 -703 -3019
rect -545 -3053 -511 -3019
rect -353 -3053 -319 -3019
rect -161 -3053 -127 -3019
rect 31 -3053 65 -3019
rect 223 -3053 257 -3019
rect 415 -3053 449 -3019
rect 607 -3053 641 -3019
rect 799 -3053 833 -3019
rect 991 -3053 1025 -3019
<< locali >>
rect -1283 3121 -1187 3155
rect 1187 3121 1283 3155
rect -1283 3059 -1249 3121
rect 1249 3059 1283 3121
rect -1137 3019 -1121 3053
rect -1087 3019 -1071 3053
rect -945 3019 -929 3053
rect -895 3019 -879 3053
rect -753 3019 -737 3053
rect -703 3019 -687 3053
rect -561 3019 -545 3053
rect -511 3019 -495 3053
rect -369 3019 -353 3053
rect -319 3019 -303 3053
rect -177 3019 -161 3053
rect -127 3019 -111 3053
rect 15 3019 31 3053
rect 65 3019 81 3053
rect 207 3019 223 3053
rect 257 3019 273 3053
rect 399 3019 415 3053
rect 449 3019 465 3053
rect 591 3019 607 3053
rect 641 3019 657 3053
rect 783 3019 799 3053
rect 833 3019 849 3053
rect 975 3019 991 3053
rect 1025 3019 1041 3053
rect -1169 2969 -1135 2985
rect -1169 2577 -1135 2593
rect -1073 2969 -1039 2985
rect -1073 2577 -1039 2593
rect -977 2969 -943 2985
rect -977 2577 -943 2593
rect -881 2969 -847 2985
rect -881 2577 -847 2593
rect -785 2969 -751 2985
rect -785 2577 -751 2593
rect -689 2969 -655 2985
rect -689 2577 -655 2593
rect -593 2969 -559 2985
rect -593 2577 -559 2593
rect -497 2969 -463 2985
rect -497 2577 -463 2593
rect -401 2969 -367 2985
rect -401 2577 -367 2593
rect -305 2969 -271 2985
rect -305 2577 -271 2593
rect -209 2969 -175 2985
rect -209 2577 -175 2593
rect -113 2969 -79 2985
rect -113 2577 -79 2593
rect -17 2969 17 2985
rect -17 2577 17 2593
rect 79 2969 113 2985
rect 79 2577 113 2593
rect 175 2969 209 2985
rect 175 2577 209 2593
rect 271 2969 305 2985
rect 271 2577 305 2593
rect 367 2969 401 2985
rect 367 2577 401 2593
rect 463 2969 497 2985
rect 463 2577 497 2593
rect 559 2969 593 2985
rect 559 2577 593 2593
rect 655 2969 689 2985
rect 655 2577 689 2593
rect 751 2969 785 2985
rect 751 2577 785 2593
rect 847 2969 881 2985
rect 847 2577 881 2593
rect 943 2969 977 2985
rect 943 2577 977 2593
rect 1039 2969 1073 2985
rect 1039 2577 1073 2593
rect 1135 2969 1169 2985
rect 1135 2577 1169 2593
rect -1041 2509 -1025 2543
rect -991 2509 -975 2543
rect -849 2509 -833 2543
rect -799 2509 -783 2543
rect -657 2509 -641 2543
rect -607 2509 -591 2543
rect -465 2509 -449 2543
rect -415 2509 -399 2543
rect -273 2509 -257 2543
rect -223 2509 -207 2543
rect -81 2509 -65 2543
rect -31 2509 -15 2543
rect 111 2509 127 2543
rect 161 2509 177 2543
rect 303 2509 319 2543
rect 353 2509 369 2543
rect 495 2509 511 2543
rect 545 2509 561 2543
rect 687 2509 703 2543
rect 737 2509 753 2543
rect 879 2509 895 2543
rect 929 2509 945 2543
rect 1071 2509 1087 2543
rect 1121 2509 1137 2543
rect -1041 2401 -1025 2435
rect -991 2401 -975 2435
rect -849 2401 -833 2435
rect -799 2401 -783 2435
rect -657 2401 -641 2435
rect -607 2401 -591 2435
rect -465 2401 -449 2435
rect -415 2401 -399 2435
rect -273 2401 -257 2435
rect -223 2401 -207 2435
rect -81 2401 -65 2435
rect -31 2401 -15 2435
rect 111 2401 127 2435
rect 161 2401 177 2435
rect 303 2401 319 2435
rect 353 2401 369 2435
rect 495 2401 511 2435
rect 545 2401 561 2435
rect 687 2401 703 2435
rect 737 2401 753 2435
rect 879 2401 895 2435
rect 929 2401 945 2435
rect 1071 2401 1087 2435
rect 1121 2401 1137 2435
rect -1169 2351 -1135 2367
rect -1169 1959 -1135 1975
rect -1073 2351 -1039 2367
rect -1073 1959 -1039 1975
rect -977 2351 -943 2367
rect -977 1959 -943 1975
rect -881 2351 -847 2367
rect -881 1959 -847 1975
rect -785 2351 -751 2367
rect -785 1959 -751 1975
rect -689 2351 -655 2367
rect -689 1959 -655 1975
rect -593 2351 -559 2367
rect -593 1959 -559 1975
rect -497 2351 -463 2367
rect -497 1959 -463 1975
rect -401 2351 -367 2367
rect -401 1959 -367 1975
rect -305 2351 -271 2367
rect -305 1959 -271 1975
rect -209 2351 -175 2367
rect -209 1959 -175 1975
rect -113 2351 -79 2367
rect -113 1959 -79 1975
rect -17 2351 17 2367
rect -17 1959 17 1975
rect 79 2351 113 2367
rect 79 1959 113 1975
rect 175 2351 209 2367
rect 175 1959 209 1975
rect 271 2351 305 2367
rect 271 1959 305 1975
rect 367 2351 401 2367
rect 367 1959 401 1975
rect 463 2351 497 2367
rect 463 1959 497 1975
rect 559 2351 593 2367
rect 559 1959 593 1975
rect 655 2351 689 2367
rect 655 1959 689 1975
rect 751 2351 785 2367
rect 751 1959 785 1975
rect 847 2351 881 2367
rect 847 1959 881 1975
rect 943 2351 977 2367
rect 943 1959 977 1975
rect 1039 2351 1073 2367
rect 1039 1959 1073 1975
rect 1135 2351 1169 2367
rect 1135 1959 1169 1975
rect -1137 1891 -1121 1925
rect -1087 1891 -1071 1925
rect -945 1891 -929 1925
rect -895 1891 -879 1925
rect -753 1891 -737 1925
rect -703 1891 -687 1925
rect -561 1891 -545 1925
rect -511 1891 -495 1925
rect -369 1891 -353 1925
rect -319 1891 -303 1925
rect -177 1891 -161 1925
rect -127 1891 -111 1925
rect 15 1891 31 1925
rect 65 1891 81 1925
rect 207 1891 223 1925
rect 257 1891 273 1925
rect 399 1891 415 1925
rect 449 1891 465 1925
rect 591 1891 607 1925
rect 641 1891 657 1925
rect 783 1891 799 1925
rect 833 1891 849 1925
rect 975 1891 991 1925
rect 1025 1891 1041 1925
rect -1137 1783 -1121 1817
rect -1087 1783 -1071 1817
rect -945 1783 -929 1817
rect -895 1783 -879 1817
rect -753 1783 -737 1817
rect -703 1783 -687 1817
rect -561 1783 -545 1817
rect -511 1783 -495 1817
rect -369 1783 -353 1817
rect -319 1783 -303 1817
rect -177 1783 -161 1817
rect -127 1783 -111 1817
rect 15 1783 31 1817
rect 65 1783 81 1817
rect 207 1783 223 1817
rect 257 1783 273 1817
rect 399 1783 415 1817
rect 449 1783 465 1817
rect 591 1783 607 1817
rect 641 1783 657 1817
rect 783 1783 799 1817
rect 833 1783 849 1817
rect 975 1783 991 1817
rect 1025 1783 1041 1817
rect -1169 1733 -1135 1749
rect -1169 1341 -1135 1357
rect -1073 1733 -1039 1749
rect -1073 1341 -1039 1357
rect -977 1733 -943 1749
rect -977 1341 -943 1357
rect -881 1733 -847 1749
rect -881 1341 -847 1357
rect -785 1733 -751 1749
rect -785 1341 -751 1357
rect -689 1733 -655 1749
rect -689 1341 -655 1357
rect -593 1733 -559 1749
rect -593 1341 -559 1357
rect -497 1733 -463 1749
rect -497 1341 -463 1357
rect -401 1733 -367 1749
rect -401 1341 -367 1357
rect -305 1733 -271 1749
rect -305 1341 -271 1357
rect -209 1733 -175 1749
rect -209 1341 -175 1357
rect -113 1733 -79 1749
rect -113 1341 -79 1357
rect -17 1733 17 1749
rect -17 1341 17 1357
rect 79 1733 113 1749
rect 79 1341 113 1357
rect 175 1733 209 1749
rect 175 1341 209 1357
rect 271 1733 305 1749
rect 271 1341 305 1357
rect 367 1733 401 1749
rect 367 1341 401 1357
rect 463 1733 497 1749
rect 463 1341 497 1357
rect 559 1733 593 1749
rect 559 1341 593 1357
rect 655 1733 689 1749
rect 655 1341 689 1357
rect 751 1733 785 1749
rect 751 1341 785 1357
rect 847 1733 881 1749
rect 847 1341 881 1357
rect 943 1733 977 1749
rect 943 1341 977 1357
rect 1039 1733 1073 1749
rect 1039 1341 1073 1357
rect 1135 1733 1169 1749
rect 1135 1341 1169 1357
rect -1041 1273 -1025 1307
rect -991 1273 -975 1307
rect -849 1273 -833 1307
rect -799 1273 -783 1307
rect -657 1273 -641 1307
rect -607 1273 -591 1307
rect -465 1273 -449 1307
rect -415 1273 -399 1307
rect -273 1273 -257 1307
rect -223 1273 -207 1307
rect -81 1273 -65 1307
rect -31 1273 -15 1307
rect 111 1273 127 1307
rect 161 1273 177 1307
rect 303 1273 319 1307
rect 353 1273 369 1307
rect 495 1273 511 1307
rect 545 1273 561 1307
rect 687 1273 703 1307
rect 737 1273 753 1307
rect 879 1273 895 1307
rect 929 1273 945 1307
rect 1071 1273 1087 1307
rect 1121 1273 1137 1307
rect -1041 1165 -1025 1199
rect -991 1165 -975 1199
rect -849 1165 -833 1199
rect -799 1165 -783 1199
rect -657 1165 -641 1199
rect -607 1165 -591 1199
rect -465 1165 -449 1199
rect -415 1165 -399 1199
rect -273 1165 -257 1199
rect -223 1165 -207 1199
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect 111 1165 127 1199
rect 161 1165 177 1199
rect 303 1165 319 1199
rect 353 1165 369 1199
rect 495 1165 511 1199
rect 545 1165 561 1199
rect 687 1165 703 1199
rect 737 1165 753 1199
rect 879 1165 895 1199
rect 929 1165 945 1199
rect 1071 1165 1087 1199
rect 1121 1165 1137 1199
rect -1169 1115 -1135 1131
rect -1169 723 -1135 739
rect -1073 1115 -1039 1131
rect -1073 723 -1039 739
rect -977 1115 -943 1131
rect -977 723 -943 739
rect -881 1115 -847 1131
rect -881 723 -847 739
rect -785 1115 -751 1131
rect -785 723 -751 739
rect -689 1115 -655 1131
rect -689 723 -655 739
rect -593 1115 -559 1131
rect -593 723 -559 739
rect -497 1115 -463 1131
rect -497 723 -463 739
rect -401 1115 -367 1131
rect -401 723 -367 739
rect -305 1115 -271 1131
rect -305 723 -271 739
rect -209 1115 -175 1131
rect -209 723 -175 739
rect -113 1115 -79 1131
rect -113 723 -79 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 79 1115 113 1131
rect 79 723 113 739
rect 175 1115 209 1131
rect 175 723 209 739
rect 271 1115 305 1131
rect 271 723 305 739
rect 367 1115 401 1131
rect 367 723 401 739
rect 463 1115 497 1131
rect 463 723 497 739
rect 559 1115 593 1131
rect 559 723 593 739
rect 655 1115 689 1131
rect 655 723 689 739
rect 751 1115 785 1131
rect 751 723 785 739
rect 847 1115 881 1131
rect 847 723 881 739
rect 943 1115 977 1131
rect 943 723 977 739
rect 1039 1115 1073 1131
rect 1039 723 1073 739
rect 1135 1115 1169 1131
rect 1135 723 1169 739
rect -1137 655 -1121 689
rect -1087 655 -1071 689
rect -945 655 -929 689
rect -895 655 -879 689
rect -753 655 -737 689
rect -703 655 -687 689
rect -561 655 -545 689
rect -511 655 -495 689
rect -369 655 -353 689
rect -319 655 -303 689
rect -177 655 -161 689
rect -127 655 -111 689
rect 15 655 31 689
rect 65 655 81 689
rect 207 655 223 689
rect 257 655 273 689
rect 399 655 415 689
rect 449 655 465 689
rect 591 655 607 689
rect 641 655 657 689
rect 783 655 799 689
rect 833 655 849 689
rect 975 655 991 689
rect 1025 655 1041 689
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -945 547 -929 581
rect -895 547 -879 581
rect -753 547 -737 581
rect -703 547 -687 581
rect -561 547 -545 581
rect -511 547 -495 581
rect -369 547 -353 581
rect -319 547 -303 581
rect -177 547 -161 581
rect -127 547 -111 581
rect 15 547 31 581
rect 65 547 81 581
rect 207 547 223 581
rect 257 547 273 581
rect 399 547 415 581
rect 449 547 465 581
rect 591 547 607 581
rect 641 547 657 581
rect 783 547 799 581
rect 833 547 849 581
rect 975 547 991 581
rect 1025 547 1041 581
rect -1169 497 -1135 513
rect -1169 105 -1135 121
rect -1073 497 -1039 513
rect -1073 105 -1039 121
rect -977 497 -943 513
rect -977 105 -943 121
rect -881 497 -847 513
rect -881 105 -847 121
rect -785 497 -751 513
rect -785 105 -751 121
rect -689 497 -655 513
rect -689 105 -655 121
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect 655 497 689 513
rect 655 105 689 121
rect 751 497 785 513
rect 751 105 785 121
rect 847 497 881 513
rect 847 105 881 121
rect 943 497 977 513
rect 943 105 977 121
rect 1039 497 1073 513
rect 1039 105 1073 121
rect 1135 497 1169 513
rect 1135 105 1169 121
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect -1169 -121 -1135 -105
rect -1169 -513 -1135 -497
rect -1073 -121 -1039 -105
rect -1073 -513 -1039 -497
rect -977 -121 -943 -105
rect -977 -513 -943 -497
rect -881 -121 -847 -105
rect -881 -513 -847 -497
rect -785 -121 -751 -105
rect -785 -513 -751 -497
rect -689 -121 -655 -105
rect -689 -513 -655 -497
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect 655 -121 689 -105
rect 655 -513 689 -497
rect 751 -121 785 -105
rect 751 -513 785 -497
rect 847 -121 881 -105
rect 847 -513 881 -497
rect 943 -121 977 -105
rect 943 -513 977 -497
rect 1039 -121 1073 -105
rect 1039 -513 1073 -497
rect 1135 -121 1169 -105
rect 1135 -513 1169 -497
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect -1137 -689 -1121 -655
rect -1087 -689 -1071 -655
rect -945 -689 -929 -655
rect -895 -689 -879 -655
rect -753 -689 -737 -655
rect -703 -689 -687 -655
rect -561 -689 -545 -655
rect -511 -689 -495 -655
rect -369 -689 -353 -655
rect -319 -689 -303 -655
rect -177 -689 -161 -655
rect -127 -689 -111 -655
rect 15 -689 31 -655
rect 65 -689 81 -655
rect 207 -689 223 -655
rect 257 -689 273 -655
rect 399 -689 415 -655
rect 449 -689 465 -655
rect 591 -689 607 -655
rect 641 -689 657 -655
rect 783 -689 799 -655
rect 833 -689 849 -655
rect 975 -689 991 -655
rect 1025 -689 1041 -655
rect -1169 -739 -1135 -723
rect -1169 -1131 -1135 -1115
rect -1073 -739 -1039 -723
rect -1073 -1131 -1039 -1115
rect -977 -739 -943 -723
rect -977 -1131 -943 -1115
rect -881 -739 -847 -723
rect -881 -1131 -847 -1115
rect -785 -739 -751 -723
rect -785 -1131 -751 -1115
rect -689 -739 -655 -723
rect -689 -1131 -655 -1115
rect -593 -739 -559 -723
rect -593 -1131 -559 -1115
rect -497 -739 -463 -723
rect -497 -1131 -463 -1115
rect -401 -739 -367 -723
rect -401 -1131 -367 -1115
rect -305 -739 -271 -723
rect -305 -1131 -271 -1115
rect -209 -739 -175 -723
rect -209 -1131 -175 -1115
rect -113 -739 -79 -723
rect -113 -1131 -79 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 79 -739 113 -723
rect 79 -1131 113 -1115
rect 175 -739 209 -723
rect 175 -1131 209 -1115
rect 271 -739 305 -723
rect 271 -1131 305 -1115
rect 367 -739 401 -723
rect 367 -1131 401 -1115
rect 463 -739 497 -723
rect 463 -1131 497 -1115
rect 559 -739 593 -723
rect 559 -1131 593 -1115
rect 655 -739 689 -723
rect 655 -1131 689 -1115
rect 751 -739 785 -723
rect 751 -1131 785 -1115
rect 847 -739 881 -723
rect 847 -1131 881 -1115
rect 943 -739 977 -723
rect 943 -1131 977 -1115
rect 1039 -739 1073 -723
rect 1039 -1131 1073 -1115
rect 1135 -739 1169 -723
rect 1135 -1131 1169 -1115
rect -1041 -1199 -1025 -1165
rect -991 -1199 -975 -1165
rect -849 -1199 -833 -1165
rect -799 -1199 -783 -1165
rect -657 -1199 -641 -1165
rect -607 -1199 -591 -1165
rect -465 -1199 -449 -1165
rect -415 -1199 -399 -1165
rect -273 -1199 -257 -1165
rect -223 -1199 -207 -1165
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect 111 -1199 127 -1165
rect 161 -1199 177 -1165
rect 303 -1199 319 -1165
rect 353 -1199 369 -1165
rect 495 -1199 511 -1165
rect 545 -1199 561 -1165
rect 687 -1199 703 -1165
rect 737 -1199 753 -1165
rect 879 -1199 895 -1165
rect 929 -1199 945 -1165
rect 1071 -1199 1087 -1165
rect 1121 -1199 1137 -1165
rect -1041 -1307 -1025 -1273
rect -991 -1307 -975 -1273
rect -849 -1307 -833 -1273
rect -799 -1307 -783 -1273
rect -657 -1307 -641 -1273
rect -607 -1307 -591 -1273
rect -465 -1307 -449 -1273
rect -415 -1307 -399 -1273
rect -273 -1307 -257 -1273
rect -223 -1307 -207 -1273
rect -81 -1307 -65 -1273
rect -31 -1307 -15 -1273
rect 111 -1307 127 -1273
rect 161 -1307 177 -1273
rect 303 -1307 319 -1273
rect 353 -1307 369 -1273
rect 495 -1307 511 -1273
rect 545 -1307 561 -1273
rect 687 -1307 703 -1273
rect 737 -1307 753 -1273
rect 879 -1307 895 -1273
rect 929 -1307 945 -1273
rect 1071 -1307 1087 -1273
rect 1121 -1307 1137 -1273
rect -1169 -1357 -1135 -1341
rect -1169 -1749 -1135 -1733
rect -1073 -1357 -1039 -1341
rect -1073 -1749 -1039 -1733
rect -977 -1357 -943 -1341
rect -977 -1749 -943 -1733
rect -881 -1357 -847 -1341
rect -881 -1749 -847 -1733
rect -785 -1357 -751 -1341
rect -785 -1749 -751 -1733
rect -689 -1357 -655 -1341
rect -689 -1749 -655 -1733
rect -593 -1357 -559 -1341
rect -593 -1749 -559 -1733
rect -497 -1357 -463 -1341
rect -497 -1749 -463 -1733
rect -401 -1357 -367 -1341
rect -401 -1749 -367 -1733
rect -305 -1357 -271 -1341
rect -305 -1749 -271 -1733
rect -209 -1357 -175 -1341
rect -209 -1749 -175 -1733
rect -113 -1357 -79 -1341
rect -113 -1749 -79 -1733
rect -17 -1357 17 -1341
rect -17 -1749 17 -1733
rect 79 -1357 113 -1341
rect 79 -1749 113 -1733
rect 175 -1357 209 -1341
rect 175 -1749 209 -1733
rect 271 -1357 305 -1341
rect 271 -1749 305 -1733
rect 367 -1357 401 -1341
rect 367 -1749 401 -1733
rect 463 -1357 497 -1341
rect 463 -1749 497 -1733
rect 559 -1357 593 -1341
rect 559 -1749 593 -1733
rect 655 -1357 689 -1341
rect 655 -1749 689 -1733
rect 751 -1357 785 -1341
rect 751 -1749 785 -1733
rect 847 -1357 881 -1341
rect 847 -1749 881 -1733
rect 943 -1357 977 -1341
rect 943 -1749 977 -1733
rect 1039 -1357 1073 -1341
rect 1039 -1749 1073 -1733
rect 1135 -1357 1169 -1341
rect 1135 -1749 1169 -1733
rect -1137 -1817 -1121 -1783
rect -1087 -1817 -1071 -1783
rect -945 -1817 -929 -1783
rect -895 -1817 -879 -1783
rect -753 -1817 -737 -1783
rect -703 -1817 -687 -1783
rect -561 -1817 -545 -1783
rect -511 -1817 -495 -1783
rect -369 -1817 -353 -1783
rect -319 -1817 -303 -1783
rect -177 -1817 -161 -1783
rect -127 -1817 -111 -1783
rect 15 -1817 31 -1783
rect 65 -1817 81 -1783
rect 207 -1817 223 -1783
rect 257 -1817 273 -1783
rect 399 -1817 415 -1783
rect 449 -1817 465 -1783
rect 591 -1817 607 -1783
rect 641 -1817 657 -1783
rect 783 -1817 799 -1783
rect 833 -1817 849 -1783
rect 975 -1817 991 -1783
rect 1025 -1817 1041 -1783
rect -1137 -1925 -1121 -1891
rect -1087 -1925 -1071 -1891
rect -945 -1925 -929 -1891
rect -895 -1925 -879 -1891
rect -753 -1925 -737 -1891
rect -703 -1925 -687 -1891
rect -561 -1925 -545 -1891
rect -511 -1925 -495 -1891
rect -369 -1925 -353 -1891
rect -319 -1925 -303 -1891
rect -177 -1925 -161 -1891
rect -127 -1925 -111 -1891
rect 15 -1925 31 -1891
rect 65 -1925 81 -1891
rect 207 -1925 223 -1891
rect 257 -1925 273 -1891
rect 399 -1925 415 -1891
rect 449 -1925 465 -1891
rect 591 -1925 607 -1891
rect 641 -1925 657 -1891
rect 783 -1925 799 -1891
rect 833 -1925 849 -1891
rect 975 -1925 991 -1891
rect 1025 -1925 1041 -1891
rect -1169 -1975 -1135 -1959
rect -1169 -2367 -1135 -2351
rect -1073 -1975 -1039 -1959
rect -1073 -2367 -1039 -2351
rect -977 -1975 -943 -1959
rect -977 -2367 -943 -2351
rect -881 -1975 -847 -1959
rect -881 -2367 -847 -2351
rect -785 -1975 -751 -1959
rect -785 -2367 -751 -2351
rect -689 -1975 -655 -1959
rect -689 -2367 -655 -2351
rect -593 -1975 -559 -1959
rect -593 -2367 -559 -2351
rect -497 -1975 -463 -1959
rect -497 -2367 -463 -2351
rect -401 -1975 -367 -1959
rect -401 -2367 -367 -2351
rect -305 -1975 -271 -1959
rect -305 -2367 -271 -2351
rect -209 -1975 -175 -1959
rect -209 -2367 -175 -2351
rect -113 -1975 -79 -1959
rect -113 -2367 -79 -2351
rect -17 -1975 17 -1959
rect -17 -2367 17 -2351
rect 79 -1975 113 -1959
rect 79 -2367 113 -2351
rect 175 -1975 209 -1959
rect 175 -2367 209 -2351
rect 271 -1975 305 -1959
rect 271 -2367 305 -2351
rect 367 -1975 401 -1959
rect 367 -2367 401 -2351
rect 463 -1975 497 -1959
rect 463 -2367 497 -2351
rect 559 -1975 593 -1959
rect 559 -2367 593 -2351
rect 655 -1975 689 -1959
rect 655 -2367 689 -2351
rect 751 -1975 785 -1959
rect 751 -2367 785 -2351
rect 847 -1975 881 -1959
rect 847 -2367 881 -2351
rect 943 -1975 977 -1959
rect 943 -2367 977 -2351
rect 1039 -1975 1073 -1959
rect 1039 -2367 1073 -2351
rect 1135 -1975 1169 -1959
rect 1135 -2367 1169 -2351
rect -1041 -2435 -1025 -2401
rect -991 -2435 -975 -2401
rect -849 -2435 -833 -2401
rect -799 -2435 -783 -2401
rect -657 -2435 -641 -2401
rect -607 -2435 -591 -2401
rect -465 -2435 -449 -2401
rect -415 -2435 -399 -2401
rect -273 -2435 -257 -2401
rect -223 -2435 -207 -2401
rect -81 -2435 -65 -2401
rect -31 -2435 -15 -2401
rect 111 -2435 127 -2401
rect 161 -2435 177 -2401
rect 303 -2435 319 -2401
rect 353 -2435 369 -2401
rect 495 -2435 511 -2401
rect 545 -2435 561 -2401
rect 687 -2435 703 -2401
rect 737 -2435 753 -2401
rect 879 -2435 895 -2401
rect 929 -2435 945 -2401
rect 1071 -2435 1087 -2401
rect 1121 -2435 1137 -2401
rect -1041 -2543 -1025 -2509
rect -991 -2543 -975 -2509
rect -849 -2543 -833 -2509
rect -799 -2543 -783 -2509
rect -657 -2543 -641 -2509
rect -607 -2543 -591 -2509
rect -465 -2543 -449 -2509
rect -415 -2543 -399 -2509
rect -273 -2543 -257 -2509
rect -223 -2543 -207 -2509
rect -81 -2543 -65 -2509
rect -31 -2543 -15 -2509
rect 111 -2543 127 -2509
rect 161 -2543 177 -2509
rect 303 -2543 319 -2509
rect 353 -2543 369 -2509
rect 495 -2543 511 -2509
rect 545 -2543 561 -2509
rect 687 -2543 703 -2509
rect 737 -2543 753 -2509
rect 879 -2543 895 -2509
rect 929 -2543 945 -2509
rect 1071 -2543 1087 -2509
rect 1121 -2543 1137 -2509
rect -1169 -2593 -1135 -2577
rect -1169 -2985 -1135 -2969
rect -1073 -2593 -1039 -2577
rect -1073 -2985 -1039 -2969
rect -977 -2593 -943 -2577
rect -977 -2985 -943 -2969
rect -881 -2593 -847 -2577
rect -881 -2985 -847 -2969
rect -785 -2593 -751 -2577
rect -785 -2985 -751 -2969
rect -689 -2593 -655 -2577
rect -689 -2985 -655 -2969
rect -593 -2593 -559 -2577
rect -593 -2985 -559 -2969
rect -497 -2593 -463 -2577
rect -497 -2985 -463 -2969
rect -401 -2593 -367 -2577
rect -401 -2985 -367 -2969
rect -305 -2593 -271 -2577
rect -305 -2985 -271 -2969
rect -209 -2593 -175 -2577
rect -209 -2985 -175 -2969
rect -113 -2593 -79 -2577
rect -113 -2985 -79 -2969
rect -17 -2593 17 -2577
rect -17 -2985 17 -2969
rect 79 -2593 113 -2577
rect 79 -2985 113 -2969
rect 175 -2593 209 -2577
rect 175 -2985 209 -2969
rect 271 -2593 305 -2577
rect 271 -2985 305 -2969
rect 367 -2593 401 -2577
rect 367 -2985 401 -2969
rect 463 -2593 497 -2577
rect 463 -2985 497 -2969
rect 559 -2593 593 -2577
rect 559 -2985 593 -2969
rect 655 -2593 689 -2577
rect 655 -2985 689 -2969
rect 751 -2593 785 -2577
rect 751 -2985 785 -2969
rect 847 -2593 881 -2577
rect 847 -2985 881 -2969
rect 943 -2593 977 -2577
rect 943 -2985 977 -2969
rect 1039 -2593 1073 -2577
rect 1039 -2985 1073 -2969
rect 1135 -2593 1169 -2577
rect 1135 -2985 1169 -2969
rect -1137 -3053 -1121 -3019
rect -1087 -3053 -1071 -3019
rect -945 -3053 -929 -3019
rect -895 -3053 -879 -3019
rect -753 -3053 -737 -3019
rect -703 -3053 -687 -3019
rect -561 -3053 -545 -3019
rect -511 -3053 -495 -3019
rect -369 -3053 -353 -3019
rect -319 -3053 -303 -3019
rect -177 -3053 -161 -3019
rect -127 -3053 -111 -3019
rect 15 -3053 31 -3019
rect 65 -3053 81 -3019
rect 207 -3053 223 -3019
rect 257 -3053 273 -3019
rect 399 -3053 415 -3019
rect 449 -3053 465 -3019
rect 591 -3053 607 -3019
rect 641 -3053 657 -3019
rect 783 -3053 799 -3019
rect 833 -3053 849 -3019
rect 975 -3053 991 -3019
rect 1025 -3053 1041 -3019
rect -1283 -3121 -1249 -3059
rect 1249 -3121 1283 -3059
rect -1283 -3155 -1187 -3121
rect 1187 -3155 1283 -3121
<< viali >>
rect -1121 3019 -1087 3053
rect -929 3019 -895 3053
rect -737 3019 -703 3053
rect -545 3019 -511 3053
rect -353 3019 -319 3053
rect -161 3019 -127 3053
rect 31 3019 65 3053
rect 223 3019 257 3053
rect 415 3019 449 3053
rect 607 3019 641 3053
rect 799 3019 833 3053
rect 991 3019 1025 3053
rect -1169 2593 -1135 2969
rect -1073 2593 -1039 2969
rect -977 2593 -943 2969
rect -881 2593 -847 2969
rect -785 2593 -751 2969
rect -689 2593 -655 2969
rect -593 2593 -559 2969
rect -497 2593 -463 2969
rect -401 2593 -367 2969
rect -305 2593 -271 2969
rect -209 2593 -175 2969
rect -113 2593 -79 2969
rect -17 2593 17 2969
rect 79 2593 113 2969
rect 175 2593 209 2969
rect 271 2593 305 2969
rect 367 2593 401 2969
rect 463 2593 497 2969
rect 559 2593 593 2969
rect 655 2593 689 2969
rect 751 2593 785 2969
rect 847 2593 881 2969
rect 943 2593 977 2969
rect 1039 2593 1073 2969
rect 1135 2593 1169 2969
rect -1025 2509 -991 2543
rect -833 2509 -799 2543
rect -641 2509 -607 2543
rect -449 2509 -415 2543
rect -257 2509 -223 2543
rect -65 2509 -31 2543
rect 127 2509 161 2543
rect 319 2509 353 2543
rect 511 2509 545 2543
rect 703 2509 737 2543
rect 895 2509 929 2543
rect 1087 2509 1121 2543
rect -1025 2401 -991 2435
rect -833 2401 -799 2435
rect -641 2401 -607 2435
rect -449 2401 -415 2435
rect -257 2401 -223 2435
rect -65 2401 -31 2435
rect 127 2401 161 2435
rect 319 2401 353 2435
rect 511 2401 545 2435
rect 703 2401 737 2435
rect 895 2401 929 2435
rect 1087 2401 1121 2435
rect -1169 1975 -1135 2351
rect -1073 1975 -1039 2351
rect -977 1975 -943 2351
rect -881 1975 -847 2351
rect -785 1975 -751 2351
rect -689 1975 -655 2351
rect -593 1975 -559 2351
rect -497 1975 -463 2351
rect -401 1975 -367 2351
rect -305 1975 -271 2351
rect -209 1975 -175 2351
rect -113 1975 -79 2351
rect -17 1975 17 2351
rect 79 1975 113 2351
rect 175 1975 209 2351
rect 271 1975 305 2351
rect 367 1975 401 2351
rect 463 1975 497 2351
rect 559 1975 593 2351
rect 655 1975 689 2351
rect 751 1975 785 2351
rect 847 1975 881 2351
rect 943 1975 977 2351
rect 1039 1975 1073 2351
rect 1135 1975 1169 2351
rect -1121 1891 -1087 1925
rect -929 1891 -895 1925
rect -737 1891 -703 1925
rect -545 1891 -511 1925
rect -353 1891 -319 1925
rect -161 1891 -127 1925
rect 31 1891 65 1925
rect 223 1891 257 1925
rect 415 1891 449 1925
rect 607 1891 641 1925
rect 799 1891 833 1925
rect 991 1891 1025 1925
rect -1121 1783 -1087 1817
rect -929 1783 -895 1817
rect -737 1783 -703 1817
rect -545 1783 -511 1817
rect -353 1783 -319 1817
rect -161 1783 -127 1817
rect 31 1783 65 1817
rect 223 1783 257 1817
rect 415 1783 449 1817
rect 607 1783 641 1817
rect 799 1783 833 1817
rect 991 1783 1025 1817
rect -1169 1357 -1135 1733
rect -1073 1357 -1039 1733
rect -977 1357 -943 1733
rect -881 1357 -847 1733
rect -785 1357 -751 1733
rect -689 1357 -655 1733
rect -593 1357 -559 1733
rect -497 1357 -463 1733
rect -401 1357 -367 1733
rect -305 1357 -271 1733
rect -209 1357 -175 1733
rect -113 1357 -79 1733
rect -17 1357 17 1733
rect 79 1357 113 1733
rect 175 1357 209 1733
rect 271 1357 305 1733
rect 367 1357 401 1733
rect 463 1357 497 1733
rect 559 1357 593 1733
rect 655 1357 689 1733
rect 751 1357 785 1733
rect 847 1357 881 1733
rect 943 1357 977 1733
rect 1039 1357 1073 1733
rect 1135 1357 1169 1733
rect -1025 1273 -991 1307
rect -833 1273 -799 1307
rect -641 1273 -607 1307
rect -449 1273 -415 1307
rect -257 1273 -223 1307
rect -65 1273 -31 1307
rect 127 1273 161 1307
rect 319 1273 353 1307
rect 511 1273 545 1307
rect 703 1273 737 1307
rect 895 1273 929 1307
rect 1087 1273 1121 1307
rect -1025 1165 -991 1199
rect -833 1165 -799 1199
rect -641 1165 -607 1199
rect -449 1165 -415 1199
rect -257 1165 -223 1199
rect -65 1165 -31 1199
rect 127 1165 161 1199
rect 319 1165 353 1199
rect 511 1165 545 1199
rect 703 1165 737 1199
rect 895 1165 929 1199
rect 1087 1165 1121 1199
rect -1169 739 -1135 1115
rect -1073 739 -1039 1115
rect -977 739 -943 1115
rect -881 739 -847 1115
rect -785 739 -751 1115
rect -689 739 -655 1115
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect 655 739 689 1115
rect 751 739 785 1115
rect 847 739 881 1115
rect 943 739 977 1115
rect 1039 739 1073 1115
rect 1135 739 1169 1115
rect -1121 655 -1087 689
rect -929 655 -895 689
rect -737 655 -703 689
rect -545 655 -511 689
rect -353 655 -319 689
rect -161 655 -127 689
rect 31 655 65 689
rect 223 655 257 689
rect 415 655 449 689
rect 607 655 641 689
rect 799 655 833 689
rect 991 655 1025 689
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect -1121 -689 -1087 -655
rect -929 -689 -895 -655
rect -737 -689 -703 -655
rect -545 -689 -511 -655
rect -353 -689 -319 -655
rect -161 -689 -127 -655
rect 31 -689 65 -655
rect 223 -689 257 -655
rect 415 -689 449 -655
rect 607 -689 641 -655
rect 799 -689 833 -655
rect 991 -689 1025 -655
rect -1169 -1115 -1135 -739
rect -1073 -1115 -1039 -739
rect -977 -1115 -943 -739
rect -881 -1115 -847 -739
rect -785 -1115 -751 -739
rect -689 -1115 -655 -739
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect 655 -1115 689 -739
rect 751 -1115 785 -739
rect 847 -1115 881 -739
rect 943 -1115 977 -739
rect 1039 -1115 1073 -739
rect 1135 -1115 1169 -739
rect -1025 -1199 -991 -1165
rect -833 -1199 -799 -1165
rect -641 -1199 -607 -1165
rect -449 -1199 -415 -1165
rect -257 -1199 -223 -1165
rect -65 -1199 -31 -1165
rect 127 -1199 161 -1165
rect 319 -1199 353 -1165
rect 511 -1199 545 -1165
rect 703 -1199 737 -1165
rect 895 -1199 929 -1165
rect 1087 -1199 1121 -1165
rect -1025 -1307 -991 -1273
rect -833 -1307 -799 -1273
rect -641 -1307 -607 -1273
rect -449 -1307 -415 -1273
rect -257 -1307 -223 -1273
rect -65 -1307 -31 -1273
rect 127 -1307 161 -1273
rect 319 -1307 353 -1273
rect 511 -1307 545 -1273
rect 703 -1307 737 -1273
rect 895 -1307 929 -1273
rect 1087 -1307 1121 -1273
rect -1169 -1733 -1135 -1357
rect -1073 -1733 -1039 -1357
rect -977 -1733 -943 -1357
rect -881 -1733 -847 -1357
rect -785 -1733 -751 -1357
rect -689 -1733 -655 -1357
rect -593 -1733 -559 -1357
rect -497 -1733 -463 -1357
rect -401 -1733 -367 -1357
rect -305 -1733 -271 -1357
rect -209 -1733 -175 -1357
rect -113 -1733 -79 -1357
rect -17 -1733 17 -1357
rect 79 -1733 113 -1357
rect 175 -1733 209 -1357
rect 271 -1733 305 -1357
rect 367 -1733 401 -1357
rect 463 -1733 497 -1357
rect 559 -1733 593 -1357
rect 655 -1733 689 -1357
rect 751 -1733 785 -1357
rect 847 -1733 881 -1357
rect 943 -1733 977 -1357
rect 1039 -1733 1073 -1357
rect 1135 -1733 1169 -1357
rect -1121 -1817 -1087 -1783
rect -929 -1817 -895 -1783
rect -737 -1817 -703 -1783
rect -545 -1817 -511 -1783
rect -353 -1817 -319 -1783
rect -161 -1817 -127 -1783
rect 31 -1817 65 -1783
rect 223 -1817 257 -1783
rect 415 -1817 449 -1783
rect 607 -1817 641 -1783
rect 799 -1817 833 -1783
rect 991 -1817 1025 -1783
rect -1121 -1925 -1087 -1891
rect -929 -1925 -895 -1891
rect -737 -1925 -703 -1891
rect -545 -1925 -511 -1891
rect -353 -1925 -319 -1891
rect -161 -1925 -127 -1891
rect 31 -1925 65 -1891
rect 223 -1925 257 -1891
rect 415 -1925 449 -1891
rect 607 -1925 641 -1891
rect 799 -1925 833 -1891
rect 991 -1925 1025 -1891
rect -1169 -2351 -1135 -1975
rect -1073 -2351 -1039 -1975
rect -977 -2351 -943 -1975
rect -881 -2351 -847 -1975
rect -785 -2351 -751 -1975
rect -689 -2351 -655 -1975
rect -593 -2351 -559 -1975
rect -497 -2351 -463 -1975
rect -401 -2351 -367 -1975
rect -305 -2351 -271 -1975
rect -209 -2351 -175 -1975
rect -113 -2351 -79 -1975
rect -17 -2351 17 -1975
rect 79 -2351 113 -1975
rect 175 -2351 209 -1975
rect 271 -2351 305 -1975
rect 367 -2351 401 -1975
rect 463 -2351 497 -1975
rect 559 -2351 593 -1975
rect 655 -2351 689 -1975
rect 751 -2351 785 -1975
rect 847 -2351 881 -1975
rect 943 -2351 977 -1975
rect 1039 -2351 1073 -1975
rect 1135 -2351 1169 -1975
rect -1025 -2435 -991 -2401
rect -833 -2435 -799 -2401
rect -641 -2435 -607 -2401
rect -449 -2435 -415 -2401
rect -257 -2435 -223 -2401
rect -65 -2435 -31 -2401
rect 127 -2435 161 -2401
rect 319 -2435 353 -2401
rect 511 -2435 545 -2401
rect 703 -2435 737 -2401
rect 895 -2435 929 -2401
rect 1087 -2435 1121 -2401
rect -1025 -2543 -991 -2509
rect -833 -2543 -799 -2509
rect -641 -2543 -607 -2509
rect -449 -2543 -415 -2509
rect -257 -2543 -223 -2509
rect -65 -2543 -31 -2509
rect 127 -2543 161 -2509
rect 319 -2543 353 -2509
rect 511 -2543 545 -2509
rect 703 -2543 737 -2509
rect 895 -2543 929 -2509
rect 1087 -2543 1121 -2509
rect -1169 -2969 -1135 -2593
rect -1073 -2969 -1039 -2593
rect -977 -2969 -943 -2593
rect -881 -2969 -847 -2593
rect -785 -2969 -751 -2593
rect -689 -2969 -655 -2593
rect -593 -2969 -559 -2593
rect -497 -2969 -463 -2593
rect -401 -2969 -367 -2593
rect -305 -2969 -271 -2593
rect -209 -2969 -175 -2593
rect -113 -2969 -79 -2593
rect -17 -2969 17 -2593
rect 79 -2969 113 -2593
rect 175 -2969 209 -2593
rect 271 -2969 305 -2593
rect 367 -2969 401 -2593
rect 463 -2969 497 -2593
rect 559 -2969 593 -2593
rect 655 -2969 689 -2593
rect 751 -2969 785 -2593
rect 847 -2969 881 -2593
rect 943 -2969 977 -2593
rect 1039 -2969 1073 -2593
rect 1135 -2969 1169 -2593
rect -1121 -3053 -1087 -3019
rect -929 -3053 -895 -3019
rect -737 -3053 -703 -3019
rect -545 -3053 -511 -3019
rect -353 -3053 -319 -3019
rect -161 -3053 -127 -3019
rect 31 -3053 65 -3019
rect 223 -3053 257 -3019
rect 415 -3053 449 -3019
rect 607 -3053 641 -3019
rect 799 -3053 833 -3019
rect 991 -3053 1025 -3019
<< metal1 >>
rect -1133 3053 -1075 3059
rect -1133 3019 -1121 3053
rect -1087 3019 -1075 3053
rect -1133 3013 -1075 3019
rect -941 3053 -883 3059
rect -941 3019 -929 3053
rect -895 3019 -883 3053
rect -941 3013 -883 3019
rect -749 3053 -691 3059
rect -749 3019 -737 3053
rect -703 3019 -691 3053
rect -749 3013 -691 3019
rect -557 3053 -499 3059
rect -557 3019 -545 3053
rect -511 3019 -499 3053
rect -557 3013 -499 3019
rect -365 3053 -307 3059
rect -365 3019 -353 3053
rect -319 3019 -307 3053
rect -365 3013 -307 3019
rect -173 3053 -115 3059
rect -173 3019 -161 3053
rect -127 3019 -115 3053
rect -173 3013 -115 3019
rect 19 3053 77 3059
rect 19 3019 31 3053
rect 65 3019 77 3053
rect 19 3013 77 3019
rect 211 3053 269 3059
rect 211 3019 223 3053
rect 257 3019 269 3053
rect 211 3013 269 3019
rect 403 3053 461 3059
rect 403 3019 415 3053
rect 449 3019 461 3053
rect 403 3013 461 3019
rect 595 3053 653 3059
rect 595 3019 607 3053
rect 641 3019 653 3053
rect 595 3013 653 3019
rect 787 3053 845 3059
rect 787 3019 799 3053
rect 833 3019 845 3053
rect 787 3013 845 3019
rect 979 3053 1037 3059
rect 979 3019 991 3053
rect 1025 3019 1037 3053
rect 979 3013 1037 3019
rect -1175 2969 -1129 2981
rect -1175 2593 -1169 2969
rect -1135 2593 -1129 2969
rect -1175 2581 -1129 2593
rect -1079 2969 -1033 2981
rect -1079 2593 -1073 2969
rect -1039 2593 -1033 2969
rect -1079 2581 -1033 2593
rect -983 2969 -937 2981
rect -983 2593 -977 2969
rect -943 2593 -937 2969
rect -983 2581 -937 2593
rect -887 2969 -841 2981
rect -887 2593 -881 2969
rect -847 2593 -841 2969
rect -887 2581 -841 2593
rect -791 2969 -745 2981
rect -791 2593 -785 2969
rect -751 2593 -745 2969
rect -791 2581 -745 2593
rect -695 2969 -649 2981
rect -695 2593 -689 2969
rect -655 2593 -649 2969
rect -695 2581 -649 2593
rect -599 2969 -553 2981
rect -599 2593 -593 2969
rect -559 2593 -553 2969
rect -599 2581 -553 2593
rect -503 2969 -457 2981
rect -503 2593 -497 2969
rect -463 2593 -457 2969
rect -503 2581 -457 2593
rect -407 2969 -361 2981
rect -407 2593 -401 2969
rect -367 2593 -361 2969
rect -407 2581 -361 2593
rect -311 2969 -265 2981
rect -311 2593 -305 2969
rect -271 2593 -265 2969
rect -311 2581 -265 2593
rect -215 2969 -169 2981
rect -215 2593 -209 2969
rect -175 2593 -169 2969
rect -215 2581 -169 2593
rect -119 2969 -73 2981
rect -119 2593 -113 2969
rect -79 2593 -73 2969
rect -119 2581 -73 2593
rect -23 2969 23 2981
rect -23 2593 -17 2969
rect 17 2593 23 2969
rect -23 2581 23 2593
rect 73 2969 119 2981
rect 73 2593 79 2969
rect 113 2593 119 2969
rect 73 2581 119 2593
rect 169 2969 215 2981
rect 169 2593 175 2969
rect 209 2593 215 2969
rect 169 2581 215 2593
rect 265 2969 311 2981
rect 265 2593 271 2969
rect 305 2593 311 2969
rect 265 2581 311 2593
rect 361 2969 407 2981
rect 361 2593 367 2969
rect 401 2593 407 2969
rect 361 2581 407 2593
rect 457 2969 503 2981
rect 457 2593 463 2969
rect 497 2593 503 2969
rect 457 2581 503 2593
rect 553 2969 599 2981
rect 553 2593 559 2969
rect 593 2593 599 2969
rect 553 2581 599 2593
rect 649 2969 695 2981
rect 649 2593 655 2969
rect 689 2593 695 2969
rect 649 2581 695 2593
rect 745 2969 791 2981
rect 745 2593 751 2969
rect 785 2593 791 2969
rect 745 2581 791 2593
rect 841 2969 887 2981
rect 841 2593 847 2969
rect 881 2593 887 2969
rect 841 2581 887 2593
rect 937 2969 983 2981
rect 937 2593 943 2969
rect 977 2593 983 2969
rect 937 2581 983 2593
rect 1033 2969 1079 2981
rect 1033 2593 1039 2969
rect 1073 2593 1079 2969
rect 1033 2581 1079 2593
rect 1129 2969 1175 2981
rect 1129 2593 1135 2969
rect 1169 2593 1175 2969
rect 1129 2581 1175 2593
rect -1037 2543 -979 2549
rect -1037 2509 -1025 2543
rect -991 2509 -979 2543
rect -1037 2503 -979 2509
rect -845 2543 -787 2549
rect -845 2509 -833 2543
rect -799 2509 -787 2543
rect -845 2503 -787 2509
rect -653 2543 -595 2549
rect -653 2509 -641 2543
rect -607 2509 -595 2543
rect -653 2503 -595 2509
rect -461 2543 -403 2549
rect -461 2509 -449 2543
rect -415 2509 -403 2543
rect -461 2503 -403 2509
rect -269 2543 -211 2549
rect -269 2509 -257 2543
rect -223 2509 -211 2543
rect -269 2503 -211 2509
rect -77 2543 -19 2549
rect -77 2509 -65 2543
rect -31 2509 -19 2543
rect -77 2503 -19 2509
rect 115 2543 173 2549
rect 115 2509 127 2543
rect 161 2509 173 2543
rect 115 2503 173 2509
rect 307 2543 365 2549
rect 307 2509 319 2543
rect 353 2509 365 2543
rect 307 2503 365 2509
rect 499 2543 557 2549
rect 499 2509 511 2543
rect 545 2509 557 2543
rect 499 2503 557 2509
rect 691 2543 749 2549
rect 691 2509 703 2543
rect 737 2509 749 2543
rect 691 2503 749 2509
rect 883 2543 941 2549
rect 883 2509 895 2543
rect 929 2509 941 2543
rect 883 2503 941 2509
rect 1075 2543 1133 2549
rect 1075 2509 1087 2543
rect 1121 2509 1133 2543
rect 1075 2503 1133 2509
rect -1037 2435 -979 2441
rect -1037 2401 -1025 2435
rect -991 2401 -979 2435
rect -1037 2395 -979 2401
rect -845 2435 -787 2441
rect -845 2401 -833 2435
rect -799 2401 -787 2435
rect -845 2395 -787 2401
rect -653 2435 -595 2441
rect -653 2401 -641 2435
rect -607 2401 -595 2435
rect -653 2395 -595 2401
rect -461 2435 -403 2441
rect -461 2401 -449 2435
rect -415 2401 -403 2435
rect -461 2395 -403 2401
rect -269 2435 -211 2441
rect -269 2401 -257 2435
rect -223 2401 -211 2435
rect -269 2395 -211 2401
rect -77 2435 -19 2441
rect -77 2401 -65 2435
rect -31 2401 -19 2435
rect -77 2395 -19 2401
rect 115 2435 173 2441
rect 115 2401 127 2435
rect 161 2401 173 2435
rect 115 2395 173 2401
rect 307 2435 365 2441
rect 307 2401 319 2435
rect 353 2401 365 2435
rect 307 2395 365 2401
rect 499 2435 557 2441
rect 499 2401 511 2435
rect 545 2401 557 2435
rect 499 2395 557 2401
rect 691 2435 749 2441
rect 691 2401 703 2435
rect 737 2401 749 2435
rect 691 2395 749 2401
rect 883 2435 941 2441
rect 883 2401 895 2435
rect 929 2401 941 2435
rect 883 2395 941 2401
rect 1075 2435 1133 2441
rect 1075 2401 1087 2435
rect 1121 2401 1133 2435
rect 1075 2395 1133 2401
rect -1175 2351 -1129 2363
rect -1175 1975 -1169 2351
rect -1135 1975 -1129 2351
rect -1175 1963 -1129 1975
rect -1079 2351 -1033 2363
rect -1079 1975 -1073 2351
rect -1039 1975 -1033 2351
rect -1079 1963 -1033 1975
rect -983 2351 -937 2363
rect -983 1975 -977 2351
rect -943 1975 -937 2351
rect -983 1963 -937 1975
rect -887 2351 -841 2363
rect -887 1975 -881 2351
rect -847 1975 -841 2351
rect -887 1963 -841 1975
rect -791 2351 -745 2363
rect -791 1975 -785 2351
rect -751 1975 -745 2351
rect -791 1963 -745 1975
rect -695 2351 -649 2363
rect -695 1975 -689 2351
rect -655 1975 -649 2351
rect -695 1963 -649 1975
rect -599 2351 -553 2363
rect -599 1975 -593 2351
rect -559 1975 -553 2351
rect -599 1963 -553 1975
rect -503 2351 -457 2363
rect -503 1975 -497 2351
rect -463 1975 -457 2351
rect -503 1963 -457 1975
rect -407 2351 -361 2363
rect -407 1975 -401 2351
rect -367 1975 -361 2351
rect -407 1963 -361 1975
rect -311 2351 -265 2363
rect -311 1975 -305 2351
rect -271 1975 -265 2351
rect -311 1963 -265 1975
rect -215 2351 -169 2363
rect -215 1975 -209 2351
rect -175 1975 -169 2351
rect -215 1963 -169 1975
rect -119 2351 -73 2363
rect -119 1975 -113 2351
rect -79 1975 -73 2351
rect -119 1963 -73 1975
rect -23 2351 23 2363
rect -23 1975 -17 2351
rect 17 1975 23 2351
rect -23 1963 23 1975
rect 73 2351 119 2363
rect 73 1975 79 2351
rect 113 1975 119 2351
rect 73 1963 119 1975
rect 169 2351 215 2363
rect 169 1975 175 2351
rect 209 1975 215 2351
rect 169 1963 215 1975
rect 265 2351 311 2363
rect 265 1975 271 2351
rect 305 1975 311 2351
rect 265 1963 311 1975
rect 361 2351 407 2363
rect 361 1975 367 2351
rect 401 1975 407 2351
rect 361 1963 407 1975
rect 457 2351 503 2363
rect 457 1975 463 2351
rect 497 1975 503 2351
rect 457 1963 503 1975
rect 553 2351 599 2363
rect 553 1975 559 2351
rect 593 1975 599 2351
rect 553 1963 599 1975
rect 649 2351 695 2363
rect 649 1975 655 2351
rect 689 1975 695 2351
rect 649 1963 695 1975
rect 745 2351 791 2363
rect 745 1975 751 2351
rect 785 1975 791 2351
rect 745 1963 791 1975
rect 841 2351 887 2363
rect 841 1975 847 2351
rect 881 1975 887 2351
rect 841 1963 887 1975
rect 937 2351 983 2363
rect 937 1975 943 2351
rect 977 1975 983 2351
rect 937 1963 983 1975
rect 1033 2351 1079 2363
rect 1033 1975 1039 2351
rect 1073 1975 1079 2351
rect 1033 1963 1079 1975
rect 1129 2351 1175 2363
rect 1129 1975 1135 2351
rect 1169 1975 1175 2351
rect 1129 1963 1175 1975
rect -1133 1925 -1075 1931
rect -1133 1891 -1121 1925
rect -1087 1891 -1075 1925
rect -1133 1885 -1075 1891
rect -941 1925 -883 1931
rect -941 1891 -929 1925
rect -895 1891 -883 1925
rect -941 1885 -883 1891
rect -749 1925 -691 1931
rect -749 1891 -737 1925
rect -703 1891 -691 1925
rect -749 1885 -691 1891
rect -557 1925 -499 1931
rect -557 1891 -545 1925
rect -511 1891 -499 1925
rect -557 1885 -499 1891
rect -365 1925 -307 1931
rect -365 1891 -353 1925
rect -319 1891 -307 1925
rect -365 1885 -307 1891
rect -173 1925 -115 1931
rect -173 1891 -161 1925
rect -127 1891 -115 1925
rect -173 1885 -115 1891
rect 19 1925 77 1931
rect 19 1891 31 1925
rect 65 1891 77 1925
rect 19 1885 77 1891
rect 211 1925 269 1931
rect 211 1891 223 1925
rect 257 1891 269 1925
rect 211 1885 269 1891
rect 403 1925 461 1931
rect 403 1891 415 1925
rect 449 1891 461 1925
rect 403 1885 461 1891
rect 595 1925 653 1931
rect 595 1891 607 1925
rect 641 1891 653 1925
rect 595 1885 653 1891
rect 787 1925 845 1931
rect 787 1891 799 1925
rect 833 1891 845 1925
rect 787 1885 845 1891
rect 979 1925 1037 1931
rect 979 1891 991 1925
rect 1025 1891 1037 1925
rect 979 1885 1037 1891
rect -1133 1817 -1075 1823
rect -1133 1783 -1121 1817
rect -1087 1783 -1075 1817
rect -1133 1777 -1075 1783
rect -941 1817 -883 1823
rect -941 1783 -929 1817
rect -895 1783 -883 1817
rect -941 1777 -883 1783
rect -749 1817 -691 1823
rect -749 1783 -737 1817
rect -703 1783 -691 1817
rect -749 1777 -691 1783
rect -557 1817 -499 1823
rect -557 1783 -545 1817
rect -511 1783 -499 1817
rect -557 1777 -499 1783
rect -365 1817 -307 1823
rect -365 1783 -353 1817
rect -319 1783 -307 1817
rect -365 1777 -307 1783
rect -173 1817 -115 1823
rect -173 1783 -161 1817
rect -127 1783 -115 1817
rect -173 1777 -115 1783
rect 19 1817 77 1823
rect 19 1783 31 1817
rect 65 1783 77 1817
rect 19 1777 77 1783
rect 211 1817 269 1823
rect 211 1783 223 1817
rect 257 1783 269 1817
rect 211 1777 269 1783
rect 403 1817 461 1823
rect 403 1783 415 1817
rect 449 1783 461 1817
rect 403 1777 461 1783
rect 595 1817 653 1823
rect 595 1783 607 1817
rect 641 1783 653 1817
rect 595 1777 653 1783
rect 787 1817 845 1823
rect 787 1783 799 1817
rect 833 1783 845 1817
rect 787 1777 845 1783
rect 979 1817 1037 1823
rect 979 1783 991 1817
rect 1025 1783 1037 1817
rect 979 1777 1037 1783
rect -1175 1733 -1129 1745
rect -1175 1357 -1169 1733
rect -1135 1357 -1129 1733
rect -1175 1345 -1129 1357
rect -1079 1733 -1033 1745
rect -1079 1357 -1073 1733
rect -1039 1357 -1033 1733
rect -1079 1345 -1033 1357
rect -983 1733 -937 1745
rect -983 1357 -977 1733
rect -943 1357 -937 1733
rect -983 1345 -937 1357
rect -887 1733 -841 1745
rect -887 1357 -881 1733
rect -847 1357 -841 1733
rect -887 1345 -841 1357
rect -791 1733 -745 1745
rect -791 1357 -785 1733
rect -751 1357 -745 1733
rect -791 1345 -745 1357
rect -695 1733 -649 1745
rect -695 1357 -689 1733
rect -655 1357 -649 1733
rect -695 1345 -649 1357
rect -599 1733 -553 1745
rect -599 1357 -593 1733
rect -559 1357 -553 1733
rect -599 1345 -553 1357
rect -503 1733 -457 1745
rect -503 1357 -497 1733
rect -463 1357 -457 1733
rect -503 1345 -457 1357
rect -407 1733 -361 1745
rect -407 1357 -401 1733
rect -367 1357 -361 1733
rect -407 1345 -361 1357
rect -311 1733 -265 1745
rect -311 1357 -305 1733
rect -271 1357 -265 1733
rect -311 1345 -265 1357
rect -215 1733 -169 1745
rect -215 1357 -209 1733
rect -175 1357 -169 1733
rect -215 1345 -169 1357
rect -119 1733 -73 1745
rect -119 1357 -113 1733
rect -79 1357 -73 1733
rect -119 1345 -73 1357
rect -23 1733 23 1745
rect -23 1357 -17 1733
rect 17 1357 23 1733
rect -23 1345 23 1357
rect 73 1733 119 1745
rect 73 1357 79 1733
rect 113 1357 119 1733
rect 73 1345 119 1357
rect 169 1733 215 1745
rect 169 1357 175 1733
rect 209 1357 215 1733
rect 169 1345 215 1357
rect 265 1733 311 1745
rect 265 1357 271 1733
rect 305 1357 311 1733
rect 265 1345 311 1357
rect 361 1733 407 1745
rect 361 1357 367 1733
rect 401 1357 407 1733
rect 361 1345 407 1357
rect 457 1733 503 1745
rect 457 1357 463 1733
rect 497 1357 503 1733
rect 457 1345 503 1357
rect 553 1733 599 1745
rect 553 1357 559 1733
rect 593 1357 599 1733
rect 553 1345 599 1357
rect 649 1733 695 1745
rect 649 1357 655 1733
rect 689 1357 695 1733
rect 649 1345 695 1357
rect 745 1733 791 1745
rect 745 1357 751 1733
rect 785 1357 791 1733
rect 745 1345 791 1357
rect 841 1733 887 1745
rect 841 1357 847 1733
rect 881 1357 887 1733
rect 841 1345 887 1357
rect 937 1733 983 1745
rect 937 1357 943 1733
rect 977 1357 983 1733
rect 937 1345 983 1357
rect 1033 1733 1079 1745
rect 1033 1357 1039 1733
rect 1073 1357 1079 1733
rect 1033 1345 1079 1357
rect 1129 1733 1175 1745
rect 1129 1357 1135 1733
rect 1169 1357 1175 1733
rect 1129 1345 1175 1357
rect -1037 1307 -979 1313
rect -1037 1273 -1025 1307
rect -991 1273 -979 1307
rect -1037 1267 -979 1273
rect -845 1307 -787 1313
rect -845 1273 -833 1307
rect -799 1273 -787 1307
rect -845 1267 -787 1273
rect -653 1307 -595 1313
rect -653 1273 -641 1307
rect -607 1273 -595 1307
rect -653 1267 -595 1273
rect -461 1307 -403 1313
rect -461 1273 -449 1307
rect -415 1273 -403 1307
rect -461 1267 -403 1273
rect -269 1307 -211 1313
rect -269 1273 -257 1307
rect -223 1273 -211 1307
rect -269 1267 -211 1273
rect -77 1307 -19 1313
rect -77 1273 -65 1307
rect -31 1273 -19 1307
rect -77 1267 -19 1273
rect 115 1307 173 1313
rect 115 1273 127 1307
rect 161 1273 173 1307
rect 115 1267 173 1273
rect 307 1307 365 1313
rect 307 1273 319 1307
rect 353 1273 365 1307
rect 307 1267 365 1273
rect 499 1307 557 1313
rect 499 1273 511 1307
rect 545 1273 557 1307
rect 499 1267 557 1273
rect 691 1307 749 1313
rect 691 1273 703 1307
rect 737 1273 749 1307
rect 691 1267 749 1273
rect 883 1307 941 1313
rect 883 1273 895 1307
rect 929 1273 941 1307
rect 883 1267 941 1273
rect 1075 1307 1133 1313
rect 1075 1273 1087 1307
rect 1121 1273 1133 1307
rect 1075 1267 1133 1273
rect -1037 1199 -979 1205
rect -1037 1165 -1025 1199
rect -991 1165 -979 1199
rect -1037 1159 -979 1165
rect -845 1199 -787 1205
rect -845 1165 -833 1199
rect -799 1165 -787 1199
rect -845 1159 -787 1165
rect -653 1199 -595 1205
rect -653 1165 -641 1199
rect -607 1165 -595 1199
rect -653 1159 -595 1165
rect -461 1199 -403 1205
rect -461 1165 -449 1199
rect -415 1165 -403 1199
rect -461 1159 -403 1165
rect -269 1199 -211 1205
rect -269 1165 -257 1199
rect -223 1165 -211 1199
rect -269 1159 -211 1165
rect -77 1199 -19 1205
rect -77 1165 -65 1199
rect -31 1165 -19 1199
rect -77 1159 -19 1165
rect 115 1199 173 1205
rect 115 1165 127 1199
rect 161 1165 173 1199
rect 115 1159 173 1165
rect 307 1199 365 1205
rect 307 1165 319 1199
rect 353 1165 365 1199
rect 307 1159 365 1165
rect 499 1199 557 1205
rect 499 1165 511 1199
rect 545 1165 557 1199
rect 499 1159 557 1165
rect 691 1199 749 1205
rect 691 1165 703 1199
rect 737 1165 749 1199
rect 691 1159 749 1165
rect 883 1199 941 1205
rect 883 1165 895 1199
rect 929 1165 941 1199
rect 883 1159 941 1165
rect 1075 1199 1133 1205
rect 1075 1165 1087 1199
rect 1121 1165 1133 1199
rect 1075 1159 1133 1165
rect -1175 1115 -1129 1127
rect -1175 739 -1169 1115
rect -1135 739 -1129 1115
rect -1175 727 -1129 739
rect -1079 1115 -1033 1127
rect -1079 739 -1073 1115
rect -1039 739 -1033 1115
rect -1079 727 -1033 739
rect -983 1115 -937 1127
rect -983 739 -977 1115
rect -943 739 -937 1115
rect -983 727 -937 739
rect -887 1115 -841 1127
rect -887 739 -881 1115
rect -847 739 -841 1115
rect -887 727 -841 739
rect -791 1115 -745 1127
rect -791 739 -785 1115
rect -751 739 -745 1115
rect -791 727 -745 739
rect -695 1115 -649 1127
rect -695 739 -689 1115
rect -655 739 -649 1115
rect -695 727 -649 739
rect -599 1115 -553 1127
rect -599 739 -593 1115
rect -559 739 -553 1115
rect -599 727 -553 739
rect -503 1115 -457 1127
rect -503 739 -497 1115
rect -463 739 -457 1115
rect -503 727 -457 739
rect -407 1115 -361 1127
rect -407 739 -401 1115
rect -367 739 -361 1115
rect -407 727 -361 739
rect -311 1115 -265 1127
rect -311 739 -305 1115
rect -271 739 -265 1115
rect -311 727 -265 739
rect -215 1115 -169 1127
rect -215 739 -209 1115
rect -175 739 -169 1115
rect -215 727 -169 739
rect -119 1115 -73 1127
rect -119 739 -113 1115
rect -79 739 -73 1115
rect -119 727 -73 739
rect -23 1115 23 1127
rect -23 739 -17 1115
rect 17 739 23 1115
rect -23 727 23 739
rect 73 1115 119 1127
rect 73 739 79 1115
rect 113 739 119 1115
rect 73 727 119 739
rect 169 1115 215 1127
rect 169 739 175 1115
rect 209 739 215 1115
rect 169 727 215 739
rect 265 1115 311 1127
rect 265 739 271 1115
rect 305 739 311 1115
rect 265 727 311 739
rect 361 1115 407 1127
rect 361 739 367 1115
rect 401 739 407 1115
rect 361 727 407 739
rect 457 1115 503 1127
rect 457 739 463 1115
rect 497 739 503 1115
rect 457 727 503 739
rect 553 1115 599 1127
rect 553 739 559 1115
rect 593 739 599 1115
rect 553 727 599 739
rect 649 1115 695 1127
rect 649 739 655 1115
rect 689 739 695 1115
rect 649 727 695 739
rect 745 1115 791 1127
rect 745 739 751 1115
rect 785 739 791 1115
rect 745 727 791 739
rect 841 1115 887 1127
rect 841 739 847 1115
rect 881 739 887 1115
rect 841 727 887 739
rect 937 1115 983 1127
rect 937 739 943 1115
rect 977 739 983 1115
rect 937 727 983 739
rect 1033 1115 1079 1127
rect 1033 739 1039 1115
rect 1073 739 1079 1115
rect 1033 727 1079 739
rect 1129 1115 1175 1127
rect 1129 739 1135 1115
rect 1169 739 1175 1115
rect 1129 727 1175 739
rect -1133 689 -1075 695
rect -1133 655 -1121 689
rect -1087 655 -1075 689
rect -1133 649 -1075 655
rect -941 689 -883 695
rect -941 655 -929 689
rect -895 655 -883 689
rect -941 649 -883 655
rect -749 689 -691 695
rect -749 655 -737 689
rect -703 655 -691 689
rect -749 649 -691 655
rect -557 689 -499 695
rect -557 655 -545 689
rect -511 655 -499 689
rect -557 649 -499 655
rect -365 689 -307 695
rect -365 655 -353 689
rect -319 655 -307 689
rect -365 649 -307 655
rect -173 689 -115 695
rect -173 655 -161 689
rect -127 655 -115 689
rect -173 649 -115 655
rect 19 689 77 695
rect 19 655 31 689
rect 65 655 77 689
rect 19 649 77 655
rect 211 689 269 695
rect 211 655 223 689
rect 257 655 269 689
rect 211 649 269 655
rect 403 689 461 695
rect 403 655 415 689
rect 449 655 461 689
rect 403 649 461 655
rect 595 689 653 695
rect 595 655 607 689
rect 641 655 653 689
rect 595 649 653 655
rect 787 689 845 695
rect 787 655 799 689
rect 833 655 845 689
rect 787 649 845 655
rect 979 689 1037 695
rect 979 655 991 689
rect 1025 655 1037 689
rect 979 649 1037 655
rect -1133 581 -1075 587
rect -1133 547 -1121 581
rect -1087 547 -1075 581
rect -1133 541 -1075 547
rect -941 581 -883 587
rect -941 547 -929 581
rect -895 547 -883 581
rect -941 541 -883 547
rect -749 581 -691 587
rect -749 547 -737 581
rect -703 547 -691 581
rect -749 541 -691 547
rect -557 581 -499 587
rect -557 547 -545 581
rect -511 547 -499 581
rect -557 541 -499 547
rect -365 581 -307 587
rect -365 547 -353 581
rect -319 547 -307 581
rect -365 541 -307 547
rect -173 581 -115 587
rect -173 547 -161 581
rect -127 547 -115 581
rect -173 541 -115 547
rect 19 581 77 587
rect 19 547 31 581
rect 65 547 77 581
rect 19 541 77 547
rect 211 581 269 587
rect 211 547 223 581
rect 257 547 269 581
rect 211 541 269 547
rect 403 581 461 587
rect 403 547 415 581
rect 449 547 461 581
rect 403 541 461 547
rect 595 581 653 587
rect 595 547 607 581
rect 641 547 653 581
rect 595 541 653 547
rect 787 581 845 587
rect 787 547 799 581
rect 833 547 845 581
rect 787 541 845 547
rect 979 581 1037 587
rect 979 547 991 581
rect 1025 547 1037 581
rect 979 541 1037 547
rect -1175 497 -1129 509
rect -1175 121 -1169 497
rect -1135 121 -1129 497
rect -1175 109 -1129 121
rect -1079 497 -1033 509
rect -1079 121 -1073 497
rect -1039 121 -1033 497
rect -1079 109 -1033 121
rect -983 497 -937 509
rect -983 121 -977 497
rect -943 121 -937 497
rect -983 109 -937 121
rect -887 497 -841 509
rect -887 121 -881 497
rect -847 121 -841 497
rect -887 109 -841 121
rect -791 497 -745 509
rect -791 121 -785 497
rect -751 121 -745 497
rect -791 109 -745 121
rect -695 497 -649 509
rect -695 121 -689 497
rect -655 121 -649 497
rect -695 109 -649 121
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect 649 497 695 509
rect 649 121 655 497
rect 689 121 695 497
rect 649 109 695 121
rect 745 497 791 509
rect 745 121 751 497
rect 785 121 791 497
rect 745 109 791 121
rect 841 497 887 509
rect 841 121 847 497
rect 881 121 887 497
rect 841 109 887 121
rect 937 497 983 509
rect 937 121 943 497
rect 977 121 983 497
rect 937 109 983 121
rect 1033 497 1079 509
rect 1033 121 1039 497
rect 1073 121 1079 497
rect 1033 109 1079 121
rect 1129 497 1175 509
rect 1129 121 1135 497
rect 1169 121 1175 497
rect 1129 109 1175 121
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect -1175 -121 -1129 -109
rect -1175 -497 -1169 -121
rect -1135 -497 -1129 -121
rect -1175 -509 -1129 -497
rect -1079 -121 -1033 -109
rect -1079 -497 -1073 -121
rect -1039 -497 -1033 -121
rect -1079 -509 -1033 -497
rect -983 -121 -937 -109
rect -983 -497 -977 -121
rect -943 -497 -937 -121
rect -983 -509 -937 -497
rect -887 -121 -841 -109
rect -887 -497 -881 -121
rect -847 -497 -841 -121
rect -887 -509 -841 -497
rect -791 -121 -745 -109
rect -791 -497 -785 -121
rect -751 -497 -745 -121
rect -791 -509 -745 -497
rect -695 -121 -649 -109
rect -695 -497 -689 -121
rect -655 -497 -649 -121
rect -695 -509 -649 -497
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect 649 -121 695 -109
rect 649 -497 655 -121
rect 689 -497 695 -121
rect 649 -509 695 -497
rect 745 -121 791 -109
rect 745 -497 751 -121
rect 785 -497 791 -121
rect 745 -509 791 -497
rect 841 -121 887 -109
rect 841 -497 847 -121
rect 881 -497 887 -121
rect 841 -509 887 -497
rect 937 -121 983 -109
rect 937 -497 943 -121
rect 977 -497 983 -121
rect 937 -509 983 -497
rect 1033 -121 1079 -109
rect 1033 -497 1039 -121
rect 1073 -497 1079 -121
rect 1033 -509 1079 -497
rect 1129 -121 1175 -109
rect 1129 -497 1135 -121
rect 1169 -497 1175 -121
rect 1129 -509 1175 -497
rect -1133 -547 -1075 -541
rect -1133 -581 -1121 -547
rect -1087 -581 -1075 -547
rect -1133 -587 -1075 -581
rect -941 -547 -883 -541
rect -941 -581 -929 -547
rect -895 -581 -883 -547
rect -941 -587 -883 -581
rect -749 -547 -691 -541
rect -749 -581 -737 -547
rect -703 -581 -691 -547
rect -749 -587 -691 -581
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
rect 595 -547 653 -541
rect 595 -581 607 -547
rect 641 -581 653 -547
rect 595 -587 653 -581
rect 787 -547 845 -541
rect 787 -581 799 -547
rect 833 -581 845 -547
rect 787 -587 845 -581
rect 979 -547 1037 -541
rect 979 -581 991 -547
rect 1025 -581 1037 -547
rect 979 -587 1037 -581
rect -1133 -655 -1075 -649
rect -1133 -689 -1121 -655
rect -1087 -689 -1075 -655
rect -1133 -695 -1075 -689
rect -941 -655 -883 -649
rect -941 -689 -929 -655
rect -895 -689 -883 -655
rect -941 -695 -883 -689
rect -749 -655 -691 -649
rect -749 -689 -737 -655
rect -703 -689 -691 -655
rect -749 -695 -691 -689
rect -557 -655 -499 -649
rect -557 -689 -545 -655
rect -511 -689 -499 -655
rect -557 -695 -499 -689
rect -365 -655 -307 -649
rect -365 -689 -353 -655
rect -319 -689 -307 -655
rect -365 -695 -307 -689
rect -173 -655 -115 -649
rect -173 -689 -161 -655
rect -127 -689 -115 -655
rect -173 -695 -115 -689
rect 19 -655 77 -649
rect 19 -689 31 -655
rect 65 -689 77 -655
rect 19 -695 77 -689
rect 211 -655 269 -649
rect 211 -689 223 -655
rect 257 -689 269 -655
rect 211 -695 269 -689
rect 403 -655 461 -649
rect 403 -689 415 -655
rect 449 -689 461 -655
rect 403 -695 461 -689
rect 595 -655 653 -649
rect 595 -689 607 -655
rect 641 -689 653 -655
rect 595 -695 653 -689
rect 787 -655 845 -649
rect 787 -689 799 -655
rect 833 -689 845 -655
rect 787 -695 845 -689
rect 979 -655 1037 -649
rect 979 -689 991 -655
rect 1025 -689 1037 -655
rect 979 -695 1037 -689
rect -1175 -739 -1129 -727
rect -1175 -1115 -1169 -739
rect -1135 -1115 -1129 -739
rect -1175 -1127 -1129 -1115
rect -1079 -739 -1033 -727
rect -1079 -1115 -1073 -739
rect -1039 -1115 -1033 -739
rect -1079 -1127 -1033 -1115
rect -983 -739 -937 -727
rect -983 -1115 -977 -739
rect -943 -1115 -937 -739
rect -983 -1127 -937 -1115
rect -887 -739 -841 -727
rect -887 -1115 -881 -739
rect -847 -1115 -841 -739
rect -887 -1127 -841 -1115
rect -791 -739 -745 -727
rect -791 -1115 -785 -739
rect -751 -1115 -745 -739
rect -791 -1127 -745 -1115
rect -695 -739 -649 -727
rect -695 -1115 -689 -739
rect -655 -1115 -649 -739
rect -695 -1127 -649 -1115
rect -599 -739 -553 -727
rect -599 -1115 -593 -739
rect -559 -1115 -553 -739
rect -599 -1127 -553 -1115
rect -503 -739 -457 -727
rect -503 -1115 -497 -739
rect -463 -1115 -457 -739
rect -503 -1127 -457 -1115
rect -407 -739 -361 -727
rect -407 -1115 -401 -739
rect -367 -1115 -361 -739
rect -407 -1127 -361 -1115
rect -311 -739 -265 -727
rect -311 -1115 -305 -739
rect -271 -1115 -265 -739
rect -311 -1127 -265 -1115
rect -215 -739 -169 -727
rect -215 -1115 -209 -739
rect -175 -1115 -169 -739
rect -215 -1127 -169 -1115
rect -119 -739 -73 -727
rect -119 -1115 -113 -739
rect -79 -1115 -73 -739
rect -119 -1127 -73 -1115
rect -23 -739 23 -727
rect -23 -1115 -17 -739
rect 17 -1115 23 -739
rect -23 -1127 23 -1115
rect 73 -739 119 -727
rect 73 -1115 79 -739
rect 113 -1115 119 -739
rect 73 -1127 119 -1115
rect 169 -739 215 -727
rect 169 -1115 175 -739
rect 209 -1115 215 -739
rect 169 -1127 215 -1115
rect 265 -739 311 -727
rect 265 -1115 271 -739
rect 305 -1115 311 -739
rect 265 -1127 311 -1115
rect 361 -739 407 -727
rect 361 -1115 367 -739
rect 401 -1115 407 -739
rect 361 -1127 407 -1115
rect 457 -739 503 -727
rect 457 -1115 463 -739
rect 497 -1115 503 -739
rect 457 -1127 503 -1115
rect 553 -739 599 -727
rect 553 -1115 559 -739
rect 593 -1115 599 -739
rect 553 -1127 599 -1115
rect 649 -739 695 -727
rect 649 -1115 655 -739
rect 689 -1115 695 -739
rect 649 -1127 695 -1115
rect 745 -739 791 -727
rect 745 -1115 751 -739
rect 785 -1115 791 -739
rect 745 -1127 791 -1115
rect 841 -739 887 -727
rect 841 -1115 847 -739
rect 881 -1115 887 -739
rect 841 -1127 887 -1115
rect 937 -739 983 -727
rect 937 -1115 943 -739
rect 977 -1115 983 -739
rect 937 -1127 983 -1115
rect 1033 -739 1079 -727
rect 1033 -1115 1039 -739
rect 1073 -1115 1079 -739
rect 1033 -1127 1079 -1115
rect 1129 -739 1175 -727
rect 1129 -1115 1135 -739
rect 1169 -1115 1175 -739
rect 1129 -1127 1175 -1115
rect -1037 -1165 -979 -1159
rect -1037 -1199 -1025 -1165
rect -991 -1199 -979 -1165
rect -1037 -1205 -979 -1199
rect -845 -1165 -787 -1159
rect -845 -1199 -833 -1165
rect -799 -1199 -787 -1165
rect -845 -1205 -787 -1199
rect -653 -1165 -595 -1159
rect -653 -1199 -641 -1165
rect -607 -1199 -595 -1165
rect -653 -1205 -595 -1199
rect -461 -1165 -403 -1159
rect -461 -1199 -449 -1165
rect -415 -1199 -403 -1165
rect -461 -1205 -403 -1199
rect -269 -1165 -211 -1159
rect -269 -1199 -257 -1165
rect -223 -1199 -211 -1165
rect -269 -1205 -211 -1199
rect -77 -1165 -19 -1159
rect -77 -1199 -65 -1165
rect -31 -1199 -19 -1165
rect -77 -1205 -19 -1199
rect 115 -1165 173 -1159
rect 115 -1199 127 -1165
rect 161 -1199 173 -1165
rect 115 -1205 173 -1199
rect 307 -1165 365 -1159
rect 307 -1199 319 -1165
rect 353 -1199 365 -1165
rect 307 -1205 365 -1199
rect 499 -1165 557 -1159
rect 499 -1199 511 -1165
rect 545 -1199 557 -1165
rect 499 -1205 557 -1199
rect 691 -1165 749 -1159
rect 691 -1199 703 -1165
rect 737 -1199 749 -1165
rect 691 -1205 749 -1199
rect 883 -1165 941 -1159
rect 883 -1199 895 -1165
rect 929 -1199 941 -1165
rect 883 -1205 941 -1199
rect 1075 -1165 1133 -1159
rect 1075 -1199 1087 -1165
rect 1121 -1199 1133 -1165
rect 1075 -1205 1133 -1199
rect -1037 -1273 -979 -1267
rect -1037 -1307 -1025 -1273
rect -991 -1307 -979 -1273
rect -1037 -1313 -979 -1307
rect -845 -1273 -787 -1267
rect -845 -1307 -833 -1273
rect -799 -1307 -787 -1273
rect -845 -1313 -787 -1307
rect -653 -1273 -595 -1267
rect -653 -1307 -641 -1273
rect -607 -1307 -595 -1273
rect -653 -1313 -595 -1307
rect -461 -1273 -403 -1267
rect -461 -1307 -449 -1273
rect -415 -1307 -403 -1273
rect -461 -1313 -403 -1307
rect -269 -1273 -211 -1267
rect -269 -1307 -257 -1273
rect -223 -1307 -211 -1273
rect -269 -1313 -211 -1307
rect -77 -1273 -19 -1267
rect -77 -1307 -65 -1273
rect -31 -1307 -19 -1273
rect -77 -1313 -19 -1307
rect 115 -1273 173 -1267
rect 115 -1307 127 -1273
rect 161 -1307 173 -1273
rect 115 -1313 173 -1307
rect 307 -1273 365 -1267
rect 307 -1307 319 -1273
rect 353 -1307 365 -1273
rect 307 -1313 365 -1307
rect 499 -1273 557 -1267
rect 499 -1307 511 -1273
rect 545 -1307 557 -1273
rect 499 -1313 557 -1307
rect 691 -1273 749 -1267
rect 691 -1307 703 -1273
rect 737 -1307 749 -1273
rect 691 -1313 749 -1307
rect 883 -1273 941 -1267
rect 883 -1307 895 -1273
rect 929 -1307 941 -1273
rect 883 -1313 941 -1307
rect 1075 -1273 1133 -1267
rect 1075 -1307 1087 -1273
rect 1121 -1307 1133 -1273
rect 1075 -1313 1133 -1307
rect -1175 -1357 -1129 -1345
rect -1175 -1733 -1169 -1357
rect -1135 -1733 -1129 -1357
rect -1175 -1745 -1129 -1733
rect -1079 -1357 -1033 -1345
rect -1079 -1733 -1073 -1357
rect -1039 -1733 -1033 -1357
rect -1079 -1745 -1033 -1733
rect -983 -1357 -937 -1345
rect -983 -1733 -977 -1357
rect -943 -1733 -937 -1357
rect -983 -1745 -937 -1733
rect -887 -1357 -841 -1345
rect -887 -1733 -881 -1357
rect -847 -1733 -841 -1357
rect -887 -1745 -841 -1733
rect -791 -1357 -745 -1345
rect -791 -1733 -785 -1357
rect -751 -1733 -745 -1357
rect -791 -1745 -745 -1733
rect -695 -1357 -649 -1345
rect -695 -1733 -689 -1357
rect -655 -1733 -649 -1357
rect -695 -1745 -649 -1733
rect -599 -1357 -553 -1345
rect -599 -1733 -593 -1357
rect -559 -1733 -553 -1357
rect -599 -1745 -553 -1733
rect -503 -1357 -457 -1345
rect -503 -1733 -497 -1357
rect -463 -1733 -457 -1357
rect -503 -1745 -457 -1733
rect -407 -1357 -361 -1345
rect -407 -1733 -401 -1357
rect -367 -1733 -361 -1357
rect -407 -1745 -361 -1733
rect -311 -1357 -265 -1345
rect -311 -1733 -305 -1357
rect -271 -1733 -265 -1357
rect -311 -1745 -265 -1733
rect -215 -1357 -169 -1345
rect -215 -1733 -209 -1357
rect -175 -1733 -169 -1357
rect -215 -1745 -169 -1733
rect -119 -1357 -73 -1345
rect -119 -1733 -113 -1357
rect -79 -1733 -73 -1357
rect -119 -1745 -73 -1733
rect -23 -1357 23 -1345
rect -23 -1733 -17 -1357
rect 17 -1733 23 -1357
rect -23 -1745 23 -1733
rect 73 -1357 119 -1345
rect 73 -1733 79 -1357
rect 113 -1733 119 -1357
rect 73 -1745 119 -1733
rect 169 -1357 215 -1345
rect 169 -1733 175 -1357
rect 209 -1733 215 -1357
rect 169 -1745 215 -1733
rect 265 -1357 311 -1345
rect 265 -1733 271 -1357
rect 305 -1733 311 -1357
rect 265 -1745 311 -1733
rect 361 -1357 407 -1345
rect 361 -1733 367 -1357
rect 401 -1733 407 -1357
rect 361 -1745 407 -1733
rect 457 -1357 503 -1345
rect 457 -1733 463 -1357
rect 497 -1733 503 -1357
rect 457 -1745 503 -1733
rect 553 -1357 599 -1345
rect 553 -1733 559 -1357
rect 593 -1733 599 -1357
rect 553 -1745 599 -1733
rect 649 -1357 695 -1345
rect 649 -1733 655 -1357
rect 689 -1733 695 -1357
rect 649 -1745 695 -1733
rect 745 -1357 791 -1345
rect 745 -1733 751 -1357
rect 785 -1733 791 -1357
rect 745 -1745 791 -1733
rect 841 -1357 887 -1345
rect 841 -1733 847 -1357
rect 881 -1733 887 -1357
rect 841 -1745 887 -1733
rect 937 -1357 983 -1345
rect 937 -1733 943 -1357
rect 977 -1733 983 -1357
rect 937 -1745 983 -1733
rect 1033 -1357 1079 -1345
rect 1033 -1733 1039 -1357
rect 1073 -1733 1079 -1357
rect 1033 -1745 1079 -1733
rect 1129 -1357 1175 -1345
rect 1129 -1733 1135 -1357
rect 1169 -1733 1175 -1357
rect 1129 -1745 1175 -1733
rect -1133 -1783 -1075 -1777
rect -1133 -1817 -1121 -1783
rect -1087 -1817 -1075 -1783
rect -1133 -1823 -1075 -1817
rect -941 -1783 -883 -1777
rect -941 -1817 -929 -1783
rect -895 -1817 -883 -1783
rect -941 -1823 -883 -1817
rect -749 -1783 -691 -1777
rect -749 -1817 -737 -1783
rect -703 -1817 -691 -1783
rect -749 -1823 -691 -1817
rect -557 -1783 -499 -1777
rect -557 -1817 -545 -1783
rect -511 -1817 -499 -1783
rect -557 -1823 -499 -1817
rect -365 -1783 -307 -1777
rect -365 -1817 -353 -1783
rect -319 -1817 -307 -1783
rect -365 -1823 -307 -1817
rect -173 -1783 -115 -1777
rect -173 -1817 -161 -1783
rect -127 -1817 -115 -1783
rect -173 -1823 -115 -1817
rect 19 -1783 77 -1777
rect 19 -1817 31 -1783
rect 65 -1817 77 -1783
rect 19 -1823 77 -1817
rect 211 -1783 269 -1777
rect 211 -1817 223 -1783
rect 257 -1817 269 -1783
rect 211 -1823 269 -1817
rect 403 -1783 461 -1777
rect 403 -1817 415 -1783
rect 449 -1817 461 -1783
rect 403 -1823 461 -1817
rect 595 -1783 653 -1777
rect 595 -1817 607 -1783
rect 641 -1817 653 -1783
rect 595 -1823 653 -1817
rect 787 -1783 845 -1777
rect 787 -1817 799 -1783
rect 833 -1817 845 -1783
rect 787 -1823 845 -1817
rect 979 -1783 1037 -1777
rect 979 -1817 991 -1783
rect 1025 -1817 1037 -1783
rect 979 -1823 1037 -1817
rect -1133 -1891 -1075 -1885
rect -1133 -1925 -1121 -1891
rect -1087 -1925 -1075 -1891
rect -1133 -1931 -1075 -1925
rect -941 -1891 -883 -1885
rect -941 -1925 -929 -1891
rect -895 -1925 -883 -1891
rect -941 -1931 -883 -1925
rect -749 -1891 -691 -1885
rect -749 -1925 -737 -1891
rect -703 -1925 -691 -1891
rect -749 -1931 -691 -1925
rect -557 -1891 -499 -1885
rect -557 -1925 -545 -1891
rect -511 -1925 -499 -1891
rect -557 -1931 -499 -1925
rect -365 -1891 -307 -1885
rect -365 -1925 -353 -1891
rect -319 -1925 -307 -1891
rect -365 -1931 -307 -1925
rect -173 -1891 -115 -1885
rect -173 -1925 -161 -1891
rect -127 -1925 -115 -1891
rect -173 -1931 -115 -1925
rect 19 -1891 77 -1885
rect 19 -1925 31 -1891
rect 65 -1925 77 -1891
rect 19 -1931 77 -1925
rect 211 -1891 269 -1885
rect 211 -1925 223 -1891
rect 257 -1925 269 -1891
rect 211 -1931 269 -1925
rect 403 -1891 461 -1885
rect 403 -1925 415 -1891
rect 449 -1925 461 -1891
rect 403 -1931 461 -1925
rect 595 -1891 653 -1885
rect 595 -1925 607 -1891
rect 641 -1925 653 -1891
rect 595 -1931 653 -1925
rect 787 -1891 845 -1885
rect 787 -1925 799 -1891
rect 833 -1925 845 -1891
rect 787 -1931 845 -1925
rect 979 -1891 1037 -1885
rect 979 -1925 991 -1891
rect 1025 -1925 1037 -1891
rect 979 -1931 1037 -1925
rect -1175 -1975 -1129 -1963
rect -1175 -2351 -1169 -1975
rect -1135 -2351 -1129 -1975
rect -1175 -2363 -1129 -2351
rect -1079 -1975 -1033 -1963
rect -1079 -2351 -1073 -1975
rect -1039 -2351 -1033 -1975
rect -1079 -2363 -1033 -2351
rect -983 -1975 -937 -1963
rect -983 -2351 -977 -1975
rect -943 -2351 -937 -1975
rect -983 -2363 -937 -2351
rect -887 -1975 -841 -1963
rect -887 -2351 -881 -1975
rect -847 -2351 -841 -1975
rect -887 -2363 -841 -2351
rect -791 -1975 -745 -1963
rect -791 -2351 -785 -1975
rect -751 -2351 -745 -1975
rect -791 -2363 -745 -2351
rect -695 -1975 -649 -1963
rect -695 -2351 -689 -1975
rect -655 -2351 -649 -1975
rect -695 -2363 -649 -2351
rect -599 -1975 -553 -1963
rect -599 -2351 -593 -1975
rect -559 -2351 -553 -1975
rect -599 -2363 -553 -2351
rect -503 -1975 -457 -1963
rect -503 -2351 -497 -1975
rect -463 -2351 -457 -1975
rect -503 -2363 -457 -2351
rect -407 -1975 -361 -1963
rect -407 -2351 -401 -1975
rect -367 -2351 -361 -1975
rect -407 -2363 -361 -2351
rect -311 -1975 -265 -1963
rect -311 -2351 -305 -1975
rect -271 -2351 -265 -1975
rect -311 -2363 -265 -2351
rect -215 -1975 -169 -1963
rect -215 -2351 -209 -1975
rect -175 -2351 -169 -1975
rect -215 -2363 -169 -2351
rect -119 -1975 -73 -1963
rect -119 -2351 -113 -1975
rect -79 -2351 -73 -1975
rect -119 -2363 -73 -2351
rect -23 -1975 23 -1963
rect -23 -2351 -17 -1975
rect 17 -2351 23 -1975
rect -23 -2363 23 -2351
rect 73 -1975 119 -1963
rect 73 -2351 79 -1975
rect 113 -2351 119 -1975
rect 73 -2363 119 -2351
rect 169 -1975 215 -1963
rect 169 -2351 175 -1975
rect 209 -2351 215 -1975
rect 169 -2363 215 -2351
rect 265 -1975 311 -1963
rect 265 -2351 271 -1975
rect 305 -2351 311 -1975
rect 265 -2363 311 -2351
rect 361 -1975 407 -1963
rect 361 -2351 367 -1975
rect 401 -2351 407 -1975
rect 361 -2363 407 -2351
rect 457 -1975 503 -1963
rect 457 -2351 463 -1975
rect 497 -2351 503 -1975
rect 457 -2363 503 -2351
rect 553 -1975 599 -1963
rect 553 -2351 559 -1975
rect 593 -2351 599 -1975
rect 553 -2363 599 -2351
rect 649 -1975 695 -1963
rect 649 -2351 655 -1975
rect 689 -2351 695 -1975
rect 649 -2363 695 -2351
rect 745 -1975 791 -1963
rect 745 -2351 751 -1975
rect 785 -2351 791 -1975
rect 745 -2363 791 -2351
rect 841 -1975 887 -1963
rect 841 -2351 847 -1975
rect 881 -2351 887 -1975
rect 841 -2363 887 -2351
rect 937 -1975 983 -1963
rect 937 -2351 943 -1975
rect 977 -2351 983 -1975
rect 937 -2363 983 -2351
rect 1033 -1975 1079 -1963
rect 1033 -2351 1039 -1975
rect 1073 -2351 1079 -1975
rect 1033 -2363 1079 -2351
rect 1129 -1975 1175 -1963
rect 1129 -2351 1135 -1975
rect 1169 -2351 1175 -1975
rect 1129 -2363 1175 -2351
rect -1037 -2401 -979 -2395
rect -1037 -2435 -1025 -2401
rect -991 -2435 -979 -2401
rect -1037 -2441 -979 -2435
rect -845 -2401 -787 -2395
rect -845 -2435 -833 -2401
rect -799 -2435 -787 -2401
rect -845 -2441 -787 -2435
rect -653 -2401 -595 -2395
rect -653 -2435 -641 -2401
rect -607 -2435 -595 -2401
rect -653 -2441 -595 -2435
rect -461 -2401 -403 -2395
rect -461 -2435 -449 -2401
rect -415 -2435 -403 -2401
rect -461 -2441 -403 -2435
rect -269 -2401 -211 -2395
rect -269 -2435 -257 -2401
rect -223 -2435 -211 -2401
rect -269 -2441 -211 -2435
rect -77 -2401 -19 -2395
rect -77 -2435 -65 -2401
rect -31 -2435 -19 -2401
rect -77 -2441 -19 -2435
rect 115 -2401 173 -2395
rect 115 -2435 127 -2401
rect 161 -2435 173 -2401
rect 115 -2441 173 -2435
rect 307 -2401 365 -2395
rect 307 -2435 319 -2401
rect 353 -2435 365 -2401
rect 307 -2441 365 -2435
rect 499 -2401 557 -2395
rect 499 -2435 511 -2401
rect 545 -2435 557 -2401
rect 499 -2441 557 -2435
rect 691 -2401 749 -2395
rect 691 -2435 703 -2401
rect 737 -2435 749 -2401
rect 691 -2441 749 -2435
rect 883 -2401 941 -2395
rect 883 -2435 895 -2401
rect 929 -2435 941 -2401
rect 883 -2441 941 -2435
rect 1075 -2401 1133 -2395
rect 1075 -2435 1087 -2401
rect 1121 -2435 1133 -2401
rect 1075 -2441 1133 -2435
rect -1037 -2509 -979 -2503
rect -1037 -2543 -1025 -2509
rect -991 -2543 -979 -2509
rect -1037 -2549 -979 -2543
rect -845 -2509 -787 -2503
rect -845 -2543 -833 -2509
rect -799 -2543 -787 -2509
rect -845 -2549 -787 -2543
rect -653 -2509 -595 -2503
rect -653 -2543 -641 -2509
rect -607 -2543 -595 -2509
rect -653 -2549 -595 -2543
rect -461 -2509 -403 -2503
rect -461 -2543 -449 -2509
rect -415 -2543 -403 -2509
rect -461 -2549 -403 -2543
rect -269 -2509 -211 -2503
rect -269 -2543 -257 -2509
rect -223 -2543 -211 -2509
rect -269 -2549 -211 -2543
rect -77 -2509 -19 -2503
rect -77 -2543 -65 -2509
rect -31 -2543 -19 -2509
rect -77 -2549 -19 -2543
rect 115 -2509 173 -2503
rect 115 -2543 127 -2509
rect 161 -2543 173 -2509
rect 115 -2549 173 -2543
rect 307 -2509 365 -2503
rect 307 -2543 319 -2509
rect 353 -2543 365 -2509
rect 307 -2549 365 -2543
rect 499 -2509 557 -2503
rect 499 -2543 511 -2509
rect 545 -2543 557 -2509
rect 499 -2549 557 -2543
rect 691 -2509 749 -2503
rect 691 -2543 703 -2509
rect 737 -2543 749 -2509
rect 691 -2549 749 -2543
rect 883 -2509 941 -2503
rect 883 -2543 895 -2509
rect 929 -2543 941 -2509
rect 883 -2549 941 -2543
rect 1075 -2509 1133 -2503
rect 1075 -2543 1087 -2509
rect 1121 -2543 1133 -2509
rect 1075 -2549 1133 -2543
rect -1175 -2593 -1129 -2581
rect -1175 -2969 -1169 -2593
rect -1135 -2969 -1129 -2593
rect -1175 -2981 -1129 -2969
rect -1079 -2593 -1033 -2581
rect -1079 -2969 -1073 -2593
rect -1039 -2969 -1033 -2593
rect -1079 -2981 -1033 -2969
rect -983 -2593 -937 -2581
rect -983 -2969 -977 -2593
rect -943 -2969 -937 -2593
rect -983 -2981 -937 -2969
rect -887 -2593 -841 -2581
rect -887 -2969 -881 -2593
rect -847 -2969 -841 -2593
rect -887 -2981 -841 -2969
rect -791 -2593 -745 -2581
rect -791 -2969 -785 -2593
rect -751 -2969 -745 -2593
rect -791 -2981 -745 -2969
rect -695 -2593 -649 -2581
rect -695 -2969 -689 -2593
rect -655 -2969 -649 -2593
rect -695 -2981 -649 -2969
rect -599 -2593 -553 -2581
rect -599 -2969 -593 -2593
rect -559 -2969 -553 -2593
rect -599 -2981 -553 -2969
rect -503 -2593 -457 -2581
rect -503 -2969 -497 -2593
rect -463 -2969 -457 -2593
rect -503 -2981 -457 -2969
rect -407 -2593 -361 -2581
rect -407 -2969 -401 -2593
rect -367 -2969 -361 -2593
rect -407 -2981 -361 -2969
rect -311 -2593 -265 -2581
rect -311 -2969 -305 -2593
rect -271 -2969 -265 -2593
rect -311 -2981 -265 -2969
rect -215 -2593 -169 -2581
rect -215 -2969 -209 -2593
rect -175 -2969 -169 -2593
rect -215 -2981 -169 -2969
rect -119 -2593 -73 -2581
rect -119 -2969 -113 -2593
rect -79 -2969 -73 -2593
rect -119 -2981 -73 -2969
rect -23 -2593 23 -2581
rect -23 -2969 -17 -2593
rect 17 -2969 23 -2593
rect -23 -2981 23 -2969
rect 73 -2593 119 -2581
rect 73 -2969 79 -2593
rect 113 -2969 119 -2593
rect 73 -2981 119 -2969
rect 169 -2593 215 -2581
rect 169 -2969 175 -2593
rect 209 -2969 215 -2593
rect 169 -2981 215 -2969
rect 265 -2593 311 -2581
rect 265 -2969 271 -2593
rect 305 -2969 311 -2593
rect 265 -2981 311 -2969
rect 361 -2593 407 -2581
rect 361 -2969 367 -2593
rect 401 -2969 407 -2593
rect 361 -2981 407 -2969
rect 457 -2593 503 -2581
rect 457 -2969 463 -2593
rect 497 -2969 503 -2593
rect 457 -2981 503 -2969
rect 553 -2593 599 -2581
rect 553 -2969 559 -2593
rect 593 -2969 599 -2593
rect 553 -2981 599 -2969
rect 649 -2593 695 -2581
rect 649 -2969 655 -2593
rect 689 -2969 695 -2593
rect 649 -2981 695 -2969
rect 745 -2593 791 -2581
rect 745 -2969 751 -2593
rect 785 -2969 791 -2593
rect 745 -2981 791 -2969
rect 841 -2593 887 -2581
rect 841 -2969 847 -2593
rect 881 -2969 887 -2593
rect 841 -2981 887 -2969
rect 937 -2593 983 -2581
rect 937 -2969 943 -2593
rect 977 -2969 983 -2593
rect 937 -2981 983 -2969
rect 1033 -2593 1079 -2581
rect 1033 -2969 1039 -2593
rect 1073 -2969 1079 -2593
rect 1033 -2981 1079 -2969
rect 1129 -2593 1175 -2581
rect 1129 -2969 1135 -2593
rect 1169 -2969 1175 -2593
rect 1129 -2981 1175 -2969
rect -1133 -3019 -1075 -3013
rect -1133 -3053 -1121 -3019
rect -1087 -3053 -1075 -3019
rect -1133 -3059 -1075 -3053
rect -941 -3019 -883 -3013
rect -941 -3053 -929 -3019
rect -895 -3053 -883 -3019
rect -941 -3059 -883 -3053
rect -749 -3019 -691 -3013
rect -749 -3053 -737 -3019
rect -703 -3053 -691 -3019
rect -749 -3059 -691 -3053
rect -557 -3019 -499 -3013
rect -557 -3053 -545 -3019
rect -511 -3053 -499 -3019
rect -557 -3059 -499 -3053
rect -365 -3019 -307 -3013
rect -365 -3053 -353 -3019
rect -319 -3053 -307 -3019
rect -365 -3059 -307 -3053
rect -173 -3019 -115 -3013
rect -173 -3053 -161 -3019
rect -127 -3053 -115 -3019
rect -173 -3059 -115 -3053
rect 19 -3019 77 -3013
rect 19 -3053 31 -3019
rect 65 -3053 77 -3019
rect 19 -3059 77 -3053
rect 211 -3019 269 -3013
rect 211 -3053 223 -3019
rect 257 -3053 269 -3019
rect 211 -3059 269 -3053
rect 403 -3019 461 -3013
rect 403 -3053 415 -3019
rect 449 -3053 461 -3019
rect 403 -3059 461 -3053
rect 595 -3019 653 -3013
rect 595 -3053 607 -3019
rect 641 -3053 653 -3019
rect 595 -3059 653 -3053
rect 787 -3019 845 -3013
rect 787 -3053 799 -3019
rect 833 -3053 845 -3019
rect 787 -3059 845 -3053
rect 979 -3019 1037 -3013
rect 979 -3053 991 -3019
rect 1025 -3053 1037 -3019
rect 979 -3059 1037 -3053
<< properties >>
string FIXED_BBOX -1266 -3138 1266 3138
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 10 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
