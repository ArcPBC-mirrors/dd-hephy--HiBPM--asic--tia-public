magic
tech sky130A
magscale 1 2
timestamp 1689856338
<< metal1 >>
rect 75393 137794 83796 137870
rect 74915 135040 74925 137794
rect 75675 137786 83796 137794
rect 75675 135040 83804 137786
rect 112630 135400 112640 135620
rect 75393 134967 83804 135040
rect 80760 134596 83804 134967
rect 112580 134940 112640 135400
rect 113480 135400 113490 135620
rect 113480 134940 113520 135400
rect 44280 134400 52420 134580
rect 42910 130220 42920 134400
rect 44820 134340 52420 134400
rect 44820 130220 50040 134340
rect 44280 130160 50040 130220
rect 53060 130160 53070 134340
rect 80760 131220 83800 134596
rect 112580 131660 113520 134940
rect 44280 130100 52420 130160
rect 80760 129580 81500 131220
rect 83680 129580 83800 131220
rect 112570 130940 112580 131660
rect 113520 130940 113530 131660
rect 80760 129520 83800 129580
rect 111200 129720 116900 129760
rect 81360 129500 83780 129520
rect 111200 129040 111260 129720
rect 112140 129040 116160 129720
rect 116860 129040 116900 129720
rect 111200 129000 116900 129040
rect 52200 126200 65800 126400
rect 52200 124200 63800 126200
rect 65800 124200 65810 126200
rect 43200 122600 53800 124200
rect 43200 111000 45000 122600
rect 48090 118380 48100 121000
rect 48580 118380 55220 121000
rect 55700 118380 56420 121000
rect 43200 110200 43600 111000
rect 43590 109000 43600 110200
rect 44600 110200 45000 111000
rect 52560 116520 53760 116560
rect 52560 115960 53620 116520
rect 53880 115960 53890 116520
rect 83710 116220 83720 116560
rect 83900 116220 83910 116560
rect 44600 109000 44610 110200
rect 52560 102680 53760 115960
rect 87200 113120 87660 113140
rect 87200 112880 87220 113120
rect 87640 112880 87660 113120
rect 83960 104540 86560 107880
rect 83960 103560 84080 104540
rect 86480 103560 86560 104540
rect 83960 103460 86560 103560
rect 52560 102620 83360 102680
rect 52560 101780 81700 102620
rect 52580 101440 81700 101780
rect 83260 101440 83360 102620
rect 52580 101360 83360 101440
rect 47610 96240 47620 100660
rect 48660 96240 55080 100660
rect 56120 96240 56140 100660
rect 87200 98940 87660 112880
rect 87110 98200 87120 98940
rect 87700 98200 87710 98940
rect 63990 70200 64000 70800
rect 55200 69200 64000 70200
rect 45480 62600 54800 62680
rect 45480 62580 53600 62600
rect 45480 61460 45600 62580
rect 45480 59040 45560 61460
rect 48720 59200 53600 62580
rect 54600 59200 54800 62600
rect 48720 59100 54800 59200
rect 48700 59040 54800 59100
rect 45480 59000 54800 59040
rect 55200 58600 56400 69200
rect 63990 68800 64000 69200
rect 66000 68800 66010 70800
rect 97920 68020 99300 68380
rect 98150 63640 98160 63920
rect 98840 63640 98850 63920
rect 58990 63200 59000 63400
rect 53400 57400 56400 58600
rect 56800 63000 59000 63200
rect 59400 63000 59410 63400
rect 56800 62800 59400 63000
rect 53400 42400 55000 57400
rect 56800 57120 57200 62800
rect 98180 62360 98840 63640
rect 84320 61980 98840 62360
rect 55560 57060 57200 57120
rect 84300 61640 98840 61980
rect 113860 62100 115660 62160
rect 84300 59680 84740 61640
rect 113860 60320 113940 62100
rect 115600 60320 115660 62100
rect 84300 57080 84860 59680
rect 113860 58540 115660 60320
rect 55550 56720 55560 57060
rect 55840 56820 57200 57060
rect 55840 56720 55850 56820
rect 84400 55260 84860 57080
rect 84970 56820 84980 57420
rect 85080 56820 85090 57420
rect 113860 56760 113940 58540
rect 115600 56760 115660 58540
rect 113860 56680 115660 56760
rect 84390 54920 84400 55260
rect 84740 54920 84860 55260
rect 84400 54900 84860 54920
rect 53400 40800 66000 42400
rect 68200 40800 68210 42400
<< via1 >>
rect 74925 135040 75675 137794
rect 112640 134940 113480 135620
rect 42920 130220 44820 134400
rect 50040 130160 53060 134340
rect 81500 129580 83680 131220
rect 112580 130940 113520 131660
rect 111260 129040 112140 129720
rect 116160 129040 116860 129720
rect 63800 124200 65800 126200
rect 48100 118380 48580 121000
rect 55220 118380 55700 121000
rect 43600 109000 44600 111000
rect 53620 115960 53880 116520
rect 83720 116220 83900 116560
rect 87220 112880 87640 113120
rect 84080 103560 86480 104540
rect 81700 101440 83260 102620
rect 47620 96240 48660 100660
rect 55080 96240 56120 100660
rect 87120 98200 87700 98940
rect 45600 61460 48720 62580
rect 45560 59100 48720 61460
rect 53600 59200 54600 62600
rect 45560 59040 48700 59100
rect 64000 68800 66000 70800
rect 98160 63640 98840 63920
rect 59000 63000 59400 63400
rect 113940 60320 115600 62100
rect 55560 56720 55840 57060
rect 84980 56820 85080 57420
rect 113940 56760 115600 58540
rect 84400 54920 84740 55260
rect 66000 40800 68200 42400
<< metal2 >>
rect 46400 140200 48600 140210
rect 48600 138400 63000 140200
rect 70800 139600 71800 139610
rect 46400 138390 48600 138400
rect 57000 136600 59000 136610
rect 44280 134410 52420 134580
rect 42920 134400 52420 134410
rect 44820 134350 52420 134400
rect 44820 134340 53060 134350
rect 44820 130220 50040 134340
rect 42920 130210 50040 130220
rect 44280 130160 50040 130210
rect 44280 130150 53060 130160
rect 57000 131400 59000 135200
rect 44280 130100 52420 130150
rect 57000 129390 59000 129400
rect 61000 131400 63000 138400
rect 61000 129390 63000 129400
rect 63800 138400 70800 139600
rect 54200 128800 56200 128810
rect 63800 128800 65800 138400
rect 70800 138390 71800 138400
rect 75393 137804 83796 137870
rect 74925 137794 83796 137804
rect 75675 137786 83796 137794
rect 75675 135040 83804 137786
rect 112640 135620 113480 135630
rect 74925 135030 83804 135040
rect 75393 134967 83804 135030
rect 80760 134596 83804 134967
rect 112580 134940 112640 135400
rect 113480 134940 113520 135400
rect 80760 131220 83780 134596
rect 80760 129580 81500 131220
rect 83680 129580 83780 131220
rect 112580 131660 113520 134940
rect 112580 130930 113520 130940
rect 80760 129520 83780 129580
rect 81360 129500 83780 129520
rect 111200 129720 116900 129760
rect 111200 129040 111260 129720
rect 112140 129040 116160 129720
rect 116860 129040 116900 129720
rect 111200 129000 116900 129040
rect 56200 126800 65800 128800
rect 54200 126790 56200 126800
rect 63800 126200 65800 126210
rect 63800 124190 65800 124200
rect 61000 123400 63000 123410
rect 40600 121400 61000 123400
rect 40600 91600 43000 121400
rect 61000 121390 63000 121400
rect 48100 121000 48580 121010
rect 55220 121000 55700 121010
rect 48580 118380 55220 121000
rect 55700 118380 57780 121000
rect 48100 118370 48580 118380
rect 55220 118370 55700 118380
rect 77326 118137 78207 118145
rect 77326 118135 78264 118137
rect 78207 117698 78264 118135
rect 77326 117688 78264 117698
rect 77757 117115 78264 117688
rect 83320 116570 83860 116580
rect 83320 116560 83900 116570
rect 53620 116520 53880 116530
rect 53880 115960 54440 116520
rect 83320 116220 83340 116560
rect 83640 116220 83720 116560
rect 83320 116210 83900 116220
rect 83320 116200 83860 116210
rect 53620 115950 53880 115960
rect 85940 113120 87660 113140
rect 85940 112880 86000 113120
rect 86260 112880 87220 113120
rect 87640 112880 87660 113120
rect 85940 112860 87660 112880
rect 61700 112600 61980 112640
rect 60500 112540 61980 112600
rect 43600 111000 44600 111010
rect 43600 108990 44600 109000
rect 43620 105960 44540 105970
rect 60500 105940 61960 112540
rect 44540 104480 61980 105940
rect 83960 104540 86560 107880
rect 43620 104470 44540 104480
rect 83960 103560 84080 104540
rect 86480 103560 86560 104540
rect 83960 103460 86560 103560
rect 81700 102620 83260 102630
rect 81700 101430 83260 101440
rect 47620 100660 48660 100670
rect 55080 100660 56120 100670
rect 48660 99240 55080 100660
rect 48760 97300 55080 99240
rect 48660 96240 55080 97300
rect 56120 99280 56140 100660
rect 56120 99200 56180 99280
rect 56140 97320 56180 99200
rect 87120 98940 87700 98950
rect 87120 98190 87700 98200
rect 56120 97260 56180 97320
rect 56120 96240 56140 97260
rect 47620 96230 48660 96240
rect 55080 96230 56120 96240
rect 43000 89400 43800 91600
rect 44600 91400 48800 91600
rect 44600 89600 45800 91400
rect 48600 89600 48800 91400
rect 44600 89400 48800 89600
rect 40600 74800 43000 89400
rect 57200 74800 59200 74810
rect 40600 72800 57200 74800
rect 57200 72790 59200 72800
rect 54400 70800 56400 70810
rect 43000 70600 54400 70800
rect 44200 68800 54400 70600
rect 54400 68790 56400 68800
rect 64000 70800 66000 70810
rect 64000 68790 66000 68800
rect 43000 68590 44200 68600
rect 57200 66800 59200 66810
rect 43000 64800 57200 66800
rect 43000 42200 44800 64800
rect 57200 64790 59200 64800
rect 98160 63920 98840 63930
rect 98160 63630 98840 63640
rect 59000 63400 59400 63410
rect 59000 62990 59400 63000
rect 45480 62600 54800 62680
rect 45480 62580 53600 62600
rect 45480 61460 45600 62580
rect 45480 59040 45560 61460
rect 48720 59200 53600 62580
rect 54600 61600 54800 62600
rect 113860 62100 115660 62160
rect 54600 59200 58600 61600
rect 48720 59100 58600 59200
rect 48700 59040 58600 59100
rect 45480 59000 58600 59040
rect 113860 60320 113940 62100
rect 115600 60320 115660 62100
rect 48800 58560 58800 58600
rect 48800 57200 48860 58560
rect 49640 57200 58800 58560
rect 113860 58540 115660 60320
rect 48860 57190 49640 57200
rect 55560 57060 55840 57070
rect 55560 56710 55840 56720
rect 57800 56800 58800 57200
rect 84980 57420 85080 57430
rect 84980 56810 85080 56820
rect 57800 52480 58860 56800
rect 113860 56760 113940 58540
rect 115600 56760 115660 58540
rect 113860 56680 115660 56760
rect 84400 55260 84740 55270
rect 84400 54910 84740 54920
rect 63120 52480 63480 54380
rect 76260 53202 76720 53220
rect 57800 52180 63480 52480
rect 57800 51480 63500 52180
rect 66400 42600 70400 42610
rect 66000 42400 66400 42410
rect 75518 42400 76720 53202
rect 43000 42010 47800 42200
rect 70400 42100 76720 42400
rect 43000 42000 48400 42010
rect 43000 40800 46600 42000
rect 46600 40790 48400 40800
rect 68200 41900 76720 42100
rect 68200 40800 76724 41900
rect 66000 40790 68200 40800
<< via2 >>
rect 46400 138400 48600 140200
rect 57000 135200 59000 136600
rect 42920 130220 44820 134400
rect 50040 130160 53060 134340
rect 57000 129400 59000 131400
rect 61000 129400 63000 131400
rect 70800 138400 71800 139600
rect 74925 135040 75675 137794
rect 112640 134940 113480 135620
rect 81500 129580 83680 131220
rect 112580 130940 113520 131660
rect 111260 129040 112140 129720
rect 116160 129040 116860 129720
rect 54200 126800 56200 128800
rect 63800 124200 65800 126200
rect 61000 121400 63000 123400
rect 48100 118380 48580 121000
rect 55220 118380 55700 121000
rect 77326 117698 78207 118135
rect 83340 116220 83640 116560
rect 86000 112880 86260 113120
rect 43600 109000 44600 111000
rect 43620 104480 44540 105960
rect 84080 103560 86480 104540
rect 81700 101440 83260 102620
rect 47620 96240 48660 100660
rect 48660 97300 48760 99240
rect 55080 96240 56120 100660
rect 56120 97320 56140 99200
rect 87120 98200 87700 98940
rect 40600 89400 43000 91600
rect 45800 89600 48600 91400
rect 57200 72800 59200 74800
rect 43000 68600 44200 70600
rect 54400 68800 56400 70800
rect 64000 68800 66000 70800
rect 57200 64800 59200 66800
rect 98160 63640 98840 63920
rect 59000 63000 59400 63400
rect 45600 61460 48720 62580
rect 45560 59100 48720 61460
rect 53600 59200 54600 62600
rect 45560 59040 48700 59100
rect 113940 60320 115600 62100
rect 48860 57200 49640 58560
rect 84980 56820 85080 57420
rect 113940 56760 115600 58540
rect 84400 54920 84740 55260
rect 66400 42400 70400 42600
rect 66400 42100 68200 42400
rect 68200 42100 70400 42400
rect 46600 40800 48400 42000
<< metal3 >>
rect 44940 140600 49940 141000
rect 65940 140600 70940 141000
rect 107940 140860 112960 141020
rect 107940 140600 110700 140860
rect 46400 140205 48600 140600
rect 46390 140200 48610 140205
rect 66300 140200 70500 140600
rect 39760 137905 43540 139740
rect 46390 138400 46400 140200
rect 48600 138400 48610 140200
rect 66390 139900 70410 140200
rect 66400 139700 70400 139900
rect 66390 139100 66400 139700
rect 70100 139100 70400 139700
rect 70790 139600 71810 139605
rect 46390 138395 48610 138400
rect 70790 138400 70800 139600
rect 71800 138400 71810 139600
rect 82100 139080 86900 140600
rect 87200 139080 91860 140520
rect 92160 139760 96940 140540
rect 70790 138395 71810 138400
rect 39760 137900 48810 137905
rect 39760 134960 42360 137900
rect 48800 137880 48820 137900
rect 48800 137794 75699 137880
rect 48800 136600 74925 137794
rect 48800 135200 57000 136600
rect 59000 135200 74925 136600
rect 48800 135040 74925 135200
rect 75675 135040 75699 137794
rect 48800 134960 75699 135040
rect 42350 134955 48820 134960
rect 40080 134580 41100 134660
rect 40080 134400 45020 134580
rect 40080 130220 42920 134400
rect 44820 130220 45020 134400
rect 40080 130080 45020 130220
rect 40080 129980 41100 130080
rect 45480 129700 48820 134955
rect 76038 134460 80857 138028
rect 84200 134560 86860 139080
rect 92160 134560 96960 139760
rect 110690 139600 110700 140600
rect 112220 140600 112960 140860
rect 112220 139600 112230 140600
rect 112630 135620 113490 135625
rect 112630 134940 112640 135620
rect 113480 134940 113490 135620
rect 112630 134935 113490 134940
rect 109460 134560 115640 134580
rect 84200 134500 115640 134560
rect 84200 134460 115700 134500
rect 52840 134380 115700 134460
rect 39800 129560 48820 129700
rect 39800 124920 45720 129560
rect 48700 124920 48820 129560
rect 39800 124900 48820 124920
rect 45480 121000 48820 124900
rect 45480 118380 48100 121000
rect 48580 118380 48820 121000
rect 39460 113200 40000 113740
rect 39460 109000 41200 113200
rect 41700 109000 41710 113200
rect 43500 111000 43800 113200
rect 44300 111040 44600 113200
rect 44300 111000 44680 111040
rect 43500 109000 43600 111000
rect 44600 109000 44680 111000
rect 39460 108740 40000 109000
rect 43500 108700 44680 109000
rect 43240 105960 44680 108700
rect 43240 104480 43620 105960
rect 44540 104480 44680 105960
rect 43240 104460 44680 104480
rect 45480 100660 48820 118380
rect 49940 134360 115700 134380
rect 49940 134340 84360 134360
rect 49940 130160 50040 134340
rect 53060 134294 84360 134340
rect 53060 132725 75776 134294
rect 77030 134241 84360 134294
rect 77030 132806 79296 134241
rect 80865 132860 84360 134241
rect 86780 134340 115700 134360
rect 86780 132860 92380 134340
rect 80865 132806 92380 132860
rect 77030 132780 92380 132806
rect 96720 132780 115700 134340
rect 77030 132725 115700 132780
rect 53060 132600 115700 132725
rect 53060 130160 53280 132600
rect 84300 132060 115700 132600
rect 109420 132040 115700 132060
rect 112570 131660 113530 131665
rect 49940 123400 53280 130160
rect 56990 131400 59010 131405
rect 56990 129400 57000 131400
rect 59000 129400 59010 131400
rect 56990 129395 59010 129400
rect 60990 131400 63010 131405
rect 60990 129400 61000 131400
rect 63000 129400 63010 131400
rect 81360 131300 86320 131320
rect 81360 131220 86340 131300
rect 81360 129580 81500 131220
rect 83680 129580 86340 131220
rect 112570 130940 112580 131660
rect 113520 130940 113530 131660
rect 112570 130935 113530 130940
rect 81360 129500 86340 129580
rect 60990 129395 63010 129400
rect 54190 128800 56210 128805
rect 54190 126800 54200 128800
rect 56200 126800 56210 128800
rect 54190 126795 56210 126800
rect 63790 126200 65810 126205
rect 63790 124200 63800 126200
rect 65800 124200 65810 126200
rect 63790 124195 65810 124200
rect 81420 124860 86340 129500
rect 111250 129720 112150 129725
rect 111250 129040 111260 129720
rect 112140 129040 112150 129720
rect 111250 129035 112150 129040
rect 60990 123400 63010 123405
rect 49940 123200 57000 123400
rect 49940 121600 50000 123200
rect 53200 121600 57000 123200
rect 49940 121400 57000 121600
rect 59000 121400 59010 123400
rect 60990 121400 61000 123400
rect 63000 121400 63010 123400
rect 49940 107900 53280 121400
rect 60990 121395 63010 121400
rect 55210 121000 55710 121005
rect 55210 118380 55220 121000
rect 55700 118380 57400 121000
rect 81420 120640 86300 124860
rect 83620 120580 86300 120640
rect 113900 118660 115700 132040
rect 118000 131705 118400 134860
rect 117510 131700 118400 131705
rect 116100 130555 118400 131700
rect 116100 130540 117520 130555
rect 116100 129720 116960 130540
rect 118000 129860 118400 130555
rect 116100 129040 116160 129720
rect 116860 129040 116960 129720
rect 116100 129000 116960 129040
rect 113900 118600 118280 118660
rect 55210 118375 55710 118380
rect 77316 118135 78217 118140
rect 77316 117698 77326 118135
rect 78207 117698 78217 118135
rect 77316 117693 78217 117698
rect 81360 116740 83660 117180
rect 83300 116560 83660 116740
rect 83300 116220 83340 116560
rect 83640 116220 83660 116560
rect 83300 116160 83660 116220
rect 83330 115700 83340 116040
rect 83620 115700 83630 116040
rect 83340 114940 83620 115700
rect 82780 114420 83620 114940
rect 113900 113960 114120 118600
rect 115660 113960 118280 118600
rect 113900 113900 118280 113960
rect 85640 113125 86100 113140
rect 85640 113120 86270 113125
rect 85640 112880 86000 113120
rect 86260 112880 86270 113120
rect 85640 112875 86270 112880
rect 85640 112860 86100 112875
rect 113900 108600 115700 113900
rect 116520 108960 117900 113540
rect 113900 108580 118220 108600
rect 49940 105520 54000 107900
rect 45480 96240 47620 100660
rect 48660 99240 48820 100660
rect 48760 97300 48820 99240
rect 48660 96240 48820 97300
rect 39466 92740 40004 92744
rect 39460 91600 40004 92740
rect 40590 91600 43010 91605
rect 39460 89400 40600 91600
rect 43000 89400 43010 91600
rect 39460 87745 40004 89400
rect 40590 89395 43010 89400
rect 45480 91400 48820 96240
rect 45480 89600 45800 91400
rect 48600 89600 48820 91400
rect 39460 87740 40000 87745
rect 39460 71000 39800 71740
rect 39460 67000 41600 71000
rect 42200 67000 42210 71000
rect 43790 70605 43800 71000
rect 42990 70600 43800 70605
rect 42990 69600 43000 70600
rect 42900 68600 43000 69600
rect 42900 67000 43800 68600
rect 44400 67000 44410 71000
rect 39460 66740 39800 67000
rect 42900 66600 44400 67000
rect 42900 58560 44340 66600
rect 45480 62580 48820 89600
rect 45480 61460 45600 62580
rect 45480 59340 45560 61460
rect 45550 59040 45560 59340
rect 48720 59340 48820 62580
rect 49960 103980 54000 105520
rect 83960 107820 85940 107880
rect 83960 104540 86560 107820
rect 49960 59920 53340 103980
rect 83960 103560 84080 104540
rect 86480 104040 86560 104540
rect 86480 103740 86540 104040
rect 113900 103940 114060 108580
rect 115600 103940 118220 108580
rect 113900 103880 118220 103940
rect 103440 103740 115700 103880
rect 86480 103600 88380 103740
rect 101360 103600 115700 103740
rect 86480 103560 115700 103600
rect 83960 103460 115700 103560
rect 81660 102620 83300 102680
rect 81660 101440 81700 102620
rect 83260 101440 83300 102620
rect 84000 101640 115700 103460
rect 81660 100760 83300 101440
rect 77940 100720 81300 100740
rect 55780 100665 81320 100720
rect 55070 100660 81320 100665
rect 55010 97320 55020 100660
rect 56540 97760 81320 100660
rect 81660 99420 112400 100760
rect 87110 98940 87710 98945
rect 87110 98200 87120 98940
rect 87700 98200 87710 98940
rect 87110 98195 87710 98200
rect 56540 97320 56550 97760
rect 55070 96240 55080 97320
rect 56120 97315 56150 97320
rect 56120 96240 56130 97315
rect 55070 96235 56130 96240
rect 77940 92840 81300 97760
rect 77940 92760 100340 92840
rect 77940 89940 86000 92760
rect 87520 92660 100340 92760
rect 87520 90200 98460 92660
rect 100060 90200 100340 92660
rect 87520 89940 100340 90200
rect 77940 89880 81300 89940
rect 70200 75580 70500 78840
rect 70200 75220 85100 75580
rect 57190 74800 59210 74805
rect 57190 72800 57200 74800
rect 59200 72800 59210 74800
rect 57190 72795 59210 72800
rect 66270 71280 66280 71880
rect 66720 71280 66730 71880
rect 83340 71840 83980 71880
rect 83340 71320 83380 71840
rect 83960 71320 83980 71840
rect 54390 70800 56410 70805
rect 54390 68800 54400 70800
rect 56400 68800 56410 70800
rect 54390 68795 56410 68800
rect 63990 70800 66010 70805
rect 63990 68800 64000 70800
rect 66000 68800 66010 70800
rect 63990 68795 66010 68800
rect 57190 66800 59210 66805
rect 57190 64800 57200 66800
rect 59200 64800 59210 66800
rect 57190 64795 59210 64800
rect 66280 63440 66720 71280
rect 59000 63405 66740 63440
rect 58990 63400 66740 63405
rect 58990 63000 59000 63400
rect 59400 63040 66740 63400
rect 59400 63000 59410 63040
rect 58990 62995 59410 63000
rect 83340 62680 83980 71320
rect 84720 67000 85100 75220
rect 97520 71960 98840 72040
rect 97520 71260 97620 71960
rect 98740 71260 98840 71960
rect 97520 71200 98840 71260
rect 97550 67760 97560 67860
rect 97500 67120 97560 67760
rect 97920 67760 97930 67860
rect 97920 67120 98020 67760
rect 97500 62680 98020 67120
rect 98160 63925 98840 71200
rect 111400 67920 112380 99420
rect 113900 95220 115700 101640
rect 113890 92560 113900 95220
rect 115640 92560 115700 95220
rect 111390 67020 111400 67920
rect 111880 67020 112380 67920
rect 111400 67000 112380 67020
rect 112660 91660 113860 91680
rect 118020 91660 118380 92860
rect 112660 90480 118380 91660
rect 98150 63920 98850 63925
rect 98150 63640 98160 63920
rect 98840 63640 98850 63920
rect 112660 63780 113860 90480
rect 98150 63635 98850 63640
rect 111760 63720 113860 63780
rect 111760 62860 111780 63720
rect 112720 62860 113860 63720
rect 111760 62800 113860 62860
rect 114420 76680 115620 90080
rect 118020 87860 118380 90480
rect 114420 71920 114440 76680
rect 115580 71920 118260 76680
rect 114420 71900 118260 71920
rect 114420 66640 115620 71900
rect 116480 66940 117900 71580
rect 114420 66560 118260 66640
rect 53590 62600 54610 62605
rect 48720 59100 48730 59340
rect 48700 59095 48730 59100
rect 48700 59040 48710 59095
rect 45550 59035 48710 59040
rect 48850 58560 49650 58565
rect 42900 57220 48860 58560
rect 43120 57200 48860 57220
rect 49640 57200 49650 58560
rect 48850 57195 49650 57200
rect 49960 55940 53360 59920
rect 53590 59200 53600 62600
rect 54600 60000 60200 62600
rect 83340 62300 98020 62680
rect 83340 62200 89980 62300
rect 114420 62200 114540 66560
rect 113860 62100 114540 62200
rect 115540 62100 118260 66560
rect 66570 60160 66580 61360
rect 69220 60160 69230 61360
rect 84950 61100 89980 61320
rect 84950 60740 88400 61100
rect 89300 60740 89980 61100
rect 54600 59200 54610 60000
rect 80410 59880 80420 60680
rect 82780 59880 82790 60680
rect 113860 60320 113940 62100
rect 115600 61860 118260 62100
rect 115600 61560 115700 61860
rect 115600 60320 115660 61560
rect 53590 59195 54610 59200
rect 112140 58680 113620 58740
rect 112140 57920 112200 58680
rect 113540 57920 113620 58680
rect 82840 57420 84760 57780
rect 84970 57420 85090 57425
rect 82840 57340 84980 57420
rect 84460 57020 84980 57340
rect 84970 56820 84980 57020
rect 85080 56820 85090 57420
rect 84970 56815 85090 56820
rect 49960 55740 53340 55940
rect 39700 55480 53340 55740
rect 39700 51280 50140 55480
rect 52920 51280 53340 55480
rect 84390 55260 84750 55265
rect 84390 54920 84400 55260
rect 84740 54920 84750 55260
rect 84390 54915 84750 54920
rect 86810 53520 86820 53700
rect 87200 53520 87210 53700
rect 39700 50960 53340 51280
rect 40540 50940 53340 50960
rect 41460 50640 48860 50660
rect 40060 50500 48860 50640
rect 40060 46180 45580 50500
rect 48780 46180 48860 50500
rect 40060 46020 48860 46180
rect 49960 47800 53340 50940
rect 112140 53420 113620 57920
rect 113860 58540 115660 60320
rect 113860 56760 113940 58540
rect 115600 56760 115660 58540
rect 113860 53780 115660 56760
rect 116300 59780 117520 59840
rect 116300 59020 116400 59780
rect 117460 59020 117520 59780
rect 49960 47400 61100 47800
rect 63680 47400 74440 47800
rect 49960 47380 74440 47400
rect 77060 47380 85640 47800
rect 40060 46000 41500 46020
rect 39700 45680 41480 45700
rect 49960 45680 85640 47380
rect 39700 45600 85640 45680
rect 39700 42500 50300 45600
rect 52660 44240 85640 45600
rect 103940 44280 111980 44320
rect 103940 44240 111240 44280
rect 52660 44140 111240 44240
rect 52660 42900 82060 44140
rect 52660 42500 65900 42900
rect 71000 42760 82060 42900
rect 86780 42760 92140 44140
rect 96860 42760 111240 44140
rect 39700 42380 65900 42500
rect 66390 42600 70410 42605
rect 39700 40900 41480 42380
rect 66390 42100 66400 42600
rect 70400 42100 70410 42600
rect 71000 42400 111240 42760
rect 111960 42400 111980 44280
rect 71000 42380 111980 42400
rect 66390 42095 70410 42100
rect 46590 42000 48410 42005
rect 46590 40800 46600 42000
rect 48400 40800 48410 42000
rect 46590 40795 48410 40800
rect 46600 40000 48400 40795
rect 66390 40300 66400 40700
rect 70400 40300 70410 40700
rect 66590 40000 70610 40300
rect 45060 39600 50080 40000
rect 66040 39600 71060 40000
rect 82040 39720 86820 42380
rect 87140 40060 91780 41480
rect 92100 39720 96880 42380
rect 112140 41940 113600 53420
rect 113860 50780 115700 53780
rect 113860 48020 115720 50780
rect 116300 50060 117520 59020
rect 118000 50060 118400 50860
rect 116300 48780 118400 50060
rect 113860 44320 115700 48020
rect 118000 45880 118400 48780
rect 113720 44300 115700 44320
rect 113720 42420 113760 44300
rect 114480 42960 115700 44300
rect 114480 42420 115620 42960
rect 113720 42380 115620 42420
rect 110380 40460 113600 41940
rect 110380 40000 112160 40460
rect 108060 39580 113060 40000
<< via3 >>
rect 66400 139100 70100 139700
rect 70800 138400 71800 139600
rect 42360 134960 48800 137900
rect 74925 135040 75675 137794
rect 42920 130220 44820 134400
rect 110700 139600 112220 140860
rect 112640 134940 113480 135620
rect 45720 124920 48700 129560
rect 48100 118380 48580 121000
rect 41200 109000 41700 113200
rect 43800 111000 44300 113200
rect 43800 109000 44300 111000
rect 50040 130160 53060 134340
rect 75776 132725 77030 134294
rect 79296 132806 80865 134241
rect 84360 132860 86780 134360
rect 92380 132780 96720 134340
rect 57000 129400 59000 131400
rect 61000 129400 63000 131400
rect 81500 129580 83680 131220
rect 112580 130940 113520 131660
rect 54200 126800 56200 128800
rect 63800 124200 65800 126200
rect 111260 129040 112140 129720
rect 50000 121600 53200 123200
rect 57000 121400 59000 123400
rect 61000 121400 63000 123400
rect 77326 117698 78207 118135
rect 83340 115700 83620 116040
rect 114120 113960 115660 118600
rect 47620 99240 48660 100660
rect 47620 97300 48760 99240
rect 47620 96240 48660 97300
rect 45800 89600 48600 91400
rect 41600 67000 42200 71000
rect 43800 70600 44400 71000
rect 43800 68600 44200 70600
rect 44200 68600 44400 70600
rect 43800 67000 44400 68600
rect 45600 61460 48720 62580
rect 45560 59100 48720 61460
rect 84080 103560 86480 104540
rect 114060 103940 115600 108580
rect 55020 97320 55080 100660
rect 55080 99200 56120 100660
rect 56120 99200 56540 100660
rect 55080 97320 56140 99200
rect 56140 97320 56540 99200
rect 87120 98200 87700 98940
rect 55080 96240 56120 97320
rect 86000 89940 87520 92760
rect 98460 90200 100060 92660
rect 57200 72800 59200 74800
rect 66280 71280 66720 71880
rect 83380 71320 83960 71840
rect 54400 68800 56400 70800
rect 64000 68800 66000 70800
rect 57200 64800 59200 66800
rect 97620 71260 98740 71960
rect 97560 67120 97920 67860
rect 113900 92560 115640 95220
rect 111400 67020 111880 67920
rect 111780 62860 112720 63720
rect 114440 71920 115580 76680
rect 45560 59040 48700 59100
rect 53600 59200 54600 62600
rect 114540 62100 115540 66560
rect 66580 60160 69220 61360
rect 80420 59880 82780 60680
rect 113940 60320 115600 62100
rect 112200 57920 113540 58680
rect 50140 51280 52920 55480
rect 84400 54920 84740 55260
rect 86820 53520 87200 53700
rect 45580 46180 48780 50500
rect 113940 56760 115600 58540
rect 116400 59020 117460 59780
rect 50300 42500 52660 45600
rect 82060 42760 86780 44140
rect 92140 42760 96860 44140
rect 66400 42100 70400 42600
rect 111240 42400 111960 44280
rect 66400 40300 70400 40700
rect 113760 42420 114480 44300
<< metal4 >>
rect 110699 140860 112221 140861
rect 66399 139700 70101 139701
rect 66399 139100 66400 139700
rect 70100 139100 70101 139700
rect 70799 139600 71801 139601
rect 66399 139099 70101 139100
rect 70600 138400 70800 139600
rect 71800 139571 71801 139600
rect 110699 139600 110700 140860
rect 112220 139600 112221 140860
rect 110699 139599 112221 139600
rect 71800 138488 78661 139571
rect 71800 138400 71801 138488
rect 70600 138399 71801 138400
rect 70600 138300 71700 138399
rect 42359 137900 48801 137901
rect 42359 134960 42360 137900
rect 48800 137880 48820 137900
rect 48800 137200 66000 137880
rect 66500 137400 71700 138300
rect 72100 137794 75699 137880
rect 72100 137200 74925 137794
rect 48800 135040 74925 137200
rect 75675 135040 75699 137794
rect 48800 134960 75699 135040
rect 42359 134959 48820 134960
rect 42919 134400 44821 134401
rect 42919 130220 42920 134400
rect 44820 130220 44821 134400
rect 42919 130219 44821 130220
rect 45480 129560 48820 134959
rect 77433 134572 78655 138488
rect 110740 135660 112160 139599
rect 110740 135620 113520 135660
rect 110740 134940 112640 135620
rect 113480 134940 113520 135620
rect 110740 134860 113520 134940
rect 49900 134340 77182 134480
rect 49900 132040 50040 134340
rect 45480 124920 45720 129560
rect 48700 124920 48820 129560
rect 45480 121000 48820 124920
rect 45480 118380 48100 121000
rect 48580 118380 48820 121000
rect 41199 113200 41701 113201
rect 43799 113200 44301 113201
rect 41199 109000 41200 113200
rect 41700 109000 41900 113200
rect 43500 109000 43800 113200
rect 44300 109000 44301 113200
rect 41199 108999 41701 109000
rect 43799 108999 44301 109000
rect 45480 100660 48820 118380
rect 49940 130160 50040 132040
rect 53060 134294 77182 134340
rect 53060 132725 75776 134294
rect 77030 132725 77182 134294
rect 53060 132500 77182 132725
rect 53060 132040 65500 132500
rect 69000 132040 77182 132500
rect 53060 130160 53280 132040
rect 77435 131708 78647 134572
rect 109460 134560 115640 134580
rect 84300 134480 115640 134560
rect 79100 134360 115640 134480
rect 79100 134241 84360 134360
rect 79100 132806 79296 134241
rect 80865 132860 84360 134241
rect 86780 134340 115640 134360
rect 86780 132860 92380 134340
rect 80865 132806 92380 132860
rect 79100 132780 92380 132806
rect 96720 132780 115640 134340
rect 79100 132040 115640 132780
rect 77431 131551 78647 131708
rect 112520 131660 113600 131740
rect 49940 123200 53280 130160
rect 56999 131400 59001 131401
rect 56999 129400 57000 131400
rect 59000 129400 59001 131400
rect 56999 129399 59001 129400
rect 60999 131400 63001 131401
rect 60999 129400 61000 131400
rect 63000 129400 63001 131400
rect 60999 129399 63001 129400
rect 54199 128800 56201 128801
rect 54199 126800 54200 128800
rect 56200 126800 56201 128800
rect 54199 126799 56201 126800
rect 63799 126200 65801 126201
rect 63799 124200 63800 126200
rect 65800 124200 65801 126200
rect 63799 124199 65801 124200
rect 49940 121600 50000 123200
rect 53200 121600 53280 123200
rect 49940 107900 53280 121600
rect 56999 123400 59001 123401
rect 56999 121400 57000 123400
rect 59000 121400 59001 123400
rect 56999 121399 59001 121400
rect 60999 123400 63001 123401
rect 60999 121400 61000 123400
rect 63000 121400 63001 123400
rect 60999 121399 63001 121400
rect 77431 118136 78633 131551
rect 81360 131300 86320 131320
rect 81360 131220 86340 131300
rect 81360 129580 81500 131220
rect 83680 129580 86340 131220
rect 112520 130940 112580 131660
rect 113520 130940 113600 131660
rect 81360 129500 86340 129580
rect 81420 124860 86340 129500
rect 111220 129720 112200 129740
rect 111220 129040 111260 129720
rect 112140 129040 112200 129720
rect 81420 120640 86300 124860
rect 83620 120580 86300 120640
rect 111220 119220 112200 129040
rect 100360 118320 112200 119220
rect 77325 118135 78633 118136
rect 77325 117698 77326 118135
rect 78207 117931 78633 118135
rect 112520 118120 113600 130940
rect 78207 117698 78208 117931
rect 77325 117697 78208 117698
rect 100340 117220 113600 118120
rect 113860 118601 115640 132040
rect 113860 118600 115661 118601
rect 81580 116320 81980 116620
rect 83339 116040 83621 116041
rect 86560 116040 87300 116060
rect 83300 115700 83340 116040
rect 83620 115860 87300 116040
rect 83620 115700 86620 115860
rect 83339 115699 83621 115700
rect 113860 113960 114120 118600
rect 115660 113960 115661 118600
rect 113860 113959 115661 113960
rect 113860 108580 115640 113959
rect 49940 107880 54000 107900
rect 49940 106520 57060 107880
rect 82280 106520 86220 107400
rect 49940 105520 86540 106520
rect 45480 96240 47620 100660
rect 48660 99240 48820 100660
rect 48760 97300 48820 99240
rect 48660 96240 48820 97300
rect 45480 91400 48820 96240
rect 45480 89600 45800 91400
rect 48600 89600 48820 91400
rect 41599 71000 42201 71001
rect 41599 67000 41600 71000
rect 42200 67000 42201 71000
rect 41599 66999 42201 67000
rect 43799 71000 44401 71001
rect 43799 67000 43800 71000
rect 44400 67000 44401 71000
rect 43799 66999 44401 67000
rect 45480 64280 48820 89600
rect 49960 104540 86540 105520
rect 49960 103560 84080 104540
rect 86480 103740 86540 104540
rect 103440 103880 109360 104840
rect 113860 103940 114060 108580
rect 115600 103940 115640 108580
rect 113860 103880 115640 103940
rect 103440 103740 115640 103880
rect 86480 103600 88380 103740
rect 101360 103600 115640 103740
rect 86480 103560 115640 103600
rect 49960 103480 115640 103560
rect 49960 78820 53340 103480
rect 84060 101660 115640 103480
rect 84340 101640 115640 101660
rect 77940 100720 81300 100740
rect 55780 100661 81320 100720
rect 55019 100660 81320 100661
rect 55019 97320 55020 100660
rect 56540 97760 81320 100660
rect 87080 98940 111820 99000
rect 87080 98200 87120 98940
rect 87700 98200 111820 98940
rect 87080 98120 111820 98200
rect 56540 97320 56541 97760
rect 55019 97319 55080 97320
rect 55079 96240 55080 97319
rect 56120 97319 56541 97320
rect 56120 96240 56121 97319
rect 75680 97280 81320 97760
rect 55079 96239 56121 96240
rect 77940 92820 81320 97280
rect 77940 92760 100340 92820
rect 77940 89940 86000 92760
rect 87520 92660 100340 92760
rect 87520 90200 98460 92660
rect 100060 90200 100340 92660
rect 87520 89940 100340 90200
rect 77940 89880 81300 89940
rect 85260 89939 87521 89940
rect 85260 85240 86440 89939
rect 99060 86460 100340 89940
rect 110980 83660 111820 98120
rect 113860 95221 115640 101640
rect 113860 95220 115641 95221
rect 113860 92560 113900 95220
rect 115640 92560 115641 95220
rect 113860 92559 115641 92560
rect 49960 75800 56440 78820
rect 49960 74400 53340 75800
rect 57199 74800 59201 74801
rect 49960 73300 52900 74400
rect 57199 74000 57200 74800
rect 56000 73600 57200 74000
rect 49960 67300 53340 73300
rect 57199 72800 57200 73600
rect 59200 72800 59201 74800
rect 61200 74000 63200 77400
rect 113860 76680 115640 92559
rect 61200 73600 64600 74000
rect 61200 72800 63200 73600
rect 57199 72799 59201 72800
rect 97520 71960 98840 72040
rect 66279 71880 66721 71881
rect 66279 71280 66280 71880
rect 66720 71840 84000 71880
rect 66720 71320 83380 71840
rect 83960 71320 84000 71840
rect 66720 71280 84000 71320
rect 66279 71279 66721 71280
rect 97520 71260 97620 71960
rect 98740 71260 98840 71960
rect 97520 71200 98840 71260
rect 113860 71920 114440 76680
rect 115580 71920 115640 76680
rect 54399 70800 56401 70801
rect 54399 68800 54400 70800
rect 56400 68800 56401 70800
rect 54399 68799 56401 68800
rect 63999 70800 66001 70801
rect 63999 68800 64000 70800
rect 66000 68800 66001 70800
rect 63999 68799 66001 68800
rect 66940 68160 83340 70300
rect 45480 62580 48840 64280
rect 45480 61460 45600 62580
rect 45480 59040 45560 61460
rect 48720 59100 48840 62580
rect 48700 59040 48840 59100
rect 45480 50500 48840 59040
rect 45480 46660 45580 50500
rect 45579 46180 45580 46660
rect 48780 46660 48840 50500
rect 49960 63300 52000 67300
rect 57199 66800 59201 66801
rect 57199 66000 57200 66800
rect 56400 65600 57200 66000
rect 57199 64800 57200 65600
rect 59200 64800 59201 66800
rect 57199 64799 59201 64800
rect 61200 66000 63200 66800
rect 66960 66400 69240 68160
rect 61200 65600 64400 66000
rect 49960 55480 53340 63300
rect 61200 62680 63200 65600
rect 67500 65300 69240 66400
rect 66960 62680 69240 65300
rect 53599 62600 54601 62601
rect 59000 62600 69260 62680
rect 53599 59200 53600 62600
rect 54600 61360 69260 62600
rect 54600 60160 66580 61360
rect 69220 60160 69260 61360
rect 54600 60080 69260 60160
rect 80180 62160 83340 68160
rect 111399 67920 111881 67921
rect 97559 67860 97921 67861
rect 97559 67120 97560 67860
rect 97920 67120 97921 67860
rect 97559 67119 97921 67120
rect 111399 67020 111400 67920
rect 111880 67020 111881 67920
rect 111399 67019 111881 67020
rect 113860 66560 115640 71920
rect 111340 63720 112740 63780
rect 111340 62860 111780 63720
rect 112720 62860 112740 63720
rect 111340 62800 112740 62860
rect 80180 60680 86500 62160
rect 54600 60000 60200 60080
rect 54600 59200 54601 60000
rect 80180 59900 80420 60680
rect 80419 59880 80420 59900
rect 82780 59900 86500 60680
rect 113860 62100 114540 66560
rect 115540 62100 115640 66560
rect 113860 60320 113940 62100
rect 115600 61780 115640 62100
rect 115600 60320 115660 61780
rect 113860 60200 115660 60320
rect 82780 59880 82781 59900
rect 80419 59879 82781 59880
rect 53599 59199 54601 59200
rect 101760 59780 117540 59840
rect 101760 59020 116400 59780
rect 117460 59020 117540 59780
rect 101760 58940 117540 59020
rect 101740 58680 113620 58740
rect 101740 57920 112200 58680
rect 113540 57920 113620 58680
rect 101740 57840 113620 57920
rect 113860 58540 115660 58640
rect 82980 56920 83380 57220
rect 113860 56760 113940 58540
rect 115600 56760 115660 58540
rect 87740 56540 88140 56640
rect 87740 56480 87860 56540
rect 84460 56340 87860 56480
rect 84460 55940 84780 56340
rect 83340 55680 84780 55940
rect 49960 51280 50140 55480
rect 52920 51280 53340 55480
rect 84399 55260 84741 55261
rect 84399 54920 84400 55260
rect 84740 54920 87160 55260
rect 84399 54919 84741 54920
rect 86780 53701 87160 54920
rect 86780 53700 87201 53701
rect 86780 53520 86820 53700
rect 87200 53520 87201 53700
rect 86780 53519 87201 53520
rect 86780 53480 87160 53519
rect 49960 47800 53340 51280
rect 113860 52320 115660 56760
rect 48780 46180 48781 46660
rect 45579 46179 48781 46180
rect 49960 45600 85640 47800
rect 49960 44320 50300 45600
rect 49900 42500 50300 44320
rect 52660 44240 85640 45600
rect 103960 44320 107720 45420
rect 113860 44320 115640 52320
rect 103940 44300 115640 44320
rect 103940 44280 113760 44300
rect 103940 44240 111240 44280
rect 52660 44140 111240 44240
rect 52660 43500 82060 44140
rect 52660 42500 65900 43500
rect 66400 42601 70400 43100
rect 71000 42760 82060 43500
rect 86780 42760 92140 44140
rect 96860 42760 111240 44140
rect 49900 42380 65900 42500
rect 66399 42600 70401 42601
rect 66399 42100 66400 42600
rect 70400 42100 70401 42600
rect 71000 42400 111240 42760
rect 111960 42420 113760 44280
rect 114480 42820 115640 44300
rect 114480 42420 115620 42820
rect 111960 42400 115620 42420
rect 71000 42380 115620 42400
rect 66399 42099 70401 42100
rect 66400 40701 70400 41600
rect 66399 40700 70401 40701
rect 66399 40300 66400 40700
rect 70400 40300 70401 40700
rect 66399 40299 70401 40300
use bias2_top  bias2_top_1 ~/code/hibpm-sky130a-tapeout/mag/bias
timestamp 1686510802
transform 1 0 85160 0 1 67000
box -160 -4200 12860 21010
use bias2_top_s  bias2_top_s_0 ~/code/hibpm-sky130a-tapeout/mag/bias
timestamp 1686327621
transform 1 0 98960 0 1 67000
box 40 -4200 12860 21010
use exp  exp_0 ~/code/hibpm-sky130a-tapeout/mag/experiment
timestamp 1689606798
transform 1 0 55624 0 1 69024
box -3224 -5024 11624 5824
use exp  exp_2
timestamp 1689606798
transform -1 0 65324 0 -1 127224
box -3224 -5024 11624 5824
use isource  isource_0 ~/code/hibpm-sky130a-tapeout/mag/isource
timestamp 1684166381
transform 1 0 55308 0 1 81700
box -308 -5900 23140 17576
use outd_50ohm_lg  outd_50ohm_lg_0 ~/code/hibpm-sky130a-tapeout/mag/outd_50Ohm
timestamp 1689672086
transform 1 0 94122 0 1 112460
box -10522 -7820 11472 8920
use outd_50ohm_lg  outd_50ohm_lg_1
timestamp 1689672086
transform 1 0 95322 0 1 53080
box -10522 -7820 11472 8920
use rm5  rm5_0
timestamp 1689607358
transform 0 -1 64724 1 0 144624
box -7224 -5724 -5376 -1676
use rm5  rm5_1
timestamp 1689607358
transform 0 1 72124 -1 0 35924
box -7224 -5724 -5376 -1676
use rm5  rm5_2
timestamp 1689607358
transform -1 0 36424 0 -1 107324
box -7224 -5724 -5376 -1676
use rm5  rm5_3
timestamp 1689607358
transform -1 0 36624 0 -1 65324
box -7224 -5724 -5376 -1676
use tia_top  tia_top_0 ~/code/hibpm-sky130a-tapeout/mag/tiaA
timestamp 1686667164
transform 1 0 58628 0 1 48680
box -3628 -4080 25704 24280
use tia_top  tia_top_1
timestamp 1686667164
transform 1 0 57228 0 1 108080
box -3628 -4080 25704 24280
<< labels >>
rlabel metal3 82360 139420 86740 140300 1 VSS
rlabel metal3 92400 139480 96780 140360 1 VSS
rlabel metal3 87460 139340 91400 140220 1 VDD
rlabel metal3 39940 135300 40880 139420 1 VDD
port 6 n
rlabel metal3 39980 125180 40920 129300 1 VDD
rlabel metal3 40240 130240 40980 134400 1 VSS
rlabel metal3 39860 51380 41320 55540 1 VSS
rlabel metal3 39920 41200 41380 45360 1 VSS
port 3 n
rlabel metal3 40280 46220 41280 50300 1 VDD
rlabel metal3 82160 39820 86760 41400 1 VSS
rlabel metal3 87260 40140 91660 41400 1 VDD
rlabel space 92520 39960 96920 41220 1 VSS
rlabel metal3 116580 61940 118060 66460 1 VSS
rlabel metal3 116620 71980 118100 76500 1 VSS
rlabel metal3 116620 67060 117740 71400 1 VDD
rlabel metal3 116540 103960 118160 108440 1 VSS
rlabel metal3 116540 108960 117800 113420 1 VDD
rlabel metal3 116620 114020 118040 118560 1 VSS
rlabel metal3 116820 90600 117840 91480 1 I_ref_out
port 1 n
rlabel metal3 118060 131800 118320 134460 1 Out_P2
port 8 n
rlabel metal3 108060 140680 110640 140940 1 Out_N2
port 9 n
rlabel metal3 118060 47560 118320 49780 1 Out_P1
port 10 n
rlabel metal3 108320 39660 112900 39920 1 Out_N1
port 11 n
rlabel metal3 80940 75300 81520 75500 1 is_out
rlabel metal3 39546 67644 40087 68765 1 In_ref1
port 4 n
rlabel metal3 67078 39687 68793 39957 1 In1
port 12 n
rlabel metal3 68074 140487 68814 140887 1 In2
port 13 n
rlabel metal3 98320 65720 98600 66080 1 bias_outd_1
rlabel metal3 111680 68620 111960 68980 1 bias_tia_2
rlabel metal4 111040 88340 111320 88700 1 bias_outd_2
rlabel metal4 64200 69000 65800 70600 1 Ex1_In
port 16 n
rlabel metal4 54600 69000 56200 70600 1 Ex1_InRef
port 15 n
rlabel metal3 39600 110000 40000 112400 1 In_ref2
port 17 n
rlabel space 64000 125600 65600 126600 1 Ex2_InRef
rlabel space 54400 126600 56000 127600 1 Ex2_In
rlabel metal3 39568 90222 40132 91116 1 Ex_com
port 18 n
rlabel metal3 47100 39950 47836 40384 1 Ex_in2
port 19 n
rlabel metal3 46926 140356 47662 140790 1 Ex_in1
port 20 n
<< end >>
