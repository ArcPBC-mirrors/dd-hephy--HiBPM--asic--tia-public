magic
tech sky130A
magscale 1 2
timestamp 1685105324
<< pwell >>
rect -2008 -1882 2008 1882
<< psubdiff >>
rect -1972 1812 -1876 1846
rect 1876 1812 1972 1846
rect -1972 1750 -1938 1812
rect 1938 1750 1972 1812
rect -1972 -1812 -1938 -1750
rect 1938 -1812 1972 -1750
rect -1972 -1846 -1876 -1812
rect 1876 -1846 1972 -1812
<< psubdiffcont >>
rect -1876 1812 1876 1846
rect -1972 -1750 -1938 1750
rect 1938 -1750 1972 1750
rect -1876 -1846 1876 -1812
<< xpolycontact >>
rect -1842 1284 -1560 1716
rect -1842 52 -1560 484
rect -1464 1284 -1182 1716
rect -1464 52 -1182 484
rect -1086 1284 -804 1716
rect -1086 52 -804 484
rect -708 1284 -426 1716
rect -708 52 -426 484
rect -330 1284 -48 1716
rect -330 52 -48 484
rect 48 1284 330 1716
rect 48 52 330 484
rect 426 1284 708 1716
rect 426 52 708 484
rect 804 1284 1086 1716
rect 804 52 1086 484
rect 1182 1284 1464 1716
rect 1182 52 1464 484
rect 1560 1284 1842 1716
rect 1560 52 1842 484
rect -1842 -484 -1560 -52
rect -1842 -1716 -1560 -1284
rect -1464 -484 -1182 -52
rect -1464 -1716 -1182 -1284
rect -1086 -484 -804 -52
rect -1086 -1716 -804 -1284
rect -708 -484 -426 -52
rect -708 -1716 -426 -1284
rect -330 -484 -48 -52
rect -330 -1716 -48 -1284
rect 48 -484 330 -52
rect 48 -1716 330 -1284
rect 426 -484 708 -52
rect 426 -1716 708 -1284
rect 804 -484 1086 -52
rect 804 -1716 1086 -1284
rect 1182 -484 1464 -52
rect 1182 -1716 1464 -1284
rect 1560 -484 1842 -52
rect 1560 -1716 1842 -1284
<< ppolyres >>
rect -1842 484 -1560 1284
rect -1464 484 -1182 1284
rect -1086 484 -804 1284
rect -708 484 -426 1284
rect -330 484 -48 1284
rect 48 484 330 1284
rect 426 484 708 1284
rect 804 484 1086 1284
rect 1182 484 1464 1284
rect 1560 484 1842 1284
rect -1842 -1284 -1560 -484
rect -1464 -1284 -1182 -484
rect -1086 -1284 -804 -484
rect -708 -1284 -426 -484
rect -330 -1284 -48 -484
rect 48 -1284 330 -484
rect 426 -1284 708 -484
rect 804 -1284 1086 -484
rect 1182 -1284 1464 -484
rect 1560 -1284 1842 -484
<< locali >>
rect -1972 1812 -1876 1846
rect 1876 1812 1972 1846
rect -1972 1750 -1938 1812
rect 1938 1750 1972 1812
rect -1972 -1812 -1938 -1750
rect 1938 -1812 1972 -1750
rect -1972 -1846 -1876 -1812
rect 1876 -1846 1972 -1812
<< viali >>
rect -1826 1301 -1576 1698
rect -1448 1301 -1198 1698
rect -1070 1301 -820 1698
rect -692 1301 -442 1698
rect -314 1301 -64 1698
rect 64 1301 314 1698
rect 442 1301 692 1698
rect 820 1301 1070 1698
rect 1198 1301 1448 1698
rect 1576 1301 1826 1698
rect -1826 70 -1576 467
rect -1448 70 -1198 467
rect -1070 70 -820 467
rect -692 70 -442 467
rect -314 70 -64 467
rect 64 70 314 467
rect 442 70 692 467
rect 820 70 1070 467
rect 1198 70 1448 467
rect 1576 70 1826 467
rect -1826 -467 -1576 -70
rect -1448 -467 -1198 -70
rect -1070 -467 -820 -70
rect -692 -467 -442 -70
rect -314 -467 -64 -70
rect 64 -467 314 -70
rect 442 -467 692 -70
rect 820 -467 1070 -70
rect 1198 -467 1448 -70
rect 1576 -467 1826 -70
rect -1826 -1698 -1576 -1301
rect -1448 -1698 -1198 -1301
rect -1070 -1698 -820 -1301
rect -692 -1698 -442 -1301
rect -314 -1698 -64 -1301
rect 64 -1698 314 -1301
rect 442 -1698 692 -1301
rect 820 -1698 1070 -1301
rect 1198 -1698 1448 -1301
rect 1576 -1698 1826 -1301
<< metal1 >>
rect -1832 1698 -1570 1710
rect -1832 1301 -1826 1698
rect -1576 1301 -1570 1698
rect -1832 1289 -1570 1301
rect -1454 1698 -1192 1710
rect -1454 1301 -1448 1698
rect -1198 1301 -1192 1698
rect -1454 1289 -1192 1301
rect -1076 1698 -814 1710
rect -1076 1301 -1070 1698
rect -820 1301 -814 1698
rect -1076 1289 -814 1301
rect -698 1698 -436 1710
rect -698 1301 -692 1698
rect -442 1301 -436 1698
rect -698 1289 -436 1301
rect -320 1698 -58 1710
rect -320 1301 -314 1698
rect -64 1301 -58 1698
rect -320 1289 -58 1301
rect 58 1698 320 1710
rect 58 1301 64 1698
rect 314 1301 320 1698
rect 58 1289 320 1301
rect 436 1698 698 1710
rect 436 1301 442 1698
rect 692 1301 698 1698
rect 436 1289 698 1301
rect 814 1698 1076 1710
rect 814 1301 820 1698
rect 1070 1301 1076 1698
rect 814 1289 1076 1301
rect 1192 1698 1454 1710
rect 1192 1301 1198 1698
rect 1448 1301 1454 1698
rect 1192 1289 1454 1301
rect 1570 1698 1832 1710
rect 1570 1301 1576 1698
rect 1826 1301 1832 1698
rect 1570 1289 1832 1301
rect -1832 467 -1570 479
rect -1832 70 -1826 467
rect -1576 70 -1570 467
rect -1832 58 -1570 70
rect -1454 467 -1192 479
rect -1454 70 -1448 467
rect -1198 70 -1192 467
rect -1454 58 -1192 70
rect -1076 467 -814 479
rect -1076 70 -1070 467
rect -820 70 -814 467
rect -1076 58 -814 70
rect -698 467 -436 479
rect -698 70 -692 467
rect -442 70 -436 467
rect -698 58 -436 70
rect -320 467 -58 479
rect -320 70 -314 467
rect -64 70 -58 467
rect -320 58 -58 70
rect 58 467 320 479
rect 58 70 64 467
rect 314 70 320 467
rect 58 58 320 70
rect 436 467 698 479
rect 436 70 442 467
rect 692 70 698 467
rect 436 58 698 70
rect 814 467 1076 479
rect 814 70 820 467
rect 1070 70 1076 467
rect 814 58 1076 70
rect 1192 467 1454 479
rect 1192 70 1198 467
rect 1448 70 1454 467
rect 1192 58 1454 70
rect 1570 467 1832 479
rect 1570 70 1576 467
rect 1826 70 1832 467
rect 1570 58 1832 70
rect -1832 -70 -1570 -58
rect -1832 -467 -1826 -70
rect -1576 -467 -1570 -70
rect -1832 -479 -1570 -467
rect -1454 -70 -1192 -58
rect -1454 -467 -1448 -70
rect -1198 -467 -1192 -70
rect -1454 -479 -1192 -467
rect -1076 -70 -814 -58
rect -1076 -467 -1070 -70
rect -820 -467 -814 -70
rect -1076 -479 -814 -467
rect -698 -70 -436 -58
rect -698 -467 -692 -70
rect -442 -467 -436 -70
rect -698 -479 -436 -467
rect -320 -70 -58 -58
rect -320 -467 -314 -70
rect -64 -467 -58 -70
rect -320 -479 -58 -467
rect 58 -70 320 -58
rect 58 -467 64 -70
rect 314 -467 320 -70
rect 58 -479 320 -467
rect 436 -70 698 -58
rect 436 -467 442 -70
rect 692 -467 698 -70
rect 436 -479 698 -467
rect 814 -70 1076 -58
rect 814 -467 820 -70
rect 1070 -467 1076 -70
rect 814 -479 1076 -467
rect 1192 -70 1454 -58
rect 1192 -467 1198 -70
rect 1448 -467 1454 -70
rect 1192 -479 1454 -467
rect 1570 -70 1832 -58
rect 1570 -467 1576 -70
rect 1826 -467 1832 -70
rect 1570 -479 1832 -467
rect -1832 -1301 -1570 -1289
rect -1832 -1698 -1826 -1301
rect -1576 -1698 -1570 -1301
rect -1832 -1710 -1570 -1698
rect -1454 -1301 -1192 -1289
rect -1454 -1698 -1448 -1301
rect -1198 -1698 -1192 -1301
rect -1454 -1710 -1192 -1698
rect -1076 -1301 -814 -1289
rect -1076 -1698 -1070 -1301
rect -820 -1698 -814 -1301
rect -1076 -1710 -814 -1698
rect -698 -1301 -436 -1289
rect -698 -1698 -692 -1301
rect -442 -1698 -436 -1301
rect -698 -1710 -436 -1698
rect -320 -1301 -58 -1289
rect -320 -1698 -314 -1301
rect -64 -1698 -58 -1301
rect -320 -1710 -58 -1698
rect 58 -1301 320 -1289
rect 58 -1698 64 -1301
rect 314 -1698 320 -1301
rect 58 -1710 320 -1698
rect 436 -1301 698 -1289
rect 436 -1698 442 -1301
rect 692 -1698 698 -1301
rect 436 -1710 698 -1698
rect 814 -1301 1076 -1289
rect 814 -1698 820 -1301
rect 1070 -1698 1076 -1301
rect 814 -1710 1076 -1698
rect 1192 -1301 1454 -1289
rect 1192 -1698 1198 -1301
rect 1448 -1698 1454 -1301
rect 1192 -1710 1454 -1698
rect 1570 -1301 1832 -1289
rect 1570 -1698 1576 -1301
rect 1826 -1698 1832 -1301
rect 1570 -1710 1832 -1698
<< res1p41 >>
rect -1844 482 -1558 1286
rect -1466 482 -1180 1286
rect -1088 482 -802 1286
rect -710 482 -424 1286
rect -332 482 -46 1286
rect 46 482 332 1286
rect 424 482 710 1286
rect 802 482 1088 1286
rect 1180 482 1466 1286
rect 1558 482 1844 1286
rect -1844 -1286 -1558 -482
rect -1466 -1286 -1180 -482
rect -1088 -1286 -802 -482
rect -710 -1286 -424 -482
rect -332 -1286 -46 -482
rect 46 -1286 332 -482
rect 424 -1286 710 -482
rect 802 -1286 1088 -482
rect 1180 -1286 1466 -482
rect 1558 -1286 1844 -482
<< properties >>
string FIXED_BBOX -1955 -1829 1955 1829
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.41 l 4.0 m 2 nx 10 wmin 1.410 lmin 0.50 rho 319.8 val 1.183k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
