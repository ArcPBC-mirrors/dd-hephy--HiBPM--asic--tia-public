magic
tech sky130A
magscale 1 2
timestamp 1683558579
<< nwell >>
rect -12473 127 -10207 709
rect -9953 127 -7687 709
rect -7433 127 -5167 709
rect -4913 127 -2647 709
rect -2393 127 -127 709
rect 127 127 2393 709
rect 2647 127 4913 709
rect 5167 127 7433 709
rect 7687 127 9953 709
rect 10207 127 12473 709
rect -12473 -709 -10207 -127
rect -9953 -709 -7687 -127
rect -7433 -709 -5167 -127
rect -4913 -709 -2647 -127
rect -2393 -709 -127 -127
rect 127 -709 2393 -127
rect 2647 -709 4913 -127
rect 5167 -709 7433 -127
rect 7687 -709 9953 -127
rect 10207 -709 12473 -127
<< pwell >>
rect -12583 709 12583 819
rect -12583 127 -12473 709
rect -10207 127 -9953 709
rect -7687 127 -7433 709
rect -5167 127 -4913 709
rect -2647 127 -2393 709
rect -127 127 127 709
rect 2393 127 2647 709
rect 4913 127 5167 709
rect 7433 127 7687 709
rect 9953 127 10207 709
rect 12473 127 12583 709
rect -12583 -127 12583 127
rect -12583 -709 -12473 -127
rect -10207 -709 -9953 -127
rect -7687 -709 -7433 -127
rect -5167 -709 -4913 -127
rect -2647 -709 -2393 -127
rect -127 -709 127 -127
rect 2393 -709 2647 -127
rect 4913 -709 5167 -127
rect 7433 -709 7687 -127
rect 9953 -709 10207 -127
rect 12473 -709 12583 -127
rect -12583 -819 12583 -709
<< varactor >>
rect -12340 218 -10340 618
rect -9820 218 -7820 618
rect -7300 218 -5300 618
rect -4780 218 -2780 618
rect -2260 218 -260 618
rect 260 218 2260 618
rect 2780 218 4780 618
rect 5300 218 7300 618
rect 7820 218 9820 618
rect 10340 218 12340 618
rect -12340 -618 -10340 -218
rect -9820 -618 -7820 -218
rect -7300 -618 -5300 -218
rect -4780 -618 -2780 -218
rect -2260 -618 -260 -218
rect 260 -618 2260 -218
rect 2780 -618 4780 -218
rect 5300 -618 7300 -218
rect 7820 -618 9820 -218
rect 10340 -618 12340 -218
<< psubdiff >>
rect -12547 749 -12451 783
rect 12451 749 12547 783
rect -12547 687 -12513 749
rect 12513 687 12547 749
rect -12547 -749 -12513 -687
rect 12513 -749 12547 -687
rect -12547 -783 -12451 -749
rect 12451 -783 12547 -749
<< nsubdiff >>
rect -12437 594 -12340 618
rect -12437 242 -12425 594
rect -12391 242 -12340 594
rect -12437 218 -12340 242
rect -10340 594 -10243 618
rect -10340 242 -10289 594
rect -10255 242 -10243 594
rect -10340 218 -10243 242
rect -9917 594 -9820 618
rect -9917 242 -9905 594
rect -9871 242 -9820 594
rect -9917 218 -9820 242
rect -7820 594 -7723 618
rect -7820 242 -7769 594
rect -7735 242 -7723 594
rect -7820 218 -7723 242
rect -7397 594 -7300 618
rect -7397 242 -7385 594
rect -7351 242 -7300 594
rect -7397 218 -7300 242
rect -5300 594 -5203 618
rect -5300 242 -5249 594
rect -5215 242 -5203 594
rect -5300 218 -5203 242
rect -4877 594 -4780 618
rect -4877 242 -4865 594
rect -4831 242 -4780 594
rect -4877 218 -4780 242
rect -2780 594 -2683 618
rect -2780 242 -2729 594
rect -2695 242 -2683 594
rect -2780 218 -2683 242
rect -2357 594 -2260 618
rect -2357 242 -2345 594
rect -2311 242 -2260 594
rect -2357 218 -2260 242
rect -260 594 -163 618
rect -260 242 -209 594
rect -175 242 -163 594
rect -260 218 -163 242
rect 163 594 260 618
rect 163 242 175 594
rect 209 242 260 594
rect 163 218 260 242
rect 2260 594 2357 618
rect 2260 242 2311 594
rect 2345 242 2357 594
rect 2260 218 2357 242
rect 2683 594 2780 618
rect 2683 242 2695 594
rect 2729 242 2780 594
rect 2683 218 2780 242
rect 4780 594 4877 618
rect 4780 242 4831 594
rect 4865 242 4877 594
rect 4780 218 4877 242
rect 5203 594 5300 618
rect 5203 242 5215 594
rect 5249 242 5300 594
rect 5203 218 5300 242
rect 7300 594 7397 618
rect 7300 242 7351 594
rect 7385 242 7397 594
rect 7300 218 7397 242
rect 7723 594 7820 618
rect 7723 242 7735 594
rect 7769 242 7820 594
rect 7723 218 7820 242
rect 9820 594 9917 618
rect 9820 242 9871 594
rect 9905 242 9917 594
rect 9820 218 9917 242
rect 10243 594 10340 618
rect 10243 242 10255 594
rect 10289 242 10340 594
rect 10243 218 10340 242
rect 12340 594 12437 618
rect 12340 242 12391 594
rect 12425 242 12437 594
rect 12340 218 12437 242
rect -12437 -242 -12340 -218
rect -12437 -594 -12425 -242
rect -12391 -594 -12340 -242
rect -12437 -618 -12340 -594
rect -10340 -242 -10243 -218
rect -10340 -594 -10289 -242
rect -10255 -594 -10243 -242
rect -10340 -618 -10243 -594
rect -9917 -242 -9820 -218
rect -9917 -594 -9905 -242
rect -9871 -594 -9820 -242
rect -9917 -618 -9820 -594
rect -7820 -242 -7723 -218
rect -7820 -594 -7769 -242
rect -7735 -594 -7723 -242
rect -7820 -618 -7723 -594
rect -7397 -242 -7300 -218
rect -7397 -594 -7385 -242
rect -7351 -594 -7300 -242
rect -7397 -618 -7300 -594
rect -5300 -242 -5203 -218
rect -5300 -594 -5249 -242
rect -5215 -594 -5203 -242
rect -5300 -618 -5203 -594
rect -4877 -242 -4780 -218
rect -4877 -594 -4865 -242
rect -4831 -594 -4780 -242
rect -4877 -618 -4780 -594
rect -2780 -242 -2683 -218
rect -2780 -594 -2729 -242
rect -2695 -594 -2683 -242
rect -2780 -618 -2683 -594
rect -2357 -242 -2260 -218
rect -2357 -594 -2345 -242
rect -2311 -594 -2260 -242
rect -2357 -618 -2260 -594
rect -260 -242 -163 -218
rect -260 -594 -209 -242
rect -175 -594 -163 -242
rect -260 -618 -163 -594
rect 163 -242 260 -218
rect 163 -594 175 -242
rect 209 -594 260 -242
rect 163 -618 260 -594
rect 2260 -242 2357 -218
rect 2260 -594 2311 -242
rect 2345 -594 2357 -242
rect 2260 -618 2357 -594
rect 2683 -242 2780 -218
rect 2683 -594 2695 -242
rect 2729 -594 2780 -242
rect 2683 -618 2780 -594
rect 4780 -242 4877 -218
rect 4780 -594 4831 -242
rect 4865 -594 4877 -242
rect 4780 -618 4877 -594
rect 5203 -242 5300 -218
rect 5203 -594 5215 -242
rect 5249 -594 5300 -242
rect 5203 -618 5300 -594
rect 7300 -242 7397 -218
rect 7300 -594 7351 -242
rect 7385 -594 7397 -242
rect 7300 -618 7397 -594
rect 7723 -242 7820 -218
rect 7723 -594 7735 -242
rect 7769 -594 7820 -242
rect 7723 -618 7820 -594
rect 9820 -242 9917 -218
rect 9820 -594 9871 -242
rect 9905 -594 9917 -242
rect 9820 -618 9917 -594
rect 10243 -242 10340 -218
rect 10243 -594 10255 -242
rect 10289 -594 10340 -242
rect 10243 -618 10340 -594
rect 12340 -242 12437 -218
rect 12340 -594 12391 -242
rect 12425 -594 12437 -242
rect 12340 -618 12437 -594
<< psubdiffcont >>
rect -12451 749 12451 783
rect -12547 -687 -12513 687
rect 12513 -687 12547 687
rect -12451 -783 12451 -749
<< nsubdiffcont >>
rect -12425 242 -12391 594
rect -10289 242 -10255 594
rect -9905 242 -9871 594
rect -7769 242 -7735 594
rect -7385 242 -7351 594
rect -5249 242 -5215 594
rect -4865 242 -4831 594
rect -2729 242 -2695 594
rect -2345 242 -2311 594
rect -209 242 -175 594
rect 175 242 209 594
rect 2311 242 2345 594
rect 2695 242 2729 594
rect 4831 242 4865 594
rect 5215 242 5249 594
rect 7351 242 7385 594
rect 7735 242 7769 594
rect 9871 242 9905 594
rect 10255 242 10289 594
rect 12391 242 12425 594
rect -12425 -594 -12391 -242
rect -10289 -594 -10255 -242
rect -9905 -594 -9871 -242
rect -7769 -594 -7735 -242
rect -7385 -594 -7351 -242
rect -5249 -594 -5215 -242
rect -4865 -594 -4831 -242
rect -2729 -594 -2695 -242
rect -2345 -594 -2311 -242
rect -209 -594 -175 -242
rect 175 -594 209 -242
rect 2311 -594 2345 -242
rect 2695 -594 2729 -242
rect 4831 -594 4865 -242
rect 5215 -594 5249 -242
rect 7351 -594 7385 -242
rect 7735 -594 7769 -242
rect 9871 -594 9905 -242
rect 10255 -594 10289 -242
rect 12391 -594 12425 -242
<< poly >>
rect -12340 690 -10340 706
rect -12340 656 -12324 690
rect -10356 656 -10340 690
rect -12340 618 -10340 656
rect -9820 690 -7820 706
rect -9820 656 -9804 690
rect -7836 656 -7820 690
rect -9820 618 -7820 656
rect -7300 690 -5300 706
rect -7300 656 -7284 690
rect -5316 656 -5300 690
rect -7300 618 -5300 656
rect -4780 690 -2780 706
rect -4780 656 -4764 690
rect -2796 656 -2780 690
rect -4780 618 -2780 656
rect -2260 690 -260 706
rect -2260 656 -2244 690
rect -276 656 -260 690
rect -2260 618 -260 656
rect 260 690 2260 706
rect 260 656 276 690
rect 2244 656 2260 690
rect 260 618 2260 656
rect 2780 690 4780 706
rect 2780 656 2796 690
rect 4764 656 4780 690
rect 2780 618 4780 656
rect 5300 690 7300 706
rect 5300 656 5316 690
rect 7284 656 7300 690
rect 5300 618 7300 656
rect 7820 690 9820 706
rect 7820 656 7836 690
rect 9804 656 9820 690
rect 7820 618 9820 656
rect 10340 690 12340 706
rect 10340 656 10356 690
rect 12324 656 12340 690
rect 10340 618 12340 656
rect -12340 180 -10340 218
rect -12340 146 -12324 180
rect -10356 146 -10340 180
rect -12340 130 -10340 146
rect -9820 180 -7820 218
rect -9820 146 -9804 180
rect -7836 146 -7820 180
rect -9820 130 -7820 146
rect -7300 180 -5300 218
rect -7300 146 -7284 180
rect -5316 146 -5300 180
rect -7300 130 -5300 146
rect -4780 180 -2780 218
rect -4780 146 -4764 180
rect -2796 146 -2780 180
rect -4780 130 -2780 146
rect -2260 180 -260 218
rect -2260 146 -2244 180
rect -276 146 -260 180
rect -2260 130 -260 146
rect 260 180 2260 218
rect 260 146 276 180
rect 2244 146 2260 180
rect 260 130 2260 146
rect 2780 180 4780 218
rect 2780 146 2796 180
rect 4764 146 4780 180
rect 2780 130 4780 146
rect 5300 180 7300 218
rect 5300 146 5316 180
rect 7284 146 7300 180
rect 5300 130 7300 146
rect 7820 180 9820 218
rect 7820 146 7836 180
rect 9804 146 9820 180
rect 7820 130 9820 146
rect 10340 180 12340 218
rect 10340 146 10356 180
rect 12324 146 12340 180
rect 10340 130 12340 146
rect -12340 -146 -10340 -130
rect -12340 -180 -12324 -146
rect -10356 -180 -10340 -146
rect -12340 -218 -10340 -180
rect -9820 -146 -7820 -130
rect -9820 -180 -9804 -146
rect -7836 -180 -7820 -146
rect -9820 -218 -7820 -180
rect -7300 -146 -5300 -130
rect -7300 -180 -7284 -146
rect -5316 -180 -5300 -146
rect -7300 -218 -5300 -180
rect -4780 -146 -2780 -130
rect -4780 -180 -4764 -146
rect -2796 -180 -2780 -146
rect -4780 -218 -2780 -180
rect -2260 -146 -260 -130
rect -2260 -180 -2244 -146
rect -276 -180 -260 -146
rect -2260 -218 -260 -180
rect 260 -146 2260 -130
rect 260 -180 276 -146
rect 2244 -180 2260 -146
rect 260 -218 2260 -180
rect 2780 -146 4780 -130
rect 2780 -180 2796 -146
rect 4764 -180 4780 -146
rect 2780 -218 4780 -180
rect 5300 -146 7300 -130
rect 5300 -180 5316 -146
rect 7284 -180 7300 -146
rect 5300 -218 7300 -180
rect 7820 -146 9820 -130
rect 7820 -180 7836 -146
rect 9804 -180 9820 -146
rect 7820 -218 9820 -180
rect 10340 -146 12340 -130
rect 10340 -180 10356 -146
rect 12324 -180 12340 -146
rect 10340 -218 12340 -180
rect -12340 -656 -10340 -618
rect -12340 -690 -12324 -656
rect -10356 -690 -10340 -656
rect -12340 -706 -10340 -690
rect -9820 -656 -7820 -618
rect -9820 -690 -9804 -656
rect -7836 -690 -7820 -656
rect -9820 -706 -7820 -690
rect -7300 -656 -5300 -618
rect -7300 -690 -7284 -656
rect -5316 -690 -5300 -656
rect -7300 -706 -5300 -690
rect -4780 -656 -2780 -618
rect -4780 -690 -4764 -656
rect -2796 -690 -2780 -656
rect -4780 -706 -2780 -690
rect -2260 -656 -260 -618
rect -2260 -690 -2244 -656
rect -276 -690 -260 -656
rect -2260 -706 -260 -690
rect 260 -656 2260 -618
rect 260 -690 276 -656
rect 2244 -690 2260 -656
rect 260 -706 2260 -690
rect 2780 -656 4780 -618
rect 2780 -690 2796 -656
rect 4764 -690 4780 -656
rect 2780 -706 4780 -690
rect 5300 -656 7300 -618
rect 5300 -690 5316 -656
rect 7284 -690 7300 -656
rect 5300 -706 7300 -690
rect 7820 -656 9820 -618
rect 7820 -690 7836 -656
rect 9804 -690 9820 -656
rect 7820 -706 9820 -690
rect 10340 -656 12340 -618
rect 10340 -690 10356 -656
rect 12324 -690 12340 -656
rect 10340 -706 12340 -690
<< polycont >>
rect -12324 656 -10356 690
rect -9804 656 -7836 690
rect -7284 656 -5316 690
rect -4764 656 -2796 690
rect -2244 656 -276 690
rect 276 656 2244 690
rect 2796 656 4764 690
rect 5316 656 7284 690
rect 7836 656 9804 690
rect 10356 656 12324 690
rect -12324 146 -10356 180
rect -9804 146 -7836 180
rect -7284 146 -5316 180
rect -4764 146 -2796 180
rect -2244 146 -276 180
rect 276 146 2244 180
rect 2796 146 4764 180
rect 5316 146 7284 180
rect 7836 146 9804 180
rect 10356 146 12324 180
rect -12324 -180 -10356 -146
rect -9804 -180 -7836 -146
rect -7284 -180 -5316 -146
rect -4764 -180 -2796 -146
rect -2244 -180 -276 -146
rect 276 -180 2244 -146
rect 2796 -180 4764 -146
rect 5316 -180 7284 -146
rect 7836 -180 9804 -146
rect 10356 -180 12324 -146
rect -12324 -690 -10356 -656
rect -9804 -690 -7836 -656
rect -7284 -690 -5316 -656
rect -4764 -690 -2796 -656
rect -2244 -690 -276 -656
rect 276 -690 2244 -656
rect 2796 -690 4764 -656
rect 5316 -690 7284 -656
rect 7836 -690 9804 -656
rect 10356 -690 12324 -656
<< locali >>
rect -12547 749 -12451 783
rect 12451 749 12547 783
rect -12547 687 -12513 749
rect -12340 656 -12324 690
rect -10356 656 -10340 690
rect -9820 656 -9804 690
rect -7836 656 -7820 690
rect -7300 656 -7284 690
rect -5316 656 -5300 690
rect -4780 656 -4764 690
rect -2796 656 -2780 690
rect -2260 656 -2244 690
rect -276 656 -260 690
rect 260 656 276 690
rect 2244 656 2260 690
rect 2780 656 2796 690
rect 4764 656 4780 690
rect 5300 656 5316 690
rect 7284 656 7300 690
rect 7820 656 7836 690
rect 9804 656 9820 690
rect 10340 656 10356 690
rect 12324 656 12340 690
rect 12513 687 12547 749
rect -12425 594 -12391 610
rect -12425 226 -12391 242
rect -10289 594 -10255 610
rect -10289 226 -10255 242
rect -9905 594 -9871 610
rect -9905 226 -9871 242
rect -7769 594 -7735 610
rect -7769 226 -7735 242
rect -7385 594 -7351 610
rect -7385 226 -7351 242
rect -5249 594 -5215 610
rect -5249 226 -5215 242
rect -4865 594 -4831 610
rect -4865 226 -4831 242
rect -2729 594 -2695 610
rect -2729 226 -2695 242
rect -2345 594 -2311 610
rect -2345 226 -2311 242
rect -209 594 -175 610
rect -209 226 -175 242
rect 175 594 209 610
rect 175 226 209 242
rect 2311 594 2345 610
rect 2311 226 2345 242
rect 2695 594 2729 610
rect 2695 226 2729 242
rect 4831 594 4865 610
rect 4831 226 4865 242
rect 5215 594 5249 610
rect 5215 226 5249 242
rect 7351 594 7385 610
rect 7351 226 7385 242
rect 7735 594 7769 610
rect 7735 226 7769 242
rect 9871 594 9905 610
rect 9871 226 9905 242
rect 10255 594 10289 610
rect 10255 226 10289 242
rect 12391 594 12425 610
rect 12391 226 12425 242
rect -12340 146 -12324 180
rect -10356 146 -10340 180
rect -9820 146 -9804 180
rect -7836 146 -7820 180
rect -7300 146 -7284 180
rect -5316 146 -5300 180
rect -4780 146 -4764 180
rect -2796 146 -2780 180
rect -2260 146 -2244 180
rect -276 146 -260 180
rect 260 146 276 180
rect 2244 146 2260 180
rect 2780 146 2796 180
rect 4764 146 4780 180
rect 5300 146 5316 180
rect 7284 146 7300 180
rect 7820 146 7836 180
rect 9804 146 9820 180
rect 10340 146 10356 180
rect 12324 146 12340 180
rect -12340 -180 -12324 -146
rect -10356 -180 -10340 -146
rect -9820 -180 -9804 -146
rect -7836 -180 -7820 -146
rect -7300 -180 -7284 -146
rect -5316 -180 -5300 -146
rect -4780 -180 -4764 -146
rect -2796 -180 -2780 -146
rect -2260 -180 -2244 -146
rect -276 -180 -260 -146
rect 260 -180 276 -146
rect 2244 -180 2260 -146
rect 2780 -180 2796 -146
rect 4764 -180 4780 -146
rect 5300 -180 5316 -146
rect 7284 -180 7300 -146
rect 7820 -180 7836 -146
rect 9804 -180 9820 -146
rect 10340 -180 10356 -146
rect 12324 -180 12340 -146
rect -12425 -242 -12391 -226
rect -12425 -610 -12391 -594
rect -10289 -242 -10255 -226
rect -10289 -610 -10255 -594
rect -9905 -242 -9871 -226
rect -9905 -610 -9871 -594
rect -7769 -242 -7735 -226
rect -7769 -610 -7735 -594
rect -7385 -242 -7351 -226
rect -7385 -610 -7351 -594
rect -5249 -242 -5215 -226
rect -5249 -610 -5215 -594
rect -4865 -242 -4831 -226
rect -4865 -610 -4831 -594
rect -2729 -242 -2695 -226
rect -2729 -610 -2695 -594
rect -2345 -242 -2311 -226
rect -2345 -610 -2311 -594
rect -209 -242 -175 -226
rect -209 -610 -175 -594
rect 175 -242 209 -226
rect 175 -610 209 -594
rect 2311 -242 2345 -226
rect 2311 -610 2345 -594
rect 2695 -242 2729 -226
rect 2695 -610 2729 -594
rect 4831 -242 4865 -226
rect 4831 -610 4865 -594
rect 5215 -242 5249 -226
rect 5215 -610 5249 -594
rect 7351 -242 7385 -226
rect 7351 -610 7385 -594
rect 7735 -242 7769 -226
rect 7735 -610 7769 -594
rect 9871 -242 9905 -226
rect 9871 -610 9905 -594
rect 10255 -242 10289 -226
rect 10255 -610 10289 -594
rect 12391 -242 12425 -226
rect 12391 -610 12425 -594
rect -12547 -749 -12513 -687
rect -12340 -690 -12324 -656
rect -10356 -690 -10340 -656
rect -9820 -690 -9804 -656
rect -7836 -690 -7820 -656
rect -7300 -690 -7284 -656
rect -5316 -690 -5300 -656
rect -4780 -690 -4764 -656
rect -2796 -690 -2780 -656
rect -2260 -690 -2244 -656
rect -276 -690 -260 -656
rect 260 -690 276 -656
rect 2244 -690 2260 -656
rect 2780 -690 2796 -656
rect 4764 -690 4780 -656
rect 5300 -690 5316 -656
rect 7284 -690 7300 -656
rect 7820 -690 7836 -656
rect 9804 -690 9820 -656
rect 10340 -690 10356 -656
rect 12324 -690 12340 -656
rect 12513 -749 12547 -687
rect -12547 -783 -12451 -749
rect 12451 -783 12547 -749
<< viali >>
rect -12324 656 -10356 690
rect -9804 656 -7836 690
rect -7284 656 -5316 690
rect -4764 656 -2796 690
rect -2244 656 -276 690
rect 276 656 2244 690
rect 2796 656 4764 690
rect 5316 656 7284 690
rect 7836 656 9804 690
rect 10356 656 12324 690
rect -12425 242 -12391 594
rect -10289 242 -10255 594
rect -9905 242 -9871 594
rect -7769 242 -7735 594
rect -7385 242 -7351 594
rect -5249 242 -5215 594
rect -4865 242 -4831 594
rect -2729 242 -2695 594
rect -2345 242 -2311 594
rect -209 242 -175 594
rect 175 242 209 594
rect 2311 242 2345 594
rect 2695 242 2729 594
rect 4831 242 4865 594
rect 5215 242 5249 594
rect 7351 242 7385 594
rect 7735 242 7769 594
rect 9871 242 9905 594
rect 10255 242 10289 594
rect 12391 242 12425 594
rect -12324 146 -10356 180
rect -9804 146 -7836 180
rect -7284 146 -5316 180
rect -4764 146 -2796 180
rect -2244 146 -276 180
rect 276 146 2244 180
rect 2796 146 4764 180
rect 5316 146 7284 180
rect 7836 146 9804 180
rect 10356 146 12324 180
rect -12324 -180 -10356 -146
rect -9804 -180 -7836 -146
rect -7284 -180 -5316 -146
rect -4764 -180 -2796 -146
rect -2244 -180 -276 -146
rect 276 -180 2244 -146
rect 2796 -180 4764 -146
rect 5316 -180 7284 -146
rect 7836 -180 9804 -146
rect 10356 -180 12324 -146
rect -12425 -594 -12391 -242
rect -10289 -594 -10255 -242
rect -9905 -594 -9871 -242
rect -7769 -594 -7735 -242
rect -7385 -594 -7351 -242
rect -5249 -594 -5215 -242
rect -4865 -594 -4831 -242
rect -2729 -594 -2695 -242
rect -2345 -594 -2311 -242
rect -209 -594 -175 -242
rect 175 -594 209 -242
rect 2311 -594 2345 -242
rect 2695 -594 2729 -242
rect 4831 -594 4865 -242
rect 5215 -594 5249 -242
rect 7351 -594 7385 -242
rect 7735 -594 7769 -242
rect 9871 -594 9905 -242
rect 10255 -594 10289 -242
rect 12391 -594 12425 -242
rect -12324 -690 -10356 -656
rect -9804 -690 -7836 -656
rect -7284 -690 -5316 -656
rect -4764 -690 -2796 -656
rect -2244 -690 -276 -656
rect 276 -690 2244 -656
rect 2796 -690 4764 -656
rect 5316 -690 7284 -656
rect 7836 -690 9804 -656
rect 10356 -690 12324 -656
<< metal1 >>
rect -12336 690 -10344 696
rect -12336 656 -12324 690
rect -10356 656 -10344 690
rect -12336 650 -10344 656
rect -9816 690 -7824 696
rect -9816 656 -9804 690
rect -7836 656 -7824 690
rect -9816 650 -7824 656
rect -7296 690 -5304 696
rect -7296 656 -7284 690
rect -5316 656 -5304 690
rect -7296 650 -5304 656
rect -4776 690 -2784 696
rect -4776 656 -4764 690
rect -2796 656 -2784 690
rect -4776 650 -2784 656
rect -2256 690 -264 696
rect -2256 656 -2244 690
rect -276 656 -264 690
rect -2256 650 -264 656
rect 264 690 2256 696
rect 264 656 276 690
rect 2244 656 2256 690
rect 264 650 2256 656
rect 2784 690 4776 696
rect 2784 656 2796 690
rect 4764 656 4776 690
rect 2784 650 4776 656
rect 5304 690 7296 696
rect 5304 656 5316 690
rect 7284 656 7296 690
rect 5304 650 7296 656
rect 7824 690 9816 696
rect 7824 656 7836 690
rect 9804 656 9816 690
rect 7824 650 9816 656
rect 10344 690 12336 696
rect 10344 656 10356 690
rect 12324 656 12336 690
rect 10344 650 12336 656
rect -12431 594 -12385 606
rect -10295 594 -10249 606
rect -12431 242 -12425 594
rect -12391 242 -10289 594
rect -10255 242 -10249 594
rect -12431 230 -12385 242
rect -10295 230 -10249 242
rect -9911 594 -9865 606
rect -7775 594 -7729 606
rect -9911 242 -9905 594
rect -9871 242 -7769 594
rect -7735 242 -7729 594
rect -9911 230 -9865 242
rect -7775 230 -7729 242
rect -7391 594 -7345 606
rect -5255 594 -5209 606
rect -7391 242 -7385 594
rect -7351 242 -5249 594
rect -5215 242 -5209 594
rect -7391 230 -7345 242
rect -5255 230 -5209 242
rect -4871 594 -4825 606
rect -2735 594 -2689 606
rect -4871 242 -4865 594
rect -4831 242 -2729 594
rect -2695 242 -2689 594
rect -4871 230 -4825 242
rect -2735 230 -2689 242
rect -2351 594 -2305 606
rect -215 594 -169 606
rect -2351 242 -2345 594
rect -2311 242 -209 594
rect -175 242 -169 594
rect -2351 230 -2305 242
rect -215 230 -169 242
rect 169 594 215 606
rect 2305 594 2351 606
rect 169 242 175 594
rect 209 242 2311 594
rect 2345 242 2351 594
rect 169 230 215 242
rect 2305 230 2351 242
rect 2689 594 2735 606
rect 4825 594 4871 606
rect 2689 242 2695 594
rect 2729 242 4831 594
rect 4865 242 4871 594
rect 2689 230 2735 242
rect 4825 230 4871 242
rect 5209 594 5255 606
rect 7345 594 7391 606
rect 5209 242 5215 594
rect 5249 242 7351 594
rect 7385 242 7391 594
rect 5209 230 5255 242
rect 7345 230 7391 242
rect 7729 594 7775 606
rect 9865 594 9911 606
rect 7729 242 7735 594
rect 7769 242 9871 594
rect 9905 242 9911 594
rect 7729 230 7775 242
rect 9865 230 9911 242
rect 10249 594 10295 606
rect 12385 594 12431 606
rect 10249 242 10255 594
rect 10289 242 12391 594
rect 12425 242 12431 594
rect 10249 230 10295 242
rect 12385 230 12431 242
rect -12336 180 -10344 186
rect -12336 146 -12324 180
rect -10356 146 -10344 180
rect -12336 140 -10344 146
rect -9816 180 -7824 186
rect -9816 146 -9804 180
rect -7836 146 -7824 180
rect -9816 140 -7824 146
rect -7296 180 -5304 186
rect -7296 146 -7284 180
rect -5316 146 -5304 180
rect -7296 140 -5304 146
rect -4776 180 -2784 186
rect -4776 146 -4764 180
rect -2796 146 -2784 180
rect -4776 140 -2784 146
rect -2256 180 -264 186
rect -2256 146 -2244 180
rect -276 146 -264 180
rect -2256 140 -264 146
rect 264 180 2256 186
rect 264 146 276 180
rect 2244 146 2256 180
rect 264 140 2256 146
rect 2784 180 4776 186
rect 2784 146 2796 180
rect 4764 146 4776 180
rect 2784 140 4776 146
rect 5304 180 7296 186
rect 5304 146 5316 180
rect 7284 146 7296 180
rect 5304 140 7296 146
rect 7824 180 9816 186
rect 7824 146 7836 180
rect 9804 146 9816 180
rect 7824 140 9816 146
rect 10344 180 12336 186
rect 10344 146 10356 180
rect 12324 146 12336 180
rect 10344 140 12336 146
rect -12336 -146 -10344 -140
rect -12336 -180 -12324 -146
rect -10356 -180 -10344 -146
rect -12336 -186 -10344 -180
rect -9816 -146 -7824 -140
rect -9816 -180 -9804 -146
rect -7836 -180 -7824 -146
rect -9816 -186 -7824 -180
rect -7296 -146 -5304 -140
rect -7296 -180 -7284 -146
rect -5316 -180 -5304 -146
rect -7296 -186 -5304 -180
rect -4776 -146 -2784 -140
rect -4776 -180 -4764 -146
rect -2796 -180 -2784 -146
rect -4776 -186 -2784 -180
rect -2256 -146 -264 -140
rect -2256 -180 -2244 -146
rect -276 -180 -264 -146
rect -2256 -186 -264 -180
rect 264 -146 2256 -140
rect 264 -180 276 -146
rect 2244 -180 2256 -146
rect 264 -186 2256 -180
rect 2784 -146 4776 -140
rect 2784 -180 2796 -146
rect 4764 -180 4776 -146
rect 2784 -186 4776 -180
rect 5304 -146 7296 -140
rect 5304 -180 5316 -146
rect 7284 -180 7296 -146
rect 5304 -186 7296 -180
rect 7824 -146 9816 -140
rect 7824 -180 7836 -146
rect 9804 -180 9816 -146
rect 7824 -186 9816 -180
rect 10344 -146 12336 -140
rect 10344 -180 10356 -146
rect 12324 -180 12336 -146
rect 10344 -186 12336 -180
rect -12431 -242 -12385 -230
rect -10295 -242 -10249 -230
rect -12431 -594 -12425 -242
rect -12391 -594 -10289 -242
rect -10255 -594 -10249 -242
rect -12431 -606 -12385 -594
rect -10295 -606 -10249 -594
rect -9911 -242 -9865 -230
rect -7775 -242 -7729 -230
rect -9911 -594 -9905 -242
rect -9871 -594 -7769 -242
rect -7735 -594 -7729 -242
rect -9911 -606 -9865 -594
rect -7775 -606 -7729 -594
rect -7391 -242 -7345 -230
rect -5255 -242 -5209 -230
rect -7391 -594 -7385 -242
rect -7351 -594 -5249 -242
rect -5215 -594 -5209 -242
rect -7391 -606 -7345 -594
rect -5255 -606 -5209 -594
rect -4871 -242 -4825 -230
rect -2735 -242 -2689 -230
rect -4871 -594 -4865 -242
rect -4831 -594 -2729 -242
rect -2695 -594 -2689 -242
rect -4871 -606 -4825 -594
rect -2735 -606 -2689 -594
rect -2351 -242 -2305 -230
rect -215 -242 -169 -230
rect -2351 -594 -2345 -242
rect -2311 -594 -209 -242
rect -175 -594 -169 -242
rect -2351 -606 -2305 -594
rect -215 -606 -169 -594
rect 169 -242 215 -230
rect 2305 -242 2351 -230
rect 169 -594 175 -242
rect 209 -594 2311 -242
rect 2345 -594 2351 -242
rect 169 -606 215 -594
rect 2305 -606 2351 -594
rect 2689 -242 2735 -230
rect 4825 -242 4871 -230
rect 2689 -594 2695 -242
rect 2729 -594 4831 -242
rect 4865 -594 4871 -242
rect 2689 -606 2735 -594
rect 4825 -606 4871 -594
rect 5209 -242 5255 -230
rect 7345 -242 7391 -230
rect 5209 -594 5215 -242
rect 5249 -594 7351 -242
rect 7385 -594 7391 -242
rect 5209 -606 5255 -594
rect 7345 -606 7391 -594
rect 7729 -242 7775 -230
rect 9865 -242 9911 -230
rect 7729 -594 7735 -242
rect 7769 -594 9871 -242
rect 9905 -594 9911 -242
rect 7729 -606 7775 -594
rect 9865 -606 9911 -594
rect 10249 -242 10295 -230
rect 12385 -242 12431 -230
rect 10249 -594 10255 -242
rect 10289 -594 12391 -242
rect 12425 -594 12431 -242
rect 10249 -606 10295 -594
rect 12385 -606 12431 -594
rect -12336 -656 -10344 -650
rect -12336 -690 -12324 -656
rect -10356 -690 -10344 -656
rect -12336 -696 -10344 -690
rect -9816 -656 -7824 -650
rect -9816 -690 -9804 -656
rect -7836 -690 -7824 -656
rect -9816 -696 -7824 -690
rect -7296 -656 -5304 -650
rect -7296 -690 -7284 -656
rect -5316 -690 -5304 -656
rect -7296 -696 -5304 -690
rect -4776 -656 -2784 -650
rect -4776 -690 -4764 -656
rect -2796 -690 -2784 -656
rect -4776 -696 -2784 -690
rect -2256 -656 -264 -650
rect -2256 -690 -2244 -656
rect -276 -690 -264 -656
rect -2256 -696 -264 -690
rect 264 -656 2256 -650
rect 264 -690 276 -656
rect 2244 -690 2256 -656
rect 264 -696 2256 -690
rect 2784 -656 4776 -650
rect 2784 -690 2796 -656
rect 4764 -690 4776 -656
rect 2784 -696 4776 -690
rect 5304 -656 7296 -650
rect 5304 -690 5316 -656
rect 7284 -690 7296 -656
rect 5304 -696 7296 -690
rect 7824 -656 9816 -650
rect 7824 -690 7836 -656
rect 9804 -690 9816 -656
rect 7824 -696 9816 -690
rect 10344 -656 12336 -650
rect 10344 -690 10356 -656
rect 12324 -690 12336 -656
rect 10344 -696 12336 -690
<< properties >>
string FIXED_BBOX -12530 -766 12530 766
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 10 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
