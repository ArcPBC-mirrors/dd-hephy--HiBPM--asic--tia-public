magic
tech sky130A
magscale 1 2
timestamp 1684829418
<< pwell >>
rect -874 -1182 874 1182
<< psubdiff >>
rect -838 1112 -742 1146
rect 742 1112 838 1146
rect -838 1050 -804 1112
rect 804 1050 838 1112
rect -838 -1112 -804 -1050
rect 804 -1112 838 -1050
rect -838 -1146 -742 -1112
rect 742 -1146 838 -1112
<< psubdiffcont >>
rect -742 1112 742 1146
rect -838 -1050 -804 1050
rect 804 -1050 838 1050
rect -742 -1146 742 -1112
<< xpolycontact >>
rect -708 584 -426 1016
rect -708 52 -426 484
rect -330 584 -48 1016
rect -330 52 -48 484
rect 48 584 330 1016
rect 48 52 330 484
rect 426 584 708 1016
rect 426 52 708 484
rect -708 -484 -426 -52
rect -708 -1016 -426 -584
rect -330 -484 -48 -52
rect -330 -1016 -48 -584
rect 48 -484 330 -52
rect 48 -1016 330 -584
rect 426 -484 708 -52
rect 426 -1016 708 -584
<< xpolyres >>
rect -708 484 -426 584
rect -330 484 -48 584
rect 48 484 330 584
rect 426 484 708 584
rect -708 -584 -426 -484
rect -330 -584 -48 -484
rect 48 -584 330 -484
rect 426 -584 708 -484
<< locali >>
rect -838 1112 -742 1146
rect 742 1112 838 1146
rect -838 1050 -804 1112
rect 804 1050 838 1112
rect -838 -1112 -804 -1050
rect 804 -1112 838 -1050
rect -838 -1146 -742 -1112
rect 742 -1146 838 -1112
<< viali >>
rect -692 601 -442 998
rect -314 601 -64 998
rect 64 601 314 998
rect 442 601 692 998
rect -692 70 -442 467
rect -314 70 -64 467
rect 64 70 314 467
rect 442 70 692 467
rect -692 -467 -442 -70
rect -314 -467 -64 -70
rect 64 -467 314 -70
rect 442 -467 692 -70
rect -692 -998 -442 -601
rect -314 -998 -64 -601
rect 64 -998 314 -601
rect 442 -998 692 -601
<< metal1 >>
rect -698 998 -436 1010
rect -698 601 -692 998
rect -442 601 -436 998
rect -698 589 -436 601
rect -320 998 -58 1010
rect -320 601 -314 998
rect -64 601 -58 998
rect -320 589 -58 601
rect 58 998 320 1010
rect 58 601 64 998
rect 314 601 320 998
rect 58 589 320 601
rect 436 998 698 1010
rect 436 601 442 998
rect 692 601 698 998
rect 436 589 698 601
rect -698 467 -436 479
rect -698 70 -692 467
rect -442 70 -436 467
rect -698 58 -436 70
rect -320 467 -58 479
rect -320 70 -314 467
rect -64 70 -58 467
rect -320 58 -58 70
rect 58 467 320 479
rect 58 70 64 467
rect 314 70 320 467
rect 58 58 320 70
rect 436 467 698 479
rect 436 70 442 467
rect 692 70 698 467
rect 436 58 698 70
rect -698 -70 -436 -58
rect -698 -467 -692 -70
rect -442 -467 -436 -70
rect -698 -479 -436 -467
rect -320 -70 -58 -58
rect -320 -467 -314 -70
rect -64 -467 -58 -70
rect -320 -479 -58 -467
rect 58 -70 320 -58
rect 58 -467 64 -70
rect 314 -467 320 -70
rect 58 -479 320 -467
rect 436 -70 698 -58
rect 436 -467 442 -70
rect 692 -467 698 -70
rect 436 -479 698 -467
rect -698 -601 -436 -589
rect -698 -998 -692 -601
rect -442 -998 -436 -601
rect -698 -1010 -436 -998
rect -320 -601 -58 -589
rect -320 -998 -314 -601
rect -64 -998 -58 -601
rect -320 -1010 -58 -998
rect 58 -601 320 -589
rect 58 -998 64 -601
rect 314 -998 320 -601
rect 58 -1010 320 -998
rect 436 -601 698 -589
rect 436 -998 442 -601
rect 692 -998 698 -601
rect 436 -1010 698 -998
<< res1p41 >>
rect -710 482 -424 586
rect -332 482 -46 586
rect 46 482 332 586
rect 424 482 710 586
rect -710 -586 -424 -482
rect -332 -586 -46 -482
rect 46 -586 332 -482
rect 424 -586 710 -482
<< properties >>
string FIXED_BBOX -821 -1129 821 1129
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 0.5 m 2 nx 4 wmin 1.410 lmin 0.50 rho 2000 val 976.17 dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
