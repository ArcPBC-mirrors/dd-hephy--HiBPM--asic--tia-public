magic
tech sky130A
timestamp 1699354420
<< end >>
