magic
tech sky130A
magscale 1 2
timestamp 1688995864
<< pwell >>
rect -941 -1646 941 1646
<< nmos >>
rect -745 1036 -545 1436
rect -487 1036 -287 1436
rect -229 1036 -29 1436
rect 29 1036 229 1436
rect 287 1036 487 1436
rect 545 1036 745 1436
rect -745 418 -545 818
rect -487 418 -287 818
rect -229 418 -29 818
rect 29 418 229 818
rect 287 418 487 818
rect 545 418 745 818
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect -745 -818 -545 -418
rect -487 -818 -287 -418
rect -229 -818 -29 -418
rect 29 -818 229 -418
rect 287 -818 487 -418
rect 545 -818 745 -418
rect -745 -1436 -545 -1036
rect -487 -1436 -287 -1036
rect -229 -1436 -29 -1036
rect 29 -1436 229 -1036
rect 287 -1436 487 -1036
rect 545 -1436 745 -1036
<< ndiff >>
rect -803 1424 -745 1436
rect -803 1048 -791 1424
rect -757 1048 -745 1424
rect -803 1036 -745 1048
rect -545 1424 -487 1436
rect -545 1048 -533 1424
rect -499 1048 -487 1424
rect -545 1036 -487 1048
rect -287 1424 -229 1436
rect -287 1048 -275 1424
rect -241 1048 -229 1424
rect -287 1036 -229 1048
rect -29 1424 29 1436
rect -29 1048 -17 1424
rect 17 1048 29 1424
rect -29 1036 29 1048
rect 229 1424 287 1436
rect 229 1048 241 1424
rect 275 1048 287 1424
rect 229 1036 287 1048
rect 487 1424 545 1436
rect 487 1048 499 1424
rect 533 1048 545 1424
rect 487 1036 545 1048
rect 745 1424 803 1436
rect 745 1048 757 1424
rect 791 1048 803 1424
rect 745 1036 803 1048
rect -803 806 -745 818
rect -803 430 -791 806
rect -757 430 -745 806
rect -803 418 -745 430
rect -545 806 -487 818
rect -545 430 -533 806
rect -499 430 -487 806
rect -545 418 -487 430
rect -287 806 -229 818
rect -287 430 -275 806
rect -241 430 -229 806
rect -287 418 -229 430
rect -29 806 29 818
rect -29 430 -17 806
rect 17 430 29 806
rect -29 418 29 430
rect 229 806 287 818
rect 229 430 241 806
rect 275 430 287 806
rect 229 418 287 430
rect 487 806 545 818
rect 487 430 499 806
rect 533 430 545 806
rect 487 418 545 430
rect 745 806 803 818
rect 745 430 757 806
rect 791 430 803 806
rect 745 418 803 430
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect -803 -430 -745 -418
rect -803 -806 -791 -430
rect -757 -806 -745 -430
rect -803 -818 -745 -806
rect -545 -430 -487 -418
rect -545 -806 -533 -430
rect -499 -806 -487 -430
rect -545 -818 -487 -806
rect -287 -430 -229 -418
rect -287 -806 -275 -430
rect -241 -806 -229 -430
rect -287 -818 -229 -806
rect -29 -430 29 -418
rect -29 -806 -17 -430
rect 17 -806 29 -430
rect -29 -818 29 -806
rect 229 -430 287 -418
rect 229 -806 241 -430
rect 275 -806 287 -430
rect 229 -818 287 -806
rect 487 -430 545 -418
rect 487 -806 499 -430
rect 533 -806 545 -430
rect 487 -818 545 -806
rect 745 -430 803 -418
rect 745 -806 757 -430
rect 791 -806 803 -430
rect 745 -818 803 -806
rect -803 -1048 -745 -1036
rect -803 -1424 -791 -1048
rect -757 -1424 -745 -1048
rect -803 -1436 -745 -1424
rect -545 -1048 -487 -1036
rect -545 -1424 -533 -1048
rect -499 -1424 -487 -1048
rect -545 -1436 -487 -1424
rect -287 -1048 -229 -1036
rect -287 -1424 -275 -1048
rect -241 -1424 -229 -1048
rect -287 -1436 -229 -1424
rect -29 -1048 29 -1036
rect -29 -1424 -17 -1048
rect 17 -1424 29 -1048
rect -29 -1436 29 -1424
rect 229 -1048 287 -1036
rect 229 -1424 241 -1048
rect 275 -1424 287 -1048
rect 229 -1436 287 -1424
rect 487 -1048 545 -1036
rect 487 -1424 499 -1048
rect 533 -1424 545 -1048
rect 487 -1436 545 -1424
rect 745 -1048 803 -1036
rect 745 -1424 757 -1048
rect 791 -1424 803 -1048
rect 745 -1436 803 -1424
<< ndiffc >>
rect -791 1048 -757 1424
rect -533 1048 -499 1424
rect -275 1048 -241 1424
rect -17 1048 17 1424
rect 241 1048 275 1424
rect 499 1048 533 1424
rect 757 1048 791 1424
rect -791 430 -757 806
rect -533 430 -499 806
rect -275 430 -241 806
rect -17 430 17 806
rect 241 430 275 806
rect 499 430 533 806
rect 757 430 791 806
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect -791 -806 -757 -430
rect -533 -806 -499 -430
rect -275 -806 -241 -430
rect -17 -806 17 -430
rect 241 -806 275 -430
rect 499 -806 533 -430
rect 757 -806 791 -430
rect -791 -1424 -757 -1048
rect -533 -1424 -499 -1048
rect -275 -1424 -241 -1048
rect -17 -1424 17 -1048
rect 241 -1424 275 -1048
rect 499 -1424 533 -1048
rect 757 -1424 791 -1048
<< psubdiff >>
rect -905 1576 -809 1610
rect 809 1576 905 1610
rect -905 1514 -871 1576
rect 871 1514 905 1576
rect -905 -1576 -871 -1514
rect 871 -1576 905 -1514
rect -905 -1610 -809 -1576
rect 809 -1610 905 -1576
<< psubdiffcont >>
rect -809 1576 809 1610
rect -905 -1514 -871 1514
rect 871 -1514 905 1514
rect -809 -1610 809 -1576
<< poly >>
rect -745 1508 -545 1524
rect -745 1474 -729 1508
rect -561 1474 -545 1508
rect -745 1436 -545 1474
rect -487 1508 -287 1524
rect -487 1474 -471 1508
rect -303 1474 -287 1508
rect -487 1436 -287 1474
rect -229 1508 -29 1524
rect -229 1474 -213 1508
rect -45 1474 -29 1508
rect -229 1436 -29 1474
rect 29 1508 229 1524
rect 29 1474 45 1508
rect 213 1474 229 1508
rect 29 1436 229 1474
rect 287 1508 487 1524
rect 287 1474 303 1508
rect 471 1474 487 1508
rect 287 1436 487 1474
rect 545 1508 745 1524
rect 545 1474 561 1508
rect 729 1474 745 1508
rect 545 1436 745 1474
rect -745 998 -545 1036
rect -745 964 -729 998
rect -561 964 -545 998
rect -745 948 -545 964
rect -487 998 -287 1036
rect -487 964 -471 998
rect -303 964 -287 998
rect -487 948 -287 964
rect -229 998 -29 1036
rect -229 964 -213 998
rect -45 964 -29 998
rect -229 948 -29 964
rect 29 998 229 1036
rect 29 964 45 998
rect 213 964 229 998
rect 29 948 229 964
rect 287 998 487 1036
rect 287 964 303 998
rect 471 964 487 998
rect 287 948 487 964
rect 545 998 745 1036
rect 545 964 561 998
rect 729 964 745 998
rect 545 948 745 964
rect -745 890 -545 906
rect -745 856 -729 890
rect -561 856 -545 890
rect -745 818 -545 856
rect -487 890 -287 906
rect -487 856 -471 890
rect -303 856 -287 890
rect -487 818 -287 856
rect -229 890 -29 906
rect -229 856 -213 890
rect -45 856 -29 890
rect -229 818 -29 856
rect 29 890 229 906
rect 29 856 45 890
rect 213 856 229 890
rect 29 818 229 856
rect 287 890 487 906
rect 287 856 303 890
rect 471 856 487 890
rect 287 818 487 856
rect 545 890 745 906
rect 545 856 561 890
rect 729 856 745 890
rect 545 818 745 856
rect -745 380 -545 418
rect -745 346 -729 380
rect -561 346 -545 380
rect -745 330 -545 346
rect -487 380 -287 418
rect -487 346 -471 380
rect -303 346 -287 380
rect -487 330 -287 346
rect -229 380 -29 418
rect -229 346 -213 380
rect -45 346 -29 380
rect -229 330 -29 346
rect 29 380 229 418
rect 29 346 45 380
rect 213 346 229 380
rect 29 330 229 346
rect 287 380 487 418
rect 287 346 303 380
rect 471 346 487 380
rect 287 330 487 346
rect 545 380 745 418
rect 545 346 561 380
rect 729 346 745 380
rect 545 330 745 346
rect -745 272 -545 288
rect -745 238 -729 272
rect -561 238 -545 272
rect -745 200 -545 238
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect 545 272 745 288
rect 545 238 561 272
rect 729 238 745 272
rect 545 200 745 238
rect -745 -238 -545 -200
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -745 -288 -545 -272
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
rect 545 -238 745 -200
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 545 -288 745 -272
rect -745 -346 -545 -330
rect -745 -380 -729 -346
rect -561 -380 -545 -346
rect -745 -418 -545 -380
rect -487 -346 -287 -330
rect -487 -380 -471 -346
rect -303 -380 -287 -346
rect -487 -418 -287 -380
rect -229 -346 -29 -330
rect -229 -380 -213 -346
rect -45 -380 -29 -346
rect -229 -418 -29 -380
rect 29 -346 229 -330
rect 29 -380 45 -346
rect 213 -380 229 -346
rect 29 -418 229 -380
rect 287 -346 487 -330
rect 287 -380 303 -346
rect 471 -380 487 -346
rect 287 -418 487 -380
rect 545 -346 745 -330
rect 545 -380 561 -346
rect 729 -380 745 -346
rect 545 -418 745 -380
rect -745 -856 -545 -818
rect -745 -890 -729 -856
rect -561 -890 -545 -856
rect -745 -906 -545 -890
rect -487 -856 -287 -818
rect -487 -890 -471 -856
rect -303 -890 -287 -856
rect -487 -906 -287 -890
rect -229 -856 -29 -818
rect -229 -890 -213 -856
rect -45 -890 -29 -856
rect -229 -906 -29 -890
rect 29 -856 229 -818
rect 29 -890 45 -856
rect 213 -890 229 -856
rect 29 -906 229 -890
rect 287 -856 487 -818
rect 287 -890 303 -856
rect 471 -890 487 -856
rect 287 -906 487 -890
rect 545 -856 745 -818
rect 545 -890 561 -856
rect 729 -890 745 -856
rect 545 -906 745 -890
rect -745 -964 -545 -948
rect -745 -998 -729 -964
rect -561 -998 -545 -964
rect -745 -1036 -545 -998
rect -487 -964 -287 -948
rect -487 -998 -471 -964
rect -303 -998 -287 -964
rect -487 -1036 -287 -998
rect -229 -964 -29 -948
rect -229 -998 -213 -964
rect -45 -998 -29 -964
rect -229 -1036 -29 -998
rect 29 -964 229 -948
rect 29 -998 45 -964
rect 213 -998 229 -964
rect 29 -1036 229 -998
rect 287 -964 487 -948
rect 287 -998 303 -964
rect 471 -998 487 -964
rect 287 -1036 487 -998
rect 545 -964 745 -948
rect 545 -998 561 -964
rect 729 -998 745 -964
rect 545 -1036 745 -998
rect -745 -1474 -545 -1436
rect -745 -1508 -729 -1474
rect -561 -1508 -545 -1474
rect -745 -1524 -545 -1508
rect -487 -1474 -287 -1436
rect -487 -1508 -471 -1474
rect -303 -1508 -287 -1474
rect -487 -1524 -287 -1508
rect -229 -1474 -29 -1436
rect -229 -1508 -213 -1474
rect -45 -1508 -29 -1474
rect -229 -1524 -29 -1508
rect 29 -1474 229 -1436
rect 29 -1508 45 -1474
rect 213 -1508 229 -1474
rect 29 -1524 229 -1508
rect 287 -1474 487 -1436
rect 287 -1508 303 -1474
rect 471 -1508 487 -1474
rect 287 -1524 487 -1508
rect 545 -1474 745 -1436
rect 545 -1508 561 -1474
rect 729 -1508 745 -1474
rect 545 -1524 745 -1508
<< polycont >>
rect -729 1474 -561 1508
rect -471 1474 -303 1508
rect -213 1474 -45 1508
rect 45 1474 213 1508
rect 303 1474 471 1508
rect 561 1474 729 1508
rect -729 964 -561 998
rect -471 964 -303 998
rect -213 964 -45 998
rect 45 964 213 998
rect 303 964 471 998
rect 561 964 729 998
rect -729 856 -561 890
rect -471 856 -303 890
rect -213 856 -45 890
rect 45 856 213 890
rect 303 856 471 890
rect 561 856 729 890
rect -729 346 -561 380
rect -471 346 -303 380
rect -213 346 -45 380
rect 45 346 213 380
rect 303 346 471 380
rect 561 346 729 380
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect -729 -380 -561 -346
rect -471 -380 -303 -346
rect -213 -380 -45 -346
rect 45 -380 213 -346
rect 303 -380 471 -346
rect 561 -380 729 -346
rect -729 -890 -561 -856
rect -471 -890 -303 -856
rect -213 -890 -45 -856
rect 45 -890 213 -856
rect 303 -890 471 -856
rect 561 -890 729 -856
rect -729 -998 -561 -964
rect -471 -998 -303 -964
rect -213 -998 -45 -964
rect 45 -998 213 -964
rect 303 -998 471 -964
rect 561 -998 729 -964
rect -729 -1508 -561 -1474
rect -471 -1508 -303 -1474
rect -213 -1508 -45 -1474
rect 45 -1508 213 -1474
rect 303 -1508 471 -1474
rect 561 -1508 729 -1474
<< locali >>
rect -905 1576 -809 1610
rect 809 1576 905 1610
rect -905 1514 -871 1576
rect 871 1514 905 1576
rect -745 1474 -729 1508
rect -561 1474 -545 1508
rect -487 1474 -471 1508
rect -303 1474 -287 1508
rect -229 1474 -213 1508
rect -45 1474 -29 1508
rect 29 1474 45 1508
rect 213 1474 229 1508
rect 287 1474 303 1508
rect 471 1474 487 1508
rect 545 1474 561 1508
rect 729 1474 745 1508
rect -791 1424 -757 1440
rect -791 1032 -757 1048
rect -533 1424 -499 1440
rect -533 1032 -499 1048
rect -275 1424 -241 1440
rect -275 1032 -241 1048
rect -17 1424 17 1440
rect -17 1032 17 1048
rect 241 1424 275 1440
rect 241 1032 275 1048
rect 499 1424 533 1440
rect 499 1032 533 1048
rect 757 1424 791 1440
rect 757 1032 791 1048
rect -745 964 -729 998
rect -561 964 -545 998
rect -487 964 -471 998
rect -303 964 -287 998
rect -229 964 -213 998
rect -45 964 -29 998
rect 29 964 45 998
rect 213 964 229 998
rect 287 964 303 998
rect 471 964 487 998
rect 545 964 561 998
rect 729 964 745 998
rect -745 856 -729 890
rect -561 856 -545 890
rect -487 856 -471 890
rect -303 856 -287 890
rect -229 856 -213 890
rect -45 856 -29 890
rect 29 856 45 890
rect 213 856 229 890
rect 287 856 303 890
rect 471 856 487 890
rect 545 856 561 890
rect 729 856 745 890
rect -791 806 -757 822
rect -791 414 -757 430
rect -533 806 -499 822
rect -533 414 -499 430
rect -275 806 -241 822
rect -275 414 -241 430
rect -17 806 17 822
rect -17 414 17 430
rect 241 806 275 822
rect 241 414 275 430
rect 499 806 533 822
rect 499 414 533 430
rect 757 806 791 822
rect 757 414 791 430
rect -745 346 -729 380
rect -561 346 -545 380
rect -487 346 -471 380
rect -303 346 -287 380
rect -229 346 -213 380
rect -45 346 -29 380
rect 29 346 45 380
rect 213 346 229 380
rect 287 346 303 380
rect 471 346 487 380
rect 545 346 561 380
rect 729 346 745 380
rect -745 238 -729 272
rect -561 238 -545 272
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect 545 238 561 272
rect 729 238 745 272
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 545 -272 561 -238
rect 729 -272 745 -238
rect -745 -380 -729 -346
rect -561 -380 -545 -346
rect -487 -380 -471 -346
rect -303 -380 -287 -346
rect -229 -380 -213 -346
rect -45 -380 -29 -346
rect 29 -380 45 -346
rect 213 -380 229 -346
rect 287 -380 303 -346
rect 471 -380 487 -346
rect 545 -380 561 -346
rect 729 -380 745 -346
rect -791 -430 -757 -414
rect -791 -822 -757 -806
rect -533 -430 -499 -414
rect -533 -822 -499 -806
rect -275 -430 -241 -414
rect -275 -822 -241 -806
rect -17 -430 17 -414
rect -17 -822 17 -806
rect 241 -430 275 -414
rect 241 -822 275 -806
rect 499 -430 533 -414
rect 499 -822 533 -806
rect 757 -430 791 -414
rect 757 -822 791 -806
rect -745 -890 -729 -856
rect -561 -890 -545 -856
rect -487 -890 -471 -856
rect -303 -890 -287 -856
rect -229 -890 -213 -856
rect -45 -890 -29 -856
rect 29 -890 45 -856
rect 213 -890 229 -856
rect 287 -890 303 -856
rect 471 -890 487 -856
rect 545 -890 561 -856
rect 729 -890 745 -856
rect -745 -998 -729 -964
rect -561 -998 -545 -964
rect -487 -998 -471 -964
rect -303 -998 -287 -964
rect -229 -998 -213 -964
rect -45 -998 -29 -964
rect 29 -998 45 -964
rect 213 -998 229 -964
rect 287 -998 303 -964
rect 471 -998 487 -964
rect 545 -998 561 -964
rect 729 -998 745 -964
rect -791 -1048 -757 -1032
rect -791 -1440 -757 -1424
rect -533 -1048 -499 -1032
rect -533 -1440 -499 -1424
rect -275 -1048 -241 -1032
rect -275 -1440 -241 -1424
rect -17 -1048 17 -1032
rect -17 -1440 17 -1424
rect 241 -1048 275 -1032
rect 241 -1440 275 -1424
rect 499 -1048 533 -1032
rect 499 -1440 533 -1424
rect 757 -1048 791 -1032
rect 757 -1440 791 -1424
rect -745 -1508 -729 -1474
rect -561 -1508 -545 -1474
rect -487 -1508 -471 -1474
rect -303 -1508 -287 -1474
rect -229 -1508 -213 -1474
rect -45 -1508 -29 -1474
rect 29 -1508 45 -1474
rect 213 -1508 229 -1474
rect 287 -1508 303 -1474
rect 471 -1508 487 -1474
rect 545 -1508 561 -1474
rect 729 -1508 745 -1474
rect -905 -1576 -871 -1514
rect 871 -1576 905 -1514
rect -905 -1610 -809 -1576
rect 809 -1610 905 -1576
<< viali >>
rect -729 1474 -561 1508
rect -471 1474 -303 1508
rect -213 1474 -45 1508
rect 45 1474 213 1508
rect 303 1474 471 1508
rect 561 1474 729 1508
rect -791 1048 -757 1424
rect -533 1048 -499 1424
rect -275 1048 -241 1424
rect -17 1048 17 1424
rect 241 1048 275 1424
rect 499 1048 533 1424
rect 757 1048 791 1424
rect -729 964 -561 998
rect -471 964 -303 998
rect -213 964 -45 998
rect 45 964 213 998
rect 303 964 471 998
rect 561 964 729 998
rect -729 856 -561 890
rect -471 856 -303 890
rect -213 856 -45 890
rect 45 856 213 890
rect 303 856 471 890
rect 561 856 729 890
rect -791 430 -757 806
rect -533 430 -499 806
rect -275 430 -241 806
rect -17 430 17 806
rect 241 430 275 806
rect 499 430 533 806
rect 757 430 791 806
rect -729 346 -561 380
rect -471 346 -303 380
rect -213 346 -45 380
rect 45 346 213 380
rect 303 346 471 380
rect 561 346 729 380
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect -729 -380 -561 -346
rect -471 -380 -303 -346
rect -213 -380 -45 -346
rect 45 -380 213 -346
rect 303 -380 471 -346
rect 561 -380 729 -346
rect -791 -806 -757 -430
rect -533 -806 -499 -430
rect -275 -806 -241 -430
rect -17 -806 17 -430
rect 241 -806 275 -430
rect 499 -806 533 -430
rect 757 -806 791 -430
rect -729 -890 -561 -856
rect -471 -890 -303 -856
rect -213 -890 -45 -856
rect 45 -890 213 -856
rect 303 -890 471 -856
rect 561 -890 729 -856
rect -729 -998 -561 -964
rect -471 -998 -303 -964
rect -213 -998 -45 -964
rect 45 -998 213 -964
rect 303 -998 471 -964
rect 561 -998 729 -964
rect -791 -1424 -757 -1048
rect -533 -1424 -499 -1048
rect -275 -1424 -241 -1048
rect -17 -1424 17 -1048
rect 241 -1424 275 -1048
rect 499 -1424 533 -1048
rect 757 -1424 791 -1048
rect -729 -1508 -561 -1474
rect -471 -1508 -303 -1474
rect -213 -1508 -45 -1474
rect 45 -1508 213 -1474
rect 303 -1508 471 -1474
rect 561 -1508 729 -1474
<< metal1 >>
rect -741 1508 -549 1514
rect -741 1474 -729 1508
rect -561 1474 -549 1508
rect -741 1468 -549 1474
rect -483 1508 -291 1514
rect -483 1474 -471 1508
rect -303 1474 -291 1508
rect -483 1468 -291 1474
rect -225 1508 -33 1514
rect -225 1474 -213 1508
rect -45 1474 -33 1508
rect -225 1468 -33 1474
rect 33 1508 225 1514
rect 33 1474 45 1508
rect 213 1474 225 1508
rect 33 1468 225 1474
rect 291 1508 483 1514
rect 291 1474 303 1508
rect 471 1474 483 1508
rect 291 1468 483 1474
rect 549 1508 741 1514
rect 549 1474 561 1508
rect 729 1474 741 1508
rect 549 1468 741 1474
rect -797 1424 -751 1436
rect -797 1048 -791 1424
rect -757 1048 -751 1424
rect -797 1036 -751 1048
rect -539 1424 -493 1436
rect -539 1048 -533 1424
rect -499 1048 -493 1424
rect -539 1036 -493 1048
rect -281 1424 -235 1436
rect -281 1048 -275 1424
rect -241 1048 -235 1424
rect -281 1036 -235 1048
rect -23 1424 23 1436
rect -23 1048 -17 1424
rect 17 1048 23 1424
rect -23 1036 23 1048
rect 235 1424 281 1436
rect 235 1048 241 1424
rect 275 1048 281 1424
rect 235 1036 281 1048
rect 493 1424 539 1436
rect 493 1048 499 1424
rect 533 1048 539 1424
rect 493 1036 539 1048
rect 751 1424 797 1436
rect 751 1048 757 1424
rect 791 1048 797 1424
rect 751 1036 797 1048
rect -741 998 -549 1004
rect -741 964 -729 998
rect -561 964 -549 998
rect -741 958 -549 964
rect -483 998 -291 1004
rect -483 964 -471 998
rect -303 964 -291 998
rect -483 958 -291 964
rect -225 998 -33 1004
rect -225 964 -213 998
rect -45 964 -33 998
rect -225 958 -33 964
rect 33 998 225 1004
rect 33 964 45 998
rect 213 964 225 998
rect 33 958 225 964
rect 291 998 483 1004
rect 291 964 303 998
rect 471 964 483 998
rect 291 958 483 964
rect 549 998 741 1004
rect 549 964 561 998
rect 729 964 741 998
rect 549 958 741 964
rect -741 890 -549 896
rect -741 856 -729 890
rect -561 856 -549 890
rect -741 850 -549 856
rect -483 890 -291 896
rect -483 856 -471 890
rect -303 856 -291 890
rect -483 850 -291 856
rect -225 890 -33 896
rect -225 856 -213 890
rect -45 856 -33 890
rect -225 850 -33 856
rect 33 890 225 896
rect 33 856 45 890
rect 213 856 225 890
rect 33 850 225 856
rect 291 890 483 896
rect 291 856 303 890
rect 471 856 483 890
rect 291 850 483 856
rect 549 890 741 896
rect 549 856 561 890
rect 729 856 741 890
rect 549 850 741 856
rect -797 806 -751 818
rect -797 430 -791 806
rect -757 430 -751 806
rect -797 418 -751 430
rect -539 806 -493 818
rect -539 430 -533 806
rect -499 430 -493 806
rect -539 418 -493 430
rect -281 806 -235 818
rect -281 430 -275 806
rect -241 430 -235 806
rect -281 418 -235 430
rect -23 806 23 818
rect -23 430 -17 806
rect 17 430 23 806
rect -23 418 23 430
rect 235 806 281 818
rect 235 430 241 806
rect 275 430 281 806
rect 235 418 281 430
rect 493 806 539 818
rect 493 430 499 806
rect 533 430 539 806
rect 493 418 539 430
rect 751 806 797 818
rect 751 430 757 806
rect 791 430 797 806
rect 751 418 797 430
rect -741 380 -549 386
rect -741 346 -729 380
rect -561 346 -549 380
rect -741 340 -549 346
rect -483 380 -291 386
rect -483 346 -471 380
rect -303 346 -291 380
rect -483 340 -291 346
rect -225 380 -33 386
rect -225 346 -213 380
rect -45 346 -33 380
rect -225 340 -33 346
rect 33 380 225 386
rect 33 346 45 380
rect 213 346 225 380
rect 33 340 225 346
rect 291 380 483 386
rect 291 346 303 380
rect 471 346 483 380
rect 291 340 483 346
rect 549 380 741 386
rect 549 346 561 380
rect 729 346 741 380
rect 549 340 741 346
rect -741 272 -549 278
rect -741 238 -729 272
rect -561 238 -549 272
rect -741 232 -549 238
rect -483 272 -291 278
rect -483 238 -471 272
rect -303 238 -291 272
rect -483 232 -291 238
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect 291 272 483 278
rect 291 238 303 272
rect 471 238 483 272
rect 291 232 483 238
rect 549 272 741 278
rect 549 238 561 272
rect 729 238 741 272
rect 549 232 741 238
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect -741 -238 -549 -232
rect -741 -272 -729 -238
rect -561 -272 -549 -238
rect -741 -278 -549 -272
rect -483 -238 -291 -232
rect -483 -272 -471 -238
rect -303 -272 -291 -238
rect -483 -278 -291 -272
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
rect 291 -238 483 -232
rect 291 -272 303 -238
rect 471 -272 483 -238
rect 291 -278 483 -272
rect 549 -238 741 -232
rect 549 -272 561 -238
rect 729 -272 741 -238
rect 549 -278 741 -272
rect -741 -346 -549 -340
rect -741 -380 -729 -346
rect -561 -380 -549 -346
rect -741 -386 -549 -380
rect -483 -346 -291 -340
rect -483 -380 -471 -346
rect -303 -380 -291 -346
rect -483 -386 -291 -380
rect -225 -346 -33 -340
rect -225 -380 -213 -346
rect -45 -380 -33 -346
rect -225 -386 -33 -380
rect 33 -346 225 -340
rect 33 -380 45 -346
rect 213 -380 225 -346
rect 33 -386 225 -380
rect 291 -346 483 -340
rect 291 -380 303 -346
rect 471 -380 483 -346
rect 291 -386 483 -380
rect 549 -346 741 -340
rect 549 -380 561 -346
rect 729 -380 741 -346
rect 549 -386 741 -380
rect -797 -430 -751 -418
rect -797 -806 -791 -430
rect -757 -806 -751 -430
rect -797 -818 -751 -806
rect -539 -430 -493 -418
rect -539 -806 -533 -430
rect -499 -806 -493 -430
rect -539 -818 -493 -806
rect -281 -430 -235 -418
rect -281 -806 -275 -430
rect -241 -806 -235 -430
rect -281 -818 -235 -806
rect -23 -430 23 -418
rect -23 -806 -17 -430
rect 17 -806 23 -430
rect -23 -818 23 -806
rect 235 -430 281 -418
rect 235 -806 241 -430
rect 275 -806 281 -430
rect 235 -818 281 -806
rect 493 -430 539 -418
rect 493 -806 499 -430
rect 533 -806 539 -430
rect 493 -818 539 -806
rect 751 -430 797 -418
rect 751 -806 757 -430
rect 791 -806 797 -430
rect 751 -818 797 -806
rect -741 -856 -549 -850
rect -741 -890 -729 -856
rect -561 -890 -549 -856
rect -741 -896 -549 -890
rect -483 -856 -291 -850
rect -483 -890 -471 -856
rect -303 -890 -291 -856
rect -483 -896 -291 -890
rect -225 -856 -33 -850
rect -225 -890 -213 -856
rect -45 -890 -33 -856
rect -225 -896 -33 -890
rect 33 -856 225 -850
rect 33 -890 45 -856
rect 213 -890 225 -856
rect 33 -896 225 -890
rect 291 -856 483 -850
rect 291 -890 303 -856
rect 471 -890 483 -856
rect 291 -896 483 -890
rect 549 -856 741 -850
rect 549 -890 561 -856
rect 729 -890 741 -856
rect 549 -896 741 -890
rect -741 -964 -549 -958
rect -741 -998 -729 -964
rect -561 -998 -549 -964
rect -741 -1004 -549 -998
rect -483 -964 -291 -958
rect -483 -998 -471 -964
rect -303 -998 -291 -964
rect -483 -1004 -291 -998
rect -225 -964 -33 -958
rect -225 -998 -213 -964
rect -45 -998 -33 -964
rect -225 -1004 -33 -998
rect 33 -964 225 -958
rect 33 -998 45 -964
rect 213 -998 225 -964
rect 33 -1004 225 -998
rect 291 -964 483 -958
rect 291 -998 303 -964
rect 471 -998 483 -964
rect 291 -1004 483 -998
rect 549 -964 741 -958
rect 549 -998 561 -964
rect 729 -998 741 -964
rect 549 -1004 741 -998
rect -797 -1048 -751 -1036
rect -797 -1424 -791 -1048
rect -757 -1424 -751 -1048
rect -797 -1436 -751 -1424
rect -539 -1048 -493 -1036
rect -539 -1424 -533 -1048
rect -499 -1424 -493 -1048
rect -539 -1436 -493 -1424
rect -281 -1048 -235 -1036
rect -281 -1424 -275 -1048
rect -241 -1424 -235 -1048
rect -281 -1436 -235 -1424
rect -23 -1048 23 -1036
rect -23 -1424 -17 -1048
rect 17 -1424 23 -1048
rect -23 -1436 23 -1424
rect 235 -1048 281 -1036
rect 235 -1424 241 -1048
rect 275 -1424 281 -1048
rect 235 -1436 281 -1424
rect 493 -1048 539 -1036
rect 493 -1424 499 -1048
rect 533 -1424 539 -1048
rect 493 -1436 539 -1424
rect 751 -1048 797 -1036
rect 751 -1424 757 -1048
rect 791 -1424 797 -1048
rect 751 -1436 797 -1424
rect -741 -1474 -549 -1468
rect -741 -1508 -729 -1474
rect -561 -1508 -549 -1474
rect -741 -1514 -549 -1508
rect -483 -1474 -291 -1468
rect -483 -1508 -471 -1474
rect -303 -1508 -291 -1474
rect -483 -1514 -291 -1508
rect -225 -1474 -33 -1468
rect -225 -1508 -213 -1474
rect -45 -1508 -33 -1474
rect -225 -1514 -33 -1508
rect 33 -1474 225 -1468
rect 33 -1508 45 -1474
rect 213 -1508 225 -1474
rect 33 -1514 225 -1508
rect 291 -1474 483 -1468
rect 291 -1508 303 -1474
rect 471 -1508 483 -1474
rect 291 -1514 483 -1508
rect 549 -1474 741 -1468
rect 549 -1508 561 -1474
rect 729 -1508 741 -1474
rect 549 -1514 741 -1508
<< properties >>
string FIXED_BBOX -888 -1593 888 1593
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 5 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
