magic
tech sky130A
magscale 1 2
timestamp 1688995864
<< error_p >>
rect 182 1918 240 1924
rect 374 1918 432 1924
rect 566 1918 624 1924
rect 758 1918 816 1924
rect 950 1918 1008 1924
rect 182 1884 194 1918
rect 374 1884 386 1918
rect 566 1884 578 1918
rect 758 1884 770 1918
rect 950 1884 962 1918
rect 182 1878 240 1884
rect 374 1878 432 1884
rect 566 1878 624 1884
rect 758 1878 816 1884
rect 950 1878 1008 1884
rect 86 1408 144 1414
rect 278 1408 336 1414
rect 470 1408 528 1414
rect 662 1408 720 1414
rect 854 1408 912 1414
rect 86 1374 98 1408
rect 278 1374 290 1408
rect 470 1374 482 1408
rect 662 1374 674 1408
rect 854 1374 866 1408
rect 86 1368 144 1374
rect 278 1368 336 1374
rect 470 1368 528 1374
rect 662 1368 720 1374
rect 854 1368 912 1374
rect 86 1300 144 1306
rect 278 1300 336 1306
rect 470 1300 528 1306
rect 662 1300 720 1306
rect 854 1300 912 1306
rect 86 1266 98 1300
rect 278 1266 290 1300
rect 470 1266 482 1300
rect 662 1266 674 1300
rect 854 1266 866 1300
rect 86 1260 144 1266
rect 278 1260 336 1266
rect 470 1260 528 1266
rect 662 1260 720 1266
rect 854 1260 912 1266
<< error_s >>
rect 182 790 240 796
rect 374 790 432 796
rect 566 790 624 796
rect 758 790 816 796
rect 950 790 1008 796
rect 182 756 194 790
rect 374 756 386 790
rect 566 756 578 790
rect 758 756 770 790
rect 950 756 962 790
rect 182 750 240 756
rect 374 750 432 756
rect 566 750 624 756
rect 758 750 816 756
rect 950 750 1008 756
rect 182 682 240 688
rect 374 682 432 688
rect 566 682 624 688
rect 758 682 816 688
rect 950 682 1008 688
rect 182 648 194 682
rect 374 648 386 682
rect 566 648 578 682
rect 758 648 770 682
rect 950 648 962 682
rect 182 642 240 648
rect 374 642 432 648
rect 566 642 624 648
rect 758 642 816 648
rect 950 642 1008 648
rect 86 172 144 178
rect 278 172 336 178
rect 470 172 528 178
rect 662 172 720 178
rect 854 172 912 178
rect 86 138 98 172
rect 278 138 290 172
rect 470 138 482 172
rect 662 138 674 172
rect 854 138 866 172
rect 86 132 144 138
rect 278 132 336 138
rect 470 132 528 138
rect 662 132 720 138
rect 854 132 912 138
use sky130_fd_pr__nfet_01v8_lvt_R2KHEY  sky130_fd_pr__nfet_01v8_lvt_R2KHEY_0
timestamp 1688995864
transform 1 0 547 0 1 1028
box -647 -1028 647 1028
use sky130_fd_pr__nfet_01v8_URJU67  sky130_fd_pr__nfet_01v8_URJU67_0
timestamp 1688995864
transform 1 0 841 0 1 -1654
box -941 -1646 941 1646
<< end >>
