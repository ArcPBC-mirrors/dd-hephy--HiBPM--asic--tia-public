magic
tech sky130A
magscale 1 2
timestamp 1683810998
<< pwell >>
rect -8457 -519 8457 519
<< nmoslvt >>
rect -8261 109 -6661 309
rect -6603 109 -5003 309
rect -4945 109 -3345 309
rect -3287 109 -1687 309
rect -1629 109 -29 309
rect 29 109 1629 309
rect 1687 109 3287 309
rect 3345 109 4945 309
rect 5003 109 6603 309
rect 6661 109 8261 309
rect -8261 -309 -6661 -109
rect -6603 -309 -5003 -109
rect -4945 -309 -3345 -109
rect -3287 -309 -1687 -109
rect -1629 -309 -29 -109
rect 29 -309 1629 -109
rect 1687 -309 3287 -109
rect 3345 -309 4945 -109
rect 5003 -309 6603 -109
rect 6661 -309 8261 -109
<< ndiff >>
rect -8319 297 -8261 309
rect -8319 121 -8307 297
rect -8273 121 -8261 297
rect -8319 109 -8261 121
rect -6661 297 -6603 309
rect -6661 121 -6649 297
rect -6615 121 -6603 297
rect -6661 109 -6603 121
rect -5003 297 -4945 309
rect -5003 121 -4991 297
rect -4957 121 -4945 297
rect -5003 109 -4945 121
rect -3345 297 -3287 309
rect -3345 121 -3333 297
rect -3299 121 -3287 297
rect -3345 109 -3287 121
rect -1687 297 -1629 309
rect -1687 121 -1675 297
rect -1641 121 -1629 297
rect -1687 109 -1629 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 1629 297 1687 309
rect 1629 121 1641 297
rect 1675 121 1687 297
rect 1629 109 1687 121
rect 3287 297 3345 309
rect 3287 121 3299 297
rect 3333 121 3345 297
rect 3287 109 3345 121
rect 4945 297 5003 309
rect 4945 121 4957 297
rect 4991 121 5003 297
rect 4945 109 5003 121
rect 6603 297 6661 309
rect 6603 121 6615 297
rect 6649 121 6661 297
rect 6603 109 6661 121
rect 8261 297 8319 309
rect 8261 121 8273 297
rect 8307 121 8319 297
rect 8261 109 8319 121
rect -8319 -121 -8261 -109
rect -8319 -297 -8307 -121
rect -8273 -297 -8261 -121
rect -8319 -309 -8261 -297
rect -6661 -121 -6603 -109
rect -6661 -297 -6649 -121
rect -6615 -297 -6603 -121
rect -6661 -309 -6603 -297
rect -5003 -121 -4945 -109
rect -5003 -297 -4991 -121
rect -4957 -297 -4945 -121
rect -5003 -309 -4945 -297
rect -3345 -121 -3287 -109
rect -3345 -297 -3333 -121
rect -3299 -297 -3287 -121
rect -3345 -309 -3287 -297
rect -1687 -121 -1629 -109
rect -1687 -297 -1675 -121
rect -1641 -297 -1629 -121
rect -1687 -309 -1629 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 1629 -121 1687 -109
rect 1629 -297 1641 -121
rect 1675 -297 1687 -121
rect 1629 -309 1687 -297
rect 3287 -121 3345 -109
rect 3287 -297 3299 -121
rect 3333 -297 3345 -121
rect 3287 -309 3345 -297
rect 4945 -121 5003 -109
rect 4945 -297 4957 -121
rect 4991 -297 5003 -121
rect 4945 -309 5003 -297
rect 6603 -121 6661 -109
rect 6603 -297 6615 -121
rect 6649 -297 6661 -121
rect 6603 -309 6661 -297
rect 8261 -121 8319 -109
rect 8261 -297 8273 -121
rect 8307 -297 8319 -121
rect 8261 -309 8319 -297
<< ndiffc >>
rect -8307 121 -8273 297
rect -6649 121 -6615 297
rect -4991 121 -4957 297
rect -3333 121 -3299 297
rect -1675 121 -1641 297
rect -17 121 17 297
rect 1641 121 1675 297
rect 3299 121 3333 297
rect 4957 121 4991 297
rect 6615 121 6649 297
rect 8273 121 8307 297
rect -8307 -297 -8273 -121
rect -6649 -297 -6615 -121
rect -4991 -297 -4957 -121
rect -3333 -297 -3299 -121
rect -1675 -297 -1641 -121
rect -17 -297 17 -121
rect 1641 -297 1675 -121
rect 3299 -297 3333 -121
rect 4957 -297 4991 -121
rect 6615 -297 6649 -121
rect 8273 -297 8307 -121
<< psubdiff >>
rect -8421 449 -8325 483
rect 8325 449 8421 483
rect -8421 387 -8387 449
rect 8387 387 8421 449
rect -8421 -449 -8387 -387
rect 8387 -449 8421 -387
rect -8421 -483 -8325 -449
rect 8325 -483 8421 -449
<< psubdiffcont >>
rect -8325 449 8325 483
rect -8421 -387 -8387 387
rect 8387 -387 8421 387
rect -8325 -483 8325 -449
<< poly >>
rect -8261 381 -6661 397
rect -8261 347 -8245 381
rect -6677 347 -6661 381
rect -8261 309 -6661 347
rect -6603 381 -5003 397
rect -6603 347 -6587 381
rect -5019 347 -5003 381
rect -6603 309 -5003 347
rect -4945 381 -3345 397
rect -4945 347 -4929 381
rect -3361 347 -3345 381
rect -4945 309 -3345 347
rect -3287 381 -1687 397
rect -3287 347 -3271 381
rect -1703 347 -1687 381
rect -3287 309 -1687 347
rect -1629 381 -29 397
rect -1629 347 -1613 381
rect -45 347 -29 381
rect -1629 309 -29 347
rect 29 381 1629 397
rect 29 347 45 381
rect 1613 347 1629 381
rect 29 309 1629 347
rect 1687 381 3287 397
rect 1687 347 1703 381
rect 3271 347 3287 381
rect 1687 309 3287 347
rect 3345 381 4945 397
rect 3345 347 3361 381
rect 4929 347 4945 381
rect 3345 309 4945 347
rect 5003 381 6603 397
rect 5003 347 5019 381
rect 6587 347 6603 381
rect 5003 309 6603 347
rect 6661 381 8261 397
rect 6661 347 6677 381
rect 8245 347 8261 381
rect 6661 309 8261 347
rect -8261 71 -6661 109
rect -8261 37 -8245 71
rect -6677 37 -6661 71
rect -8261 21 -6661 37
rect -6603 71 -5003 109
rect -6603 37 -6587 71
rect -5019 37 -5003 71
rect -6603 21 -5003 37
rect -4945 71 -3345 109
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -4945 21 -3345 37
rect -3287 71 -1687 109
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -3287 21 -1687 37
rect -1629 71 -29 109
rect -1629 37 -1613 71
rect -45 37 -29 71
rect -1629 21 -29 37
rect 29 71 1629 109
rect 29 37 45 71
rect 1613 37 1629 71
rect 29 21 1629 37
rect 1687 71 3287 109
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 1687 21 3287 37
rect 3345 71 4945 109
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 3345 21 4945 37
rect 5003 71 6603 109
rect 5003 37 5019 71
rect 6587 37 6603 71
rect 5003 21 6603 37
rect 6661 71 8261 109
rect 6661 37 6677 71
rect 8245 37 8261 71
rect 6661 21 8261 37
rect -8261 -37 -6661 -21
rect -8261 -71 -8245 -37
rect -6677 -71 -6661 -37
rect -8261 -109 -6661 -71
rect -6603 -37 -5003 -21
rect -6603 -71 -6587 -37
rect -5019 -71 -5003 -37
rect -6603 -109 -5003 -71
rect -4945 -37 -3345 -21
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -4945 -109 -3345 -71
rect -3287 -37 -1687 -21
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -3287 -109 -1687 -71
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -109 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -109 1629 -71
rect 1687 -37 3287 -21
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 1687 -109 3287 -71
rect 3345 -37 4945 -21
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 3345 -109 4945 -71
rect 5003 -37 6603 -21
rect 5003 -71 5019 -37
rect 6587 -71 6603 -37
rect 5003 -109 6603 -71
rect 6661 -37 8261 -21
rect 6661 -71 6677 -37
rect 8245 -71 8261 -37
rect 6661 -109 8261 -71
rect -8261 -347 -6661 -309
rect -8261 -381 -8245 -347
rect -6677 -381 -6661 -347
rect -8261 -397 -6661 -381
rect -6603 -347 -5003 -309
rect -6603 -381 -6587 -347
rect -5019 -381 -5003 -347
rect -6603 -397 -5003 -381
rect -4945 -347 -3345 -309
rect -4945 -381 -4929 -347
rect -3361 -381 -3345 -347
rect -4945 -397 -3345 -381
rect -3287 -347 -1687 -309
rect -3287 -381 -3271 -347
rect -1703 -381 -1687 -347
rect -3287 -397 -1687 -381
rect -1629 -347 -29 -309
rect -1629 -381 -1613 -347
rect -45 -381 -29 -347
rect -1629 -397 -29 -381
rect 29 -347 1629 -309
rect 29 -381 45 -347
rect 1613 -381 1629 -347
rect 29 -397 1629 -381
rect 1687 -347 3287 -309
rect 1687 -381 1703 -347
rect 3271 -381 3287 -347
rect 1687 -397 3287 -381
rect 3345 -347 4945 -309
rect 3345 -381 3361 -347
rect 4929 -381 4945 -347
rect 3345 -397 4945 -381
rect 5003 -347 6603 -309
rect 5003 -381 5019 -347
rect 6587 -381 6603 -347
rect 5003 -397 6603 -381
rect 6661 -347 8261 -309
rect 6661 -381 6677 -347
rect 8245 -381 8261 -347
rect 6661 -397 8261 -381
<< polycont >>
rect -8245 347 -6677 381
rect -6587 347 -5019 381
rect -4929 347 -3361 381
rect -3271 347 -1703 381
rect -1613 347 -45 381
rect 45 347 1613 381
rect 1703 347 3271 381
rect 3361 347 4929 381
rect 5019 347 6587 381
rect 6677 347 8245 381
rect -8245 37 -6677 71
rect -6587 37 -5019 71
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect 5019 37 6587 71
rect 6677 37 8245 71
rect -8245 -71 -6677 -37
rect -6587 -71 -5019 -37
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect 5019 -71 6587 -37
rect 6677 -71 8245 -37
rect -8245 -381 -6677 -347
rect -6587 -381 -5019 -347
rect -4929 -381 -3361 -347
rect -3271 -381 -1703 -347
rect -1613 -381 -45 -347
rect 45 -381 1613 -347
rect 1703 -381 3271 -347
rect 3361 -381 4929 -347
rect 5019 -381 6587 -347
rect 6677 -381 8245 -347
<< locali >>
rect -8421 449 -8325 483
rect 8325 449 8421 483
rect -8421 387 -8387 449
rect 8387 387 8421 449
rect -8261 347 -8245 381
rect -6677 347 -6661 381
rect -6603 347 -6587 381
rect -5019 347 -5003 381
rect -4945 347 -4929 381
rect -3361 347 -3345 381
rect -3287 347 -3271 381
rect -1703 347 -1687 381
rect -1629 347 -1613 381
rect -45 347 -29 381
rect 29 347 45 381
rect 1613 347 1629 381
rect 1687 347 1703 381
rect 3271 347 3287 381
rect 3345 347 3361 381
rect 4929 347 4945 381
rect 5003 347 5019 381
rect 6587 347 6603 381
rect 6661 347 6677 381
rect 8245 347 8261 381
rect -8307 297 -8273 313
rect -8307 105 -8273 121
rect -6649 297 -6615 313
rect -6649 105 -6615 121
rect -4991 297 -4957 313
rect -4991 105 -4957 121
rect -3333 297 -3299 313
rect -3333 105 -3299 121
rect -1675 297 -1641 313
rect -1675 105 -1641 121
rect -17 297 17 313
rect -17 105 17 121
rect 1641 297 1675 313
rect 1641 105 1675 121
rect 3299 297 3333 313
rect 3299 105 3333 121
rect 4957 297 4991 313
rect 4957 105 4991 121
rect 6615 297 6649 313
rect 6615 105 6649 121
rect 8273 297 8307 313
rect 8273 105 8307 121
rect -8261 37 -8245 71
rect -6677 37 -6661 71
rect -6603 37 -6587 71
rect -5019 37 -5003 71
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -1629 37 -1613 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1613 37 1629 71
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 5003 37 5019 71
rect 6587 37 6603 71
rect 6661 37 6677 71
rect 8245 37 8261 71
rect -8261 -71 -8245 -37
rect -6677 -71 -6661 -37
rect -6603 -71 -6587 -37
rect -5019 -71 -5003 -37
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 5003 -71 5019 -37
rect 6587 -71 6603 -37
rect 6661 -71 6677 -37
rect 8245 -71 8261 -37
rect -8307 -121 -8273 -105
rect -8307 -313 -8273 -297
rect -6649 -121 -6615 -105
rect -6649 -313 -6615 -297
rect -4991 -121 -4957 -105
rect -4991 -313 -4957 -297
rect -3333 -121 -3299 -105
rect -3333 -313 -3299 -297
rect -1675 -121 -1641 -105
rect -1675 -313 -1641 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 1641 -121 1675 -105
rect 1641 -313 1675 -297
rect 3299 -121 3333 -105
rect 3299 -313 3333 -297
rect 4957 -121 4991 -105
rect 4957 -313 4991 -297
rect 6615 -121 6649 -105
rect 6615 -313 6649 -297
rect 8273 -121 8307 -105
rect 8273 -313 8307 -297
rect -8261 -381 -8245 -347
rect -6677 -381 -6661 -347
rect -6603 -381 -6587 -347
rect -5019 -381 -5003 -347
rect -4945 -381 -4929 -347
rect -3361 -381 -3345 -347
rect -3287 -381 -3271 -347
rect -1703 -381 -1687 -347
rect -1629 -381 -1613 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 1613 -381 1629 -347
rect 1687 -381 1703 -347
rect 3271 -381 3287 -347
rect 3345 -381 3361 -347
rect 4929 -381 4945 -347
rect 5003 -381 5019 -347
rect 6587 -381 6603 -347
rect 6661 -381 6677 -347
rect 8245 -381 8261 -347
rect -8421 -449 -8387 -387
rect 8387 -449 8421 -387
rect -8421 -483 -8325 -449
rect 8325 -483 8421 -449
<< viali >>
rect -8245 347 -6677 381
rect -6587 347 -5019 381
rect -4929 347 -3361 381
rect -3271 347 -1703 381
rect -1613 347 -45 381
rect 45 347 1613 381
rect 1703 347 3271 381
rect 3361 347 4929 381
rect 5019 347 6587 381
rect 6677 347 8245 381
rect -8307 121 -8273 297
rect -6649 121 -6615 297
rect -4991 121 -4957 297
rect -3333 121 -3299 297
rect -1675 121 -1641 297
rect -17 121 17 297
rect 1641 121 1675 297
rect 3299 121 3333 297
rect 4957 121 4991 297
rect 6615 121 6649 297
rect 8273 121 8307 297
rect -8245 37 -6677 71
rect -6587 37 -5019 71
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect 5019 37 6587 71
rect 6677 37 8245 71
rect -8245 -71 -6677 -37
rect -6587 -71 -5019 -37
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect 5019 -71 6587 -37
rect 6677 -71 8245 -37
rect -8307 -297 -8273 -121
rect -6649 -297 -6615 -121
rect -4991 -297 -4957 -121
rect -3333 -297 -3299 -121
rect -1675 -297 -1641 -121
rect -17 -297 17 -121
rect 1641 -297 1675 -121
rect 3299 -297 3333 -121
rect 4957 -297 4991 -121
rect 6615 -297 6649 -121
rect 8273 -297 8307 -121
rect -8245 -381 -6677 -347
rect -6587 -381 -5019 -347
rect -4929 -381 -3361 -347
rect -3271 -381 -1703 -347
rect -1613 -381 -45 -347
rect 45 -381 1613 -347
rect 1703 -381 3271 -347
rect 3361 -381 4929 -347
rect 5019 -381 6587 -347
rect 6677 -381 8245 -347
<< metal1 >>
rect -8257 381 -6665 387
rect -8257 347 -8245 381
rect -6677 347 -6665 381
rect -8257 341 -6665 347
rect -6599 381 -5007 387
rect -6599 347 -6587 381
rect -5019 347 -5007 381
rect -6599 341 -5007 347
rect -4941 381 -3349 387
rect -4941 347 -4929 381
rect -3361 347 -3349 381
rect -4941 341 -3349 347
rect -3283 381 -1691 387
rect -3283 347 -3271 381
rect -1703 347 -1691 381
rect -3283 341 -1691 347
rect -1625 381 -33 387
rect -1625 347 -1613 381
rect -45 347 -33 381
rect -1625 341 -33 347
rect 33 381 1625 387
rect 33 347 45 381
rect 1613 347 1625 381
rect 33 341 1625 347
rect 1691 381 3283 387
rect 1691 347 1703 381
rect 3271 347 3283 381
rect 1691 341 3283 347
rect 3349 381 4941 387
rect 3349 347 3361 381
rect 4929 347 4941 381
rect 3349 341 4941 347
rect 5007 381 6599 387
rect 5007 347 5019 381
rect 6587 347 6599 381
rect 5007 341 6599 347
rect 6665 381 8257 387
rect 6665 347 6677 381
rect 8245 347 8257 381
rect 6665 341 8257 347
rect -8313 297 -8267 309
rect -8313 121 -8307 297
rect -8273 121 -8267 297
rect -8313 109 -8267 121
rect -6655 297 -6609 309
rect -6655 121 -6649 297
rect -6615 121 -6609 297
rect -6655 109 -6609 121
rect -4997 297 -4951 309
rect -4997 121 -4991 297
rect -4957 121 -4951 297
rect -4997 109 -4951 121
rect -3339 297 -3293 309
rect -3339 121 -3333 297
rect -3299 121 -3293 297
rect -3339 109 -3293 121
rect -1681 297 -1635 309
rect -1681 121 -1675 297
rect -1641 121 -1635 297
rect -1681 109 -1635 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 1635 297 1681 309
rect 1635 121 1641 297
rect 1675 121 1681 297
rect 1635 109 1681 121
rect 3293 297 3339 309
rect 3293 121 3299 297
rect 3333 121 3339 297
rect 3293 109 3339 121
rect 4951 297 4997 309
rect 4951 121 4957 297
rect 4991 121 4997 297
rect 4951 109 4997 121
rect 6609 297 6655 309
rect 6609 121 6615 297
rect 6649 121 6655 297
rect 6609 109 6655 121
rect 8267 297 8313 309
rect 8267 121 8273 297
rect 8307 121 8313 297
rect 8267 109 8313 121
rect -8257 71 -6665 77
rect -8257 37 -8245 71
rect -6677 37 -6665 71
rect -8257 31 -6665 37
rect -6599 71 -5007 77
rect -6599 37 -6587 71
rect -5019 37 -5007 71
rect -6599 31 -5007 37
rect -4941 71 -3349 77
rect -4941 37 -4929 71
rect -3361 37 -3349 71
rect -4941 31 -3349 37
rect -3283 71 -1691 77
rect -3283 37 -3271 71
rect -1703 37 -1691 71
rect -3283 31 -1691 37
rect -1625 71 -33 77
rect -1625 37 -1613 71
rect -45 37 -33 71
rect -1625 31 -33 37
rect 33 71 1625 77
rect 33 37 45 71
rect 1613 37 1625 71
rect 33 31 1625 37
rect 1691 71 3283 77
rect 1691 37 1703 71
rect 3271 37 3283 71
rect 1691 31 3283 37
rect 3349 71 4941 77
rect 3349 37 3361 71
rect 4929 37 4941 71
rect 3349 31 4941 37
rect 5007 71 6599 77
rect 5007 37 5019 71
rect 6587 37 6599 71
rect 5007 31 6599 37
rect 6665 71 8257 77
rect 6665 37 6677 71
rect 8245 37 8257 71
rect 6665 31 8257 37
rect -8257 -37 -6665 -31
rect -8257 -71 -8245 -37
rect -6677 -71 -6665 -37
rect -8257 -77 -6665 -71
rect -6599 -37 -5007 -31
rect -6599 -71 -6587 -37
rect -5019 -71 -5007 -37
rect -6599 -77 -5007 -71
rect -4941 -37 -3349 -31
rect -4941 -71 -4929 -37
rect -3361 -71 -3349 -37
rect -4941 -77 -3349 -71
rect -3283 -37 -1691 -31
rect -3283 -71 -3271 -37
rect -1703 -71 -1691 -37
rect -3283 -77 -1691 -71
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect 1691 -37 3283 -31
rect 1691 -71 1703 -37
rect 3271 -71 3283 -37
rect 1691 -77 3283 -71
rect 3349 -37 4941 -31
rect 3349 -71 3361 -37
rect 4929 -71 4941 -37
rect 3349 -77 4941 -71
rect 5007 -37 6599 -31
rect 5007 -71 5019 -37
rect 6587 -71 6599 -37
rect 5007 -77 6599 -71
rect 6665 -37 8257 -31
rect 6665 -71 6677 -37
rect 8245 -71 8257 -37
rect 6665 -77 8257 -71
rect -8313 -121 -8267 -109
rect -8313 -297 -8307 -121
rect -8273 -297 -8267 -121
rect -8313 -309 -8267 -297
rect -6655 -121 -6609 -109
rect -6655 -297 -6649 -121
rect -6615 -297 -6609 -121
rect -6655 -309 -6609 -297
rect -4997 -121 -4951 -109
rect -4997 -297 -4991 -121
rect -4957 -297 -4951 -121
rect -4997 -309 -4951 -297
rect -3339 -121 -3293 -109
rect -3339 -297 -3333 -121
rect -3299 -297 -3293 -121
rect -3339 -309 -3293 -297
rect -1681 -121 -1635 -109
rect -1681 -297 -1675 -121
rect -1641 -297 -1635 -121
rect -1681 -309 -1635 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 1635 -121 1681 -109
rect 1635 -297 1641 -121
rect 1675 -297 1681 -121
rect 1635 -309 1681 -297
rect 3293 -121 3339 -109
rect 3293 -297 3299 -121
rect 3333 -297 3339 -121
rect 3293 -309 3339 -297
rect 4951 -121 4997 -109
rect 4951 -297 4957 -121
rect 4991 -297 4997 -121
rect 4951 -309 4997 -297
rect 6609 -121 6655 -109
rect 6609 -297 6615 -121
rect 6649 -297 6655 -121
rect 6609 -309 6655 -297
rect 8267 -121 8313 -109
rect 8267 -297 8273 -121
rect 8307 -297 8313 -121
rect 8267 -309 8313 -297
rect -8257 -347 -6665 -341
rect -8257 -381 -8245 -347
rect -6677 -381 -6665 -347
rect -8257 -387 -6665 -381
rect -6599 -347 -5007 -341
rect -6599 -381 -6587 -347
rect -5019 -381 -5007 -347
rect -6599 -387 -5007 -381
rect -4941 -347 -3349 -341
rect -4941 -381 -4929 -347
rect -3361 -381 -3349 -347
rect -4941 -387 -3349 -381
rect -3283 -347 -1691 -341
rect -3283 -381 -3271 -347
rect -1703 -381 -1691 -347
rect -3283 -387 -1691 -381
rect -1625 -347 -33 -341
rect -1625 -381 -1613 -347
rect -45 -381 -33 -347
rect -1625 -387 -33 -381
rect 33 -347 1625 -341
rect 33 -381 45 -347
rect 1613 -381 1625 -347
rect 33 -387 1625 -381
rect 1691 -347 3283 -341
rect 1691 -381 1703 -347
rect 3271 -381 3283 -347
rect 1691 -387 3283 -381
rect 3349 -347 4941 -341
rect 3349 -381 3361 -347
rect 4929 -381 4941 -347
rect 3349 -387 4941 -381
rect 5007 -347 6599 -341
rect 5007 -381 5019 -347
rect 6587 -381 6599 -347
rect 5007 -387 6599 -381
rect 6665 -347 8257 -341
rect 6665 -381 6677 -347
rect 8245 -381 8257 -347
rect 6665 -387 8257 -381
<< properties >>
string FIXED_BBOX -8404 -466 8404 466
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 8 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
