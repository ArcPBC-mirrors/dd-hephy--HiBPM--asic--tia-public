magic
tech sky130A
magscale 1 2
timestamp 1685110944
<< metal3 >>
rect -11410 8492 -7038 8520
rect -11410 4468 -7122 8492
rect -7058 4468 -7038 8492
rect -11410 4440 -7038 4468
rect -6798 8492 -2426 8520
rect -6798 4468 -2510 8492
rect -2446 4468 -2426 8492
rect -6798 4440 -2426 4468
rect -2186 8492 2186 8520
rect -2186 4468 2102 8492
rect 2166 4468 2186 8492
rect -2186 4440 2186 4468
rect 2426 8492 6798 8520
rect 2426 4468 6714 8492
rect 6778 4468 6798 8492
rect 2426 4440 6798 4468
rect 7038 8492 11410 8520
rect 7038 4468 11326 8492
rect 11390 4468 11410 8492
rect 7038 4440 11410 4468
rect -11410 4172 -7038 4200
rect -11410 148 -7122 4172
rect -7058 148 -7038 4172
rect -11410 120 -7038 148
rect -6798 4172 -2426 4200
rect -6798 148 -2510 4172
rect -2446 148 -2426 4172
rect -6798 120 -2426 148
rect -2186 4172 2186 4200
rect -2186 148 2102 4172
rect 2166 148 2186 4172
rect -2186 120 2186 148
rect 2426 4172 6798 4200
rect 2426 148 6714 4172
rect 6778 148 6798 4172
rect 2426 120 6798 148
rect 7038 4172 11410 4200
rect 7038 148 11326 4172
rect 11390 148 11410 4172
rect 7038 120 11410 148
rect -11410 -148 -7038 -120
rect -11410 -4172 -7122 -148
rect -7058 -4172 -7038 -148
rect -11410 -4200 -7038 -4172
rect -6798 -148 -2426 -120
rect -6798 -4172 -2510 -148
rect -2446 -4172 -2426 -148
rect -6798 -4200 -2426 -4172
rect -2186 -148 2186 -120
rect -2186 -4172 2102 -148
rect 2166 -4172 2186 -148
rect -2186 -4200 2186 -4172
rect 2426 -148 6798 -120
rect 2426 -4172 6714 -148
rect 6778 -4172 6798 -148
rect 2426 -4200 6798 -4172
rect 7038 -148 11410 -120
rect 7038 -4172 11326 -148
rect 11390 -4172 11410 -148
rect 7038 -4200 11410 -4172
rect -11410 -4468 -7038 -4440
rect -11410 -8492 -7122 -4468
rect -7058 -8492 -7038 -4468
rect -11410 -8520 -7038 -8492
rect -6798 -4468 -2426 -4440
rect -6798 -8492 -2510 -4468
rect -2446 -8492 -2426 -4468
rect -6798 -8520 -2426 -8492
rect -2186 -4468 2186 -4440
rect -2186 -8492 2102 -4468
rect 2166 -8492 2186 -4468
rect -2186 -8520 2186 -8492
rect 2426 -4468 6798 -4440
rect 2426 -8492 6714 -4468
rect 6778 -8492 6798 -4468
rect 2426 -8520 6798 -8492
rect 7038 -4468 11410 -4440
rect 7038 -8492 11326 -4468
rect 11390 -8492 11410 -4468
rect 7038 -8520 11410 -8492
<< via3 >>
rect -7122 4468 -7058 8492
rect -2510 4468 -2446 8492
rect 2102 4468 2166 8492
rect 6714 4468 6778 8492
rect 11326 4468 11390 8492
rect -7122 148 -7058 4172
rect -2510 148 -2446 4172
rect 2102 148 2166 4172
rect 6714 148 6778 4172
rect 11326 148 11390 4172
rect -7122 -4172 -7058 -148
rect -2510 -4172 -2446 -148
rect 2102 -4172 2166 -148
rect 6714 -4172 6778 -148
rect 11326 -4172 11390 -148
rect -7122 -8492 -7058 -4468
rect -2510 -8492 -2446 -4468
rect 2102 -8492 2166 -4468
rect 6714 -8492 6778 -4468
rect 11326 -8492 11390 -4468
<< mimcap >>
rect -11370 8440 -7370 8480
rect -11370 4520 -11330 8440
rect -7410 4520 -7370 8440
rect -11370 4480 -7370 4520
rect -6758 8440 -2758 8480
rect -6758 4520 -6718 8440
rect -2798 4520 -2758 8440
rect -6758 4480 -2758 4520
rect -2146 8440 1854 8480
rect -2146 4520 -2106 8440
rect 1814 4520 1854 8440
rect -2146 4480 1854 4520
rect 2466 8440 6466 8480
rect 2466 4520 2506 8440
rect 6426 4520 6466 8440
rect 2466 4480 6466 4520
rect 7078 8440 11078 8480
rect 7078 4520 7118 8440
rect 11038 4520 11078 8440
rect 7078 4480 11078 4520
rect -11370 4120 -7370 4160
rect -11370 200 -11330 4120
rect -7410 200 -7370 4120
rect -11370 160 -7370 200
rect -6758 4120 -2758 4160
rect -6758 200 -6718 4120
rect -2798 200 -2758 4120
rect -6758 160 -2758 200
rect -2146 4120 1854 4160
rect -2146 200 -2106 4120
rect 1814 200 1854 4120
rect -2146 160 1854 200
rect 2466 4120 6466 4160
rect 2466 200 2506 4120
rect 6426 200 6466 4120
rect 2466 160 6466 200
rect 7078 4120 11078 4160
rect 7078 200 7118 4120
rect 11038 200 11078 4120
rect 7078 160 11078 200
rect -11370 -200 -7370 -160
rect -11370 -4120 -11330 -200
rect -7410 -4120 -7370 -200
rect -11370 -4160 -7370 -4120
rect -6758 -200 -2758 -160
rect -6758 -4120 -6718 -200
rect -2798 -4120 -2758 -200
rect -6758 -4160 -2758 -4120
rect -2146 -200 1854 -160
rect -2146 -4120 -2106 -200
rect 1814 -4120 1854 -200
rect -2146 -4160 1854 -4120
rect 2466 -200 6466 -160
rect 2466 -4120 2506 -200
rect 6426 -4120 6466 -200
rect 2466 -4160 6466 -4120
rect 7078 -200 11078 -160
rect 7078 -4120 7118 -200
rect 11038 -4120 11078 -200
rect 7078 -4160 11078 -4120
rect -11370 -4520 -7370 -4480
rect -11370 -8440 -11330 -4520
rect -7410 -8440 -7370 -4520
rect -11370 -8480 -7370 -8440
rect -6758 -4520 -2758 -4480
rect -6758 -8440 -6718 -4520
rect -2798 -8440 -2758 -4520
rect -6758 -8480 -2758 -8440
rect -2146 -4520 1854 -4480
rect -2146 -8440 -2106 -4520
rect 1814 -8440 1854 -4520
rect -2146 -8480 1854 -8440
rect 2466 -4520 6466 -4480
rect 2466 -8440 2506 -4520
rect 6426 -8440 6466 -4520
rect 2466 -8480 6466 -8440
rect 7078 -4520 11078 -4480
rect 7078 -8440 7118 -4520
rect 11038 -8440 11078 -4520
rect 7078 -8480 11078 -8440
<< mimcapcontact >>
rect -11330 4520 -7410 8440
rect -6718 4520 -2798 8440
rect -2106 4520 1814 8440
rect 2506 4520 6426 8440
rect 7118 4520 11038 8440
rect -11330 200 -7410 4120
rect -6718 200 -2798 4120
rect -2106 200 1814 4120
rect 2506 200 6426 4120
rect 7118 200 11038 4120
rect -11330 -4120 -7410 -200
rect -6718 -4120 -2798 -200
rect -2106 -4120 1814 -200
rect 2506 -4120 6426 -200
rect 7118 -4120 11038 -200
rect -11330 -8440 -7410 -4520
rect -6718 -8440 -2798 -4520
rect -2106 -8440 1814 -4520
rect 2506 -8440 6426 -4520
rect 7118 -8440 11038 -4520
<< metal4 >>
rect -9422 8441 -9318 8640
rect -7142 8492 -7038 8640
rect -11331 8440 -7409 8441
rect -11331 4520 -11330 8440
rect -7410 4520 -7409 8440
rect -11331 4519 -7409 4520
rect -9422 4121 -9318 4519
rect -7142 4468 -7122 8492
rect -7058 4468 -7038 8492
rect -4810 8441 -4706 8640
rect -2530 8492 -2426 8640
rect -6719 8440 -2797 8441
rect -6719 4520 -6718 8440
rect -2798 4520 -2797 8440
rect -6719 4519 -2797 4520
rect -7142 4172 -7038 4468
rect -11331 4120 -7409 4121
rect -11331 200 -11330 4120
rect -7410 200 -7409 4120
rect -11331 199 -7409 200
rect -9422 -199 -9318 199
rect -7142 148 -7122 4172
rect -7058 148 -7038 4172
rect -4810 4121 -4706 4519
rect -2530 4468 -2510 8492
rect -2446 4468 -2426 8492
rect -198 8441 -94 8640
rect 2082 8492 2186 8640
rect -2107 8440 1815 8441
rect -2107 4520 -2106 8440
rect 1814 4520 1815 8440
rect -2107 4519 1815 4520
rect -2530 4172 -2426 4468
rect -6719 4120 -2797 4121
rect -6719 200 -6718 4120
rect -2798 200 -2797 4120
rect -6719 199 -2797 200
rect -7142 -148 -7038 148
rect -11331 -200 -7409 -199
rect -11331 -4120 -11330 -200
rect -7410 -4120 -7409 -200
rect -11331 -4121 -7409 -4120
rect -9422 -4519 -9318 -4121
rect -7142 -4172 -7122 -148
rect -7058 -4172 -7038 -148
rect -4810 -199 -4706 199
rect -2530 148 -2510 4172
rect -2446 148 -2426 4172
rect -198 4121 -94 4519
rect 2082 4468 2102 8492
rect 2166 4468 2186 8492
rect 4414 8441 4518 8640
rect 6694 8492 6798 8640
rect 2505 8440 6427 8441
rect 2505 4520 2506 8440
rect 6426 4520 6427 8440
rect 2505 4519 6427 4520
rect 2082 4172 2186 4468
rect -2107 4120 1815 4121
rect -2107 200 -2106 4120
rect 1814 200 1815 4120
rect -2107 199 1815 200
rect -2530 -148 -2426 148
rect -6719 -200 -2797 -199
rect -6719 -4120 -6718 -200
rect -2798 -4120 -2797 -200
rect -6719 -4121 -2797 -4120
rect -7142 -4468 -7038 -4172
rect -11331 -4520 -7409 -4519
rect -11331 -8440 -11330 -4520
rect -7410 -8440 -7409 -4520
rect -11331 -8441 -7409 -8440
rect -9422 -8640 -9318 -8441
rect -7142 -8492 -7122 -4468
rect -7058 -8492 -7038 -4468
rect -4810 -4519 -4706 -4121
rect -2530 -4172 -2510 -148
rect -2446 -4172 -2426 -148
rect -198 -199 -94 199
rect 2082 148 2102 4172
rect 2166 148 2186 4172
rect 4414 4121 4518 4519
rect 6694 4468 6714 8492
rect 6778 4468 6798 8492
rect 9026 8441 9130 8640
rect 11306 8492 11410 8640
rect 7117 8440 11039 8441
rect 7117 4520 7118 8440
rect 11038 4520 11039 8440
rect 7117 4519 11039 4520
rect 6694 4172 6798 4468
rect 2505 4120 6427 4121
rect 2505 200 2506 4120
rect 6426 200 6427 4120
rect 2505 199 6427 200
rect 2082 -148 2186 148
rect -2107 -200 1815 -199
rect -2107 -4120 -2106 -200
rect 1814 -4120 1815 -200
rect -2107 -4121 1815 -4120
rect -2530 -4468 -2426 -4172
rect -6719 -4520 -2797 -4519
rect -6719 -8440 -6718 -4520
rect -2798 -8440 -2797 -4520
rect -6719 -8441 -2797 -8440
rect -7142 -8640 -7038 -8492
rect -4810 -8640 -4706 -8441
rect -2530 -8492 -2510 -4468
rect -2446 -8492 -2426 -4468
rect -198 -4519 -94 -4121
rect 2082 -4172 2102 -148
rect 2166 -4172 2186 -148
rect 4414 -199 4518 199
rect 6694 148 6714 4172
rect 6778 148 6798 4172
rect 9026 4121 9130 4519
rect 11306 4468 11326 8492
rect 11390 4468 11410 8492
rect 11306 4172 11410 4468
rect 7117 4120 11039 4121
rect 7117 200 7118 4120
rect 11038 200 11039 4120
rect 7117 199 11039 200
rect 6694 -148 6798 148
rect 2505 -200 6427 -199
rect 2505 -4120 2506 -200
rect 6426 -4120 6427 -200
rect 2505 -4121 6427 -4120
rect 2082 -4468 2186 -4172
rect -2107 -4520 1815 -4519
rect -2107 -8440 -2106 -4520
rect 1814 -8440 1815 -4520
rect -2107 -8441 1815 -8440
rect -2530 -8640 -2426 -8492
rect -198 -8640 -94 -8441
rect 2082 -8492 2102 -4468
rect 2166 -8492 2186 -4468
rect 4414 -4519 4518 -4121
rect 6694 -4172 6714 -148
rect 6778 -4172 6798 -148
rect 9026 -199 9130 199
rect 11306 148 11326 4172
rect 11390 148 11410 4172
rect 11306 -148 11410 148
rect 7117 -200 11039 -199
rect 7117 -4120 7118 -200
rect 11038 -4120 11039 -200
rect 7117 -4121 11039 -4120
rect 6694 -4468 6798 -4172
rect 2505 -4520 6427 -4519
rect 2505 -8440 2506 -4520
rect 6426 -8440 6427 -4520
rect 2505 -8441 6427 -8440
rect 2082 -8640 2186 -8492
rect 4414 -8640 4518 -8441
rect 6694 -8492 6714 -4468
rect 6778 -8492 6798 -4468
rect 9026 -4519 9130 -4121
rect 11306 -4172 11326 -148
rect 11390 -4172 11410 -148
rect 11306 -4468 11410 -4172
rect 7117 -4520 11039 -4519
rect 7117 -8440 7118 -4520
rect 11038 -8440 11039 -4520
rect 7117 -8441 11039 -8440
rect 6694 -8640 6798 -8492
rect 9026 -8640 9130 -8441
rect 11306 -8492 11326 -4468
rect 11390 -8492 11410 -4468
rect 11306 -8640 11410 -8492
<< properties >>
string FIXED_BBOX 7038 4440 11118 8520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 5 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
