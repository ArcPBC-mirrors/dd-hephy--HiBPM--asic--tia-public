magic
tech sky130A
magscale 1 2
timestamp 1687117224
<< error_p >>
rect -1325 272 -1267 278
rect -1133 272 -1075 278
rect -941 272 -883 278
rect -749 272 -691 278
rect -557 272 -499 278
rect -365 272 -307 278
rect -173 272 -115 278
rect 19 272 77 278
rect 211 272 269 278
rect 403 272 461 278
rect 595 272 653 278
rect 787 272 845 278
rect 979 272 1037 278
rect 1171 272 1229 278
rect 1363 272 1421 278
rect -1325 238 -1313 272
rect -1133 238 -1121 272
rect -941 238 -929 272
rect -749 238 -737 272
rect -557 238 -545 272
rect -365 238 -353 272
rect -173 238 -161 272
rect 19 238 31 272
rect 211 238 223 272
rect 403 238 415 272
rect 595 238 607 272
rect 787 238 799 272
rect 979 238 991 272
rect 1171 238 1183 272
rect 1363 238 1375 272
rect -1325 232 -1267 238
rect -1133 232 -1075 238
rect -941 232 -883 238
rect -749 232 -691 238
rect -557 232 -499 238
rect -365 232 -307 238
rect -173 232 -115 238
rect 19 232 77 238
rect 211 232 269 238
rect 403 232 461 238
rect 595 232 653 238
rect 787 232 845 238
rect 979 232 1037 238
rect 1171 232 1229 238
rect 1363 232 1421 238
rect -1421 -238 -1363 -232
rect -1229 -238 -1171 -232
rect -1037 -238 -979 -232
rect -845 -238 -787 -232
rect -653 -238 -595 -232
rect -461 -238 -403 -232
rect -269 -238 -211 -232
rect -77 -238 -19 -232
rect 115 -238 173 -232
rect 307 -238 365 -232
rect 499 -238 557 -232
rect 691 -238 749 -232
rect 883 -238 941 -232
rect 1075 -238 1133 -232
rect 1267 -238 1325 -232
rect -1421 -272 -1409 -238
rect -1229 -272 -1217 -238
rect -1037 -272 -1025 -238
rect -845 -272 -833 -238
rect -653 -272 -641 -238
rect -461 -272 -449 -238
rect -269 -272 -257 -238
rect -77 -272 -65 -238
rect 115 -272 127 -238
rect 307 -272 319 -238
rect 499 -272 511 -238
rect 691 -272 703 -238
rect 883 -272 895 -238
rect 1075 -272 1087 -238
rect 1267 -272 1279 -238
rect -1421 -278 -1363 -272
rect -1229 -278 -1171 -272
rect -1037 -278 -979 -272
rect -845 -278 -787 -272
rect -653 -278 -595 -272
rect -461 -278 -403 -272
rect -269 -278 -211 -272
rect -77 -278 -19 -272
rect 115 -278 173 -272
rect 307 -278 365 -272
rect 499 -278 557 -272
rect 691 -278 749 -272
rect 883 -278 941 -272
rect 1075 -278 1133 -272
rect 1267 -278 1325 -272
<< pwell >>
rect -1607 -410 1607 410
<< nmoslvt >>
rect -1407 -200 -1377 200
rect -1311 -200 -1281 200
rect -1215 -200 -1185 200
rect -1119 -200 -1089 200
rect -1023 -200 -993 200
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
rect 993 -200 1023 200
rect 1089 -200 1119 200
rect 1185 -200 1215 200
rect 1281 -200 1311 200
rect 1377 -200 1407 200
<< ndiff >>
rect -1469 188 -1407 200
rect -1469 -188 -1457 188
rect -1423 -188 -1407 188
rect -1469 -200 -1407 -188
rect -1377 188 -1311 200
rect -1377 -188 -1361 188
rect -1327 -188 -1311 188
rect -1377 -200 -1311 -188
rect -1281 188 -1215 200
rect -1281 -188 -1265 188
rect -1231 -188 -1215 188
rect -1281 -200 -1215 -188
rect -1185 188 -1119 200
rect -1185 -188 -1169 188
rect -1135 -188 -1119 188
rect -1185 -200 -1119 -188
rect -1089 188 -1023 200
rect -1089 -188 -1073 188
rect -1039 -188 -1023 188
rect -1089 -200 -1023 -188
rect -993 188 -927 200
rect -993 -188 -977 188
rect -943 -188 -927 188
rect -993 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 993 200
rect 927 -188 943 188
rect 977 -188 993 188
rect 927 -200 993 -188
rect 1023 188 1089 200
rect 1023 -188 1039 188
rect 1073 -188 1089 188
rect 1023 -200 1089 -188
rect 1119 188 1185 200
rect 1119 -188 1135 188
rect 1169 -188 1185 188
rect 1119 -200 1185 -188
rect 1215 188 1281 200
rect 1215 -188 1231 188
rect 1265 -188 1281 188
rect 1215 -200 1281 -188
rect 1311 188 1377 200
rect 1311 -188 1327 188
rect 1361 -188 1377 188
rect 1311 -200 1377 -188
rect 1407 188 1469 200
rect 1407 -188 1423 188
rect 1457 -188 1469 188
rect 1407 -200 1469 -188
<< ndiffc >>
rect -1457 -188 -1423 188
rect -1361 -188 -1327 188
rect -1265 -188 -1231 188
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect 1231 -188 1265 188
rect 1327 -188 1361 188
rect 1423 -188 1457 188
<< psubdiff >>
rect -1571 340 -1475 374
rect 1475 340 1571 374
rect -1571 278 -1537 340
rect 1537 278 1571 340
rect -1571 -340 -1537 -278
rect 1537 -340 1571 -278
rect -1571 -374 -1475 -340
rect 1475 -374 1571 -340
<< psubdiffcont >>
rect -1475 340 1475 374
rect -1571 -278 -1537 278
rect 1537 -278 1571 278
rect -1475 -374 1475 -340
<< poly >>
rect -1329 272 -1263 288
rect -1329 238 -1313 272
rect -1279 238 -1263 272
rect -1407 200 -1377 226
rect -1329 222 -1263 238
rect -1137 272 -1071 288
rect -1137 238 -1121 272
rect -1087 238 -1071 272
rect -1311 200 -1281 222
rect -1215 200 -1185 226
rect -1137 222 -1071 238
rect -945 272 -879 288
rect -945 238 -929 272
rect -895 238 -879 272
rect -1119 200 -1089 222
rect -1023 200 -993 226
rect -945 222 -879 238
rect -753 272 -687 288
rect -753 238 -737 272
rect -703 238 -687 272
rect -927 200 -897 222
rect -831 200 -801 226
rect -753 222 -687 238
rect -561 272 -495 288
rect -561 238 -545 272
rect -511 238 -495 272
rect -735 200 -705 222
rect -639 200 -609 226
rect -561 222 -495 238
rect -369 272 -303 288
rect -369 238 -353 272
rect -319 238 -303 272
rect -543 200 -513 222
rect -447 200 -417 226
rect -369 222 -303 238
rect -177 272 -111 288
rect -177 238 -161 272
rect -127 238 -111 272
rect -351 200 -321 222
rect -255 200 -225 226
rect -177 222 -111 238
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -159 200 -129 222
rect -63 200 -33 226
rect 15 222 81 238
rect 207 272 273 288
rect 207 238 223 272
rect 257 238 273 272
rect 33 200 63 222
rect 129 200 159 226
rect 207 222 273 238
rect 399 272 465 288
rect 399 238 415 272
rect 449 238 465 272
rect 225 200 255 222
rect 321 200 351 226
rect 399 222 465 238
rect 591 272 657 288
rect 591 238 607 272
rect 641 238 657 272
rect 417 200 447 222
rect 513 200 543 226
rect 591 222 657 238
rect 783 272 849 288
rect 783 238 799 272
rect 833 238 849 272
rect 609 200 639 222
rect 705 200 735 226
rect 783 222 849 238
rect 975 272 1041 288
rect 975 238 991 272
rect 1025 238 1041 272
rect 801 200 831 222
rect 897 200 927 226
rect 975 222 1041 238
rect 1167 272 1233 288
rect 1167 238 1183 272
rect 1217 238 1233 272
rect 993 200 1023 222
rect 1089 200 1119 226
rect 1167 222 1233 238
rect 1359 272 1425 288
rect 1359 238 1375 272
rect 1409 238 1425 272
rect 1185 200 1215 222
rect 1281 200 1311 226
rect 1359 222 1425 238
rect 1377 200 1407 222
rect -1407 -222 -1377 -200
rect -1425 -238 -1359 -222
rect -1311 -226 -1281 -200
rect -1215 -222 -1185 -200
rect -1425 -272 -1409 -238
rect -1375 -272 -1359 -238
rect -1425 -288 -1359 -272
rect -1233 -238 -1167 -222
rect -1119 -226 -1089 -200
rect -1023 -222 -993 -200
rect -1233 -272 -1217 -238
rect -1183 -272 -1167 -238
rect -1233 -288 -1167 -272
rect -1041 -238 -975 -222
rect -927 -226 -897 -200
rect -831 -222 -801 -200
rect -1041 -272 -1025 -238
rect -991 -272 -975 -238
rect -1041 -288 -975 -272
rect -849 -238 -783 -222
rect -735 -226 -705 -200
rect -639 -222 -609 -200
rect -849 -272 -833 -238
rect -799 -272 -783 -238
rect -849 -288 -783 -272
rect -657 -238 -591 -222
rect -543 -226 -513 -200
rect -447 -222 -417 -200
rect -657 -272 -641 -238
rect -607 -272 -591 -238
rect -657 -288 -591 -272
rect -465 -238 -399 -222
rect -351 -226 -321 -200
rect -255 -222 -225 -200
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -465 -288 -399 -272
rect -273 -238 -207 -222
rect -159 -226 -129 -200
rect -63 -222 -33 -200
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -273 -288 -207 -272
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect 129 -222 159 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
rect 111 -238 177 -222
rect 225 -226 255 -200
rect 321 -222 351 -200
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 111 -288 177 -272
rect 303 -238 369 -222
rect 417 -226 447 -200
rect 513 -222 543 -200
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 303 -288 369 -272
rect 495 -238 561 -222
rect 609 -226 639 -200
rect 705 -222 735 -200
rect 495 -272 511 -238
rect 545 -272 561 -238
rect 495 -288 561 -272
rect 687 -238 753 -222
rect 801 -226 831 -200
rect 897 -222 927 -200
rect 687 -272 703 -238
rect 737 -272 753 -238
rect 687 -288 753 -272
rect 879 -238 945 -222
rect 993 -226 1023 -200
rect 1089 -222 1119 -200
rect 879 -272 895 -238
rect 929 -272 945 -238
rect 879 -288 945 -272
rect 1071 -238 1137 -222
rect 1185 -226 1215 -200
rect 1281 -222 1311 -200
rect 1071 -272 1087 -238
rect 1121 -272 1137 -238
rect 1071 -288 1137 -272
rect 1263 -238 1329 -222
rect 1377 -226 1407 -200
rect 1263 -272 1279 -238
rect 1313 -272 1329 -238
rect 1263 -288 1329 -272
<< polycont >>
rect -1313 238 -1279 272
rect -1121 238 -1087 272
rect -929 238 -895 272
rect -737 238 -703 272
rect -545 238 -511 272
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect 607 238 641 272
rect 799 238 833 272
rect 991 238 1025 272
rect 1183 238 1217 272
rect 1375 238 1409 272
rect -1409 -272 -1375 -238
rect -1217 -272 -1183 -238
rect -1025 -272 -991 -238
rect -833 -272 -799 -238
rect -641 -272 -607 -238
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect 511 -272 545 -238
rect 703 -272 737 -238
rect 895 -272 929 -238
rect 1087 -272 1121 -238
rect 1279 -272 1313 -238
<< locali >>
rect -1571 340 -1475 374
rect 1475 340 1571 374
rect -1571 278 -1537 340
rect 1537 278 1571 340
rect -1329 238 -1313 272
rect -1279 238 -1263 272
rect -1137 238 -1121 272
rect -1087 238 -1071 272
rect -945 238 -929 272
rect -895 238 -879 272
rect -753 238 -737 272
rect -703 238 -687 272
rect -561 238 -545 272
rect -511 238 -495 272
rect -369 238 -353 272
rect -319 238 -303 272
rect -177 238 -161 272
rect -127 238 -111 272
rect 15 238 31 272
rect 65 238 81 272
rect 207 238 223 272
rect 257 238 273 272
rect 399 238 415 272
rect 449 238 465 272
rect 591 238 607 272
rect 641 238 657 272
rect 783 238 799 272
rect 833 238 849 272
rect 975 238 991 272
rect 1025 238 1041 272
rect 1167 238 1183 272
rect 1217 238 1233 272
rect 1359 238 1375 272
rect 1409 238 1425 272
rect -1457 188 -1423 204
rect -1457 -204 -1423 -188
rect -1361 188 -1327 204
rect -1361 -204 -1327 -188
rect -1265 188 -1231 204
rect -1265 -204 -1231 -188
rect -1169 188 -1135 204
rect -1169 -204 -1135 -188
rect -1073 188 -1039 204
rect -1073 -204 -1039 -188
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect 1039 188 1073 204
rect 1039 -204 1073 -188
rect 1135 188 1169 204
rect 1135 -204 1169 -188
rect 1231 188 1265 204
rect 1231 -204 1265 -188
rect 1327 188 1361 204
rect 1327 -204 1361 -188
rect 1423 188 1457 204
rect 1423 -204 1457 -188
rect -1425 -272 -1409 -238
rect -1375 -272 -1359 -238
rect -1233 -272 -1217 -238
rect -1183 -272 -1167 -238
rect -1041 -272 -1025 -238
rect -991 -272 -975 -238
rect -849 -272 -833 -238
rect -799 -272 -783 -238
rect -657 -272 -641 -238
rect -607 -272 -591 -238
rect -465 -272 -449 -238
rect -415 -272 -399 -238
rect -273 -272 -257 -238
rect -223 -272 -207 -238
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect 111 -272 127 -238
rect 161 -272 177 -238
rect 303 -272 319 -238
rect 353 -272 369 -238
rect 495 -272 511 -238
rect 545 -272 561 -238
rect 687 -272 703 -238
rect 737 -272 753 -238
rect 879 -272 895 -238
rect 929 -272 945 -238
rect 1071 -272 1087 -238
rect 1121 -272 1137 -238
rect 1263 -272 1279 -238
rect 1313 -272 1329 -238
rect -1571 -340 -1537 -278
rect 1537 -340 1571 -278
rect -1571 -374 -1475 -340
rect 1475 -374 1571 -340
<< viali >>
rect -1313 238 -1279 272
rect -1121 238 -1087 272
rect -929 238 -895 272
rect -737 238 -703 272
rect -545 238 -511 272
rect -353 238 -319 272
rect -161 238 -127 272
rect 31 238 65 272
rect 223 238 257 272
rect 415 238 449 272
rect 607 238 641 272
rect 799 238 833 272
rect 991 238 1025 272
rect 1183 238 1217 272
rect 1375 238 1409 272
rect -1457 -188 -1423 188
rect -1361 -188 -1327 188
rect -1265 -188 -1231 188
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect 1231 -188 1265 188
rect 1327 -188 1361 188
rect 1423 -188 1457 188
rect -1409 -272 -1375 -238
rect -1217 -272 -1183 -238
rect -1025 -272 -991 -238
rect -833 -272 -799 -238
rect -641 -272 -607 -238
rect -449 -272 -415 -238
rect -257 -272 -223 -238
rect -65 -272 -31 -238
rect 127 -272 161 -238
rect 319 -272 353 -238
rect 511 -272 545 -238
rect 703 -272 737 -238
rect 895 -272 929 -238
rect 1087 -272 1121 -238
rect 1279 -272 1313 -238
<< metal1 >>
rect -1325 272 -1267 278
rect -1325 238 -1313 272
rect -1279 238 -1267 272
rect -1325 232 -1267 238
rect -1133 272 -1075 278
rect -1133 238 -1121 272
rect -1087 238 -1075 272
rect -1133 232 -1075 238
rect -941 272 -883 278
rect -941 238 -929 272
rect -895 238 -883 272
rect -941 232 -883 238
rect -749 272 -691 278
rect -749 238 -737 272
rect -703 238 -691 272
rect -749 232 -691 238
rect -557 272 -499 278
rect -557 238 -545 272
rect -511 238 -499 272
rect -557 232 -499 238
rect -365 272 -307 278
rect -365 238 -353 272
rect -319 238 -307 272
rect -365 232 -307 238
rect -173 272 -115 278
rect -173 238 -161 272
rect -127 238 -115 272
rect -173 232 -115 238
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect 211 272 269 278
rect 211 238 223 272
rect 257 238 269 272
rect 211 232 269 238
rect 403 272 461 278
rect 403 238 415 272
rect 449 238 461 272
rect 403 232 461 238
rect 595 272 653 278
rect 595 238 607 272
rect 641 238 653 272
rect 595 232 653 238
rect 787 272 845 278
rect 787 238 799 272
rect 833 238 845 272
rect 787 232 845 238
rect 979 272 1037 278
rect 979 238 991 272
rect 1025 238 1037 272
rect 979 232 1037 238
rect 1171 272 1229 278
rect 1171 238 1183 272
rect 1217 238 1229 272
rect 1171 232 1229 238
rect 1363 272 1421 278
rect 1363 238 1375 272
rect 1409 238 1421 272
rect 1363 232 1421 238
rect -1463 188 -1417 200
rect -1463 -188 -1457 188
rect -1423 -188 -1417 188
rect -1463 -200 -1417 -188
rect -1367 188 -1321 200
rect -1367 -188 -1361 188
rect -1327 -188 -1321 188
rect -1367 -200 -1321 -188
rect -1271 188 -1225 200
rect -1271 -188 -1265 188
rect -1231 -188 -1225 188
rect -1271 -200 -1225 -188
rect -1175 188 -1129 200
rect -1175 -188 -1169 188
rect -1135 -188 -1129 188
rect -1175 -200 -1129 -188
rect -1079 188 -1033 200
rect -1079 -188 -1073 188
rect -1039 -188 -1033 188
rect -1079 -200 -1033 -188
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect 1033 188 1079 200
rect 1033 -188 1039 188
rect 1073 -188 1079 188
rect 1033 -200 1079 -188
rect 1129 188 1175 200
rect 1129 -188 1135 188
rect 1169 -188 1175 188
rect 1129 -200 1175 -188
rect 1225 188 1271 200
rect 1225 -188 1231 188
rect 1265 -188 1271 188
rect 1225 -200 1271 -188
rect 1321 188 1367 200
rect 1321 -188 1327 188
rect 1361 -188 1367 188
rect 1321 -200 1367 -188
rect 1417 188 1463 200
rect 1417 -188 1423 188
rect 1457 -188 1463 188
rect 1417 -200 1463 -188
rect -1421 -238 -1363 -232
rect -1421 -272 -1409 -238
rect -1375 -272 -1363 -238
rect -1421 -278 -1363 -272
rect -1229 -238 -1171 -232
rect -1229 -272 -1217 -238
rect -1183 -272 -1171 -238
rect -1229 -278 -1171 -272
rect -1037 -238 -979 -232
rect -1037 -272 -1025 -238
rect -991 -272 -979 -238
rect -1037 -278 -979 -272
rect -845 -238 -787 -232
rect -845 -272 -833 -238
rect -799 -272 -787 -238
rect -845 -278 -787 -272
rect -653 -238 -595 -232
rect -653 -272 -641 -238
rect -607 -272 -595 -238
rect -653 -278 -595 -272
rect -461 -238 -403 -232
rect -461 -272 -449 -238
rect -415 -272 -403 -238
rect -461 -278 -403 -272
rect -269 -238 -211 -232
rect -269 -272 -257 -238
rect -223 -272 -211 -238
rect -269 -278 -211 -272
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
rect 115 -238 173 -232
rect 115 -272 127 -238
rect 161 -272 173 -238
rect 115 -278 173 -272
rect 307 -238 365 -232
rect 307 -272 319 -238
rect 353 -272 365 -238
rect 307 -278 365 -272
rect 499 -238 557 -232
rect 499 -272 511 -238
rect 545 -272 557 -238
rect 499 -278 557 -272
rect 691 -238 749 -232
rect 691 -272 703 -238
rect 737 -272 749 -238
rect 691 -278 749 -272
rect 883 -238 941 -232
rect 883 -272 895 -238
rect 929 -272 941 -238
rect 883 -278 941 -272
rect 1075 -238 1133 -232
rect 1075 -272 1087 -238
rect 1121 -272 1133 -238
rect 1075 -278 1133 -272
rect 1267 -238 1325 -232
rect 1267 -272 1279 -238
rect 1313 -272 1325 -238
rect 1267 -278 1325 -272
<< properties >>
string FIXED_BBOX -1554 -357 1554 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
