magic
tech sky130A
magscale 1 2
timestamp 1689778135
<< error_p >>
rect -514156 1655671 -514154 1655796
rect -428682 1655712 -428680 1655796
rect -428598 1655671 -428596 1655712
rect -467904 1652732 -467870 1652820
rect -467174 1652732 -467140 1652820
rect -455460 1652732 -455454 1652820
rect -454118 1652732 -454112 1652820
rect -467904 1651572 -467870 1651660
rect -467174 1651572 -467140 1651660
rect -455460 1651572 -455454 1651660
rect -454118 1651572 -454112 1651660
rect 625740 1543178 625744 1543194
rect 646740 1543178 646744 1543194
rect 667740 1543180 667742 1543194
rect 667742 1543178 667744 1543180
rect 688740 1543178 688744 1543194
rect 799740 1543178 799744 1543194
rect 820740 1543178 820744 1543194
rect 841740 1543180 841742 1543194
rect 841742 1543178 841744 1543180
rect 862740 1543178 862744 1543194
rect 625744 1542958 625747 1543178
rect 646744 1542958 646747 1543178
rect 667744 1543137 667747 1543178
rect 688744 1542958 688747 1543178
rect 799744 1542958 799747 1543178
rect 820744 1542958 820747 1543178
rect 841744 1543137 841747 1543178
rect 862744 1542958 862747 1543178
rect 612987 1542909 613215 1542925
rect 633987 1542909 634215 1542925
rect 654987 1542909 655215 1542925
rect 675987 1542909 676215 1542925
rect 786987 1542909 787215 1542925
rect 807987 1542909 808215 1542925
rect 828987 1542909 829215 1542925
rect 849987 1542909 850215 1542925
rect 612984 1542898 612987 1542909
rect 633984 1542898 633987 1542909
rect 654984 1542898 654987 1542909
rect 675984 1542898 675987 1542909
rect 786984 1542898 786987 1542909
rect 807984 1542898 807987 1542909
rect 828984 1542898 828987 1542909
rect 849984 1542898 849987 1542909
rect 275740 1542178 275744 1542194
rect 296740 1542178 296744 1542194
rect 317740 1542178 317744 1542194
rect 338740 1542178 338744 1542194
rect 449740 1542178 449744 1542194
rect 470740 1542178 470744 1542194
rect 491740 1542178 491744 1542194
rect 512740 1542178 512744 1542194
rect 275744 1541958 275747 1542178
rect 296744 1541958 296747 1542178
rect 317744 1541958 317747 1542178
rect 338744 1541958 338747 1542178
rect 449744 1541958 449747 1542178
rect 470744 1541958 470747 1542178
rect 491744 1541958 491747 1542178
rect 512744 1541958 512747 1542178
rect 262987 1541909 263215 1541925
rect 283987 1541909 284215 1541925
rect 304987 1541909 305215 1541925
rect 325987 1541909 326215 1541925
rect 436987 1541909 437215 1541925
rect 457987 1541909 458215 1541925
rect 478987 1541909 479215 1541925
rect 499987 1541909 500215 1541925
rect 262984 1541898 262987 1541909
rect 283984 1541898 283987 1541909
rect 304984 1541898 304987 1541909
rect 325984 1541898 325987 1541909
rect 436984 1541898 436987 1541909
rect 457984 1541898 457987 1541909
rect 478984 1541898 478987 1541909
rect 499984 1541898 499987 1541909
rect 626004 1530442 626016 1530462
rect 647004 1530442 647016 1530462
rect 668004 1530442 668016 1530462
rect 689004 1530442 689016 1530462
rect 800004 1530442 800016 1530462
rect 821004 1530442 821016 1530462
rect 842004 1530442 842016 1530462
rect 863004 1530442 863016 1530462
rect 625780 1530435 626004 1530442
rect 646780 1530435 647004 1530442
rect 667780 1530435 668004 1530442
rect 688780 1530435 689004 1530442
rect 799780 1530435 800004 1530442
rect 820780 1530435 821004 1530442
rect 841780 1530435 842004 1530442
rect 862780 1530435 863004 1530442
rect 613253 1530182 613256 1530190
rect 634253 1530182 634256 1530190
rect 655253 1530182 655256 1530190
rect 676253 1530182 676256 1530190
rect 787253 1530182 787256 1530190
rect 808253 1530182 808256 1530190
rect 829253 1530182 829256 1530190
rect 850253 1530182 850256 1530190
rect 613256 1530166 613260 1530182
rect 634256 1530166 634260 1530182
rect 655256 1530166 655260 1530182
rect 676256 1530166 676260 1530182
rect 787256 1530166 787260 1530182
rect 808256 1530166 808260 1530182
rect 829256 1530166 829260 1530182
rect 850256 1530166 850260 1530182
rect 276004 1529442 276016 1529462
rect 297004 1529442 297016 1529462
rect 318004 1529442 318016 1529462
rect 339004 1529442 339016 1529462
rect 450004 1529442 450016 1529462
rect 471004 1529442 471016 1529462
rect 492004 1529442 492016 1529462
rect 513004 1529442 513016 1529462
rect 275780 1529435 276004 1529442
rect 296780 1529435 297004 1529442
rect 317780 1529435 318004 1529442
rect 338780 1529435 339004 1529442
rect 449780 1529435 450004 1529442
rect 470780 1529435 471004 1529442
rect 491780 1529435 492004 1529442
rect 512780 1529435 513004 1529442
rect 263253 1529182 263256 1529190
rect 284253 1529182 284256 1529190
rect 305253 1529182 305256 1529402
rect 326253 1529182 326256 1529190
rect 437253 1529182 437256 1529190
rect 458253 1529182 458256 1529190
rect 479253 1529182 479256 1529402
rect 500253 1529182 500256 1529190
rect 263256 1529166 263260 1529182
rect 284256 1529166 284260 1529182
rect 305256 1529166 305260 1529182
rect 326256 1529166 326260 1529182
rect 437256 1529166 437260 1529182
rect 458256 1529166 458260 1529182
rect 479256 1529166 479260 1529182
rect 500256 1529166 500260 1529182
rect 608178 1518213 608180 1518297
rect 608262 1518172 608264 1518213
rect 693820 1518172 693822 1518297
rect 782178 1518213 782180 1518297
rect 782262 1518172 782264 1518213
rect 867820 1518172 867822 1518297
rect 258178 1517213 258180 1517297
rect 258262 1517172 258264 1517213
rect 343820 1517172 343822 1517297
rect 432178 1517213 432180 1517297
rect 432262 1517172 432264 1517213
rect 517820 1517172 517822 1517297
rect 591138 1507804 591158 1507816
rect 723298 1507813 723309 1507816
rect 591158 1507580 591165 1507804
rect 723309 1507585 723325 1507813
rect 765138 1507804 765158 1507816
rect 897298 1507813 897309 1507816
rect 765158 1507580 765165 1507804
rect 897309 1507585 897325 1507813
rect 578422 1507544 578642 1507547
rect 710582 1507544 710802 1507547
rect 752422 1507544 752642 1507547
rect 884582 1507544 884802 1507547
rect 578406 1507540 578422 1507544
rect 710566 1507540 710582 1507544
rect 752406 1507540 752422 1507544
rect 884566 1507540 884582 1507544
rect 241138 1506804 241158 1506816
rect 373298 1506813 373309 1506816
rect 241158 1506580 241165 1506804
rect 373309 1506585 373325 1506813
rect 415138 1506804 415158 1506816
rect 547298 1506813 547309 1506816
rect 415158 1506580 415165 1506804
rect 547309 1506585 547325 1506813
rect 228422 1506544 228642 1506547
rect 360582 1506544 360802 1506547
rect 402422 1506544 402642 1506547
rect 534582 1506544 534802 1506547
rect 228406 1506540 228422 1506544
rect 360566 1506540 360582 1506544
rect 402406 1506540 402422 1506544
rect 534566 1506540 534582 1506544
rect 787220 1498962 787825 1498967
rect 591418 1495056 591434 1495060
rect 723578 1495056 723594 1495060
rect 765418 1495056 765434 1495060
rect 897578 1495056 897594 1495060
rect 591198 1495053 591418 1495056
rect 723358 1495053 723578 1495056
rect 765198 1495053 765418 1495056
rect 897358 1495053 897578 1495056
rect 578675 1494787 578691 1495015
rect 710835 1494796 710842 1495020
rect 578691 1494784 578702 1494787
rect 710842 1494784 710862 1494796
rect 752675 1494787 752691 1495015
rect 884835 1494796 884842 1495020
rect 752691 1494784 752702 1494787
rect 884842 1494784 884862 1494796
rect 241418 1494056 241434 1494060
rect 373578 1494056 373594 1494060
rect 415418 1494056 415434 1494060
rect 547578 1494056 547594 1494060
rect 241198 1494053 241418 1494056
rect 373358 1494053 373578 1494056
rect 415198 1494053 415418 1494056
rect 547358 1494053 547578 1494056
rect 228675 1493787 228691 1494015
rect 360835 1493796 360842 1494020
rect 228691 1493784 228702 1493787
rect 360842 1493784 360862 1493796
rect 402675 1493787 402691 1494015
rect 534835 1493796 534842 1494020
rect 402691 1493784 402702 1493787
rect 534842 1493784 534862 1493796
rect 591138 1487804 591158 1487816
rect 723298 1487813 723309 1487816
rect 591158 1487580 591165 1487804
rect 723309 1487585 723325 1487813
rect 765138 1487804 765158 1487816
rect 897298 1487813 897309 1487816
rect 765158 1487580 765165 1487804
rect 897309 1487585 897325 1487813
rect 578422 1487544 578642 1487547
rect 710582 1487544 710802 1487547
rect 752422 1487544 752642 1487547
rect 884582 1487544 884802 1487547
rect 578406 1487540 578422 1487544
rect 710566 1487540 710582 1487544
rect 752406 1487540 752422 1487544
rect 884566 1487540 884582 1487544
rect 241138 1485804 241158 1485816
rect 373298 1485813 373309 1485816
rect 241158 1485580 241165 1485804
rect 373309 1485585 373325 1485813
rect 415138 1485804 415158 1485816
rect 547298 1485813 547309 1485816
rect 415158 1485580 415165 1485804
rect 547309 1485585 547325 1485813
rect 228422 1485544 228642 1485547
rect 360582 1485544 360802 1485547
rect 402422 1485544 402642 1485547
rect 534582 1485544 534802 1485547
rect 228406 1485540 228422 1485544
rect 360566 1485540 360582 1485544
rect 402406 1485540 402422 1485544
rect 534566 1485540 534582 1485544
rect 785940 1483722 786000 1483744
rect 786020 1483722 786080 1483762
rect 591418 1475056 591434 1475060
rect 723578 1475056 723594 1475060
rect 765418 1475056 765434 1475060
rect 897578 1475056 897594 1475060
rect 591198 1475053 591418 1475056
rect 723358 1475053 723578 1475056
rect 765198 1475053 765418 1475056
rect 897358 1475053 897578 1475056
rect 578675 1474787 578691 1475015
rect 710835 1474796 710842 1475020
rect 578691 1474784 578702 1474787
rect 710842 1474784 710862 1474796
rect 752675 1474787 752691 1475015
rect 884835 1474796 884842 1475020
rect 752691 1474784 752702 1474787
rect 884842 1474784 884862 1474796
rect 241418 1473056 241434 1473060
rect 373578 1473056 373594 1473060
rect 415418 1473056 415434 1473060
rect 547578 1473056 547594 1473060
rect 241198 1473053 241418 1473056
rect 373358 1473053 373578 1473056
rect 415198 1473053 415418 1473056
rect 547358 1473053 547578 1473056
rect 228675 1472787 228691 1473015
rect 360835 1472796 360842 1473020
rect 228691 1472784 228702 1472787
rect 360842 1472784 360862 1472796
rect 402675 1472787 402691 1473015
rect 534835 1472796 534842 1473020
rect 402691 1472784 402702 1472787
rect 534842 1472784 534862 1472796
rect 591138 1467804 591158 1467816
rect 723298 1467813 723309 1467816
rect 591158 1467580 591165 1467804
rect 723309 1467585 723325 1467813
rect 765138 1467804 765158 1467816
rect 897298 1467813 897309 1467816
rect 765158 1467580 765165 1467804
rect 897309 1467585 897325 1467813
rect 578422 1467544 578642 1467547
rect 710582 1467544 710802 1467547
rect 752422 1467544 752642 1467547
rect 884582 1467544 884802 1467547
rect 578406 1467540 578422 1467544
rect 710566 1467540 710582 1467544
rect 752406 1467540 752422 1467544
rect 884566 1467540 884582 1467544
rect 229583 1464800 230483 1465115
rect 241138 1464804 241158 1464816
rect 373298 1464813 373309 1464816
rect 241158 1464580 241165 1464804
rect 373309 1464585 373325 1464813
rect 403583 1464800 404483 1465115
rect 415138 1464804 415158 1464816
rect 547298 1464813 547309 1464816
rect 415158 1464580 415165 1464804
rect 547309 1464585 547325 1464813
rect 228422 1464544 228642 1464547
rect 360582 1464544 360802 1464547
rect 402422 1464544 402642 1464547
rect 534582 1464544 534802 1464547
rect 228406 1464311 228422 1464544
rect 241252 1464490 241472 1464493
rect 241472 1464257 241488 1464490
rect 360566 1464311 360582 1464544
rect 373537 1464490 373632 1464493
rect 373632 1464257 373648 1464490
rect 402406 1464311 402422 1464544
rect 415252 1464490 415472 1464493
rect 415472 1464257 415488 1464490
rect 534566 1464311 534582 1464544
rect 547537 1464490 547632 1464493
rect 547632 1464257 547648 1464490
rect 228102 1464224 228322 1464227
rect 228086 1463991 228102 1464224
rect 360256 1464218 360482 1464227
rect 402102 1464224 402322 1464227
rect 241572 1464160 241802 1464173
rect 241802 1463937 241808 1464160
rect 360246 1463991 360256 1464218
rect 373732 1464170 373952 1464173
rect 373952 1464053 373968 1464170
rect 402086 1463991 402102 1464224
rect 534256 1464218 534482 1464227
rect 415572 1464160 415802 1464173
rect 415802 1463937 415808 1464160
rect 534246 1463991 534256 1464218
rect 547732 1464170 547952 1464173
rect 547952 1464053 547968 1464170
rect 227782 1463904 228002 1463907
rect 359942 1463904 360162 1463907
rect 401782 1463904 402002 1463907
rect 533942 1463904 534162 1463907
rect 227766 1463774 227782 1463904
rect 241892 1463850 242112 1463853
rect 242112 1463617 242128 1463850
rect 359926 1463671 359942 1463904
rect 374069 1463850 374272 1463853
rect 374272 1463784 374288 1463850
rect 401766 1463774 401782 1463904
rect 415892 1463850 416112 1463853
rect 416112 1463617 416128 1463850
rect 533926 1463671 533942 1463904
rect 548069 1463850 548272 1463853
rect 548272 1463784 548288 1463850
rect 227420 1463542 227640 1463545
rect 359580 1463542 359800 1463545
rect 401420 1463542 401640 1463545
rect 533580 1463542 533800 1463545
rect 227404 1463518 227420 1463542
rect 242200 1463518 242436 1463531
rect 359564 1463518 359580 1463542
rect 374360 1463518 374596 1463531
rect 401404 1463518 401420 1463542
rect 416200 1463518 416436 1463531
rect 533564 1463518 533580 1463542
rect 548360 1463518 548596 1463531
rect 231275 1463323 231309 1463357
rect 234297 1463323 234331 1463357
rect 367669 1463323 367703 1463357
rect 370691 1463323 370725 1463357
rect 405275 1463323 405309 1463357
rect 408297 1463323 408331 1463357
rect 541669 1463323 541703 1463357
rect 544691 1463323 544725 1463357
rect 231275 1463285 231347 1463321
rect 234259 1463285 234331 1463321
rect 367669 1463285 367741 1463321
rect 370653 1463285 370725 1463321
rect 405275 1463285 405347 1463321
rect 408259 1463285 408331 1463321
rect 541669 1463285 541741 1463321
rect 544653 1463285 544725 1463321
rect 785960 1458902 786000 1459122
rect 786020 1458962 786080 1459122
rect 591418 1455056 591434 1455060
rect 723578 1455056 723594 1455060
rect 765418 1455056 765434 1455060
rect 897578 1455056 897594 1455060
rect 591198 1455053 591418 1455056
rect 723358 1455053 723578 1455056
rect 765198 1455053 765418 1455056
rect 897358 1455053 897578 1455056
rect 578675 1454787 578691 1455015
rect 710835 1454796 710842 1455020
rect 578691 1454784 578702 1454787
rect 710842 1454784 710862 1454796
rect 752675 1454787 752691 1455015
rect 884835 1454796 884842 1455020
rect 752691 1454784 752702 1454787
rect 884842 1454784 884862 1454796
rect 231275 1453279 231347 1453315
rect 234259 1453279 234331 1453315
rect 367669 1453279 367741 1453315
rect 370653 1453279 370725 1453315
rect 405275 1453279 405347 1453315
rect 408259 1453279 408331 1453315
rect 541669 1453279 541741 1453315
rect 544653 1453279 544725 1453315
rect 231275 1453243 231309 1453277
rect 234297 1453243 234331 1453277
rect 367669 1453243 367703 1453277
rect 370691 1453243 370725 1453277
rect 405275 1453243 405309 1453277
rect 408297 1453243 408331 1453277
rect 541669 1453243 541703 1453277
rect 544691 1453243 544725 1453277
rect 227404 1453069 227640 1453082
rect 242420 1453058 242436 1453082
rect 359564 1453069 359800 1453082
rect 374580 1453058 374596 1453082
rect 401404 1453069 401640 1453082
rect 416420 1453058 416436 1453082
rect 533564 1453069 533800 1453082
rect 548580 1453058 548596 1453082
rect 242200 1453055 242420 1453058
rect 374360 1453055 374580 1453058
rect 416200 1453055 416420 1453058
rect 548360 1453055 548580 1453058
rect 227712 1452750 227728 1452816
rect 227728 1452747 227931 1452750
rect 242058 1452696 242074 1452929
rect 359872 1452750 359888 1452983
rect 359888 1452747 360108 1452750
rect 374218 1452696 374234 1452826
rect 401712 1452750 401728 1452816
rect 401728 1452747 401931 1452750
rect 416058 1452696 416074 1452929
rect 533872 1452750 533888 1452983
rect 533888 1452747 534108 1452750
rect 548218 1452696 548234 1452826
rect 241838 1452693 242058 1452696
rect 373998 1452693 374218 1452696
rect 415838 1452693 416058 1452696
rect 547998 1452693 548218 1452696
rect 228032 1452430 228048 1452547
rect 228048 1452427 228268 1452430
rect 241744 1452382 241754 1452609
rect 360192 1452440 360198 1452663
rect 360198 1452427 360428 1452440
rect 241518 1452373 241744 1452382
rect 373898 1452376 373914 1452609
rect 402032 1452430 402048 1452547
rect 402048 1452427 402268 1452430
rect 415744 1452382 415754 1452609
rect 534192 1452440 534198 1452663
rect 534198 1452427 534428 1452440
rect 373678 1452373 373898 1452376
rect 415518 1452373 415744 1452382
rect 547898 1452376 547914 1452609
rect 547678 1452373 547898 1452376
rect 228352 1452110 228368 1452343
rect 228368 1452107 228463 1452110
rect 241418 1452056 241434 1452289
rect 360512 1452110 360528 1452343
rect 360528 1452107 360748 1452110
rect 373578 1452056 373594 1452289
rect 402352 1452110 402368 1452343
rect 402368 1452107 402463 1452110
rect 415418 1452056 415434 1452289
rect 534512 1452110 534528 1452343
rect 534528 1452107 534748 1452110
rect 547578 1452056 547594 1452289
rect 241198 1452053 241418 1452056
rect 373358 1452053 373578 1452056
rect 415198 1452053 415418 1452056
rect 547358 1452053 547578 1452056
rect 228675 1451787 228691 1452015
rect 360835 1451796 360842 1452020
rect 228691 1451784 228702 1451787
rect 360842 1451784 360862 1451796
rect 402675 1451787 402691 1452015
rect 534835 1451796 534842 1452020
rect 402691 1451784 402702 1451787
rect 534842 1451784 534862 1451796
rect 591138 1447804 591158 1447816
rect 723298 1447813 723309 1447816
rect 591158 1447580 591165 1447804
rect 723309 1447585 723325 1447813
rect 765138 1447804 765158 1447816
rect 897298 1447813 897309 1447816
rect 765158 1447580 765165 1447804
rect 897309 1447585 897325 1447813
rect 578422 1447544 578642 1447547
rect 710582 1447544 710802 1447547
rect 752422 1447544 752642 1447547
rect 884582 1447544 884802 1447547
rect 578406 1447540 578422 1447544
rect 710566 1447540 710582 1447544
rect 752406 1447540 752422 1447544
rect 884566 1447540 884582 1447544
rect 241138 1443804 241158 1443816
rect 373298 1443813 373309 1443816
rect 241158 1443580 241165 1443804
rect 373309 1443585 373325 1443813
rect 415138 1443804 415158 1443816
rect 547298 1443813 547309 1443816
rect 415158 1443580 415165 1443804
rect 547309 1443585 547325 1443813
rect 228422 1443544 228642 1443547
rect 360582 1443544 360802 1443547
rect 402422 1443544 402642 1443547
rect 534582 1443544 534802 1443547
rect 228406 1443311 228422 1443544
rect 241252 1443490 241472 1443493
rect 241472 1443257 241488 1443490
rect 360566 1443311 360582 1443544
rect 373537 1443490 373632 1443493
rect 373632 1443257 373648 1443490
rect 402406 1443311 402422 1443544
rect 415252 1443490 415472 1443493
rect 415472 1443257 415488 1443490
rect 534566 1443311 534582 1443544
rect 547537 1443490 547632 1443493
rect 547632 1443257 547648 1443490
rect 228102 1443224 228322 1443227
rect 228086 1442991 228102 1443224
rect 360256 1443218 360482 1443227
rect 402102 1443224 402322 1443227
rect 241572 1443160 241802 1443173
rect 241802 1442937 241808 1443160
rect 360246 1442991 360256 1443218
rect 373732 1443170 373952 1443173
rect 373952 1443053 373968 1443170
rect 402086 1442991 402102 1443224
rect 534256 1443218 534482 1443227
rect 415572 1443160 415802 1443173
rect 415802 1442937 415808 1443160
rect 534246 1442991 534256 1443218
rect 547732 1443170 547952 1443173
rect 547952 1443053 547968 1443170
rect 227782 1442904 228002 1442907
rect 359942 1442904 360162 1442907
rect 401782 1442904 402002 1442907
rect 533942 1442904 534162 1442907
rect 227766 1442774 227782 1442904
rect 241892 1442850 242112 1442853
rect 242112 1442617 242128 1442850
rect 359926 1442671 359942 1442904
rect 374069 1442850 374272 1442853
rect 374272 1442617 374288 1442850
rect 401766 1442774 401782 1442904
rect 415892 1442850 416112 1442853
rect 416112 1442617 416128 1442850
rect 533926 1442671 533942 1442904
rect 548069 1442850 548272 1442853
rect 548272 1442617 548288 1442850
rect 227420 1442542 227640 1442545
rect 359580 1442542 359800 1442545
rect 401420 1442542 401640 1442545
rect 533580 1442542 533800 1442545
rect 227404 1442518 227420 1442542
rect 242200 1442518 242436 1442531
rect 359564 1442518 359580 1442542
rect 374360 1442518 374596 1442531
rect 401404 1442518 401420 1442542
rect 416200 1442518 416436 1442531
rect 533564 1442518 533580 1442542
rect 548360 1442518 548596 1442531
rect 231275 1442323 231309 1442357
rect 234297 1442323 234331 1442357
rect 405275 1442323 405309 1442357
rect 408297 1442323 408331 1442357
rect 231275 1442285 231347 1442321
rect 234259 1442285 234331 1442321
rect 405275 1442285 405347 1442321
rect 408259 1442285 408331 1442321
rect 591418 1435056 591434 1435060
rect 723578 1435056 723594 1435060
rect 765418 1435056 765434 1435060
rect 897578 1435056 897594 1435060
rect 591198 1435053 591418 1435056
rect 723358 1435053 723578 1435056
rect 765198 1435053 765418 1435056
rect 897358 1435053 897578 1435056
rect 578675 1434787 578691 1435015
rect 710835 1434796 710842 1435020
rect 578691 1434784 578702 1434787
rect 710842 1434784 710862 1434796
rect 752675 1434787 752691 1435015
rect 884835 1434796 884842 1435020
rect 752691 1434784 752702 1434787
rect 884842 1434784 884862 1434796
rect 231275 1432279 231347 1432315
rect 234259 1432279 234331 1432315
rect 405275 1432279 405347 1432315
rect 408259 1432279 408331 1432315
rect 231275 1432243 231309 1432277
rect 234297 1432243 234331 1432277
rect 405275 1432243 405309 1432277
rect 408297 1432243 408331 1432277
rect 227404 1432069 227640 1432082
rect 242420 1432058 242436 1432082
rect 359564 1432069 359800 1432082
rect 374580 1432058 374596 1432082
rect 401404 1432069 401640 1432082
rect 416420 1432058 416436 1432082
rect 533564 1432069 533800 1432082
rect 548580 1432058 548596 1432082
rect 242200 1432055 242420 1432058
rect 374360 1432055 374580 1432058
rect 416200 1432055 416420 1432058
rect 548360 1432055 548580 1432058
rect 227712 1431750 227728 1431816
rect 227728 1431747 227931 1431750
rect 242058 1431696 242074 1431929
rect 359872 1431750 359888 1431983
rect 359888 1431747 360108 1431750
rect 374218 1431696 374234 1431929
rect 401712 1431750 401728 1431816
rect 401728 1431747 401931 1431750
rect 416058 1431696 416074 1431929
rect 533872 1431750 533888 1431983
rect 533888 1431747 534108 1431750
rect 548218 1431696 548234 1431929
rect 241838 1431693 242058 1431696
rect 373998 1431693 374218 1431696
rect 415838 1431693 416058 1431696
rect 547998 1431693 548218 1431696
rect 228032 1431430 228048 1431547
rect 228048 1431427 228268 1431430
rect 241744 1431382 241754 1431609
rect 360192 1431440 360198 1431663
rect 360198 1431427 360428 1431440
rect 241518 1431373 241744 1431382
rect 373898 1431376 373914 1431609
rect 402032 1431430 402048 1431547
rect 402048 1431427 402268 1431430
rect 415744 1431382 415754 1431609
rect 534192 1431440 534198 1431663
rect 534198 1431427 534428 1431440
rect 373678 1431373 373898 1431376
rect 415518 1431373 415744 1431382
rect 547898 1431376 547914 1431609
rect 547678 1431373 547898 1431376
rect 228352 1431110 228368 1431343
rect 228368 1431107 228463 1431110
rect 241418 1431056 241434 1431289
rect 360512 1431110 360528 1431343
rect 360528 1431107 360748 1431110
rect 373578 1431056 373594 1431289
rect 402352 1431110 402368 1431343
rect 402368 1431107 402463 1431110
rect 415418 1431056 415434 1431289
rect 534512 1431110 534528 1431343
rect 534528 1431107 534748 1431110
rect 547578 1431056 547594 1431289
rect 241198 1431053 241418 1431056
rect 373358 1431053 373578 1431056
rect 415198 1431053 415418 1431056
rect 547358 1431053 547578 1431056
rect 228675 1430787 228691 1431015
rect 360835 1430796 360842 1431020
rect 228691 1430784 228702 1430787
rect 360842 1430784 360862 1430796
rect 402675 1430787 402691 1431015
rect 534835 1430796 534842 1431020
rect 402691 1430784 402702 1430787
rect 534842 1430784 534862 1430796
rect 591138 1427804 591158 1427816
rect 723298 1427813 723309 1427816
rect 591158 1427580 591165 1427804
rect 723309 1427585 723325 1427813
rect 765138 1427804 765158 1427816
rect 897298 1427813 897309 1427816
rect 765158 1427580 765165 1427804
rect 897309 1427585 897325 1427813
rect 578422 1427544 578642 1427547
rect 710582 1427544 710802 1427547
rect 752422 1427544 752642 1427547
rect 884582 1427544 884802 1427547
rect 578406 1427540 578422 1427544
rect 710566 1427540 710582 1427544
rect 752406 1427540 752422 1427544
rect 884566 1427540 884582 1427544
rect 241138 1422804 241158 1422816
rect 373298 1422813 373309 1422816
rect 241158 1422580 241165 1422804
rect 373309 1422585 373325 1422813
rect 415138 1422804 415158 1422816
rect 547298 1422813 547309 1422816
rect 415158 1422580 415165 1422804
rect 547309 1422585 547325 1422813
rect 228422 1422544 228642 1422547
rect 360582 1422544 360802 1422547
rect 402422 1422544 402642 1422547
rect 534582 1422544 534802 1422547
rect 228406 1422311 228422 1422544
rect 241252 1422490 241472 1422493
rect 241472 1422257 241488 1422490
rect 360566 1422311 360582 1422544
rect 373537 1422490 373632 1422493
rect 373632 1422257 373648 1422490
rect 402406 1422311 402422 1422544
rect 415252 1422490 415472 1422493
rect 415472 1422257 415488 1422490
rect 534566 1422311 534582 1422544
rect 547537 1422490 547632 1422493
rect 547632 1422257 547648 1422490
rect 228102 1422224 228322 1422227
rect 228086 1421991 228102 1422224
rect 360256 1422218 360482 1422227
rect 402102 1422224 402322 1422227
rect 241572 1422160 241802 1422173
rect 241802 1421937 241808 1422160
rect 360246 1421991 360256 1422218
rect 373732 1422170 373952 1422173
rect 373952 1422053 373968 1422170
rect 402086 1421991 402102 1422224
rect 534256 1422218 534482 1422227
rect 415572 1422160 415802 1422173
rect 415802 1421937 415808 1422160
rect 534246 1421991 534256 1422218
rect 547732 1422170 547952 1422173
rect 547952 1422053 547968 1422170
rect 227782 1421904 228002 1421907
rect 359942 1421904 360162 1421907
rect 401782 1421904 402002 1421907
rect 533942 1421904 534162 1421907
rect 227766 1421671 227782 1421904
rect 241892 1421850 242112 1421853
rect 242112 1421617 242128 1421850
rect 359926 1421671 359942 1421904
rect 374069 1421850 374272 1421853
rect 374272 1421784 374288 1421850
rect 401766 1421671 401782 1421904
rect 415892 1421850 416112 1421853
rect 416112 1421617 416128 1421850
rect 533926 1421671 533942 1421904
rect 548069 1421850 548272 1421853
rect 548272 1421784 548288 1421850
rect 227420 1421542 227640 1421545
rect 359580 1421542 359800 1421545
rect 401420 1421542 401640 1421545
rect 533580 1421542 533800 1421545
rect 227404 1421518 227420 1421542
rect 242200 1421518 242436 1421531
rect 359564 1421518 359580 1421542
rect 374360 1421518 374596 1421531
rect 401404 1421518 401420 1421542
rect 416200 1421518 416436 1421531
rect 533564 1421518 533580 1421542
rect 548360 1421518 548596 1421531
rect 367669 1421323 367703 1421357
rect 370691 1421323 370725 1421357
rect 541669 1421323 541703 1421357
rect 544691 1421323 544725 1421357
rect 367669 1421285 367741 1421321
rect 370653 1421285 370725 1421321
rect 541669 1421285 541741 1421321
rect 544653 1421285 544725 1421321
rect 785940 1419162 786000 1423642
rect 785960 1418902 786000 1419162
rect 786020 1418962 786080 1423562
rect 591418 1415056 591434 1415060
rect 723578 1415056 723594 1415060
rect 765418 1415056 765434 1415060
rect 897578 1415056 897594 1415060
rect 591198 1415053 591418 1415056
rect 723358 1415053 723578 1415056
rect 765198 1415053 765418 1415056
rect 897358 1415053 897578 1415056
rect 578675 1414787 578691 1415015
rect 710835 1414796 710842 1415020
rect 578691 1414784 578702 1414787
rect 710842 1414784 710862 1414796
rect 752675 1414787 752691 1415015
rect 884835 1414796 884842 1415020
rect 752691 1414784 752702 1414787
rect 884842 1414784 884862 1414796
rect 367669 1411279 367741 1411315
rect 370653 1411279 370725 1411315
rect 541669 1411279 541741 1411315
rect 544653 1411279 544725 1411315
rect 367669 1411243 367703 1411277
rect 370691 1411243 370725 1411277
rect 541669 1411243 541703 1411277
rect 544691 1411243 544725 1411277
rect 227404 1411069 227640 1411082
rect 242420 1411058 242436 1411082
rect 359564 1411069 359800 1411082
rect 374580 1411058 374596 1411082
rect 401404 1411069 401640 1411082
rect 416420 1411058 416436 1411082
rect 533564 1411069 533800 1411082
rect 548580 1411058 548596 1411082
rect 242200 1411055 242420 1411058
rect 374360 1411055 374580 1411058
rect 416200 1411055 416420 1411058
rect 548360 1411055 548580 1411058
rect 227712 1410750 227728 1410983
rect 227728 1410747 227931 1410750
rect 242058 1410696 242074 1410929
rect 359872 1410750 359888 1410983
rect 359888 1410747 360108 1410750
rect 374218 1410696 374234 1410826
rect 401712 1410750 401728 1410983
rect 401728 1410747 401931 1410750
rect 416058 1410696 416074 1410929
rect 533872 1410750 533888 1410983
rect 533888 1410747 534108 1410750
rect 548218 1410696 548234 1410826
rect 241838 1410693 242058 1410696
rect 373998 1410693 374218 1410696
rect 415838 1410693 416058 1410696
rect 547998 1410693 548218 1410696
rect 228032 1410430 228048 1410547
rect 228048 1410427 228268 1410430
rect 241744 1410382 241754 1410609
rect 360192 1410440 360198 1410663
rect 360198 1410427 360428 1410440
rect 241518 1410373 241744 1410382
rect 373898 1410376 373914 1410609
rect 402032 1410430 402048 1410547
rect 402048 1410427 402268 1410430
rect 415744 1410382 415754 1410609
rect 534192 1410440 534198 1410663
rect 534198 1410427 534428 1410440
rect 373678 1410373 373898 1410376
rect 415518 1410373 415744 1410382
rect 547898 1410376 547914 1410609
rect 547678 1410373 547898 1410376
rect 228352 1410110 228368 1410343
rect 228368 1410107 228463 1410110
rect 241418 1410056 241434 1410289
rect 360512 1410110 360528 1410343
rect 360528 1410107 360748 1410110
rect 373578 1410056 373594 1410289
rect 402352 1410110 402368 1410343
rect 402368 1410107 402463 1410110
rect 415418 1410056 415434 1410289
rect 534512 1410110 534528 1410343
rect 534528 1410107 534748 1410110
rect 547578 1410056 547594 1410289
rect 241198 1410053 241418 1410056
rect 373358 1410053 373578 1410056
rect 415198 1410053 415418 1410056
rect 547358 1410053 547578 1410056
rect 228675 1409787 228691 1410015
rect 360835 1409796 360842 1410020
rect 228691 1409784 228702 1409787
rect 360842 1409784 360862 1409796
rect 402675 1409787 402691 1410015
rect 534835 1409796 534842 1410020
rect 402691 1409784 402702 1409787
rect 534842 1409784 534862 1409796
rect 591138 1407804 591158 1407816
rect 723298 1407813 723309 1407816
rect 591158 1407580 591165 1407804
rect 723309 1407585 723325 1407813
rect 765138 1407804 765158 1407816
rect 897298 1407813 897309 1407816
rect 765158 1407580 765165 1407804
rect 897309 1407585 897325 1407813
rect 578422 1407544 578642 1407547
rect 710582 1407544 710802 1407547
rect 752422 1407544 752642 1407547
rect 884582 1407544 884802 1407547
rect 578406 1407540 578422 1407544
rect 710566 1407540 710582 1407544
rect 752406 1407540 752422 1407544
rect 884566 1407540 884582 1407544
rect 787220 1399000 787825 1399005
rect 591418 1395056 591434 1395060
rect 723578 1395056 723594 1395060
rect 765418 1395056 765434 1395060
rect 897578 1395056 897594 1395060
rect 591198 1395053 591418 1395056
rect 723358 1395053 723578 1395056
rect 765198 1395053 765418 1395056
rect 897358 1395053 897578 1395056
rect 578675 1394787 578691 1395015
rect 710835 1394796 710842 1395020
rect 578691 1394784 578702 1394787
rect 710842 1394784 710862 1394796
rect 752675 1394787 752691 1395015
rect 884835 1394796 884842 1395020
rect 752691 1394784 752702 1394787
rect 884842 1394784 884862 1394796
rect 591138 1387804 591158 1387816
rect 723298 1387813 723309 1387816
rect 591158 1387580 591165 1387804
rect 723309 1387585 723325 1387813
rect 765138 1387804 765158 1387816
rect 897298 1387813 897309 1387816
rect 765158 1387580 765165 1387804
rect 897309 1387585 897325 1387813
rect 578422 1387544 578642 1387547
rect 710582 1387544 710802 1387547
rect 752422 1387544 752642 1387547
rect 884582 1387544 884802 1387547
rect 578406 1387540 578422 1387544
rect 710566 1387540 710582 1387544
rect 752406 1387540 752422 1387544
rect 884566 1387540 884582 1387544
rect 275740 1387418 275744 1387434
rect 296740 1387418 296744 1387434
rect 317540 1387418 317744 1387434
rect 338740 1387418 338744 1387434
rect 449740 1387418 449744 1387434
rect 470740 1387418 470744 1387434
rect 491540 1387418 491744 1387434
rect 512740 1387418 512744 1387434
rect 275744 1387410 275747 1387418
rect 296744 1387410 296747 1387418
rect 317744 1387198 317747 1387418
rect 338744 1387410 338747 1387418
rect 449744 1387410 449747 1387418
rect 470744 1387410 470747 1387418
rect 491744 1387198 491747 1387418
rect 512744 1387410 512747 1387418
rect 262996 1387158 263220 1387165
rect 283996 1387158 284220 1387165
rect 304996 1387158 305220 1387165
rect 325996 1387158 326220 1387165
rect 436996 1387158 437220 1387165
rect 457996 1387158 458220 1387165
rect 478996 1387158 479220 1387165
rect 499996 1387158 500220 1387165
rect 262984 1387138 262996 1387158
rect 283984 1387138 283996 1387158
rect 304984 1387138 304996 1387158
rect 325984 1387138 325996 1387158
rect 436984 1387138 436996 1387158
rect 457984 1387138 457996 1387158
rect 478984 1387138 478996 1387158
rect 499984 1387138 499996 1387158
rect 591418 1375056 591434 1375060
rect 723578 1375056 723594 1375060
rect 765418 1375056 765434 1375060
rect 897578 1375056 897594 1375060
rect 591198 1375053 591418 1375056
rect 723358 1375053 723578 1375056
rect 765198 1375053 765418 1375056
rect 897358 1375053 897578 1375056
rect 578675 1374787 578691 1375015
rect 710835 1374796 710842 1375020
rect 578691 1374784 578702 1374787
rect 710842 1374784 710862 1374796
rect 752675 1374787 752691 1375015
rect 884835 1374796 884842 1375020
rect 752691 1374784 752702 1374787
rect 884842 1374784 884862 1374796
rect 276013 1374691 276016 1374702
rect 297013 1374691 297016 1374702
rect 318013 1374691 318016 1374702
rect 339013 1374691 339016 1374702
rect 450013 1374691 450016 1374702
rect 471013 1374691 471016 1374702
rect 492013 1374691 492016 1374702
rect 513013 1374691 513016 1374702
rect 275785 1374675 276013 1374691
rect 296785 1374675 297013 1374691
rect 317785 1374675 318013 1374691
rect 338785 1374675 339013 1374691
rect 449785 1374675 450013 1374691
rect 470785 1374675 471013 1374691
rect 491785 1374675 492013 1374691
rect 512785 1374675 513013 1374691
rect 263253 1374422 263256 1374642
rect 284253 1374422 284256 1374463
rect 305253 1374422 305256 1374642
rect 263256 1374406 263260 1374422
rect 284256 1374420 284258 1374422
rect 284258 1374406 284260 1374420
rect 305256 1374406 305260 1374422
rect 317690 1374368 317693 1374463
rect 326253 1374422 326256 1374642
rect 437253 1374422 437256 1374642
rect 458253 1374422 458256 1374463
rect 479253 1374422 479256 1374642
rect 326256 1374406 326260 1374422
rect 437256 1374406 437260 1374422
rect 458256 1374420 458258 1374422
rect 458258 1374406 458260 1374420
rect 479256 1374406 479260 1374422
rect 491690 1374368 491693 1374463
rect 500253 1374422 500256 1374642
rect 500256 1374406 500260 1374422
rect 317540 1374352 317690 1374368
rect 491540 1374352 491690 1374368
rect 591138 1367804 591158 1367816
rect 723298 1367813 723309 1367816
rect 591158 1367580 591165 1367804
rect 723309 1367585 723325 1367813
rect 765138 1367804 765158 1367816
rect 897298 1367813 897309 1367816
rect 765158 1367580 765165 1367804
rect 897309 1367585 897325 1367813
rect 578422 1367544 578642 1367547
rect 710582 1367544 710802 1367547
rect 752422 1367544 752642 1367547
rect 884582 1367544 884802 1367547
rect 578406 1367540 578422 1367544
rect 710566 1367540 710582 1367544
rect 752406 1367540 752422 1367544
rect 884566 1367540 884582 1367544
rect 785960 1358940 786000 1359160
rect 786020 1359000 786080 1359160
rect 591418 1355056 591434 1355060
rect 723578 1355056 723594 1355060
rect 765418 1355056 765434 1355060
rect 897578 1355056 897594 1355060
rect 591198 1355053 591418 1355056
rect 723358 1355053 723578 1355056
rect 765198 1355053 765418 1355056
rect 897358 1355053 897578 1355056
rect 578675 1354787 578691 1355015
rect 710835 1354796 710842 1355020
rect 578691 1354784 578702 1354787
rect 710842 1354784 710862 1354796
rect 752675 1354787 752691 1355015
rect 884835 1354796 884842 1355020
rect 752691 1354784 752702 1354787
rect 884842 1354784 884862 1354796
rect 591138 1347804 591158 1347816
rect 723298 1347813 723309 1347816
rect 591158 1347580 591165 1347804
rect 723309 1347585 723325 1347813
rect 765138 1347804 765158 1347816
rect 897298 1347813 897309 1347816
rect 765158 1347580 765165 1347804
rect 897309 1347585 897325 1347813
rect 578422 1347544 578642 1347547
rect 710582 1347544 710802 1347547
rect 752422 1347544 752642 1347547
rect 884582 1347544 884802 1347547
rect 578406 1347540 578422 1347544
rect 710566 1347540 710582 1347544
rect 752406 1347540 752422 1347544
rect 884566 1347540 884582 1347544
rect 275740 1342178 275744 1342194
rect 296740 1342178 296744 1342194
rect 317740 1342178 317744 1342194
rect 338740 1342178 338744 1342194
rect 449740 1342178 449744 1342194
rect 470740 1342178 470744 1342194
rect 491740 1342178 491744 1342194
rect 512740 1342178 512744 1342194
rect 275744 1341958 275747 1342178
rect 296744 1341958 296747 1342178
rect 317744 1341958 317747 1342178
rect 338744 1341958 338747 1342178
rect 449744 1341958 449747 1342178
rect 470744 1341958 470747 1342178
rect 491744 1341958 491747 1342178
rect 512744 1341958 512747 1342178
rect 262987 1341909 263215 1341925
rect 283987 1341909 284215 1341925
rect 304987 1341909 305215 1341925
rect 325987 1341909 326215 1341925
rect 436987 1341909 437215 1341925
rect 457987 1341909 458215 1341925
rect 478987 1341909 479215 1341925
rect 499987 1341909 500215 1341925
rect 262984 1341898 262987 1341909
rect 283984 1341898 283987 1341909
rect 304984 1341898 304987 1341909
rect 325984 1341898 325987 1341909
rect 436984 1341898 436987 1341909
rect 457984 1341898 457987 1341909
rect 478984 1341898 478987 1341909
rect 499984 1341898 499987 1341909
rect 591418 1335056 591434 1335060
rect 723578 1335056 723594 1335060
rect 765418 1335056 765434 1335060
rect 897578 1335056 897594 1335060
rect 591198 1335053 591418 1335056
rect 723358 1335053 723578 1335056
rect 765198 1335053 765418 1335056
rect 897358 1335053 897578 1335056
rect 578675 1334787 578691 1335015
rect 710835 1334796 710842 1335020
rect 578691 1334784 578702 1334787
rect 710842 1334784 710862 1334796
rect 752675 1334787 752691 1335015
rect 884835 1334796 884842 1335020
rect 752691 1334784 752702 1334787
rect 884842 1334784 884862 1334796
rect 276004 1329442 276016 1329462
rect 297004 1329442 297016 1329462
rect 318004 1329442 318016 1329462
rect 339004 1329442 339016 1329462
rect 450004 1329442 450016 1329462
rect 471004 1329442 471016 1329462
rect 492004 1329442 492016 1329462
rect 513004 1329442 513016 1329462
rect 275780 1329435 276004 1329442
rect 296780 1329435 297004 1329442
rect 317780 1329435 318004 1329442
rect 338780 1329435 339004 1329442
rect 449780 1329435 450004 1329442
rect 470780 1329435 471004 1329442
rect 491780 1329435 492004 1329442
rect 512780 1329435 513004 1329442
rect 263253 1329182 263256 1329190
rect 284253 1329182 284256 1329190
rect 305253 1329182 305256 1329402
rect 326253 1329182 326256 1329190
rect 437253 1329182 437256 1329190
rect 458253 1329182 458256 1329190
rect 479253 1329182 479256 1329402
rect 500253 1329182 500256 1329190
rect 263256 1329166 263260 1329182
rect 284256 1329166 284260 1329182
rect 305256 1329166 305260 1329182
rect 326256 1329166 326260 1329182
rect 437256 1329166 437260 1329182
rect 458256 1329166 458260 1329182
rect 479256 1329166 479260 1329182
rect 500256 1329166 500260 1329182
rect 591138 1327804 591158 1327816
rect 723298 1327813 723309 1327816
rect 591158 1327580 591165 1327804
rect 723309 1327585 723325 1327813
rect 765138 1327804 765158 1327816
rect 897298 1327813 897309 1327816
rect 765158 1327580 765165 1327804
rect 897309 1327585 897325 1327813
rect 578422 1327544 578642 1327547
rect 710582 1327544 710802 1327547
rect 752422 1327544 752642 1327547
rect 884582 1327544 884802 1327547
rect 578406 1327540 578422 1327544
rect 710566 1327540 710582 1327544
rect 752406 1327540 752422 1327544
rect 884566 1327540 884582 1327544
rect 785940 1319200 786000 1323680
rect 785960 1318940 786000 1319200
rect 786020 1319000 786080 1323600
rect 258178 1317213 258180 1317297
rect 258262 1317172 258264 1317213
rect 343820 1317172 343822 1317297
rect 432178 1317213 432180 1317297
rect 432262 1317172 432264 1317213
rect 517820 1317172 517822 1317297
rect 591418 1315056 591434 1315060
rect 723578 1315056 723594 1315060
rect 765418 1315056 765434 1315060
rect 897578 1315056 897594 1315060
rect 591198 1315053 591418 1315056
rect 723358 1315053 723578 1315056
rect 765198 1315053 765418 1315056
rect 897358 1315053 897578 1315056
rect 578675 1314787 578691 1315015
rect 710835 1314796 710842 1315020
rect 578691 1314784 578702 1314787
rect 710842 1314784 710862 1314796
rect 752675 1314787 752691 1315015
rect 884835 1314796 884842 1315020
rect 752691 1314784 752702 1314787
rect 884842 1314784 884862 1314796
rect 591138 1307804 591158 1307816
rect 723298 1307813 723309 1307816
rect 591158 1307580 591165 1307804
rect 723309 1307585 723325 1307813
rect 765138 1307804 765158 1307816
rect 897298 1307813 897309 1307816
rect 765158 1307580 765165 1307804
rect 897309 1307585 897325 1307813
rect 578422 1307544 578642 1307547
rect 710582 1307544 710802 1307547
rect 752422 1307544 752642 1307547
rect 884582 1307544 884802 1307547
rect 578406 1307540 578422 1307544
rect 710566 1307540 710582 1307544
rect 752406 1307540 752422 1307544
rect 884566 1307540 884582 1307544
rect 241138 1306804 241158 1306816
rect 373298 1306813 373309 1306816
rect 241158 1306580 241165 1306804
rect 373309 1306585 373325 1306813
rect 415138 1306804 415158 1306816
rect 547298 1306813 547309 1306816
rect 415158 1306580 415165 1306804
rect 547309 1306585 547325 1306813
rect 228422 1306544 228642 1306547
rect 360582 1306544 360802 1306547
rect 402422 1306544 402642 1306547
rect 534582 1306544 534802 1306547
rect 228406 1306540 228422 1306544
rect 360566 1306540 360582 1306544
rect 402406 1306540 402422 1306544
rect 534566 1306540 534582 1306544
rect 787220 1299000 787825 1299005
rect 591418 1295056 591434 1295060
rect 723578 1295056 723594 1295060
rect 765418 1295056 765434 1295060
rect 897578 1295056 897594 1295060
rect 591198 1295053 591418 1295056
rect 723358 1295053 723578 1295056
rect 765198 1295053 765418 1295056
rect 897358 1295053 897578 1295056
rect 578675 1294787 578691 1295015
rect 710835 1294796 710842 1295020
rect 578691 1294784 578702 1294787
rect 710842 1294784 710862 1294796
rect 752675 1294787 752691 1295015
rect 884835 1294796 884842 1295020
rect 752691 1294784 752702 1294787
rect 884842 1294784 884862 1294796
rect 241418 1294056 241434 1294060
rect 373578 1294056 373594 1294060
rect 415418 1294056 415434 1294060
rect 547578 1294056 547594 1294060
rect 241198 1294053 241418 1294056
rect 373358 1294053 373578 1294056
rect 415198 1294053 415418 1294056
rect 547358 1294053 547578 1294056
rect 228675 1293787 228691 1294015
rect 360835 1293796 360842 1294020
rect 228691 1293784 228702 1293787
rect 360842 1293784 360862 1293796
rect 402675 1293787 402691 1294015
rect 534835 1293796 534842 1294020
rect 402691 1293784 402702 1293787
rect 534842 1293784 534862 1293796
rect 591138 1287804 591158 1287816
rect 723298 1287813 723309 1287816
rect 591158 1287580 591165 1287804
rect 723309 1287585 723325 1287813
rect 765138 1287804 765158 1287816
rect 897298 1287813 897309 1287816
rect 765158 1287580 765165 1287804
rect 897309 1287585 897325 1287813
rect 578422 1287544 578642 1287547
rect 710582 1287544 710802 1287547
rect 752422 1287544 752642 1287547
rect 884582 1287544 884802 1287547
rect 578406 1287540 578422 1287544
rect 710566 1287540 710582 1287544
rect 752406 1287540 752422 1287544
rect 884566 1287540 884582 1287544
rect 241138 1285804 241158 1285816
rect 373298 1285813 373309 1285816
rect 241158 1285580 241165 1285804
rect 373309 1285585 373325 1285813
rect 415138 1285804 415158 1285816
rect 547298 1285813 547309 1285816
rect 415158 1285580 415165 1285804
rect 547309 1285585 547325 1285813
rect 228422 1285544 228642 1285547
rect 360582 1285544 360802 1285547
rect 402422 1285544 402642 1285547
rect 534582 1285544 534802 1285547
rect 228406 1285540 228422 1285544
rect 360566 1285540 360582 1285544
rect 402406 1285540 402422 1285544
rect 534566 1285540 534582 1285544
rect 591418 1275056 591434 1275060
rect 723578 1275056 723594 1275060
rect 765418 1275056 765434 1275060
rect 897578 1275056 897594 1275060
rect 591198 1275053 591418 1275056
rect 723358 1275053 723578 1275056
rect 765198 1275053 765418 1275056
rect 897358 1275053 897578 1275056
rect 578675 1274787 578691 1275015
rect 710835 1274796 710842 1275020
rect 578691 1274784 578702 1274787
rect 710842 1274784 710862 1274796
rect 752675 1274787 752691 1275015
rect 884835 1274796 884842 1275020
rect 752691 1274784 752702 1274787
rect 884842 1274784 884862 1274796
rect 241418 1273056 241434 1273060
rect 373578 1273056 373594 1273060
rect 415418 1273056 415434 1273060
rect 547578 1273056 547594 1273060
rect 241198 1273053 241418 1273056
rect 373358 1273053 373578 1273056
rect 415198 1273053 415418 1273056
rect 547358 1273053 547578 1273056
rect 228675 1272787 228691 1273015
rect 360835 1272796 360842 1273020
rect 228691 1272784 228702 1272787
rect 360842 1272784 360862 1272796
rect 402675 1272787 402691 1273015
rect 534835 1272796 534842 1273020
rect 402691 1272784 402702 1272787
rect 534842 1272784 534862 1272796
rect 591138 1267804 591158 1267816
rect 723298 1267813 723309 1267816
rect 591158 1267580 591165 1267804
rect 723309 1267585 723325 1267813
rect 765138 1267804 765158 1267816
rect 897298 1267813 897309 1267816
rect 765158 1267580 765165 1267804
rect 897309 1267585 897325 1267813
rect 578422 1267544 578642 1267547
rect 710582 1267544 710802 1267547
rect 752422 1267544 752642 1267547
rect 884582 1267544 884802 1267547
rect 578406 1267540 578422 1267544
rect 710566 1267540 710582 1267544
rect 752406 1267540 752422 1267544
rect 884566 1267540 884582 1267544
rect 229583 1264800 230483 1265115
rect 241138 1264804 241158 1264816
rect 373298 1264813 373309 1264816
rect 241158 1264580 241165 1264804
rect 373309 1264585 373325 1264813
rect 403583 1264800 404483 1265115
rect 415138 1264804 415158 1264816
rect 547298 1264813 547309 1264816
rect 415158 1264580 415165 1264804
rect 547309 1264585 547325 1264813
rect 228422 1264544 228642 1264547
rect 360582 1264544 360802 1264547
rect 402422 1264544 402642 1264547
rect 534582 1264544 534802 1264547
rect 228406 1264311 228422 1264544
rect 241252 1264490 241472 1264493
rect 241472 1264257 241488 1264490
rect 360566 1264311 360582 1264544
rect 373537 1264490 373632 1264493
rect 373632 1264257 373648 1264490
rect 402406 1264311 402422 1264544
rect 415252 1264490 415472 1264493
rect 415472 1264257 415488 1264490
rect 534566 1264311 534582 1264544
rect 547537 1264490 547632 1264493
rect 547632 1264257 547648 1264490
rect 228102 1264224 228322 1264227
rect 228086 1263991 228102 1264224
rect 360256 1264218 360482 1264227
rect 402102 1264224 402322 1264227
rect 241572 1264160 241802 1264173
rect 241802 1263937 241808 1264160
rect 360246 1263991 360256 1264218
rect 373732 1264170 373952 1264173
rect 373952 1264053 373968 1264170
rect 402086 1263991 402102 1264224
rect 534256 1264218 534482 1264227
rect 415572 1264160 415802 1264173
rect 415802 1263937 415808 1264160
rect 534246 1263991 534256 1264218
rect 547732 1264170 547952 1264173
rect 547952 1264053 547968 1264170
rect 227782 1263904 228002 1263907
rect 359942 1263904 360162 1263907
rect 401782 1263904 402002 1263907
rect 533942 1263904 534162 1263907
rect 227766 1263774 227782 1263904
rect 241892 1263850 242112 1263853
rect 242112 1263617 242128 1263850
rect 359926 1263671 359942 1263904
rect 374069 1263850 374272 1263853
rect 374272 1263784 374288 1263850
rect 401766 1263774 401782 1263904
rect 415892 1263850 416112 1263853
rect 416112 1263617 416128 1263850
rect 533926 1263671 533942 1263904
rect 548069 1263850 548272 1263853
rect 548272 1263784 548288 1263850
rect 227420 1263542 227640 1263545
rect 359580 1263542 359800 1263545
rect 401420 1263542 401640 1263545
rect 533580 1263542 533800 1263545
rect 227404 1263518 227420 1263542
rect 242200 1263518 242436 1263531
rect 359564 1263518 359580 1263542
rect 374360 1263518 374596 1263531
rect 401404 1263518 401420 1263542
rect 416200 1263518 416436 1263531
rect 533564 1263518 533580 1263542
rect 548360 1263518 548596 1263531
rect 231275 1263323 231309 1263357
rect 234297 1263323 234331 1263357
rect 367669 1263323 367703 1263357
rect 370691 1263323 370725 1263357
rect 405275 1263323 405309 1263357
rect 408297 1263323 408331 1263357
rect 541669 1263323 541703 1263357
rect 544691 1263323 544725 1263357
rect 231275 1263285 231347 1263321
rect 234259 1263285 234331 1263321
rect 367669 1263285 367741 1263321
rect 370653 1263285 370725 1263321
rect 405275 1263285 405347 1263321
rect 408259 1263285 408331 1263321
rect 541669 1263285 541741 1263321
rect 544653 1263285 544725 1263321
rect 785960 1258940 786000 1259160
rect 786020 1259000 786080 1259160
rect 591418 1255056 591434 1255060
rect 723578 1255056 723594 1255060
rect 765418 1255056 765434 1255060
rect 897578 1255056 897594 1255060
rect 591198 1255053 591418 1255056
rect 723358 1255053 723578 1255056
rect 765198 1255053 765418 1255056
rect 897358 1255053 897578 1255056
rect 578675 1254787 578691 1255015
rect 710835 1254796 710842 1255020
rect 578691 1254784 578702 1254787
rect 710842 1254784 710862 1254796
rect 752675 1254787 752691 1255015
rect 884835 1254796 884842 1255020
rect 752691 1254784 752702 1254787
rect 884842 1254784 884862 1254796
rect 231275 1253279 231347 1253315
rect 234259 1253279 234331 1253315
rect 367669 1253279 367741 1253315
rect 370653 1253279 370725 1253315
rect 405275 1253279 405347 1253315
rect 408259 1253279 408331 1253315
rect 541669 1253279 541741 1253315
rect 544653 1253279 544725 1253315
rect 231275 1253243 231309 1253277
rect 234297 1253243 234331 1253277
rect 367669 1253243 367703 1253277
rect 370691 1253243 370725 1253277
rect 405275 1253243 405309 1253277
rect 408297 1253243 408331 1253277
rect 541669 1253243 541703 1253277
rect 544691 1253243 544725 1253277
rect 227404 1253069 227640 1253082
rect 242420 1253058 242436 1253082
rect 359564 1253069 359800 1253082
rect 374580 1253058 374596 1253082
rect 401404 1253069 401640 1253082
rect 416420 1253058 416436 1253082
rect 533564 1253069 533800 1253082
rect 548580 1253058 548596 1253082
rect 242200 1253055 242420 1253058
rect 374360 1253055 374580 1253058
rect 416200 1253055 416420 1253058
rect 548360 1253055 548580 1253058
rect 227712 1252750 227728 1252816
rect 227728 1252747 227931 1252750
rect 242058 1252696 242074 1252929
rect 359872 1252750 359888 1252983
rect 359888 1252747 360108 1252750
rect 374218 1252696 374234 1252826
rect 401712 1252750 401728 1252816
rect 401728 1252747 401931 1252750
rect 416058 1252696 416074 1252929
rect 533872 1252750 533888 1252983
rect 533888 1252747 534108 1252750
rect 548218 1252696 548234 1252826
rect 241838 1252693 242058 1252696
rect 373998 1252693 374218 1252696
rect 415838 1252693 416058 1252696
rect 547998 1252693 548218 1252696
rect 228032 1252430 228048 1252547
rect 228048 1252427 228268 1252430
rect 241744 1252382 241754 1252609
rect 360192 1252440 360198 1252663
rect 360198 1252427 360428 1252440
rect 241518 1252373 241744 1252382
rect 373898 1252376 373914 1252609
rect 402032 1252430 402048 1252547
rect 402048 1252427 402268 1252430
rect 415744 1252382 415754 1252609
rect 534192 1252440 534198 1252663
rect 534198 1252427 534428 1252440
rect 373678 1252373 373898 1252376
rect 415518 1252373 415744 1252382
rect 547898 1252376 547914 1252609
rect 547678 1252373 547898 1252376
rect 228352 1252110 228368 1252343
rect 228368 1252107 228463 1252110
rect 241418 1252056 241434 1252289
rect 360512 1252110 360528 1252343
rect 360528 1252107 360748 1252110
rect 373578 1252056 373594 1252289
rect 402352 1252110 402368 1252343
rect 402368 1252107 402463 1252110
rect 415418 1252056 415434 1252289
rect 534512 1252110 534528 1252343
rect 534528 1252107 534748 1252110
rect 547578 1252056 547594 1252289
rect 241198 1252053 241418 1252056
rect 373358 1252053 373578 1252056
rect 415198 1252053 415418 1252056
rect 547358 1252053 547578 1252056
rect 228675 1251787 228691 1252015
rect 360835 1251796 360842 1252020
rect 228691 1251784 228702 1251787
rect 360842 1251784 360862 1251796
rect 402675 1251787 402691 1252015
rect 534835 1251796 534842 1252020
rect 402691 1251784 402702 1251787
rect 534842 1251784 534862 1251796
rect 591138 1247804 591158 1247816
rect 723298 1247813 723309 1247816
rect 591158 1247580 591165 1247804
rect 723309 1247585 723325 1247813
rect 765138 1247804 765158 1247816
rect 897298 1247813 897309 1247816
rect 765158 1247580 765165 1247804
rect 897309 1247585 897325 1247813
rect 578422 1247544 578642 1247547
rect 710582 1247544 710802 1247547
rect 752422 1247544 752642 1247547
rect 884582 1247544 884802 1247547
rect 578406 1247540 578422 1247544
rect 710566 1247540 710582 1247544
rect 752406 1247540 752422 1247544
rect 884566 1247540 884582 1247544
rect 241138 1243804 241158 1243816
rect 373298 1243813 373309 1243816
rect 241158 1243580 241165 1243804
rect 373309 1243585 373325 1243813
rect 415138 1243804 415158 1243816
rect 547298 1243813 547309 1243816
rect 415158 1243580 415165 1243804
rect 547309 1243585 547325 1243813
rect 228422 1243544 228642 1243547
rect 360582 1243544 360802 1243547
rect 402422 1243544 402642 1243547
rect 534582 1243544 534802 1243547
rect 228406 1243311 228422 1243544
rect 241252 1243490 241472 1243493
rect 241472 1243257 241488 1243490
rect 360566 1243311 360582 1243544
rect 373537 1243490 373632 1243493
rect 373632 1243257 373648 1243490
rect 402406 1243311 402422 1243544
rect 415252 1243490 415472 1243493
rect 415472 1243257 415488 1243490
rect 534566 1243311 534582 1243544
rect 547537 1243490 547632 1243493
rect 547632 1243257 547648 1243490
rect 228102 1243224 228322 1243227
rect 228086 1242991 228102 1243224
rect 360256 1243218 360482 1243227
rect 402102 1243224 402322 1243227
rect 241572 1243160 241802 1243173
rect 241802 1242937 241808 1243160
rect 360246 1242991 360256 1243218
rect 373732 1243170 373952 1243173
rect 373952 1243053 373968 1243170
rect 402086 1242991 402102 1243224
rect 534256 1243218 534482 1243227
rect 415572 1243160 415802 1243173
rect 415802 1242937 415808 1243160
rect 534246 1242991 534256 1243218
rect 547732 1243170 547952 1243173
rect 547952 1243053 547968 1243170
rect 227782 1242904 228002 1242907
rect 359942 1242904 360162 1242907
rect 401782 1242904 402002 1242907
rect 533942 1242904 534162 1242907
rect 227766 1242774 227782 1242904
rect 241892 1242850 242112 1242853
rect 242112 1242617 242128 1242850
rect 359926 1242671 359942 1242904
rect 374069 1242850 374272 1242853
rect 374272 1242617 374288 1242850
rect 401766 1242774 401782 1242904
rect 415892 1242850 416112 1242853
rect 416112 1242617 416128 1242850
rect 533926 1242671 533942 1242904
rect 548069 1242850 548272 1242853
rect 548272 1242617 548288 1242850
rect 227420 1242542 227640 1242545
rect 359580 1242542 359800 1242545
rect 401420 1242542 401640 1242545
rect 533580 1242542 533800 1242545
rect 227404 1242518 227420 1242542
rect 242200 1242518 242436 1242531
rect 359564 1242518 359580 1242542
rect 374360 1242518 374596 1242531
rect 401404 1242518 401420 1242542
rect 416200 1242518 416436 1242531
rect 533564 1242518 533580 1242542
rect 548360 1242518 548596 1242531
rect 231275 1242323 231309 1242357
rect 234297 1242323 234331 1242357
rect 405275 1242323 405309 1242357
rect 408297 1242323 408331 1242357
rect 231275 1242285 231347 1242321
rect 234259 1242285 234331 1242321
rect 405275 1242285 405347 1242321
rect 408259 1242285 408331 1242321
rect 591418 1235056 591434 1235060
rect 723578 1235056 723594 1235060
rect 765418 1235056 765434 1235060
rect 897578 1235056 897594 1235060
rect 591198 1235053 591418 1235056
rect 723358 1235053 723578 1235056
rect 765198 1235053 765418 1235056
rect 897358 1235053 897578 1235056
rect 578675 1234787 578691 1235015
rect 710835 1234796 710842 1235020
rect 578691 1234784 578702 1234787
rect 710842 1234784 710862 1234796
rect 752675 1234787 752691 1235015
rect 884835 1234796 884842 1235020
rect 752691 1234784 752702 1234787
rect 884842 1234784 884862 1234796
rect 231275 1232279 231347 1232315
rect 234259 1232279 234331 1232315
rect 405275 1232279 405347 1232315
rect 408259 1232279 408331 1232315
rect 231275 1232243 231309 1232277
rect 234297 1232243 234331 1232277
rect 405275 1232243 405309 1232277
rect 408297 1232243 408331 1232277
rect 227404 1232069 227640 1232082
rect 242420 1232058 242436 1232082
rect 359564 1232069 359800 1232082
rect 374580 1232058 374596 1232082
rect 401404 1232069 401640 1232082
rect 416420 1232058 416436 1232082
rect 533564 1232069 533800 1232082
rect 548580 1232058 548596 1232082
rect 242200 1232055 242420 1232058
rect 374360 1232055 374580 1232058
rect 416200 1232055 416420 1232058
rect 548360 1232055 548580 1232058
rect 227712 1231750 227728 1231816
rect 227728 1231747 227931 1231750
rect 242058 1231696 242074 1231929
rect 359872 1231750 359888 1231983
rect 359888 1231747 360108 1231750
rect 374218 1231696 374234 1231929
rect 401712 1231750 401728 1231816
rect 401728 1231747 401931 1231750
rect 416058 1231696 416074 1231929
rect 533872 1231750 533888 1231983
rect 533888 1231747 534108 1231750
rect 548218 1231696 548234 1231929
rect 241838 1231693 242058 1231696
rect 373998 1231693 374218 1231696
rect 415838 1231693 416058 1231696
rect 547998 1231693 548218 1231696
rect 228032 1231430 228048 1231547
rect 228048 1231427 228268 1231430
rect 241744 1231382 241754 1231609
rect 360192 1231440 360198 1231663
rect 360198 1231427 360428 1231440
rect 241518 1231373 241744 1231382
rect 373898 1231376 373914 1231609
rect 402032 1231430 402048 1231547
rect 402048 1231427 402268 1231430
rect 415744 1231382 415754 1231609
rect 534192 1231440 534198 1231663
rect 534198 1231427 534428 1231440
rect 373678 1231373 373898 1231376
rect 415518 1231373 415744 1231382
rect 547898 1231376 547914 1231609
rect 547678 1231373 547898 1231376
rect 228352 1231110 228368 1231343
rect 228368 1231107 228463 1231110
rect 241418 1231056 241434 1231289
rect 360512 1231110 360528 1231343
rect 360528 1231107 360748 1231110
rect 373578 1231056 373594 1231289
rect 402352 1231110 402368 1231343
rect 402368 1231107 402463 1231110
rect 415418 1231056 415434 1231289
rect 534512 1231110 534528 1231343
rect 534528 1231107 534748 1231110
rect 547578 1231056 547594 1231289
rect 241198 1231053 241418 1231056
rect 373358 1231053 373578 1231056
rect 415198 1231053 415418 1231056
rect 547358 1231053 547578 1231056
rect 228675 1230787 228691 1231015
rect 360835 1230796 360842 1231020
rect 228691 1230784 228702 1230787
rect 360842 1230784 360862 1230796
rect 402675 1230787 402691 1231015
rect 534835 1230796 534842 1231020
rect 402691 1230784 402702 1230787
rect 534842 1230784 534862 1230796
rect 591138 1227804 591158 1227816
rect 723298 1227813 723309 1227816
rect 591158 1227580 591165 1227804
rect 723309 1227585 723325 1227813
rect 765138 1227804 765158 1227816
rect 897298 1227813 897309 1227816
rect 765158 1227580 765165 1227804
rect 897309 1227585 897325 1227813
rect 578422 1227544 578642 1227547
rect 710582 1227544 710802 1227547
rect 752422 1227544 752642 1227547
rect 884582 1227544 884802 1227547
rect 578406 1227540 578422 1227544
rect 710566 1227540 710582 1227544
rect 752406 1227540 752422 1227544
rect 884566 1227540 884582 1227544
rect 241138 1222804 241158 1222816
rect 373298 1222813 373309 1222816
rect 241158 1222580 241165 1222804
rect 373309 1222585 373325 1222813
rect 415138 1222804 415158 1222816
rect 547298 1222813 547309 1222816
rect 415158 1222580 415165 1222804
rect 547309 1222585 547325 1222813
rect 228422 1222544 228642 1222547
rect 360582 1222544 360802 1222547
rect 402422 1222544 402642 1222547
rect 534582 1222544 534802 1222547
rect 228406 1222311 228422 1222544
rect 241252 1222490 241472 1222493
rect 241472 1222257 241488 1222490
rect 360566 1222311 360582 1222544
rect 373537 1222490 373632 1222493
rect 373632 1222257 373648 1222490
rect 402406 1222311 402422 1222544
rect 415252 1222490 415472 1222493
rect 415472 1222257 415488 1222490
rect 534566 1222311 534582 1222544
rect 547537 1222490 547632 1222493
rect 547632 1222257 547648 1222490
rect 228102 1222224 228322 1222227
rect 228086 1221991 228102 1222224
rect 360256 1222218 360482 1222227
rect 402102 1222224 402322 1222227
rect 241572 1222160 241802 1222173
rect 241802 1221937 241808 1222160
rect 360246 1221991 360256 1222218
rect 373732 1222170 373952 1222173
rect 373952 1222053 373968 1222170
rect 402086 1221991 402102 1222224
rect 534256 1222218 534482 1222227
rect 415572 1222160 415802 1222173
rect 415802 1221937 415808 1222160
rect 534246 1221991 534256 1222218
rect 547732 1222170 547952 1222173
rect 547952 1222053 547968 1222170
rect 227782 1221904 228002 1221907
rect 359942 1221904 360162 1221907
rect 401782 1221904 402002 1221907
rect 533942 1221904 534162 1221907
rect 227766 1221671 227782 1221904
rect 241892 1221850 242112 1221853
rect 242112 1221617 242128 1221850
rect 359926 1221671 359942 1221904
rect 374069 1221850 374272 1221853
rect 374272 1221784 374288 1221850
rect 401766 1221671 401782 1221904
rect 415892 1221850 416112 1221853
rect 416112 1221617 416128 1221850
rect 533926 1221671 533942 1221904
rect 548069 1221850 548272 1221853
rect 548272 1221784 548288 1221850
rect 227420 1221542 227640 1221545
rect 359580 1221542 359800 1221545
rect 401420 1221542 401640 1221545
rect 533580 1221542 533800 1221545
rect 227404 1221518 227420 1221542
rect 242200 1221518 242436 1221531
rect 359564 1221518 359580 1221542
rect 374360 1221518 374596 1221531
rect 401404 1221518 401420 1221542
rect 416200 1221518 416436 1221531
rect 533564 1221518 533580 1221542
rect 548360 1221518 548596 1221531
rect 367669 1221323 367703 1221357
rect 370691 1221323 370725 1221357
rect 541669 1221323 541703 1221357
rect 544691 1221323 544725 1221357
rect 367669 1221285 367741 1221321
rect 370653 1221285 370725 1221321
rect 541669 1221285 541741 1221321
rect 544653 1221285 544725 1221321
rect 785940 1219200 786000 1223680
rect 785960 1218940 786000 1219200
rect 786020 1219000 786080 1223600
rect 591418 1215056 591434 1215060
rect 723578 1215056 723594 1215060
rect 765418 1215056 765434 1215060
rect 897578 1215056 897594 1215060
rect 591198 1215053 591418 1215056
rect 723358 1215053 723578 1215056
rect 765198 1215053 765418 1215056
rect 897358 1215053 897578 1215056
rect 578675 1214787 578691 1215015
rect 710835 1214796 710842 1215020
rect 578691 1214784 578702 1214787
rect 710842 1214784 710862 1214796
rect 752675 1214787 752691 1215015
rect 884835 1214796 884842 1215020
rect 752691 1214784 752702 1214787
rect 884842 1214784 884862 1214796
rect 367669 1211279 367741 1211315
rect 370653 1211279 370725 1211315
rect 541669 1211279 541741 1211315
rect 544653 1211279 544725 1211315
rect 367669 1211243 367703 1211277
rect 370691 1211243 370725 1211277
rect 541669 1211243 541703 1211277
rect 544691 1211243 544725 1211277
rect 227404 1211069 227640 1211082
rect 242420 1211058 242436 1211082
rect 359564 1211069 359800 1211082
rect 374580 1211058 374596 1211082
rect 401404 1211069 401640 1211082
rect 416420 1211058 416436 1211082
rect 533564 1211069 533800 1211082
rect 548580 1211058 548596 1211082
rect 242200 1211055 242420 1211058
rect 374360 1211055 374580 1211058
rect 416200 1211055 416420 1211058
rect 548360 1211055 548580 1211058
rect 227712 1210750 227728 1210983
rect 227728 1210747 227931 1210750
rect 242058 1210696 242074 1210929
rect 359872 1210750 359888 1210983
rect 359888 1210747 360108 1210750
rect 374218 1210696 374234 1210826
rect 401712 1210750 401728 1210983
rect 401728 1210747 401931 1210750
rect 416058 1210696 416074 1210929
rect 533872 1210750 533888 1210983
rect 533888 1210747 534108 1210750
rect 548218 1210696 548234 1210826
rect 241838 1210693 242058 1210696
rect 373998 1210693 374218 1210696
rect 415838 1210693 416058 1210696
rect 547998 1210693 548218 1210696
rect 228032 1210430 228048 1210547
rect 228048 1210427 228268 1210430
rect 241744 1210382 241754 1210609
rect 360192 1210440 360198 1210663
rect 360198 1210427 360428 1210440
rect 241518 1210373 241744 1210382
rect 373898 1210376 373914 1210609
rect 402032 1210430 402048 1210547
rect 402048 1210427 402268 1210430
rect 415744 1210382 415754 1210609
rect 534192 1210440 534198 1210663
rect 534198 1210427 534428 1210440
rect 373678 1210373 373898 1210376
rect 415518 1210373 415744 1210382
rect 547898 1210376 547914 1210609
rect 547678 1210373 547898 1210376
rect 228352 1210110 228368 1210343
rect 228368 1210107 228463 1210110
rect 241418 1210056 241434 1210289
rect 360512 1210110 360528 1210343
rect 360528 1210107 360748 1210110
rect 373578 1210056 373594 1210289
rect 402352 1210110 402368 1210343
rect 402368 1210107 402463 1210110
rect 415418 1210056 415434 1210289
rect 534512 1210110 534528 1210343
rect 534528 1210107 534748 1210110
rect 547578 1210056 547594 1210289
rect 241198 1210053 241418 1210056
rect 373358 1210053 373578 1210056
rect 415198 1210053 415418 1210056
rect 547358 1210053 547578 1210056
rect 228675 1209787 228691 1210015
rect 360835 1209796 360842 1210020
rect 228691 1209784 228702 1209787
rect 360842 1209784 360862 1209796
rect 402675 1209787 402691 1210015
rect 534835 1209796 534842 1210020
rect 402691 1209784 402702 1209787
rect 534842 1209784 534862 1209796
rect 591138 1207804 591158 1207816
rect 723298 1207813 723309 1207816
rect 591158 1207580 591165 1207804
rect 723309 1207585 723325 1207813
rect 765138 1207804 765158 1207816
rect 897298 1207813 897309 1207816
rect 765158 1207580 765165 1207804
rect 897309 1207585 897325 1207813
rect 578422 1207544 578642 1207547
rect 710582 1207544 710802 1207547
rect 752422 1207544 752642 1207547
rect 884582 1207544 884802 1207547
rect 578406 1207540 578422 1207544
rect 710566 1207540 710582 1207544
rect 752406 1207540 752422 1207544
rect 884566 1207540 884582 1207544
rect 611080 1203720 611680 1203731
rect 611000 1203640 611600 1203651
rect 787220 1198800 787825 1198805
rect 591418 1195056 591434 1195060
rect 723578 1195056 723594 1195060
rect 765418 1195056 765434 1195060
rect 897578 1195056 897594 1195060
rect 591198 1195053 591418 1195056
rect 723358 1195053 723578 1195056
rect 765198 1195053 765418 1195056
rect 897358 1195053 897578 1195056
rect 578675 1194787 578691 1195015
rect 710835 1194796 710842 1195020
rect 578691 1194784 578702 1194787
rect 710842 1194784 710862 1194796
rect 752675 1194787 752691 1195015
rect 884835 1194796 884842 1195020
rect 752691 1194784 752702 1194787
rect 884842 1194784 884862 1194796
rect 591138 1187804 591158 1187816
rect 723298 1187813 723309 1187816
rect 591158 1187580 591165 1187804
rect 723309 1187585 723325 1187813
rect 765138 1187804 765158 1187816
rect 897298 1187813 897309 1187816
rect 765158 1187580 765165 1187804
rect 897309 1187585 897325 1187813
rect 578422 1187544 578642 1187547
rect 710582 1187544 710802 1187547
rect 752422 1187544 752642 1187547
rect 884582 1187544 884802 1187547
rect 578406 1187540 578422 1187544
rect 710566 1187540 710582 1187544
rect 752406 1187540 752422 1187544
rect 884566 1187540 884582 1187544
rect 275740 1187418 275744 1187434
rect 296740 1187418 296744 1187434
rect 317540 1187418 317744 1187434
rect 338740 1187418 338744 1187434
rect 449740 1187418 449744 1187434
rect 470740 1187418 470744 1187434
rect 491540 1187418 491744 1187434
rect 512740 1187418 512744 1187434
rect 275744 1187410 275747 1187418
rect 296744 1187410 296747 1187418
rect 317744 1187198 317747 1187418
rect 338744 1187410 338747 1187418
rect 449744 1187410 449747 1187418
rect 470744 1187410 470747 1187418
rect 491744 1187198 491747 1187418
rect 512744 1187410 512747 1187418
rect 262996 1187158 263220 1187165
rect 283996 1187158 284220 1187165
rect 304996 1187158 305220 1187165
rect 325996 1187158 326220 1187165
rect 436996 1187158 437220 1187165
rect 457996 1187158 458220 1187165
rect 478996 1187158 479220 1187165
rect 499996 1187158 500220 1187165
rect 262984 1187138 262996 1187158
rect 283984 1187138 283996 1187158
rect 304984 1187138 304996 1187158
rect 325984 1187138 325996 1187158
rect 436984 1187138 436996 1187158
rect 457984 1187138 457996 1187158
rect 478984 1187138 478996 1187158
rect 499984 1187138 499996 1187158
rect 785940 1183560 786000 1183680
rect 786020 1183560 786080 1183600
rect 591418 1175056 591434 1175060
rect 723578 1175056 723594 1175060
rect 765418 1175056 765434 1175060
rect 897578 1175056 897594 1175060
rect 591198 1175053 591418 1175056
rect 723358 1175053 723578 1175056
rect 765198 1175053 765418 1175056
rect 897358 1175053 897578 1175056
rect 578675 1174787 578691 1175015
rect 710835 1174796 710842 1175020
rect 578691 1174784 578702 1174787
rect 710842 1174784 710862 1174796
rect 752675 1174787 752691 1175015
rect 884835 1174796 884842 1175020
rect 752691 1174784 752702 1174787
rect 884842 1174784 884862 1174796
rect 276013 1174691 276016 1174702
rect 297013 1174691 297016 1174702
rect 318013 1174691 318016 1174702
rect 339013 1174691 339016 1174702
rect 450013 1174691 450016 1174702
rect 471013 1174691 471016 1174702
rect 492013 1174691 492016 1174702
rect 513013 1174691 513016 1174702
rect 275785 1174675 276013 1174691
rect 296785 1174675 297013 1174691
rect 317785 1174675 318013 1174691
rect 338785 1174675 339013 1174691
rect 449785 1174675 450013 1174691
rect 470785 1174675 471013 1174691
rect 491785 1174675 492013 1174691
rect 512785 1174675 513013 1174691
rect 263253 1174422 263256 1174642
rect 284253 1174422 284256 1174463
rect 305253 1174422 305256 1174642
rect 263256 1174406 263260 1174422
rect 284256 1174420 284258 1174422
rect 284258 1174406 284260 1174420
rect 305256 1174406 305260 1174422
rect 317690 1174368 317693 1174463
rect 326253 1174422 326256 1174642
rect 437253 1174422 437256 1174642
rect 458253 1174422 458256 1174463
rect 479253 1174422 479256 1174642
rect 326256 1174406 326260 1174422
rect 437256 1174406 437260 1174422
rect 458256 1174420 458258 1174422
rect 458258 1174406 458260 1174420
rect 479256 1174406 479260 1174422
rect 491690 1174368 491693 1174463
rect 500253 1174422 500256 1174642
rect 500256 1174406 500260 1174422
rect 317540 1174352 317690 1174368
rect 491540 1174352 491690 1174368
rect 591138 1167804 591158 1167816
rect 723298 1167813 723309 1167816
rect 591158 1167580 591165 1167804
rect 723309 1167585 723325 1167813
rect 765138 1167804 765158 1167816
rect 897298 1167813 897309 1167816
rect 765158 1167580 765165 1167804
rect 897309 1167585 897325 1167813
rect 578422 1167544 578642 1167547
rect 710582 1167544 710802 1167547
rect 752422 1167544 752642 1167547
rect 884582 1167544 884802 1167547
rect 578406 1167540 578422 1167544
rect 710566 1167540 710582 1167544
rect 752406 1167540 752422 1167544
rect 884566 1167540 884582 1167544
rect 785960 1158744 786000 1158960
rect 786020 1158800 786080 1158960
rect 591418 1155056 591434 1155060
rect 723578 1155056 723594 1155060
rect 765418 1155056 765434 1155060
rect 897578 1155056 897594 1155060
rect 591198 1155053 591418 1155056
rect 723358 1155053 723578 1155056
rect 765198 1155053 765418 1155056
rect 897358 1155053 897578 1155056
rect 578675 1154787 578691 1155015
rect 710835 1154796 710842 1155020
rect 578691 1154784 578702 1154787
rect 710842 1154784 710862 1154796
rect 752675 1154787 752691 1155015
rect 884835 1154796 884842 1155020
rect 752691 1154784 752702 1154787
rect 884842 1154784 884862 1154796
rect 591138 1147804 591158 1147816
rect 723298 1147813 723309 1147816
rect 591158 1147580 591165 1147804
rect 723309 1147585 723325 1147813
rect 765138 1147804 765158 1147816
rect 897298 1147813 897309 1147816
rect 765158 1147580 765165 1147804
rect 897309 1147585 897325 1147813
rect 578422 1147544 578642 1147547
rect 710582 1147544 710802 1147547
rect 752422 1147544 752642 1147547
rect 884582 1147544 884802 1147547
rect 578406 1147540 578422 1147544
rect 710566 1147540 710582 1147544
rect 752406 1147540 752422 1147544
rect 884566 1147540 884582 1147544
rect 275740 1142178 275744 1142194
rect 296740 1142178 296744 1142194
rect 317740 1142178 317744 1142194
rect 338740 1142178 338744 1142194
rect 449740 1142178 449744 1142194
rect 470740 1142178 470744 1142194
rect 491740 1142178 491744 1142194
rect 512740 1142178 512744 1142194
rect 275744 1141958 275747 1142178
rect 296744 1141958 296747 1142178
rect 317744 1141958 317747 1142178
rect 338744 1141958 338747 1142178
rect 449744 1141958 449747 1142178
rect 470744 1141958 470747 1142178
rect 491744 1141958 491747 1142178
rect 512744 1141958 512747 1142178
rect 262987 1141909 263215 1141925
rect 283987 1141909 284215 1141925
rect 304987 1141909 305215 1141925
rect 325987 1141909 326215 1141925
rect 436987 1141909 437215 1141925
rect 457987 1141909 458215 1141925
rect 478987 1141909 479215 1141925
rect 499987 1141909 500215 1141925
rect 262984 1141898 262987 1141909
rect 283984 1141898 283987 1141909
rect 304984 1141898 304987 1141909
rect 325984 1141898 325987 1141909
rect 436984 1141898 436987 1141909
rect 457984 1141898 457987 1141909
rect 478984 1141898 478987 1141909
rect 499984 1141898 499987 1141909
rect 591418 1135056 591434 1135060
rect 723578 1135056 723594 1135060
rect 765418 1135056 765434 1135060
rect 897578 1135056 897594 1135060
rect 591198 1135053 591418 1135056
rect 723358 1135053 723578 1135056
rect 765198 1135053 765418 1135056
rect 897358 1135053 897578 1135056
rect 578675 1134787 578691 1135015
rect 710835 1134796 710842 1135020
rect 578691 1134784 578702 1134787
rect 710842 1134784 710862 1134796
rect 752675 1134787 752691 1135015
rect 884835 1134796 884842 1135020
rect 752691 1134784 752702 1134787
rect 884842 1134784 884862 1134796
rect 276004 1129442 276016 1129462
rect 297004 1129442 297016 1129462
rect 318004 1129442 318016 1129462
rect 339004 1129442 339016 1129462
rect 450004 1129442 450016 1129462
rect 471004 1129442 471016 1129462
rect 492004 1129442 492016 1129462
rect 513004 1129442 513016 1129462
rect 275780 1129435 276004 1129442
rect 296780 1129435 297004 1129442
rect 317780 1129435 318004 1129442
rect 338780 1129435 339004 1129442
rect 449780 1129435 450004 1129442
rect 470780 1129435 471004 1129442
rect 491780 1129435 492004 1129442
rect 512780 1129435 513004 1129442
rect 263253 1129182 263256 1129190
rect 284253 1129182 284256 1129190
rect 305253 1129182 305256 1129402
rect 326253 1129182 326256 1129190
rect 437253 1129182 437256 1129190
rect 458253 1129182 458256 1129190
rect 479253 1129182 479256 1129402
rect 500253 1129182 500256 1129190
rect 263256 1129166 263260 1129182
rect 284256 1129166 284260 1129182
rect 305256 1129166 305260 1129182
rect 326256 1129166 326260 1129182
rect 437256 1129166 437260 1129182
rect 458256 1129166 458260 1129182
rect 479256 1129166 479260 1129182
rect 500256 1129166 500260 1129182
rect 591138 1127804 591158 1127816
rect 723298 1127813 723309 1127816
rect 591158 1127580 591165 1127804
rect 723309 1127585 723325 1127813
rect 765138 1127804 765158 1127816
rect 897298 1127813 897309 1127816
rect 765158 1127580 765165 1127804
rect 897309 1127585 897325 1127813
rect 578422 1127544 578642 1127547
rect 710582 1127544 710802 1127547
rect 752422 1127544 752642 1127547
rect 884582 1127544 884802 1127547
rect 578406 1127540 578422 1127544
rect 710566 1127540 710582 1127544
rect 752406 1127540 752422 1127544
rect 884566 1127540 884582 1127544
rect 785940 1119000 786000 1123480
rect 785960 1118744 786000 1119000
rect 786020 1118800 786080 1123400
rect 258178 1117213 258180 1117297
rect 258262 1117172 258264 1117213
rect 343820 1117172 343822 1117297
rect 432178 1117213 432180 1117297
rect 432262 1117172 432264 1117213
rect 517820 1117172 517822 1117297
rect 591418 1115056 591434 1115060
rect 723578 1115056 723594 1115060
rect 765418 1115056 765434 1115060
rect 897578 1115056 897594 1115060
rect 591198 1115053 591418 1115056
rect 723358 1115053 723578 1115056
rect 765198 1115053 765418 1115056
rect 897358 1115053 897578 1115056
rect 578675 1114787 578691 1115015
rect 710835 1114796 710842 1115020
rect 578691 1114784 578702 1114787
rect 710842 1114784 710862 1114796
rect 752675 1114787 752691 1115015
rect 884835 1114796 884842 1115020
rect 752691 1114784 752702 1114787
rect 884842 1114784 884862 1114796
rect 591138 1107804 591158 1107816
rect 723298 1107813 723309 1107816
rect 591158 1107580 591165 1107804
rect 723309 1107585 723325 1107813
rect 765138 1107804 765158 1107816
rect 897298 1107813 897309 1107816
rect 765158 1107580 765165 1107804
rect 897309 1107585 897325 1107813
rect 578422 1107544 578642 1107547
rect 710582 1107544 710802 1107547
rect 752422 1107544 752642 1107547
rect 884582 1107544 884802 1107547
rect 578406 1107540 578422 1107544
rect 710566 1107540 710582 1107544
rect 752406 1107540 752422 1107544
rect 884566 1107540 884582 1107544
rect 241138 1106804 241158 1106816
rect 373298 1106813 373309 1106816
rect 241158 1106580 241165 1106804
rect 373309 1106585 373325 1106813
rect 415138 1106804 415158 1106816
rect 547298 1106813 547309 1106816
rect 415158 1106580 415165 1106804
rect 547309 1106585 547325 1106813
rect 228422 1106544 228642 1106547
rect 360582 1106544 360802 1106547
rect 402422 1106544 402642 1106547
rect 534582 1106544 534802 1106547
rect 228406 1106540 228422 1106544
rect 360566 1106540 360582 1106544
rect 402406 1106540 402422 1106544
rect 534566 1106540 534582 1106544
rect 611080 1103720 611680 1103731
rect 611000 1103640 611600 1103651
rect 787220 1098800 787825 1098805
rect 591418 1095056 591434 1095060
rect 723578 1095056 723594 1095060
rect 765418 1095056 765434 1095060
rect 897578 1095056 897594 1095060
rect 591198 1095053 591418 1095056
rect 723358 1095053 723578 1095056
rect 765198 1095053 765418 1095056
rect 897358 1095053 897578 1095056
rect 578675 1094787 578691 1095015
rect 710835 1094796 710842 1095020
rect 578691 1094784 578702 1094787
rect 710842 1094784 710862 1094796
rect 752675 1094787 752691 1095015
rect 884835 1094796 884842 1095020
rect 752691 1094784 752702 1094787
rect 884842 1094784 884862 1094796
rect 241418 1094056 241434 1094060
rect 373578 1094056 373594 1094060
rect 415418 1094056 415434 1094060
rect 547578 1094056 547594 1094060
rect 241198 1094053 241418 1094056
rect 373358 1094053 373578 1094056
rect 415198 1094053 415418 1094056
rect 547358 1094053 547578 1094056
rect 228675 1093787 228691 1094015
rect 360835 1093796 360842 1094020
rect 228691 1093784 228702 1093787
rect 360842 1093784 360862 1093796
rect 402675 1093787 402691 1094015
rect 534835 1093796 534842 1094020
rect 402691 1093784 402702 1093787
rect 534842 1093784 534862 1093796
rect 591138 1087804 591158 1087816
rect 723298 1087813 723309 1087816
rect 591158 1087580 591165 1087804
rect 723309 1087585 723325 1087813
rect 765138 1087804 765158 1087816
rect 897298 1087813 897309 1087816
rect 765158 1087580 765165 1087804
rect 897309 1087585 897325 1087813
rect 578422 1087544 578642 1087547
rect 710582 1087544 710802 1087547
rect 752422 1087544 752642 1087547
rect 884582 1087544 884802 1087547
rect 578406 1087540 578422 1087544
rect 710566 1087540 710582 1087544
rect 752406 1087540 752422 1087544
rect 884566 1087540 884582 1087544
rect 241138 1085804 241158 1085816
rect 373298 1085813 373309 1085816
rect 241158 1085580 241165 1085804
rect 373309 1085585 373325 1085813
rect 415138 1085804 415158 1085816
rect 547298 1085813 547309 1085816
rect 415158 1085580 415165 1085804
rect 547309 1085585 547325 1085813
rect 228422 1085544 228642 1085547
rect 360582 1085544 360802 1085547
rect 402422 1085544 402642 1085547
rect 534582 1085544 534802 1085547
rect 228406 1085540 228422 1085544
rect 360566 1085540 360582 1085544
rect 402406 1085540 402422 1085544
rect 534566 1085540 534582 1085544
rect 785940 1083560 786000 1083680
rect 786020 1083560 786080 1083600
rect 591418 1075056 591434 1075060
rect 723578 1075056 723594 1075060
rect 765418 1075056 765434 1075060
rect 897578 1075056 897594 1075060
rect 591198 1075053 591418 1075056
rect 723358 1075053 723578 1075056
rect 765198 1075053 765418 1075056
rect 897358 1075053 897578 1075056
rect 578675 1074787 578691 1075015
rect 710835 1074796 710842 1075020
rect 578691 1074784 578702 1074787
rect 710842 1074784 710862 1074796
rect 752675 1074787 752691 1075015
rect 884835 1074796 884842 1075020
rect 752691 1074784 752702 1074787
rect 884842 1074784 884862 1074796
rect 241418 1073056 241434 1073060
rect 373578 1073056 373594 1073060
rect 415418 1073056 415434 1073060
rect 547578 1073056 547594 1073060
rect 241198 1073053 241418 1073056
rect 373358 1073053 373578 1073056
rect 415198 1073053 415418 1073056
rect 547358 1073053 547578 1073056
rect 228675 1072787 228691 1073015
rect 360835 1072796 360842 1073020
rect 228691 1072784 228702 1072787
rect 360842 1072784 360862 1072796
rect 402675 1072787 402691 1073015
rect 534835 1072796 534842 1073020
rect 402691 1072784 402702 1072787
rect 534842 1072784 534862 1072796
rect 591138 1067804 591158 1067816
rect 723298 1067813 723309 1067816
rect 591158 1067580 591165 1067804
rect 723309 1067585 723325 1067813
rect 765138 1067804 765158 1067816
rect 897298 1067813 897309 1067816
rect 765158 1067580 765165 1067804
rect 897309 1067585 897325 1067813
rect 578422 1067544 578642 1067547
rect 710582 1067544 710802 1067547
rect 752422 1067544 752642 1067547
rect 884582 1067544 884802 1067547
rect 578406 1067540 578422 1067544
rect 710566 1067540 710582 1067544
rect 752406 1067540 752422 1067544
rect 884566 1067540 884582 1067544
rect 229583 1064800 230483 1065115
rect 241138 1064804 241158 1064816
rect 373298 1064813 373309 1064816
rect 241158 1064580 241165 1064804
rect 373309 1064585 373325 1064813
rect 403583 1064800 404483 1065115
rect 415138 1064804 415158 1064816
rect 547298 1064813 547309 1064816
rect 415158 1064580 415165 1064804
rect 547309 1064585 547325 1064813
rect 228422 1064544 228642 1064547
rect 360582 1064544 360802 1064547
rect 402422 1064544 402642 1064547
rect 534582 1064544 534802 1064547
rect 228406 1064311 228422 1064544
rect 241252 1064490 241472 1064493
rect 241472 1064257 241488 1064490
rect 360566 1064311 360582 1064544
rect 373537 1064490 373632 1064493
rect 373632 1064257 373648 1064490
rect 402406 1064311 402422 1064544
rect 415252 1064490 415472 1064493
rect 415472 1064257 415488 1064490
rect 534566 1064311 534582 1064544
rect 547537 1064490 547632 1064493
rect 547632 1064257 547648 1064490
rect 228102 1064224 228322 1064227
rect 228086 1063991 228102 1064224
rect 360256 1064218 360482 1064227
rect 402102 1064224 402322 1064227
rect 241572 1064160 241802 1064173
rect 241802 1063937 241808 1064160
rect 360246 1063991 360256 1064218
rect 373732 1064170 373952 1064173
rect 373952 1064053 373968 1064170
rect 402086 1063991 402102 1064224
rect 534256 1064218 534482 1064227
rect 415572 1064160 415802 1064173
rect 415802 1063937 415808 1064160
rect 534246 1063991 534256 1064218
rect 547732 1064170 547952 1064173
rect 547952 1064053 547968 1064170
rect 227782 1063904 228002 1063907
rect 359942 1063904 360162 1063907
rect 401782 1063904 402002 1063907
rect 533942 1063904 534162 1063907
rect 227766 1063774 227782 1063904
rect 241892 1063850 242112 1063853
rect 242112 1063617 242128 1063850
rect 359926 1063671 359942 1063904
rect 374069 1063850 374272 1063853
rect 374272 1063784 374288 1063850
rect 401766 1063774 401782 1063904
rect 415892 1063850 416112 1063853
rect 416112 1063617 416128 1063850
rect 533926 1063671 533942 1063904
rect 548069 1063850 548272 1063853
rect 548272 1063784 548288 1063850
rect 227420 1063542 227640 1063545
rect 359580 1063542 359800 1063545
rect 401420 1063542 401640 1063545
rect 533580 1063542 533800 1063545
rect 227404 1063518 227420 1063542
rect 242200 1063518 242436 1063531
rect 359564 1063518 359580 1063542
rect 374360 1063518 374596 1063531
rect 401404 1063518 401420 1063542
rect 416200 1063518 416436 1063531
rect 533564 1063518 533580 1063542
rect 548360 1063518 548596 1063531
rect 231275 1063323 231309 1063357
rect 234297 1063323 234331 1063357
rect 367669 1063323 367703 1063357
rect 370691 1063323 370725 1063357
rect 405275 1063323 405309 1063357
rect 408297 1063323 408331 1063357
rect 541669 1063323 541703 1063357
rect 544691 1063323 544725 1063357
rect 231275 1063285 231347 1063321
rect 234259 1063285 234331 1063321
rect 367669 1063285 367741 1063321
rect 370653 1063285 370725 1063321
rect 405275 1063285 405347 1063321
rect 408259 1063285 408331 1063321
rect 541669 1063285 541741 1063321
rect 544653 1063285 544725 1063321
rect 785960 1058744 786000 1058960
rect 786020 1058800 786080 1058960
rect 591418 1055056 591434 1055060
rect 723578 1055056 723594 1055060
rect 765418 1055056 765434 1055060
rect 897578 1055056 897594 1055060
rect 591198 1055053 591418 1055056
rect 723358 1055053 723578 1055056
rect 765198 1055053 765418 1055056
rect 897358 1055053 897578 1055056
rect 578675 1054787 578691 1055015
rect 710835 1054796 710842 1055020
rect 578691 1054784 578702 1054787
rect 710842 1054784 710862 1054796
rect 752675 1054787 752691 1055015
rect 884835 1054796 884842 1055020
rect 752691 1054784 752702 1054787
rect 884842 1054784 884862 1054796
rect 231275 1053279 231347 1053315
rect 234259 1053279 234331 1053315
rect 367669 1053279 367741 1053315
rect 370653 1053279 370725 1053315
rect 405275 1053279 405347 1053315
rect 408259 1053279 408331 1053315
rect 541669 1053279 541741 1053315
rect 544653 1053279 544725 1053315
rect 231275 1053243 231309 1053277
rect 234297 1053243 234331 1053277
rect 367669 1053243 367703 1053277
rect 370691 1053243 370725 1053277
rect 405275 1053243 405309 1053277
rect 408297 1053243 408331 1053277
rect 541669 1053243 541703 1053277
rect 544691 1053243 544725 1053277
rect 227404 1053069 227640 1053082
rect 242420 1053058 242436 1053082
rect 359564 1053069 359800 1053082
rect 374580 1053058 374596 1053082
rect 401404 1053069 401640 1053082
rect 416420 1053058 416436 1053082
rect 533564 1053069 533800 1053082
rect 548580 1053058 548596 1053082
rect 242200 1053055 242420 1053058
rect 374360 1053055 374580 1053058
rect 416200 1053055 416420 1053058
rect 548360 1053055 548580 1053058
rect 227712 1052750 227728 1052816
rect 227728 1052747 227931 1052750
rect 242058 1052696 242074 1052929
rect 359872 1052750 359888 1052983
rect 359888 1052747 360108 1052750
rect 374218 1052696 374234 1052826
rect 401712 1052750 401728 1052816
rect 401728 1052747 401931 1052750
rect 416058 1052696 416074 1052929
rect 533872 1052750 533888 1052983
rect 533888 1052747 534108 1052750
rect 548218 1052696 548234 1052826
rect 241838 1052693 242058 1052696
rect 373998 1052693 374218 1052696
rect 415838 1052693 416058 1052696
rect 547998 1052693 548218 1052696
rect 228032 1052430 228048 1052547
rect 228048 1052427 228268 1052430
rect 241744 1052382 241754 1052609
rect 360192 1052440 360198 1052663
rect 360198 1052427 360428 1052440
rect 241518 1052373 241744 1052382
rect 373898 1052376 373914 1052609
rect 402032 1052430 402048 1052547
rect 402048 1052427 402268 1052430
rect 415744 1052382 415754 1052609
rect 534192 1052440 534198 1052663
rect 534198 1052427 534428 1052440
rect 373678 1052373 373898 1052376
rect 415518 1052373 415744 1052382
rect 547898 1052376 547914 1052609
rect 547678 1052373 547898 1052376
rect 228352 1052110 228368 1052343
rect 228368 1052107 228463 1052110
rect 241418 1052056 241434 1052289
rect 360512 1052110 360528 1052343
rect 360528 1052107 360748 1052110
rect 373578 1052056 373594 1052289
rect 402352 1052110 402368 1052343
rect 402368 1052107 402463 1052110
rect 415418 1052056 415434 1052289
rect 534512 1052110 534528 1052343
rect 534528 1052107 534748 1052110
rect 547578 1052056 547594 1052289
rect 241198 1052053 241418 1052056
rect 373358 1052053 373578 1052056
rect 415198 1052053 415418 1052056
rect 547358 1052053 547578 1052056
rect 228675 1051787 228691 1052015
rect 360835 1051796 360842 1052020
rect 228691 1051784 228702 1051787
rect 360842 1051784 360862 1051796
rect 402675 1051787 402691 1052015
rect 534835 1051796 534842 1052020
rect 402691 1051784 402702 1051787
rect 534842 1051784 534862 1051796
rect 591138 1047804 591158 1047816
rect 723298 1047813 723309 1047816
rect 591158 1047580 591165 1047804
rect 723309 1047585 723325 1047813
rect 765138 1047804 765158 1047816
rect 897298 1047813 897309 1047816
rect 765158 1047580 765165 1047804
rect 897309 1047585 897325 1047813
rect 578422 1047544 578642 1047547
rect 710582 1047544 710802 1047547
rect 752422 1047544 752642 1047547
rect 884582 1047544 884802 1047547
rect 578406 1047540 578422 1047544
rect 710566 1047540 710582 1047544
rect 752406 1047540 752422 1047544
rect 884566 1047540 884582 1047544
rect 241138 1043804 241158 1043816
rect 373298 1043813 373309 1043816
rect 241158 1043580 241165 1043804
rect 373309 1043585 373325 1043813
rect 415138 1043804 415158 1043816
rect 547298 1043813 547309 1043816
rect 415158 1043580 415165 1043804
rect 547309 1043585 547325 1043813
rect 228422 1043544 228642 1043547
rect 360582 1043544 360802 1043547
rect 402422 1043544 402642 1043547
rect 534582 1043544 534802 1043547
rect 228406 1043311 228422 1043544
rect 241252 1043490 241472 1043493
rect 241472 1043257 241488 1043490
rect 360566 1043311 360582 1043544
rect 373537 1043490 373632 1043493
rect 373632 1043257 373648 1043490
rect 402406 1043311 402422 1043544
rect 415252 1043490 415472 1043493
rect 415472 1043257 415488 1043490
rect 534566 1043311 534582 1043544
rect 547537 1043490 547632 1043493
rect 547632 1043257 547648 1043490
rect 228102 1043224 228322 1043227
rect 228086 1042991 228102 1043224
rect 360256 1043218 360482 1043227
rect 402102 1043224 402322 1043227
rect 241572 1043160 241802 1043173
rect 241802 1042937 241808 1043160
rect 360246 1042991 360256 1043218
rect 373732 1043170 373952 1043173
rect 373952 1043053 373968 1043170
rect 402086 1042991 402102 1043224
rect 534256 1043218 534482 1043227
rect 415572 1043160 415802 1043173
rect 415802 1042937 415808 1043160
rect 534246 1042991 534256 1043218
rect 547732 1043170 547952 1043173
rect 547952 1043053 547968 1043170
rect 227782 1042904 228002 1042907
rect 359942 1042904 360162 1042907
rect 401782 1042904 402002 1042907
rect 533942 1042904 534162 1042907
rect 227766 1042774 227782 1042904
rect 241892 1042850 242112 1042853
rect 242112 1042617 242128 1042850
rect 359926 1042671 359942 1042904
rect 374069 1042850 374272 1042853
rect 374272 1042617 374288 1042850
rect 401766 1042774 401782 1042904
rect 415892 1042850 416112 1042853
rect 416112 1042617 416128 1042850
rect 533926 1042671 533942 1042904
rect 548069 1042850 548272 1042853
rect 548272 1042617 548288 1042850
rect 227420 1042542 227640 1042545
rect 359580 1042542 359800 1042545
rect 401420 1042542 401640 1042545
rect 533580 1042542 533800 1042545
rect 227404 1042518 227420 1042542
rect 242200 1042518 242436 1042531
rect 359564 1042518 359580 1042542
rect 374360 1042518 374596 1042531
rect 401404 1042518 401420 1042542
rect 416200 1042518 416436 1042531
rect 533564 1042518 533580 1042542
rect 548360 1042518 548596 1042531
rect 231275 1042323 231309 1042357
rect 234297 1042323 234331 1042357
rect 405275 1042323 405309 1042357
rect 408297 1042323 408331 1042357
rect 231275 1042285 231347 1042321
rect 234259 1042285 234331 1042321
rect 405275 1042285 405347 1042321
rect 408259 1042285 408331 1042321
rect 591418 1035056 591434 1035060
rect 723578 1035056 723594 1035060
rect 765418 1035056 765434 1035060
rect 897578 1035056 897594 1035060
rect 591198 1035053 591418 1035056
rect 723358 1035053 723578 1035056
rect 765198 1035053 765418 1035056
rect 897358 1035053 897578 1035056
rect 578675 1034787 578691 1035015
rect 710835 1034796 710842 1035020
rect 578691 1034784 578702 1034787
rect 710842 1034784 710862 1034796
rect 752675 1034787 752691 1035015
rect 884835 1034796 884842 1035020
rect 752691 1034784 752702 1034787
rect 884842 1034784 884862 1034796
rect 231275 1032279 231347 1032315
rect 234259 1032279 234331 1032315
rect 405275 1032279 405347 1032315
rect 408259 1032279 408331 1032315
rect 231275 1032243 231309 1032277
rect 234297 1032243 234331 1032277
rect 405275 1032243 405309 1032277
rect 408297 1032243 408331 1032277
rect 227404 1032069 227640 1032082
rect 242420 1032058 242436 1032082
rect 359564 1032069 359800 1032082
rect 374580 1032058 374596 1032082
rect 401404 1032069 401640 1032082
rect 416420 1032058 416436 1032082
rect 533564 1032069 533800 1032082
rect 548580 1032058 548596 1032082
rect 242200 1032055 242420 1032058
rect 374360 1032055 374580 1032058
rect 416200 1032055 416420 1032058
rect 548360 1032055 548580 1032058
rect 227712 1031750 227728 1031816
rect 227728 1031747 227931 1031750
rect 242058 1031696 242074 1031929
rect 359872 1031750 359888 1031983
rect 359888 1031747 360108 1031750
rect 374218 1031696 374234 1031929
rect 401712 1031750 401728 1031816
rect 401728 1031747 401931 1031750
rect 416058 1031696 416074 1031929
rect 533872 1031750 533888 1031983
rect 533888 1031747 534108 1031750
rect 548218 1031696 548234 1031929
rect 241838 1031693 242058 1031696
rect 373998 1031693 374218 1031696
rect 415838 1031693 416058 1031696
rect 547998 1031693 548218 1031696
rect 228032 1031430 228048 1031547
rect 228048 1031427 228268 1031430
rect 241744 1031382 241754 1031609
rect 360192 1031440 360198 1031663
rect 360198 1031427 360428 1031440
rect 241518 1031373 241744 1031382
rect 373898 1031376 373914 1031609
rect 402032 1031430 402048 1031547
rect 402048 1031427 402268 1031430
rect 415744 1031382 415754 1031609
rect 534192 1031440 534198 1031663
rect 534198 1031427 534428 1031440
rect 373678 1031373 373898 1031376
rect 415518 1031373 415744 1031382
rect 547898 1031376 547914 1031609
rect 547678 1031373 547898 1031376
rect 228352 1031110 228368 1031343
rect 228368 1031107 228463 1031110
rect 241418 1031056 241434 1031289
rect 360512 1031110 360528 1031343
rect 360528 1031107 360748 1031110
rect 373578 1031056 373594 1031289
rect 402352 1031110 402368 1031343
rect 402368 1031107 402463 1031110
rect 415418 1031056 415434 1031289
rect 534512 1031110 534528 1031343
rect 534528 1031107 534748 1031110
rect 547578 1031056 547594 1031289
rect 241198 1031053 241418 1031056
rect 373358 1031053 373578 1031056
rect 415198 1031053 415418 1031056
rect 547358 1031053 547578 1031056
rect 228675 1030787 228691 1031015
rect 360835 1030796 360842 1031020
rect 228691 1030784 228702 1030787
rect 360842 1030784 360862 1030796
rect 402675 1030787 402691 1031015
rect 534835 1030796 534842 1031020
rect 402691 1030784 402702 1030787
rect 534842 1030784 534862 1030796
rect 591138 1027804 591158 1027816
rect 723298 1027813 723309 1027816
rect 591158 1027580 591165 1027804
rect 723309 1027585 723325 1027813
rect 765138 1027804 765158 1027816
rect 897298 1027813 897309 1027816
rect 765158 1027580 765165 1027804
rect 897309 1027585 897325 1027813
rect 578422 1027544 578642 1027547
rect 710582 1027544 710802 1027547
rect 752422 1027544 752642 1027547
rect 884582 1027544 884802 1027547
rect 578406 1027540 578422 1027544
rect 710566 1027540 710582 1027544
rect 752406 1027540 752422 1027544
rect 884566 1027540 884582 1027544
rect 241138 1022804 241158 1022816
rect 373298 1022813 373309 1022816
rect 241158 1022580 241165 1022804
rect 373309 1022585 373325 1022813
rect 415138 1022804 415158 1022816
rect 547298 1022813 547309 1022816
rect 415158 1022580 415165 1022804
rect 547309 1022585 547325 1022813
rect 228422 1022544 228642 1022547
rect 360582 1022544 360802 1022547
rect 402422 1022544 402642 1022547
rect 534582 1022544 534802 1022547
rect 228406 1022311 228422 1022544
rect 241252 1022490 241472 1022493
rect 241472 1022257 241488 1022490
rect 360566 1022311 360582 1022544
rect 373537 1022490 373632 1022493
rect 373632 1022257 373648 1022490
rect 402406 1022311 402422 1022544
rect 415252 1022490 415472 1022493
rect 415472 1022257 415488 1022490
rect 534566 1022311 534582 1022544
rect 547537 1022490 547632 1022493
rect 547632 1022257 547648 1022490
rect 228102 1022224 228322 1022227
rect 228086 1021991 228102 1022224
rect 360256 1022218 360482 1022227
rect 402102 1022224 402322 1022227
rect 241572 1022160 241802 1022173
rect 241802 1021937 241808 1022160
rect 360246 1021991 360256 1022218
rect 373732 1022170 373952 1022173
rect 373952 1022053 373968 1022170
rect 402086 1021991 402102 1022224
rect 534256 1022218 534482 1022227
rect 415572 1022160 415802 1022173
rect 415802 1021937 415808 1022160
rect 534246 1021991 534256 1022218
rect 547732 1022170 547952 1022173
rect 547952 1022053 547968 1022170
rect 227782 1021904 228002 1021907
rect 359942 1021904 360162 1021907
rect 401782 1021904 402002 1021907
rect 533942 1021904 534162 1021907
rect 227766 1021671 227782 1021904
rect 241892 1021850 242112 1021853
rect 242112 1021617 242128 1021850
rect 359926 1021671 359942 1021904
rect 374069 1021850 374272 1021853
rect 374272 1021784 374288 1021850
rect 401766 1021671 401782 1021904
rect 415892 1021850 416112 1021853
rect 416112 1021617 416128 1021850
rect 533926 1021671 533942 1021904
rect 548069 1021850 548272 1021853
rect 548272 1021784 548288 1021850
rect 227420 1021542 227640 1021545
rect 359580 1021542 359800 1021545
rect 401420 1021542 401640 1021545
rect 533580 1021542 533800 1021545
rect 227404 1021518 227420 1021542
rect 242200 1021518 242436 1021531
rect 359564 1021518 359580 1021542
rect 374360 1021518 374596 1021531
rect 401404 1021518 401420 1021542
rect 416200 1021518 416436 1021531
rect 533564 1021518 533580 1021542
rect 548360 1021518 548596 1021531
rect 367669 1021323 367703 1021357
rect 370691 1021323 370725 1021357
rect 541669 1021323 541703 1021357
rect 544691 1021323 544725 1021357
rect 367669 1021285 367741 1021321
rect 370653 1021285 370725 1021321
rect 541669 1021285 541741 1021321
rect 544653 1021285 544725 1021321
rect 785940 1019000 786000 1023480
rect 785960 1018744 786000 1019000
rect 786020 1018800 786080 1023400
rect 591418 1015056 591434 1015060
rect 723578 1015056 723594 1015060
rect 765418 1015056 765434 1015060
rect 897578 1015056 897594 1015060
rect 591198 1015053 591418 1015056
rect 723358 1015053 723578 1015056
rect 765198 1015053 765418 1015056
rect 897358 1015053 897578 1015056
rect 578675 1014787 578691 1015015
rect 710835 1014796 710842 1015020
rect 578691 1014784 578702 1014787
rect 710842 1014784 710862 1014796
rect 752675 1014787 752691 1015015
rect 884835 1014796 884842 1015020
rect 752691 1014784 752702 1014787
rect 884842 1014784 884862 1014796
rect 367669 1011279 367741 1011315
rect 370653 1011279 370725 1011315
rect 541669 1011279 541741 1011315
rect 544653 1011279 544725 1011315
rect 367669 1011243 367703 1011277
rect 370691 1011243 370725 1011277
rect 541669 1011243 541703 1011277
rect 544691 1011243 544725 1011277
rect 227404 1011069 227640 1011082
rect 242420 1011058 242436 1011082
rect 359564 1011069 359800 1011082
rect 374580 1011058 374596 1011082
rect 401404 1011069 401640 1011082
rect 416420 1011058 416436 1011082
rect 533564 1011069 533800 1011082
rect 548580 1011058 548596 1011082
rect 242200 1011055 242420 1011058
rect 374360 1011055 374580 1011058
rect 416200 1011055 416420 1011058
rect 548360 1011055 548580 1011058
rect 227712 1010750 227728 1010983
rect 227728 1010747 227931 1010750
rect 242058 1010696 242074 1010929
rect 359872 1010750 359888 1010983
rect 359888 1010747 360108 1010750
rect 374218 1010696 374234 1010826
rect 401712 1010750 401728 1010983
rect 401728 1010747 401931 1010750
rect 416058 1010696 416074 1010929
rect 533872 1010750 533888 1010983
rect 533888 1010747 534108 1010750
rect 548218 1010696 548234 1010826
rect 241838 1010693 242058 1010696
rect 373998 1010693 374218 1010696
rect 415838 1010693 416058 1010696
rect 547998 1010693 548218 1010696
rect 228032 1010430 228048 1010547
rect 228048 1010427 228268 1010430
rect 241744 1010382 241754 1010609
rect 360192 1010440 360198 1010663
rect 360198 1010427 360428 1010440
rect 241518 1010373 241744 1010382
rect 373898 1010376 373914 1010609
rect 402032 1010430 402048 1010547
rect 402048 1010427 402268 1010430
rect 415744 1010382 415754 1010609
rect 534192 1010440 534198 1010663
rect 534198 1010427 534428 1010440
rect 373678 1010373 373898 1010376
rect 415518 1010373 415744 1010382
rect 547898 1010376 547914 1010609
rect 547678 1010373 547898 1010376
rect 228352 1010110 228368 1010343
rect 228368 1010107 228463 1010110
rect 241418 1010056 241434 1010289
rect 360512 1010110 360528 1010343
rect 360528 1010107 360748 1010110
rect 373578 1010056 373594 1010289
rect 402352 1010110 402368 1010343
rect 402368 1010107 402463 1010110
rect 415418 1010056 415434 1010289
rect 534512 1010110 534528 1010343
rect 534528 1010107 534748 1010110
rect 547578 1010056 547594 1010289
rect 241198 1010053 241418 1010056
rect 373358 1010053 373578 1010056
rect 415198 1010053 415418 1010056
rect 547358 1010053 547578 1010056
rect 228675 1009787 228691 1010015
rect 360835 1009796 360842 1010020
rect 228691 1009784 228702 1009787
rect 360842 1009784 360862 1009796
rect 402675 1009787 402691 1010015
rect 534835 1009796 534842 1010020
rect 402691 1009784 402702 1009787
rect 534842 1009784 534862 1009796
rect 591138 1007804 591158 1007816
rect 723298 1007813 723309 1007816
rect 591158 1007580 591165 1007804
rect 723309 1007585 723325 1007813
rect 765138 1007804 765158 1007816
rect 897298 1007813 897309 1007816
rect 765158 1007580 765165 1007804
rect 897309 1007585 897325 1007813
rect 578422 1007544 578642 1007547
rect 710582 1007544 710802 1007547
rect 752422 1007544 752642 1007547
rect 884582 1007544 884802 1007547
rect 578406 1007540 578422 1007544
rect 710566 1007540 710582 1007544
rect 752406 1007540 752422 1007544
rect 884566 1007540 884582 1007544
rect 787220 997000 787825 997005
rect 591418 995056 591434 995060
rect 723578 995056 723594 995060
rect 765418 995056 765434 995060
rect 897578 995056 897594 995060
rect 591198 995053 591418 995056
rect 723358 995053 723578 995056
rect 765198 995053 765418 995056
rect 897358 995053 897578 995056
rect 578675 994787 578691 995015
rect 710835 994796 710842 995020
rect 578691 994784 578702 994787
rect 710842 994784 710862 994796
rect 752675 994787 752691 995015
rect 884835 994796 884842 995020
rect 752691 994784 752702 994787
rect 884842 994784 884862 994796
rect 591138 987804 591158 987816
rect 723298 987813 723309 987816
rect 591158 987580 591165 987804
rect 723309 987585 723325 987813
rect 765138 987804 765158 987816
rect 897298 987813 897309 987816
rect 765158 987580 765165 987804
rect 897309 987585 897325 987813
rect 578422 987544 578642 987547
rect 710582 987544 710802 987547
rect 752422 987544 752642 987547
rect 884582 987544 884802 987547
rect 578406 987540 578422 987544
rect 710566 987540 710582 987544
rect 752406 987540 752422 987544
rect 884566 987540 884582 987544
rect 275740 987418 275744 987434
rect 296740 987418 296744 987434
rect 317540 987418 317744 987434
rect 338740 987418 338744 987434
rect 449740 987418 449744 987434
rect 470740 987418 470744 987434
rect 491540 987418 491744 987434
rect 512740 987418 512744 987434
rect 275744 987410 275747 987418
rect 296744 987410 296747 987418
rect 317744 987198 317747 987418
rect 338744 987410 338747 987418
rect 449744 987410 449747 987418
rect 470744 987410 470747 987418
rect 491744 987198 491747 987418
rect 512744 987410 512747 987418
rect 262996 987158 263220 987165
rect 283996 987158 284220 987165
rect 304996 987158 305220 987165
rect 325996 987158 326220 987165
rect 436996 987158 437220 987165
rect 457996 987158 458220 987165
rect 478996 987158 479220 987165
rect 499996 987158 500220 987165
rect 262984 987138 262996 987158
rect 283984 987138 283996 987158
rect 304984 987138 304996 987158
rect 325984 987138 325996 987158
rect 436984 987138 436996 987158
rect 457984 987138 457996 987158
rect 478984 987138 478996 987158
rect 499984 987138 499996 987158
rect 785940 981760 786000 981880
rect 786020 981760 786080 981800
rect 591418 975056 591434 975060
rect 723578 975056 723594 975060
rect 765418 975056 765434 975060
rect 897578 975056 897594 975060
rect 591198 975053 591418 975056
rect 723358 975053 723578 975056
rect 765198 975053 765418 975056
rect 897358 975053 897578 975056
rect 578675 974787 578691 975015
rect 710835 974796 710842 975020
rect 578691 974784 578702 974787
rect 710842 974784 710862 974796
rect 752675 974787 752691 975015
rect 884835 974796 884842 975020
rect 752691 974784 752702 974787
rect 884842 974784 884862 974796
rect 276013 974691 276016 974702
rect 297013 974691 297016 974702
rect 318013 974691 318016 974702
rect 339013 974691 339016 974702
rect 450013 974691 450016 974702
rect 471013 974691 471016 974702
rect 492013 974691 492016 974702
rect 513013 974691 513016 974702
rect 275785 974675 276013 974691
rect 296785 974675 297013 974691
rect 317785 974675 318013 974691
rect 338785 974675 339013 974691
rect 449785 974675 450013 974691
rect 470785 974675 471013 974691
rect 491785 974675 492013 974691
rect 512785 974675 513013 974691
rect 263253 974422 263256 974642
rect 284253 974422 284256 974463
rect 305253 974422 305256 974642
rect 263256 974406 263260 974422
rect 284256 974420 284258 974422
rect 284258 974406 284260 974420
rect 305256 974406 305260 974422
rect 317690 974368 317693 974463
rect 326253 974422 326256 974642
rect 437253 974422 437256 974642
rect 458253 974422 458256 974463
rect 479253 974422 479256 974642
rect 326256 974406 326260 974422
rect 437256 974406 437260 974422
rect 458256 974420 458258 974422
rect 458258 974406 458260 974420
rect 479256 974406 479260 974422
rect 491690 974368 491693 974463
rect 500253 974422 500256 974642
rect 500256 974406 500260 974422
rect 317540 974352 317690 974368
rect 491540 974352 491690 974368
rect 591138 967804 591158 967816
rect 723298 967813 723309 967816
rect 591158 967580 591165 967804
rect 723309 967585 723325 967813
rect 765138 967804 765158 967816
rect 897298 967813 897309 967816
rect 765158 967580 765165 967804
rect 897309 967585 897325 967813
rect 578422 967544 578642 967547
rect 710582 967544 710802 967547
rect 752422 967544 752642 967547
rect 884582 967544 884802 967547
rect 578406 967540 578422 967544
rect 710566 967540 710582 967544
rect 752406 967540 752422 967544
rect 884566 967540 884582 967544
rect 591418 955056 591434 955060
rect 723578 955056 723594 955060
rect 765418 955056 765434 955060
rect 897578 955056 897594 955060
rect 591198 955053 591418 955056
rect 723358 955053 723578 955056
rect 765198 955053 765418 955056
rect 897358 955053 897578 955056
rect 578675 954787 578691 955015
rect 710835 954796 710842 955020
rect 578691 954784 578702 954787
rect 710842 954784 710862 954796
rect 752675 954787 752691 955015
rect 884835 954796 884842 955020
rect 752691 954784 752702 954787
rect 884842 954784 884862 954796
rect 591138 947804 591158 947816
rect 723298 947813 723309 947816
rect 591158 947580 591165 947804
rect 723309 947585 723325 947813
rect 765138 947804 765158 947816
rect 897298 947813 897309 947816
rect 765158 947580 765165 947804
rect 897309 947585 897325 947813
rect 578422 947544 578642 947547
rect 710582 947544 710802 947547
rect 752422 947544 752642 947547
rect 884582 947544 884802 947547
rect 578406 947540 578422 947544
rect 710566 947540 710582 947544
rect 752406 947540 752422 947544
rect 884566 947540 884582 947544
rect 275740 942178 275744 942194
rect 296740 942178 296744 942194
rect 317740 942178 317744 942194
rect 338740 942178 338744 942194
rect 449740 942178 449744 942194
rect 470740 942178 470744 942194
rect 491740 942178 491744 942194
rect 512740 942178 512744 942194
rect 275744 941958 275747 942178
rect 296744 941958 296747 942178
rect 317744 941958 317747 942178
rect 338744 941958 338747 942178
rect 449744 941958 449747 942178
rect 470744 941958 470747 942178
rect 491744 941958 491747 942178
rect 512744 941958 512747 942178
rect 262987 941909 263215 941925
rect 283987 941909 284215 941925
rect 304987 941909 305215 941925
rect 325987 941909 326215 941925
rect 436987 941909 437215 941925
rect 457987 941909 458215 941925
rect 478987 941909 479215 941925
rect 499987 941909 500215 941925
rect 262984 941898 262987 941909
rect 283984 941898 283987 941909
rect 304984 941898 304987 941909
rect 325984 941898 325987 941909
rect 436984 941898 436987 941909
rect 457984 941898 457987 941909
rect 478984 941898 478987 941909
rect 499984 941898 499987 941909
rect 591418 935056 591434 935060
rect 723578 935056 723594 935060
rect 765418 935056 765434 935060
rect 897578 935056 897594 935060
rect 591198 935053 591418 935056
rect 723358 935053 723578 935056
rect 765198 935053 765418 935056
rect 897358 935053 897578 935056
rect 578675 934787 578691 935015
rect 710835 934796 710842 935020
rect 578691 934784 578702 934787
rect 710842 934784 710862 934796
rect 752675 934787 752691 935015
rect 884835 934796 884842 935020
rect 752691 934784 752702 934787
rect 884842 934784 884862 934796
rect 276004 929442 276016 929462
rect 297004 929442 297016 929462
rect 318004 929442 318016 929462
rect 339004 929442 339016 929462
rect 450004 929442 450016 929462
rect 471004 929442 471016 929462
rect 492004 929442 492016 929462
rect 513004 929442 513016 929462
rect 275780 929435 276004 929442
rect 296780 929435 297004 929442
rect 317780 929435 318004 929442
rect 338780 929435 339004 929442
rect 449780 929435 450004 929442
rect 470780 929435 471004 929442
rect 491780 929435 492004 929442
rect 512780 929435 513004 929442
rect 263253 929182 263256 929190
rect 284253 929182 284256 929190
rect 305253 929182 305256 929402
rect 326253 929182 326256 929190
rect 437253 929182 437256 929190
rect 458253 929182 458256 929190
rect 479253 929182 479256 929402
rect 500253 929182 500256 929190
rect 263256 929166 263260 929182
rect 284256 929166 284260 929182
rect 305256 929166 305260 929182
rect 326256 929166 326260 929182
rect 437256 929166 437260 929182
rect 458256 929166 458260 929182
rect 479256 929166 479260 929182
rect 500256 929166 500260 929182
rect 591138 927804 591158 927816
rect 723298 927813 723309 927816
rect 591158 927580 591165 927804
rect 723309 927585 723325 927813
rect 765138 927804 765158 927816
rect 897298 927813 897309 927816
rect 765158 927580 765165 927804
rect 897309 927585 897325 927813
rect 578422 927544 578642 927547
rect 710582 927544 710802 927547
rect 752422 927544 752642 927547
rect 884582 927544 884802 927547
rect 578406 927540 578422 927544
rect 710566 927540 710582 927544
rect 752406 927540 752422 927544
rect 884566 927540 884582 927544
rect 785940 918744 786000 921680
rect 786020 918664 786080 921600
rect 258178 917213 258180 917297
rect 258262 917172 258264 917213
rect 343820 917172 343822 917297
rect 432178 917213 432180 917297
rect 432262 917172 432264 917213
rect 517820 917172 517822 917297
rect 591418 915056 591434 915060
rect 723578 915056 723594 915060
rect 765418 915056 765434 915060
rect 897578 915056 897594 915060
rect 591198 915053 591418 915056
rect 723358 915053 723578 915056
rect 765198 915053 765418 915056
rect 897358 915053 897578 915056
rect 578675 914787 578691 915015
rect 710835 914796 710842 915020
rect 578691 914784 578702 914787
rect 710842 914784 710862 914796
rect 752675 914787 752691 915015
rect 884835 914796 884842 915020
rect 752691 914784 752702 914787
rect 884842 914784 884862 914796
rect 591138 907804 591158 907816
rect 723298 907813 723309 907816
rect 591158 907580 591165 907804
rect 723309 907585 723325 907813
rect 765138 907804 765158 907816
rect 897298 907813 897309 907816
rect 765158 907580 765165 907804
rect 897309 907585 897325 907813
rect 578422 907544 578642 907547
rect 710582 907544 710802 907547
rect 752422 907544 752642 907547
rect 884582 907544 884802 907547
rect 578406 907540 578422 907544
rect 710566 907540 710582 907544
rect 752406 907540 752422 907544
rect 884566 907540 884582 907544
rect 241138 906804 241158 906816
rect 373298 906813 373309 906816
rect 241158 906580 241165 906804
rect 373309 906585 373325 906813
rect 415138 906804 415158 906816
rect 547298 906813 547309 906816
rect 415158 906580 415165 906804
rect 547309 906585 547325 906813
rect 228422 906544 228642 906547
rect 360582 906544 360802 906547
rect 402422 906544 402642 906547
rect 534582 906544 534802 906547
rect 228406 906540 228422 906544
rect 360566 906540 360582 906544
rect 402406 906540 402422 906544
rect 534566 906540 534582 906544
rect 787220 899000 787825 899005
rect 591418 895056 591434 895060
rect 723578 895056 723594 895060
rect 765418 895056 765434 895060
rect 897578 895056 897594 895060
rect 591198 895053 591418 895056
rect 723358 895053 723578 895056
rect 765198 895053 765418 895056
rect 897358 895053 897578 895056
rect 578675 894787 578691 895015
rect 710835 894796 710842 895020
rect 578691 894784 578702 894787
rect 710842 894784 710862 894796
rect 752675 894787 752691 895015
rect 884835 894796 884842 895020
rect 752691 894784 752702 894787
rect 884842 894784 884862 894796
rect 241418 894056 241434 894060
rect 373578 894056 373594 894060
rect 415418 894056 415434 894060
rect 547578 894056 547594 894060
rect 241198 894053 241418 894056
rect 373358 894053 373578 894056
rect 415198 894053 415418 894056
rect 547358 894053 547578 894056
rect 228675 893787 228691 894015
rect 360835 893796 360842 894020
rect 228691 893784 228702 893787
rect 360842 893784 360862 893796
rect 402675 893787 402691 894015
rect 534835 893796 534842 894020
rect 402691 893784 402702 893787
rect 534842 893784 534862 893796
rect 591138 887804 591158 887816
rect 723298 887813 723309 887816
rect 591158 887580 591165 887804
rect 723309 887585 723325 887813
rect 765138 887804 765158 887816
rect 897298 887813 897309 887816
rect 765158 887580 765165 887804
rect 897309 887585 897325 887813
rect 578422 887544 578642 887547
rect 710582 887544 710802 887547
rect 752422 887544 752642 887547
rect 884582 887544 884802 887547
rect 578406 887540 578422 887544
rect 710566 887540 710582 887544
rect 752406 887540 752422 887544
rect 884566 887540 884582 887544
rect 241138 885804 241158 885816
rect 373298 885813 373309 885816
rect 241158 885580 241165 885804
rect 373309 885585 373325 885813
rect 415138 885804 415158 885816
rect 547298 885813 547309 885816
rect 415158 885580 415165 885804
rect 547309 885585 547325 885813
rect 228422 885544 228642 885547
rect 360582 885544 360802 885547
rect 402422 885544 402642 885547
rect 534582 885544 534802 885547
rect 228406 885540 228422 885544
rect 360566 885540 360582 885544
rect 402406 885540 402422 885544
rect 534566 885540 534582 885544
rect 591418 875056 591434 875060
rect 723578 875056 723594 875060
rect 765418 875056 765434 875060
rect 897578 875056 897594 875060
rect 591198 875053 591418 875056
rect 723358 875053 723578 875056
rect 765198 875053 765418 875056
rect 897358 875053 897578 875056
rect 578675 874787 578691 875015
rect 710835 874796 710842 875020
rect 578691 874784 578702 874787
rect 710842 874784 710862 874796
rect 752675 874787 752691 875015
rect 884835 874796 884842 875020
rect 752691 874784 752702 874787
rect 884842 874784 884862 874796
rect 241418 873056 241434 873060
rect 373578 873056 373594 873060
rect 415418 873056 415434 873060
rect 547578 873056 547594 873060
rect 241198 873053 241418 873056
rect 373358 873053 373578 873056
rect 415198 873053 415418 873056
rect 547358 873053 547578 873056
rect 228675 872787 228691 873015
rect 360835 872796 360842 873020
rect 228691 872784 228702 872787
rect 360842 872784 360862 872796
rect 402675 872787 402691 873015
rect 534835 872796 534842 873020
rect 402691 872784 402702 872787
rect 534842 872784 534862 872796
rect 591138 867804 591158 867816
rect 723298 867813 723309 867816
rect 591158 867580 591165 867804
rect 723309 867585 723325 867813
rect 765138 867804 765158 867816
rect 897298 867813 897309 867816
rect 765158 867580 765165 867804
rect 897309 867585 897325 867813
rect 578422 867544 578642 867547
rect 710582 867544 710802 867547
rect 752422 867544 752642 867547
rect 884582 867544 884802 867547
rect 578406 867540 578422 867544
rect 710566 867540 710582 867544
rect 752406 867540 752422 867544
rect 884566 867540 884582 867544
rect 229583 864800 230483 865115
rect 241138 864804 241158 864816
rect 373298 864813 373309 864816
rect 241158 864580 241165 864804
rect 373309 864585 373325 864813
rect 403583 864800 404483 865115
rect 415138 864804 415158 864816
rect 547298 864813 547309 864816
rect 415158 864580 415165 864804
rect 547309 864585 547325 864813
rect 228422 864544 228642 864547
rect 360582 864544 360802 864547
rect 402422 864544 402642 864547
rect 534582 864544 534802 864547
rect 228406 864311 228422 864544
rect 241252 864490 241472 864493
rect 241472 864257 241488 864490
rect 360566 864311 360582 864544
rect 373537 864490 373632 864493
rect 373632 864257 373648 864490
rect 402406 864311 402422 864544
rect 415252 864490 415472 864493
rect 415472 864257 415488 864490
rect 534566 864311 534582 864544
rect 547537 864490 547632 864493
rect 547632 864257 547648 864490
rect 228102 864224 228322 864227
rect 228086 863991 228102 864224
rect 360256 864218 360482 864227
rect 402102 864224 402322 864227
rect 241572 864160 241802 864173
rect 241802 863937 241808 864160
rect 360246 863991 360256 864218
rect 373732 864170 373952 864173
rect 373952 864053 373968 864170
rect 402086 863991 402102 864224
rect 534256 864218 534482 864227
rect 415572 864160 415802 864173
rect 415802 863937 415808 864160
rect 534246 863991 534256 864218
rect 547732 864170 547952 864173
rect 547952 864053 547968 864170
rect 227782 863904 228002 863907
rect 359942 863904 360162 863907
rect 401782 863904 402002 863907
rect 533942 863904 534162 863907
rect 227766 863774 227782 863904
rect 241892 863850 242112 863853
rect 242112 863617 242128 863850
rect 359926 863671 359942 863904
rect 374069 863850 374272 863853
rect 374272 863784 374288 863850
rect 401766 863774 401782 863904
rect 415892 863850 416112 863853
rect 416112 863617 416128 863850
rect 533926 863671 533942 863904
rect 548069 863850 548272 863853
rect 548272 863784 548288 863850
rect 227420 863542 227640 863545
rect 359580 863542 359800 863545
rect 401420 863542 401640 863545
rect 533580 863542 533800 863545
rect 227404 863518 227420 863542
rect 242200 863518 242436 863531
rect 359564 863518 359580 863542
rect 374360 863518 374596 863531
rect 401404 863518 401420 863542
rect 416200 863518 416436 863531
rect 533564 863518 533580 863542
rect 548360 863518 548596 863531
rect 231275 863323 231309 863357
rect 234297 863323 234331 863357
rect 367669 863323 367703 863357
rect 370691 863323 370725 863357
rect 405275 863323 405309 863357
rect 408297 863323 408331 863357
rect 541669 863323 541703 863357
rect 544691 863323 544725 863357
rect 231275 863285 231347 863321
rect 234259 863285 234331 863321
rect 367669 863285 367741 863321
rect 370653 863285 370725 863321
rect 405275 863285 405347 863321
rect 408259 863285 408331 863321
rect 541669 863285 541741 863321
rect 544653 863285 544725 863321
rect 785960 858940 786000 859160
rect 786020 859000 786080 859160
rect 591418 855056 591434 855060
rect 723578 855056 723594 855060
rect 765418 855056 765434 855060
rect 897578 855056 897594 855060
rect 591198 855053 591418 855056
rect 723358 855053 723578 855056
rect 765198 855053 765418 855056
rect 897358 855053 897578 855056
rect 578675 854787 578691 855015
rect 710835 854796 710842 855020
rect 578691 854784 578702 854787
rect 710842 854784 710862 854796
rect 752675 854787 752691 855015
rect 884835 854796 884842 855020
rect 752691 854784 752702 854787
rect 884842 854784 884862 854796
rect 231275 853279 231347 853315
rect 234259 853279 234331 853315
rect 367669 853279 367741 853315
rect 370653 853279 370725 853315
rect 405275 853279 405347 853315
rect 408259 853279 408331 853315
rect 541669 853279 541741 853315
rect 544653 853279 544725 853315
rect 231275 853243 231309 853277
rect 234297 853243 234331 853277
rect 367669 853243 367703 853277
rect 370691 853243 370725 853277
rect 405275 853243 405309 853277
rect 408297 853243 408331 853277
rect 541669 853243 541703 853277
rect 544691 853243 544725 853277
rect 227404 853069 227640 853082
rect 242420 853058 242436 853082
rect 359564 853069 359800 853082
rect 374580 853058 374596 853082
rect 401404 853069 401640 853082
rect 416420 853058 416436 853082
rect 533564 853069 533800 853082
rect 548580 853058 548596 853082
rect 242200 853055 242420 853058
rect 374360 853055 374580 853058
rect 416200 853055 416420 853058
rect 548360 853055 548580 853058
rect 227712 852750 227728 852816
rect 227728 852747 227931 852750
rect 242058 852696 242074 852929
rect 359872 852750 359888 852983
rect 359888 852747 360108 852750
rect 374218 852696 374234 852826
rect 401712 852750 401728 852816
rect 401728 852747 401931 852750
rect 416058 852696 416074 852929
rect 533872 852750 533888 852983
rect 533888 852747 534108 852750
rect 548218 852696 548234 852826
rect 241838 852693 242058 852696
rect 373998 852693 374218 852696
rect 415838 852693 416058 852696
rect 547998 852693 548218 852696
rect 228032 852430 228048 852547
rect 228048 852427 228268 852430
rect 241744 852382 241754 852609
rect 360192 852440 360198 852663
rect 360198 852427 360428 852440
rect 241518 852373 241744 852382
rect 373898 852376 373914 852609
rect 402032 852430 402048 852547
rect 402048 852427 402268 852430
rect 415744 852382 415754 852609
rect 534192 852440 534198 852663
rect 534198 852427 534428 852440
rect 373678 852373 373898 852376
rect 415518 852373 415744 852382
rect 547898 852376 547914 852609
rect 547678 852373 547898 852376
rect 228352 852110 228368 852343
rect 228368 852107 228463 852110
rect 241418 852056 241434 852289
rect 360512 852110 360528 852343
rect 360528 852107 360748 852110
rect 373578 852056 373594 852289
rect 402352 852110 402368 852343
rect 402368 852107 402463 852110
rect 415418 852056 415434 852289
rect 534512 852110 534528 852343
rect 534528 852107 534748 852110
rect 547578 852056 547594 852289
rect 241198 852053 241418 852056
rect 373358 852053 373578 852056
rect 415198 852053 415418 852056
rect 547358 852053 547578 852056
rect 228675 851787 228691 852015
rect 360835 851796 360842 852020
rect 228691 851784 228702 851787
rect 360842 851784 360862 851796
rect 402675 851787 402691 852015
rect 534835 851796 534842 852020
rect 402691 851784 402702 851787
rect 534842 851784 534862 851796
rect 591138 847804 591158 847816
rect 723298 847813 723309 847816
rect 591158 847580 591165 847804
rect 723309 847585 723325 847813
rect 765138 847804 765158 847816
rect 897298 847813 897309 847816
rect 765158 847580 765165 847804
rect 897309 847585 897325 847813
rect 578422 847544 578642 847547
rect 710582 847544 710802 847547
rect 752422 847544 752642 847547
rect 884582 847544 884802 847547
rect 578406 847540 578422 847544
rect 710566 847540 710582 847544
rect 752406 847540 752422 847544
rect 884566 847540 884582 847544
rect 241138 843804 241158 843816
rect 373298 843813 373309 843816
rect 241158 843580 241165 843804
rect 373309 843585 373325 843813
rect 415138 843804 415158 843816
rect 547298 843813 547309 843816
rect 415158 843580 415165 843804
rect 547309 843585 547325 843813
rect 228422 843544 228642 843547
rect 360582 843544 360802 843547
rect 402422 843544 402642 843547
rect 534582 843544 534802 843547
rect 228406 843311 228422 843544
rect 241252 843490 241472 843493
rect 241472 843257 241488 843490
rect 360566 843311 360582 843544
rect 373537 843490 373632 843493
rect 373632 843257 373648 843490
rect 402406 843311 402422 843544
rect 415252 843490 415472 843493
rect 415472 843257 415488 843490
rect 534566 843311 534582 843544
rect 547537 843490 547632 843493
rect 547632 843257 547648 843490
rect 228102 843224 228322 843227
rect 228086 842991 228102 843224
rect 360256 843218 360482 843227
rect 402102 843224 402322 843227
rect 241572 843160 241802 843173
rect 241802 842937 241808 843160
rect 360246 842991 360256 843218
rect 373732 843170 373952 843173
rect 373952 843053 373968 843170
rect 402086 842991 402102 843224
rect 534256 843218 534482 843227
rect 415572 843160 415802 843173
rect 415802 842937 415808 843160
rect 534246 842991 534256 843218
rect 547732 843170 547952 843173
rect 547952 843053 547968 843170
rect 227782 842904 228002 842907
rect 359942 842904 360162 842907
rect 401782 842904 402002 842907
rect 533942 842904 534162 842907
rect 227766 842774 227782 842904
rect 241892 842850 242112 842853
rect 242112 842617 242128 842850
rect 359926 842671 359942 842904
rect 374069 842850 374272 842853
rect 374272 842617 374288 842850
rect 401766 842774 401782 842904
rect 415892 842850 416112 842853
rect 416112 842617 416128 842850
rect 533926 842671 533942 842904
rect 548069 842850 548272 842853
rect 548272 842617 548288 842850
rect 227420 842542 227640 842545
rect 359580 842542 359800 842545
rect 401420 842542 401640 842545
rect 533580 842542 533800 842545
rect 227404 842518 227420 842542
rect 242200 842518 242436 842531
rect 359564 842518 359580 842542
rect 374360 842518 374596 842531
rect 401404 842518 401420 842542
rect 416200 842518 416436 842531
rect 533564 842518 533580 842542
rect 548360 842518 548596 842531
rect 231275 842323 231309 842357
rect 234297 842323 234331 842357
rect 405275 842323 405309 842357
rect 408297 842323 408331 842357
rect 231275 842285 231347 842321
rect 234259 842285 234331 842321
rect 405275 842285 405347 842321
rect 408259 842285 408331 842321
rect 591418 835056 591434 835060
rect 723578 835056 723594 835060
rect 765418 835056 765434 835060
rect 897578 835056 897594 835060
rect 591198 835053 591418 835056
rect 723358 835053 723578 835056
rect 765198 835053 765418 835056
rect 897358 835053 897578 835056
rect 578675 834787 578691 835015
rect 710835 834796 710842 835020
rect 578691 834784 578702 834787
rect 710842 834784 710862 834796
rect 752675 834787 752691 835015
rect 884835 834796 884842 835020
rect 752691 834784 752702 834787
rect 884842 834784 884862 834796
rect 231275 832279 231347 832315
rect 234259 832279 234331 832315
rect 405275 832279 405347 832315
rect 408259 832279 408331 832315
rect 231275 832243 231309 832277
rect 234297 832243 234331 832277
rect 405275 832243 405309 832277
rect 408297 832243 408331 832277
rect 227404 832069 227640 832082
rect 242420 832058 242436 832082
rect 359564 832069 359800 832082
rect 374580 832058 374596 832082
rect 401404 832069 401640 832082
rect 416420 832058 416436 832082
rect 533564 832069 533800 832082
rect 548580 832058 548596 832082
rect 242200 832055 242420 832058
rect 374360 832055 374580 832058
rect 416200 832055 416420 832058
rect 548360 832055 548580 832058
rect 227712 831750 227728 831816
rect 227728 831747 227931 831750
rect 242058 831696 242074 831929
rect 359872 831750 359888 831983
rect 359888 831747 360108 831750
rect 374218 831696 374234 831929
rect 401712 831750 401728 831816
rect 401728 831747 401931 831750
rect 416058 831696 416074 831929
rect 533872 831750 533888 831983
rect 533888 831747 534108 831750
rect 548218 831696 548234 831929
rect 241838 831693 242058 831696
rect 373998 831693 374218 831696
rect 415838 831693 416058 831696
rect 547998 831693 548218 831696
rect 228032 831430 228048 831547
rect 228048 831427 228268 831430
rect 241744 831382 241754 831609
rect 360192 831440 360198 831663
rect 360198 831427 360428 831440
rect 241518 831373 241744 831382
rect 373898 831376 373914 831609
rect 402032 831430 402048 831547
rect 402048 831427 402268 831430
rect 415744 831382 415754 831609
rect 534192 831440 534198 831663
rect 534198 831427 534428 831440
rect 373678 831373 373898 831376
rect 415518 831373 415744 831382
rect 547898 831376 547914 831609
rect 547678 831373 547898 831376
rect 228352 831110 228368 831343
rect 228368 831107 228463 831110
rect 241418 831056 241434 831289
rect 360512 831110 360528 831343
rect 360528 831107 360748 831110
rect 373578 831056 373594 831289
rect 402352 831110 402368 831343
rect 402368 831107 402463 831110
rect 415418 831056 415434 831289
rect 534512 831110 534528 831343
rect 534528 831107 534748 831110
rect 547578 831056 547594 831289
rect 241198 831053 241418 831056
rect 373358 831053 373578 831056
rect 415198 831053 415418 831056
rect 547358 831053 547578 831056
rect 228675 830787 228691 831015
rect 360835 830796 360842 831020
rect 228691 830784 228702 830787
rect 360842 830784 360862 830796
rect 402675 830787 402691 831015
rect 534835 830796 534842 831020
rect 402691 830784 402702 830787
rect 534842 830784 534862 830796
rect 591138 827804 591158 827816
rect 723298 827813 723309 827816
rect 591158 827580 591165 827804
rect 723309 827585 723325 827813
rect 765138 827804 765158 827816
rect 897298 827813 897309 827816
rect 765158 827580 765165 827804
rect 897309 827585 897325 827813
rect 578422 827544 578642 827547
rect 710582 827544 710802 827547
rect 752422 827544 752642 827547
rect 884582 827544 884802 827547
rect 578406 827540 578422 827544
rect 710566 827540 710582 827544
rect 752406 827540 752422 827544
rect 884566 827540 884582 827544
rect 241138 822804 241158 822816
rect 373298 822813 373309 822816
rect 241158 822580 241165 822804
rect 373309 822585 373325 822813
rect 415138 822804 415158 822816
rect 547298 822813 547309 822816
rect 415158 822580 415165 822804
rect 547309 822585 547325 822813
rect 228422 822544 228642 822547
rect 360582 822544 360802 822547
rect 402422 822544 402642 822547
rect 534582 822544 534802 822547
rect 228406 822311 228422 822544
rect 241252 822490 241472 822493
rect 241472 822257 241488 822490
rect 360566 822311 360582 822544
rect 373537 822490 373632 822493
rect 373632 822257 373648 822490
rect 402406 822311 402422 822544
rect 415252 822490 415472 822493
rect 415472 822257 415488 822490
rect 534566 822311 534582 822544
rect 547537 822490 547632 822493
rect 547632 822257 547648 822490
rect 228102 822224 228322 822227
rect 228086 821991 228102 822224
rect 360256 822218 360482 822227
rect 402102 822224 402322 822227
rect 241572 822160 241802 822173
rect 241802 821937 241808 822160
rect 360246 821991 360256 822218
rect 373732 822170 373952 822173
rect 373952 822053 373968 822170
rect 402086 821991 402102 822224
rect 534256 822218 534482 822227
rect 415572 822160 415802 822173
rect 415802 821937 415808 822160
rect 534246 821991 534256 822218
rect 547732 822170 547952 822173
rect 547952 822053 547968 822170
rect 227782 821904 228002 821907
rect 359942 821904 360162 821907
rect 401782 821904 402002 821907
rect 533942 821904 534162 821907
rect 227766 821671 227782 821904
rect 241892 821850 242112 821853
rect 242112 821617 242128 821850
rect 359926 821671 359942 821904
rect 374069 821850 374272 821853
rect 374272 821784 374288 821850
rect 401766 821671 401782 821904
rect 415892 821850 416112 821853
rect 416112 821617 416128 821850
rect 533926 821671 533942 821904
rect 548069 821850 548272 821853
rect 548272 821784 548288 821850
rect 227420 821542 227640 821545
rect 359580 821542 359800 821545
rect 401420 821542 401640 821545
rect 533580 821542 533800 821545
rect 227404 821518 227420 821542
rect 242200 821518 242436 821531
rect 359564 821518 359580 821542
rect 374360 821518 374596 821531
rect 401404 821518 401420 821542
rect 416200 821518 416436 821531
rect 533564 821518 533580 821542
rect 548360 821518 548596 821531
rect 367669 821323 367703 821357
rect 370691 821323 370725 821357
rect 541669 821323 541703 821357
rect 544691 821323 544725 821357
rect 367669 821285 367741 821321
rect 370653 821285 370725 821321
rect 541669 821285 541741 821321
rect 544653 821285 544725 821321
rect 785940 819200 786000 823680
rect 785960 818940 786000 819200
rect 786020 819000 786080 823600
rect 591418 815056 591434 815060
rect 723578 815056 723594 815060
rect 765418 815056 765434 815060
rect 897578 815056 897594 815060
rect 591198 815053 591418 815056
rect 723358 815053 723578 815056
rect 765198 815053 765418 815056
rect 897358 815053 897578 815056
rect 578675 814787 578691 815015
rect 710835 814796 710842 815020
rect 578691 814784 578702 814787
rect 710842 814784 710862 814796
rect 752675 814787 752691 815015
rect 884835 814796 884842 815020
rect 752691 814784 752702 814787
rect 884842 814784 884862 814796
rect 367669 811279 367741 811315
rect 370653 811279 370725 811315
rect 541669 811279 541741 811315
rect 544653 811279 544725 811315
rect 367669 811243 367703 811277
rect 370691 811243 370725 811277
rect 541669 811243 541703 811277
rect 544691 811243 544725 811277
rect 227404 811069 227640 811082
rect 242420 811058 242436 811082
rect 359564 811069 359800 811082
rect 374580 811058 374596 811082
rect 401404 811069 401640 811082
rect 416420 811058 416436 811082
rect 533564 811069 533800 811082
rect 548580 811058 548596 811082
rect 242200 811055 242420 811058
rect 374360 811055 374580 811058
rect 416200 811055 416420 811058
rect 548360 811055 548580 811058
rect 227712 810750 227728 810983
rect 227728 810747 227931 810750
rect 242058 810696 242074 810929
rect 359872 810750 359888 810983
rect 359888 810747 360108 810750
rect 374218 810696 374234 810826
rect 401712 810750 401728 810983
rect 401728 810747 401931 810750
rect 416058 810696 416074 810929
rect 533872 810750 533888 810983
rect 533888 810747 534108 810750
rect 548218 810696 548234 810826
rect 241838 810693 242058 810696
rect 373998 810693 374218 810696
rect 415838 810693 416058 810696
rect 547998 810693 548218 810696
rect 228032 810430 228048 810547
rect 228048 810427 228268 810430
rect 241744 810382 241754 810609
rect 360192 810440 360198 810663
rect 360198 810427 360428 810440
rect 241518 810373 241744 810382
rect 373898 810376 373914 810609
rect 402032 810430 402048 810547
rect 402048 810427 402268 810430
rect 415744 810382 415754 810609
rect 534192 810440 534198 810663
rect 534198 810427 534428 810440
rect 373678 810373 373898 810376
rect 415518 810373 415744 810382
rect 547898 810376 547914 810609
rect 547678 810373 547898 810376
rect 228352 810110 228368 810343
rect 228368 810107 228463 810110
rect 241418 810056 241434 810289
rect 360512 810110 360528 810343
rect 360528 810107 360748 810110
rect 373578 810056 373594 810289
rect 402352 810110 402368 810343
rect 402368 810107 402463 810110
rect 415418 810056 415434 810289
rect 534512 810110 534528 810343
rect 534528 810107 534748 810110
rect 547578 810056 547594 810289
rect 241198 810053 241418 810056
rect 373358 810053 373578 810056
rect 415198 810053 415418 810056
rect 547358 810053 547578 810056
rect 228675 809787 228691 810015
rect 360835 809796 360842 810020
rect 228691 809784 228702 809787
rect 360842 809784 360862 809796
rect 402675 809787 402691 810015
rect 534835 809796 534842 810020
rect 402691 809784 402702 809787
rect 534842 809784 534862 809796
rect 591138 807804 591158 807816
rect 723298 807813 723309 807816
rect 591158 807580 591165 807804
rect 723309 807585 723325 807813
rect 765138 807804 765158 807816
rect 897298 807813 897309 807816
rect 765158 807580 765165 807804
rect 897309 807585 897325 807813
rect 578422 807544 578642 807547
rect 710582 807544 710802 807547
rect 752422 807544 752642 807547
rect 884582 807544 884802 807547
rect 578406 807540 578422 807544
rect 710566 807540 710582 807544
rect 752406 807540 752422 807544
rect 884566 807540 884582 807544
rect 787220 799000 787825 799005
rect 591418 795056 591434 795060
rect 723578 795056 723594 795060
rect 765418 795056 765434 795060
rect 897578 795056 897594 795060
rect 591198 795053 591418 795056
rect 723358 795053 723578 795056
rect 765198 795053 765418 795056
rect 897358 795053 897578 795056
rect 578675 794787 578691 795015
rect 710835 794796 710842 795020
rect 578691 794784 578702 794787
rect 710842 794784 710862 794796
rect 752675 794787 752691 795015
rect 884835 794796 884842 795020
rect 752691 794784 752702 794787
rect 884842 794784 884862 794796
rect 591138 787804 591158 787816
rect 723298 787813 723309 787816
rect 591158 787580 591165 787804
rect 723309 787585 723325 787813
rect 765138 787804 765158 787816
rect 897298 787813 897309 787816
rect 765158 787580 765165 787804
rect 897309 787585 897325 787813
rect 578422 787544 578642 787547
rect 710582 787544 710802 787547
rect 752422 787544 752642 787547
rect 884582 787544 884802 787547
rect 578406 787540 578422 787544
rect 710566 787540 710582 787544
rect 752406 787540 752422 787544
rect 884566 787540 884582 787544
rect 275740 787418 275744 787434
rect 296740 787418 296744 787434
rect 317540 787418 317744 787434
rect 338740 787418 338744 787434
rect 449740 787418 449744 787434
rect 470740 787418 470744 787434
rect 491540 787418 491744 787434
rect 512740 787418 512744 787434
rect 275744 787410 275747 787418
rect 296744 787410 296747 787418
rect 317744 787198 317747 787418
rect 338744 787410 338747 787418
rect 449744 787410 449747 787418
rect 470744 787410 470747 787418
rect 491744 787198 491747 787418
rect 512744 787410 512747 787418
rect 262996 787158 263220 787165
rect 283996 787158 284220 787165
rect 304996 787158 305220 787165
rect 325996 787158 326220 787165
rect 436996 787158 437220 787165
rect 457996 787158 458220 787165
rect 478996 787158 479220 787165
rect 499996 787158 500220 787165
rect 262984 787138 262996 787158
rect 283984 787138 283996 787158
rect 304984 787138 304996 787158
rect 325984 787138 325996 787158
rect 436984 787138 436996 787158
rect 457984 787138 457996 787158
rect 478984 787138 478996 787158
rect 499984 787138 499996 787158
rect 591418 775056 591434 775060
rect 723578 775056 723594 775060
rect 765418 775056 765434 775060
rect 897578 775056 897594 775060
rect 591198 775053 591418 775056
rect 723358 775053 723578 775056
rect 765198 775053 765418 775056
rect 897358 775053 897578 775056
rect 578675 774787 578691 775015
rect 710835 774796 710842 775020
rect 578691 774784 578702 774787
rect 710842 774784 710862 774796
rect 752675 774787 752691 775015
rect 884835 774796 884842 775020
rect 752691 774784 752702 774787
rect 884842 774784 884862 774796
rect 276013 774691 276016 774702
rect 297013 774691 297016 774702
rect 318013 774691 318016 774702
rect 339013 774691 339016 774702
rect 450013 774691 450016 774702
rect 471013 774691 471016 774702
rect 492013 774691 492016 774702
rect 513013 774691 513016 774702
rect 275785 774675 276013 774691
rect 296785 774675 297013 774691
rect 317785 774675 318013 774691
rect 338785 774675 339013 774691
rect 449785 774675 450013 774691
rect 470785 774675 471013 774691
rect 491785 774675 492013 774691
rect 512785 774675 513013 774691
rect 263253 774422 263256 774642
rect 284253 774422 284256 774463
rect 305253 774422 305256 774642
rect 263256 774406 263260 774422
rect 284256 774420 284258 774422
rect 284258 774406 284260 774420
rect 305256 774406 305260 774422
rect 317690 774368 317693 774463
rect 326253 774422 326256 774642
rect 437253 774422 437256 774642
rect 458253 774422 458256 774463
rect 479253 774422 479256 774642
rect 326256 774406 326260 774422
rect 437256 774406 437260 774422
rect 458256 774420 458258 774422
rect 458258 774406 458260 774420
rect 479256 774406 479260 774422
rect 491690 774368 491693 774463
rect 500253 774422 500256 774642
rect 500256 774406 500260 774422
rect 317540 774352 317690 774368
rect 491540 774352 491690 774368
rect 591138 767804 591158 767816
rect 723298 767813 723309 767816
rect 591158 767580 591165 767804
rect 723309 767585 723325 767813
rect 765138 767804 765158 767816
rect 897298 767813 897309 767816
rect 765158 767580 765165 767804
rect 897309 767585 897325 767813
rect 578422 767544 578642 767547
rect 710582 767544 710802 767547
rect 752422 767544 752642 767547
rect 884582 767544 884802 767547
rect 578406 767540 578422 767544
rect 710566 767540 710582 767544
rect 752406 767540 752422 767544
rect 884566 767540 884582 767544
rect 785960 758940 786000 759160
rect 786020 759000 786080 759160
rect 591418 755056 591434 755060
rect 723578 755056 723594 755060
rect 765418 755056 765434 755060
rect 897578 755056 897594 755060
rect 591198 755053 591418 755056
rect 723358 755053 723578 755056
rect 765198 755053 765418 755056
rect 897358 755053 897578 755056
rect 578675 754787 578691 755015
rect 710835 754796 710842 755020
rect 578691 754784 578702 754787
rect 710842 754784 710862 754796
rect 752675 754787 752691 755015
rect 884835 754796 884842 755020
rect 752691 754784 752702 754787
rect 884842 754784 884862 754796
rect 591138 747804 591158 747816
rect 723298 747813 723309 747816
rect 591158 747580 591165 747804
rect 723309 747585 723325 747813
rect 765138 747804 765158 747816
rect 897298 747813 897309 747816
rect 765158 747580 765165 747804
rect 897309 747585 897325 747813
rect 578422 747544 578642 747547
rect 710582 747544 710802 747547
rect 752422 747544 752642 747547
rect 884582 747544 884802 747547
rect 578406 747540 578422 747544
rect 710566 747540 710582 747544
rect 752406 747540 752422 747544
rect 884566 747540 884582 747544
rect 275740 742178 275744 742194
rect 296740 742178 296744 742194
rect 317740 742178 317744 742194
rect 338740 742178 338744 742194
rect 449740 742178 449744 742194
rect 470740 742178 470744 742194
rect 491740 742178 491744 742194
rect 512740 742178 512744 742194
rect 275744 741958 275747 742178
rect 296744 741958 296747 742178
rect 317744 741958 317747 742178
rect 338744 741958 338747 742178
rect 449744 741958 449747 742178
rect 470744 741958 470747 742178
rect 491744 741958 491747 742178
rect 512744 741958 512747 742178
rect 262987 741909 263215 741925
rect 283987 741909 284215 741925
rect 304987 741909 305215 741925
rect 325987 741909 326215 741925
rect 436987 741909 437215 741925
rect 457987 741909 458215 741925
rect 478987 741909 479215 741925
rect 499987 741909 500215 741925
rect 262984 741898 262987 741909
rect 283984 741898 283987 741909
rect 304984 741898 304987 741909
rect 325984 741898 325987 741909
rect 436984 741898 436987 741909
rect 457984 741898 457987 741909
rect 478984 741898 478987 741909
rect 499984 741898 499987 741909
rect 591418 735056 591434 735060
rect 723578 735056 723594 735060
rect 765418 735056 765434 735060
rect 897578 735056 897594 735060
rect 591198 735053 591418 735056
rect 723358 735053 723578 735056
rect 765198 735053 765418 735056
rect 897358 735053 897578 735056
rect 578675 734787 578691 735015
rect 710835 734796 710842 735020
rect 578691 734784 578702 734787
rect 710842 734784 710862 734796
rect 752675 734787 752691 735015
rect 884835 734796 884842 735020
rect 752691 734784 752702 734787
rect 884842 734784 884862 734796
rect 276004 729442 276016 729462
rect 297004 729442 297016 729462
rect 318004 729442 318016 729462
rect 339004 729442 339016 729462
rect 450004 729442 450016 729462
rect 471004 729442 471016 729462
rect 492004 729442 492016 729462
rect 513004 729442 513016 729462
rect 275780 729435 276004 729442
rect 296780 729435 297004 729442
rect 317780 729435 318004 729442
rect 338780 729435 339004 729442
rect 449780 729435 450004 729442
rect 470780 729435 471004 729442
rect 491780 729435 492004 729442
rect 512780 729435 513004 729442
rect 263253 729182 263256 729190
rect 284253 729182 284256 729190
rect 305253 729182 305256 729402
rect 326253 729182 326256 729190
rect 437253 729182 437256 729190
rect 458253 729182 458256 729190
rect 479253 729182 479256 729402
rect 500253 729182 500256 729190
rect 263256 729166 263260 729182
rect 284256 729166 284260 729182
rect 305256 729166 305260 729182
rect 326256 729166 326260 729182
rect 437256 729166 437260 729182
rect 458256 729166 458260 729182
rect 479256 729166 479260 729182
rect 500256 729166 500260 729182
rect 591138 727804 591158 727816
rect 723298 727813 723309 727816
rect 591158 727580 591165 727804
rect 723309 727585 723325 727813
rect 765138 727804 765158 727816
rect 897298 727813 897309 727816
rect 765158 727580 765165 727804
rect 897309 727585 897325 727813
rect 578422 727544 578642 727547
rect 710582 727544 710802 727547
rect 752422 727544 752642 727547
rect 884582 727544 884802 727547
rect 578406 727540 578422 727544
rect 710566 727540 710582 727544
rect 752406 727540 752422 727544
rect 884566 727540 884582 727544
rect 785940 719200 786000 723680
rect 785960 718940 786000 719200
rect 786020 719000 786080 723600
rect 258178 717213 258180 717297
rect 258262 717172 258264 717213
rect 343820 717172 343822 717297
rect 432178 717213 432180 717297
rect 432262 717172 432264 717213
rect 517820 717172 517822 717297
rect 591418 715056 591434 715060
rect 723578 715056 723594 715060
rect 765418 715056 765434 715060
rect 897578 715056 897594 715060
rect 591198 715053 591418 715056
rect 723358 715053 723578 715056
rect 765198 715053 765418 715056
rect 897358 715053 897578 715056
rect 578675 714787 578691 715015
rect 710835 714796 710842 715020
rect 578691 714784 578702 714787
rect 710842 714784 710862 714796
rect 752675 714787 752691 715015
rect 884835 714796 884842 715020
rect 752691 714784 752702 714787
rect 884842 714784 884862 714796
rect 591138 707804 591158 707816
rect 723298 707813 723309 707816
rect 591158 707580 591165 707804
rect 723309 707585 723325 707813
rect 765138 707804 765158 707816
rect 897298 707813 897309 707816
rect 765158 707580 765165 707804
rect 897309 707585 897325 707813
rect 578422 707544 578642 707547
rect 710582 707544 710802 707547
rect 752422 707544 752642 707547
rect 884582 707544 884802 707547
rect 578406 707540 578422 707544
rect 710566 707540 710582 707544
rect 752406 707540 752422 707544
rect 884566 707540 884582 707544
rect 241138 706804 241158 706816
rect 373298 706813 373309 706816
rect 241158 706580 241165 706804
rect 373309 706585 373325 706813
rect 415138 706804 415158 706816
rect 547298 706813 547309 706816
rect 415158 706580 415165 706804
rect 547309 706585 547325 706813
rect 228422 706544 228642 706547
rect 360582 706544 360802 706547
rect 402422 706544 402642 706547
rect 534582 706544 534802 706547
rect 228406 706540 228422 706544
rect 360566 706540 360582 706544
rect 402406 706540 402422 706544
rect 534566 706540 534582 706544
rect 787220 699000 787825 699005
rect 591418 695056 591434 695060
rect 723578 695056 723594 695060
rect 765418 695056 765434 695060
rect 897578 695056 897594 695060
rect 591198 695053 591418 695056
rect 723358 695053 723578 695056
rect 765198 695053 765418 695056
rect 897358 695053 897578 695056
rect 578675 694787 578691 695015
rect 710835 694796 710842 695020
rect 578691 694784 578702 694787
rect 710842 694784 710862 694796
rect 752675 694787 752691 695015
rect 884835 694796 884842 695020
rect 752691 694784 752702 694787
rect 884842 694784 884862 694796
rect 241418 694056 241434 694060
rect 373578 694056 373594 694060
rect 415418 694056 415434 694060
rect 547578 694056 547594 694060
rect 241198 694053 241418 694056
rect 373358 694053 373578 694056
rect 415198 694053 415418 694056
rect 547358 694053 547578 694056
rect 228675 693787 228691 694015
rect 360835 693796 360842 694020
rect 228691 693784 228702 693787
rect 360842 693784 360862 693796
rect 402675 693787 402691 694015
rect 534835 693796 534842 694020
rect 402691 693784 402702 693787
rect 534842 693784 534862 693796
rect 591138 687804 591158 687816
rect 723298 687813 723309 687816
rect 591158 687580 591165 687804
rect 723309 687585 723325 687813
rect 765138 687804 765158 687816
rect 897298 687813 897309 687816
rect 765158 687580 765165 687804
rect 897309 687585 897325 687813
rect 578422 687544 578642 687547
rect 710582 687544 710802 687547
rect 752422 687544 752642 687547
rect 884582 687544 884802 687547
rect 578406 687540 578422 687544
rect 710566 687540 710582 687544
rect 752406 687540 752422 687544
rect 884566 687540 884582 687544
rect 241138 685804 241158 685816
rect 373298 685813 373309 685816
rect 241158 685580 241165 685804
rect 373309 685585 373325 685813
rect 415138 685804 415158 685816
rect 547298 685813 547309 685816
rect 415158 685580 415165 685804
rect 547309 685585 547325 685813
rect 228422 685544 228642 685547
rect 360582 685544 360802 685547
rect 402422 685544 402642 685547
rect 534582 685544 534802 685547
rect 228406 685540 228422 685544
rect 360566 685540 360582 685544
rect 402406 685540 402422 685544
rect 534566 685540 534582 685544
rect 591418 675056 591434 675060
rect 723578 675056 723594 675060
rect 765418 675056 765434 675060
rect 897578 675056 897594 675060
rect 591198 675053 591418 675056
rect 723358 675053 723578 675056
rect 765198 675053 765418 675056
rect 897358 675053 897578 675056
rect 578675 674787 578691 675015
rect 710835 674796 710842 675020
rect 578691 674784 578702 674787
rect 710842 674784 710862 674796
rect 752675 674787 752691 675015
rect 884835 674796 884842 675020
rect 752691 674784 752702 674787
rect 884842 674784 884862 674796
rect 241418 673056 241434 673060
rect 373578 673056 373594 673060
rect 415418 673056 415434 673060
rect 547578 673056 547594 673060
rect 241198 673053 241418 673056
rect 373358 673053 373578 673056
rect 415198 673053 415418 673056
rect 547358 673053 547578 673056
rect 228675 672787 228691 673015
rect 360835 672796 360842 673020
rect 228691 672784 228702 672787
rect 360842 672784 360862 672796
rect 402675 672787 402691 673015
rect 534835 672796 534842 673020
rect 402691 672784 402702 672787
rect 534842 672784 534862 672796
rect 591138 667804 591158 667816
rect 723298 667813 723309 667816
rect 591158 667580 591165 667804
rect 723309 667585 723325 667813
rect 765138 667804 765158 667816
rect 897298 667813 897309 667816
rect 765158 667580 765165 667804
rect 897309 667585 897325 667813
rect 578422 667544 578642 667547
rect 710582 667544 710802 667547
rect 752422 667544 752642 667547
rect 884582 667544 884802 667547
rect 578406 667540 578422 667544
rect 710566 667540 710582 667544
rect 752406 667540 752422 667544
rect 884566 667540 884582 667544
rect 229583 664800 230483 665115
rect 241138 664804 241158 664816
rect 373298 664813 373309 664816
rect 241158 664580 241165 664804
rect 373309 664585 373325 664813
rect 403583 664800 404483 665115
rect 415138 664804 415158 664816
rect 547298 664813 547309 664816
rect 415158 664580 415165 664804
rect 547309 664585 547325 664813
rect 228422 664544 228642 664547
rect 360582 664544 360802 664547
rect 402422 664544 402642 664547
rect 534582 664544 534802 664547
rect 228406 664311 228422 664544
rect 241252 664490 241472 664493
rect 241472 664257 241488 664490
rect 360566 664311 360582 664544
rect 373537 664490 373632 664493
rect 373632 664257 373648 664490
rect 402406 664311 402422 664544
rect 415252 664490 415472 664493
rect 415472 664257 415488 664490
rect 534566 664311 534582 664544
rect 547537 664490 547632 664493
rect 547632 664257 547648 664490
rect 228102 664224 228322 664227
rect 228086 663991 228102 664224
rect 360256 664218 360482 664227
rect 402102 664224 402322 664227
rect 241572 664160 241802 664173
rect 241802 663937 241808 664160
rect 360246 663991 360256 664218
rect 373732 664170 373952 664173
rect 373952 664053 373968 664170
rect 402086 663991 402102 664224
rect 534256 664218 534482 664227
rect 415572 664160 415802 664173
rect 415802 663937 415808 664160
rect 534246 663991 534256 664218
rect 547732 664170 547952 664173
rect 547952 664053 547968 664170
rect 227782 663904 228002 663907
rect 359942 663904 360162 663907
rect 401782 663904 402002 663907
rect 533942 663904 534162 663907
rect 227766 663774 227782 663904
rect 241892 663850 242112 663853
rect 242112 663617 242128 663850
rect 359926 663671 359942 663904
rect 374069 663850 374272 663853
rect 374272 663784 374288 663850
rect 401766 663774 401782 663904
rect 415892 663850 416112 663853
rect 416112 663617 416128 663850
rect 533926 663671 533942 663904
rect 548069 663850 548272 663853
rect 548272 663784 548288 663850
rect 227420 663542 227640 663545
rect 359580 663542 359800 663545
rect 401420 663542 401640 663545
rect 533580 663542 533800 663545
rect 227404 663518 227420 663542
rect 242200 663518 242436 663531
rect 359564 663518 359580 663542
rect 374360 663518 374596 663531
rect 401404 663518 401420 663542
rect 416200 663518 416436 663531
rect 533564 663518 533580 663542
rect 548360 663518 548596 663531
rect 231275 663323 231309 663357
rect 234297 663323 234331 663357
rect 367669 663323 367703 663357
rect 370691 663323 370725 663357
rect 405275 663323 405309 663357
rect 408297 663323 408331 663357
rect 541669 663323 541703 663357
rect 544691 663323 544725 663357
rect 231275 663285 231347 663321
rect 234259 663285 234331 663321
rect 367669 663285 367741 663321
rect 370653 663285 370725 663321
rect 405275 663285 405347 663321
rect 408259 663285 408331 663321
rect 541669 663285 541741 663321
rect 544653 663285 544725 663321
rect 785960 658940 786000 659160
rect 786020 659000 786080 659160
rect 591418 655056 591434 655060
rect 723578 655056 723594 655060
rect 765418 655056 765434 655060
rect 897578 655056 897594 655060
rect 591198 655053 591418 655056
rect 723358 655053 723578 655056
rect 765198 655053 765418 655056
rect 897358 655053 897578 655056
rect 578675 654787 578691 655015
rect 710835 654796 710842 655020
rect 578691 654784 578702 654787
rect 710842 654784 710862 654796
rect 752675 654787 752691 655015
rect 884835 654796 884842 655020
rect 752691 654784 752702 654787
rect 884842 654784 884862 654796
rect 231275 653279 231347 653315
rect 234259 653279 234331 653315
rect 367669 653279 367741 653315
rect 370653 653279 370725 653315
rect 405275 653279 405347 653315
rect 408259 653279 408331 653315
rect 541669 653279 541741 653315
rect 544653 653279 544725 653315
rect 231275 653243 231309 653277
rect 234297 653243 234331 653277
rect 367669 653243 367703 653277
rect 370691 653243 370725 653277
rect 405275 653243 405309 653277
rect 408297 653243 408331 653277
rect 541669 653243 541703 653277
rect 544691 653243 544725 653277
rect 227404 653069 227640 653082
rect 242420 653058 242436 653082
rect 359564 653069 359800 653082
rect 374580 653058 374596 653082
rect 401404 653069 401640 653082
rect 416420 653058 416436 653082
rect 533564 653069 533800 653082
rect 548580 653058 548596 653082
rect 242200 653055 242420 653058
rect 374360 653055 374580 653058
rect 416200 653055 416420 653058
rect 548360 653055 548580 653058
rect 227712 652750 227728 652816
rect 227728 652747 227931 652750
rect 242058 652696 242074 652929
rect 359872 652750 359888 652983
rect 359888 652747 360108 652750
rect 374218 652696 374234 652826
rect 401712 652750 401728 652816
rect 401728 652747 401931 652750
rect 416058 652696 416074 652929
rect 533872 652750 533888 652983
rect 533888 652747 534108 652750
rect 548218 652696 548234 652826
rect 241838 652693 242058 652696
rect 373998 652693 374218 652696
rect 415838 652693 416058 652696
rect 547998 652693 548218 652696
rect 228032 652430 228048 652547
rect 228048 652427 228268 652430
rect 241744 652382 241754 652609
rect 360192 652440 360198 652663
rect 360198 652427 360428 652440
rect 241518 652373 241744 652382
rect 373898 652376 373914 652609
rect 402032 652430 402048 652547
rect 402048 652427 402268 652430
rect 415744 652382 415754 652609
rect 534192 652440 534198 652663
rect 534198 652427 534428 652440
rect 373678 652373 373898 652376
rect 415518 652373 415744 652382
rect 547898 652376 547914 652609
rect 547678 652373 547898 652376
rect 228352 652110 228368 652343
rect 228368 652107 228463 652110
rect 241418 652056 241434 652289
rect 360512 652110 360528 652343
rect 360528 652107 360748 652110
rect 373578 652056 373594 652289
rect 402352 652110 402368 652343
rect 402368 652107 402463 652110
rect 415418 652056 415434 652289
rect 534512 652110 534528 652343
rect 534528 652107 534748 652110
rect 547578 652056 547594 652289
rect 241198 652053 241418 652056
rect 373358 652053 373578 652056
rect 415198 652053 415418 652056
rect 547358 652053 547578 652056
rect 228675 651787 228691 652015
rect 360835 651796 360842 652020
rect 228691 651784 228702 651787
rect 360842 651784 360862 651796
rect 402675 651787 402691 652015
rect 534835 651796 534842 652020
rect 402691 651784 402702 651787
rect 534842 651784 534862 651796
rect 591138 647804 591158 647816
rect 723298 647813 723309 647816
rect 591158 647580 591165 647804
rect 723309 647585 723325 647813
rect 765138 647804 765158 647816
rect 897298 647813 897309 647816
rect 765158 647580 765165 647804
rect 897309 647585 897325 647813
rect 578422 647544 578642 647547
rect 710582 647544 710802 647547
rect 752422 647544 752642 647547
rect 884582 647544 884802 647547
rect 578406 647540 578422 647544
rect 710566 647540 710582 647544
rect 752406 647540 752422 647544
rect 884566 647540 884582 647544
rect 241138 643804 241158 643816
rect 373298 643813 373309 643816
rect 241158 643580 241165 643804
rect 373309 643585 373325 643813
rect 415138 643804 415158 643816
rect 547298 643813 547309 643816
rect 415158 643580 415165 643804
rect 547309 643585 547325 643813
rect 228422 643544 228642 643547
rect 360582 643544 360802 643547
rect 402422 643544 402642 643547
rect 534582 643544 534802 643547
rect 228406 643311 228422 643544
rect 241252 643490 241472 643493
rect 241472 643257 241488 643490
rect 360566 643311 360582 643544
rect 373537 643490 373632 643493
rect 373632 643257 373648 643490
rect 402406 643311 402422 643544
rect 415252 643490 415472 643493
rect 415472 643257 415488 643490
rect 534566 643311 534582 643544
rect 547537 643490 547632 643493
rect 547632 643257 547648 643490
rect 228102 643224 228322 643227
rect 228086 642991 228102 643224
rect 360256 643218 360482 643227
rect 402102 643224 402322 643227
rect 241572 643160 241802 643173
rect 241802 642937 241808 643160
rect 360246 642991 360256 643218
rect 373732 643170 373952 643173
rect 373952 643053 373968 643170
rect 402086 642991 402102 643224
rect 534256 643218 534482 643227
rect 415572 643160 415802 643173
rect 415802 642937 415808 643160
rect 534246 642991 534256 643218
rect 547732 643170 547952 643173
rect 547952 643053 547968 643170
rect 227782 642904 228002 642907
rect 359942 642904 360162 642907
rect 401782 642904 402002 642907
rect 533942 642904 534162 642907
rect 227766 642774 227782 642904
rect 241892 642850 242112 642853
rect 242112 642617 242128 642850
rect 359926 642671 359942 642904
rect 374069 642850 374272 642853
rect 374272 642617 374288 642850
rect 401766 642774 401782 642904
rect 415892 642850 416112 642853
rect 416112 642617 416128 642850
rect 533926 642671 533942 642904
rect 548069 642850 548272 642853
rect 548272 642617 548288 642850
rect 227420 642542 227640 642545
rect 359580 642542 359800 642545
rect 401420 642542 401640 642545
rect 533580 642542 533800 642545
rect 227404 642518 227420 642542
rect 242200 642518 242436 642531
rect 359564 642518 359580 642542
rect 374360 642518 374596 642531
rect 401404 642518 401420 642542
rect 416200 642518 416436 642531
rect 533564 642518 533580 642542
rect 548360 642518 548596 642531
rect 231275 642323 231309 642357
rect 234297 642323 234331 642357
rect 405275 642323 405309 642357
rect 408297 642323 408331 642357
rect 231275 642285 231347 642321
rect 234259 642285 234331 642321
rect 405275 642285 405347 642321
rect 408259 642285 408331 642321
rect 591418 635056 591434 635060
rect 723578 635056 723594 635060
rect 765418 635056 765434 635060
rect 897578 635056 897594 635060
rect 591198 635053 591418 635056
rect 723358 635053 723578 635056
rect 765198 635053 765418 635056
rect 897358 635053 897578 635056
rect 578675 634787 578691 635015
rect 710835 634796 710842 635020
rect 578691 634784 578702 634787
rect 710842 634784 710862 634796
rect 752675 634787 752691 635015
rect 884835 634796 884842 635020
rect 752691 634784 752702 634787
rect 884842 634784 884862 634796
rect 231275 632279 231347 632315
rect 234259 632279 234331 632315
rect 405275 632279 405347 632315
rect 408259 632279 408331 632315
rect 231275 632243 231309 632277
rect 234297 632243 234331 632277
rect 405275 632243 405309 632277
rect 408297 632243 408331 632277
rect 227404 632069 227640 632082
rect 242420 632058 242436 632082
rect 359564 632069 359800 632082
rect 374580 632058 374596 632082
rect 401404 632069 401640 632082
rect 416420 632058 416436 632082
rect 533564 632069 533800 632082
rect 548580 632058 548596 632082
rect 242200 632055 242420 632058
rect 374360 632055 374580 632058
rect 416200 632055 416420 632058
rect 548360 632055 548580 632058
rect 227712 631750 227728 631816
rect 227728 631747 227931 631750
rect 242058 631696 242074 631929
rect 359872 631750 359888 631983
rect 359888 631747 360108 631750
rect 374218 631696 374234 631929
rect 401712 631750 401728 631816
rect 401728 631747 401931 631750
rect 416058 631696 416074 631929
rect 533872 631750 533888 631983
rect 533888 631747 534108 631750
rect 548218 631696 548234 631929
rect 241838 631693 242058 631696
rect 373998 631693 374218 631696
rect 415838 631693 416058 631696
rect 547998 631693 548218 631696
rect 228032 631430 228048 631547
rect 228048 631427 228268 631430
rect 241744 631382 241754 631609
rect 360192 631440 360198 631663
rect 360198 631427 360428 631440
rect 241518 631373 241744 631382
rect 373898 631376 373914 631609
rect 402032 631430 402048 631547
rect 402048 631427 402268 631430
rect 415744 631382 415754 631609
rect 534192 631440 534198 631663
rect 534198 631427 534428 631440
rect 373678 631373 373898 631376
rect 415518 631373 415744 631382
rect 547898 631376 547914 631609
rect 547678 631373 547898 631376
rect 228352 631110 228368 631343
rect 228368 631107 228463 631110
rect 241418 631056 241434 631289
rect 360512 631110 360528 631343
rect 360528 631107 360748 631110
rect 373578 631056 373594 631289
rect 402352 631110 402368 631343
rect 402368 631107 402463 631110
rect 415418 631056 415434 631289
rect 534512 631110 534528 631343
rect 534528 631107 534748 631110
rect 547578 631056 547594 631289
rect 241198 631053 241418 631056
rect 373358 631053 373578 631056
rect 415198 631053 415418 631056
rect 547358 631053 547578 631056
rect 228675 630787 228691 631015
rect 360835 630796 360842 631020
rect 228691 630784 228702 630787
rect 360842 630784 360862 630796
rect 402675 630787 402691 631015
rect 534835 630796 534842 631020
rect 402691 630784 402702 630787
rect 534842 630784 534862 630796
rect 591138 627804 591158 627816
rect 723298 627813 723309 627816
rect 591158 627580 591165 627804
rect 723309 627585 723325 627813
rect 765138 627804 765158 627816
rect 897298 627813 897309 627816
rect 765158 627580 765165 627804
rect 897309 627585 897325 627813
rect 578422 627544 578642 627547
rect 710582 627544 710802 627547
rect 752422 627544 752642 627547
rect 884582 627544 884802 627547
rect 578406 627540 578422 627544
rect 710566 627540 710582 627544
rect 752406 627540 752422 627544
rect 884566 627540 884582 627544
rect 241138 622804 241158 622816
rect 373298 622813 373309 622816
rect 241158 622580 241165 622804
rect 373309 622585 373325 622813
rect 415138 622804 415158 622816
rect 547298 622813 547309 622816
rect 415158 622580 415165 622804
rect 547309 622585 547325 622813
rect 228422 622544 228642 622547
rect 360582 622544 360802 622547
rect 402422 622544 402642 622547
rect 534582 622544 534802 622547
rect 228406 622311 228422 622544
rect 241252 622490 241472 622493
rect 241472 622257 241488 622490
rect 360566 622311 360582 622544
rect 373537 622490 373632 622493
rect 373632 622257 373648 622490
rect 402406 622311 402422 622544
rect 415252 622490 415472 622493
rect 415472 622257 415488 622490
rect 534566 622311 534582 622544
rect 547537 622490 547632 622493
rect 547632 622257 547648 622490
rect 228102 622224 228322 622227
rect 228086 621991 228102 622224
rect 360256 622218 360482 622227
rect 402102 622224 402322 622227
rect 241572 622160 241802 622173
rect 241802 621937 241808 622160
rect 360246 621991 360256 622218
rect 373732 622170 373952 622173
rect 373952 622053 373968 622170
rect 402086 621991 402102 622224
rect 534256 622218 534482 622227
rect 415572 622160 415802 622173
rect 415802 621937 415808 622160
rect 534246 621991 534256 622218
rect 547732 622170 547952 622173
rect 547952 622053 547968 622170
rect 227782 621904 228002 621907
rect 359942 621904 360162 621907
rect 401782 621904 402002 621907
rect 533942 621904 534162 621907
rect 227766 621671 227782 621904
rect 241892 621850 242112 621853
rect 242112 621617 242128 621850
rect 359926 621671 359942 621904
rect 374069 621850 374272 621853
rect 374272 621784 374288 621850
rect 401766 621671 401782 621904
rect 415892 621850 416112 621853
rect 416112 621617 416128 621850
rect 533926 621671 533942 621904
rect 548069 621850 548272 621853
rect 548272 621784 548288 621850
rect 227420 621542 227640 621545
rect 359580 621542 359800 621545
rect 401420 621542 401640 621545
rect 533580 621542 533800 621545
rect 227404 621518 227420 621542
rect 242200 621518 242436 621531
rect 359564 621518 359580 621542
rect 374360 621518 374596 621531
rect 401404 621518 401420 621542
rect 416200 621518 416436 621531
rect 533564 621518 533580 621542
rect 548360 621518 548596 621531
rect 367669 621323 367703 621357
rect 370691 621323 370725 621357
rect 541669 621323 541703 621357
rect 544691 621323 544725 621357
rect 367669 621285 367741 621321
rect 370653 621285 370725 621321
rect 541669 621285 541741 621321
rect 544653 621285 544725 621321
rect 785940 619200 786000 623680
rect 785960 618940 786000 619200
rect 786020 619000 786080 623600
rect 591418 615056 591434 615060
rect 723578 615056 723594 615060
rect 765418 615056 765434 615060
rect 897578 615056 897594 615060
rect 591198 615053 591418 615056
rect 723358 615053 723578 615056
rect 765198 615053 765418 615056
rect 897358 615053 897578 615056
rect 578675 614787 578691 615015
rect 710835 614796 710842 615020
rect 578691 614784 578702 614787
rect 710842 614784 710862 614796
rect 752675 614787 752691 615015
rect 884835 614796 884842 615020
rect 752691 614784 752702 614787
rect 884842 614784 884862 614796
rect 367669 611279 367741 611315
rect 370653 611279 370725 611315
rect 541669 611279 541741 611315
rect 544653 611279 544725 611315
rect 367669 611243 367703 611277
rect 370691 611243 370725 611277
rect 541669 611243 541703 611277
rect 544691 611243 544725 611277
rect 227404 611069 227640 611082
rect 242420 611058 242436 611082
rect 359564 611069 359800 611082
rect 374580 611058 374596 611082
rect 401404 611069 401640 611082
rect 416420 611058 416436 611082
rect 533564 611069 533800 611082
rect 548580 611058 548596 611082
rect 242200 611055 242420 611058
rect 374360 611055 374580 611058
rect 416200 611055 416420 611058
rect 548360 611055 548580 611058
rect 227712 610750 227728 610983
rect 227728 610747 227931 610750
rect 242058 610696 242074 610929
rect 359872 610750 359888 610983
rect 359888 610747 360108 610750
rect 374218 610696 374234 610826
rect 401712 610750 401728 610983
rect 401728 610747 401931 610750
rect 416058 610696 416074 610929
rect 533872 610750 533888 610983
rect 533888 610747 534108 610750
rect 548218 610696 548234 610826
rect 241838 610693 242058 610696
rect 373998 610693 374218 610696
rect 415838 610693 416058 610696
rect 547998 610693 548218 610696
rect 228032 610430 228048 610547
rect 228048 610427 228268 610430
rect 241744 610382 241754 610609
rect 360192 610440 360198 610663
rect 360198 610427 360428 610440
rect 241518 610373 241744 610382
rect 373898 610376 373914 610609
rect 402032 610430 402048 610547
rect 402048 610427 402268 610430
rect 415744 610382 415754 610609
rect 534192 610440 534198 610663
rect 534198 610427 534428 610440
rect 373678 610373 373898 610376
rect 415518 610373 415744 610382
rect 547898 610376 547914 610609
rect 547678 610373 547898 610376
rect 228352 610110 228368 610343
rect 228368 610107 228463 610110
rect 241418 610056 241434 610289
rect 360512 610110 360528 610343
rect 360528 610107 360748 610110
rect 373578 610056 373594 610289
rect 402352 610110 402368 610343
rect 402368 610107 402463 610110
rect 415418 610056 415434 610289
rect 534512 610110 534528 610343
rect 534528 610107 534748 610110
rect 547578 610056 547594 610289
rect 241198 610053 241418 610056
rect 373358 610053 373578 610056
rect 415198 610053 415418 610056
rect 547358 610053 547578 610056
rect 228675 609787 228691 610015
rect 360835 609796 360842 610020
rect 228691 609784 228702 609787
rect 360842 609784 360862 609796
rect 402675 609787 402691 610015
rect 534835 609796 534842 610020
rect 402691 609784 402702 609787
rect 534842 609784 534862 609796
rect 608262 599387 608264 599512
rect 693736 599428 693738 599512
rect 693820 599387 693822 599428
rect 782262 599387 782264 599512
rect 867736 599428 867738 599512
rect 867820 599387 867822 599428
rect 275740 587418 275744 587434
rect 296740 587418 296744 587434
rect 317540 587418 317744 587434
rect 338740 587418 338744 587434
rect 449740 587418 449744 587434
rect 470740 587418 470744 587434
rect 491540 587418 491744 587434
rect 512740 587418 512744 587434
rect 625740 587418 625744 587434
rect 646740 587418 646744 587434
rect 667740 587418 667744 587434
rect 688740 587418 688744 587434
rect 799740 587418 799744 587434
rect 820740 587418 820744 587434
rect 841740 587418 841744 587434
rect 862740 587418 862744 587434
rect 275744 587410 275747 587418
rect 296744 587410 296747 587418
rect 317744 587198 317747 587418
rect 338744 587410 338747 587418
rect 449744 587410 449747 587418
rect 470744 587410 470747 587418
rect 491744 587198 491747 587418
rect 512744 587410 512747 587418
rect 625744 587410 625747 587418
rect 646744 587410 646747 587418
rect 667744 587410 667747 587418
rect 688744 587410 688747 587418
rect 799744 587410 799747 587418
rect 820744 587410 820747 587418
rect 841744 587410 841747 587418
rect 862744 587410 862747 587418
rect 262996 587158 263220 587165
rect 283996 587158 284220 587165
rect 304996 587158 305220 587165
rect 325996 587158 326220 587165
rect 436996 587158 437220 587165
rect 457996 587158 458220 587165
rect 478996 587158 479220 587165
rect 499996 587158 500220 587165
rect 612996 587158 613220 587165
rect 633996 587158 634220 587165
rect 654996 587158 655220 587165
rect 675996 587158 676220 587165
rect 786996 587158 787220 587165
rect 807996 587158 808220 587165
rect 828996 587158 829220 587165
rect 849996 587158 850220 587165
rect 262984 587138 262996 587158
rect 283984 587138 283996 587158
rect 304984 587138 304996 587158
rect 325984 587138 325996 587158
rect 436984 587138 436996 587158
rect 457984 587138 457996 587158
rect 478984 587138 478996 587158
rect 499984 587138 499996 587158
rect 612984 587138 612996 587158
rect 633984 587138 633996 587158
rect 654984 587138 654996 587158
rect 675984 587138 675996 587158
rect 786984 587138 786996 587158
rect 807984 587138 807996 587158
rect 828984 587138 828996 587158
rect 849984 587138 849996 587158
rect 276013 574691 276016 574702
rect 297013 574691 297016 574702
rect 318013 574691 318016 574702
rect 339013 574691 339016 574702
rect 450013 574691 450016 574702
rect 471013 574691 471016 574702
rect 492013 574691 492016 574702
rect 513013 574691 513016 574702
rect 626013 574691 626016 574702
rect 647013 574691 647016 574702
rect 668013 574691 668016 574702
rect 689013 574691 689016 574702
rect 800013 574691 800016 574702
rect 821013 574691 821016 574702
rect 842013 574691 842016 574702
rect 863013 574691 863016 574702
rect 275785 574675 276013 574691
rect 296785 574675 297013 574691
rect 317785 574675 318013 574691
rect 338785 574675 339013 574691
rect 449785 574675 450013 574691
rect 470785 574675 471013 574691
rect 491785 574675 492013 574691
rect 512785 574675 513013 574691
rect 625785 574675 626013 574691
rect 646785 574675 647013 574691
rect 667785 574675 668013 574691
rect 688785 574675 689013 574691
rect 799785 574675 800013 574691
rect 820785 574675 821013 574691
rect 841785 574675 842013 574691
rect 862785 574675 863013 574691
rect 263253 574422 263256 574642
rect 284253 574422 284256 574463
rect 305253 574422 305256 574642
rect 263256 574406 263260 574422
rect 284256 574420 284258 574422
rect 284258 574406 284260 574420
rect 305256 574406 305260 574422
rect 317690 574368 317693 574463
rect 326253 574422 326256 574642
rect 437253 574422 437256 574642
rect 458253 574422 458256 574463
rect 479253 574422 479256 574642
rect 326256 574406 326260 574422
rect 437256 574406 437260 574422
rect 458256 574420 458258 574422
rect 458258 574406 458260 574420
rect 479256 574406 479260 574422
rect 491690 574368 491693 574463
rect 500253 574422 500256 574642
rect 613253 574422 613256 574642
rect 634253 574422 634256 574463
rect 655253 574422 655256 574463
rect 676253 574422 676256 574642
rect 787253 574422 787256 574642
rect 808253 574422 808256 574463
rect 829253 574422 829256 574463
rect 850253 574422 850256 574642
rect 500256 574406 500260 574422
rect 613256 574406 613260 574422
rect 634256 574420 634258 574422
rect 655256 574420 655258 574422
rect 634258 574406 634260 574420
rect 655258 574406 655260 574420
rect 676256 574406 676260 574422
rect 787256 574406 787260 574422
rect 808256 574420 808258 574422
rect 829256 574420 829258 574422
rect 808258 574406 808260 574420
rect 829258 574406 829260 574420
rect 850256 574406 850260 574422
rect 317540 574352 317690 574368
rect 491540 574352 491690 574368
use one_padframe_var1  one_padframe_var1_0
timestamp 1689778135
transform 1 0 222000 0 1 568000
box 0 0 158000 180600
use one_padframe_var1  one_padframe_var1_1
timestamp 1689778135
transform 1 0 222000 0 1 768000
box 0 0 158000 180600
use one_padframe_var1  one_padframe_var1_2
timestamp 1689778135
transform 1 0 222000 0 1 968000
box 0 0 158000 180600
use one_padframe_var1  one_padframe_var1_3
timestamp 1689778135
transform 1 0 222000 0 1 1168000
box 0 0 158000 180600
use one_padframe_var1B  one_padframe_var1B_0
timestamp 1689778135
transform 1 0 222000 0 1 1368000
box 0 0 158000 180600
use one_padframe_var2  one_padframe_var2_0
timestamp 1689778135
transform 1 0 396000 0 1 568000
box 0 0 158000 180600
use one_padframe_var2  one_padframe_var2_1
timestamp 1689778135
transform 1 0 396000 0 1 768000
box 0 0 158000 180600
use one_padframe_var2  one_padframe_var2_2
timestamp 1689778135
transform 1 0 396000 0 1 968000
box 0 0 158000 180600
use one_padframe_var2  one_padframe_var2_3
timestamp 1689778135
transform 1 0 396000 0 1 1168000
box 0 0 158000 180600
use one_padframe_var2B  one_padframe_var2B_0
timestamp 1689778135
transform 1 0 396000 0 1 1368000
box 0 0 158000 180600
use one_padframe_var3  one_padframe_var3_0
timestamp 1689778135
transform 1 0 572000 0 1 427000
box 0 141000 158000 1122600
use one_padframe_var4  one_padframe_var4_0
timestamp 1689778135
transform 1 0 746000 0 1 427000
box 0 141000 158000 1122600
<< end >>
