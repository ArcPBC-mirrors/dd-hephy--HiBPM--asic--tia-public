magic
tech sky130A
magscale 1 2
timestamp 1699354420
<< error_p >>
rect 55542 94254 55779 94278
rect 55542 94217 55562 94254
rect 55539 94208 55542 94217
rect 55564 94210 55584 94254
rect 55629 94217 55779 94254
rect 55402 94201 55539 94208
rect 55561 94201 55564 94210
rect 55402 93785 55561 94201
rect 55629 94197 55770 94217
rect 55779 94208 55798 94217
rect 55769 94187 55788 94196
rect 55798 94188 56771 94208
rect 55302 93778 55402 93785
rect 55424 93778 55561 93785
rect 55789 93785 56771 94188
rect 55302 93638 55424 93778
rect 55789 93765 56762 93785
rect 56771 93765 57110 93785
rect 56762 93638 57110 93765
rect 55302 93478 55402 93638
rect 56762 93618 57101 93638
rect 57110 93618 57399 93638
rect 57101 93512 57399 93618
rect 57101 93507 57390 93512
rect 57399 93507 57410 93512
rect 57101 93492 57478 93507
rect 57386 93483 57478 93492
rect 55227 93471 55302 93478
rect 55324 93471 55424 93478
rect 55227 93402 55324 93471
rect 57403 93458 57478 93483
rect 57454 93412 57478 93458
rect 55227 93246 55302 93402
rect 57390 93281 57478 93412
rect 57378 93271 57390 93280
rect 57411 93271 57478 93281
rect 57378 93269 57411 93271
rect 57374 93267 57411 93269
rect 57373 93252 57411 93267
rect 57340 93247 57411 93252
rect 54175 93239 55227 93246
rect 55249 93239 55324 93246
rect 57340 93245 57399 93247
rect 57340 93243 57398 93245
rect 54175 93170 55249 93239
rect 57340 93180 57397 93243
rect 57259 93170 57340 93180
rect 57361 93170 57397 93180
rect 54175 90008 55227 93170
rect 57259 93021 57361 93170
rect 55617 93011 57259 93020
rect 57280 93011 57361 93021
rect 55617 93010 57280 93011
rect 55638 90008 57280 93010
rect 53985 90001 54175 90008
rect 54197 90001 55249 90008
rect 53985 89772 54197 90001
rect 55617 89782 57280 90008
rect 55321 89772 55617 89782
rect 55638 89772 57280 89782
rect 53985 89423 54175 89772
rect 53960 89416 53985 89423
rect 54007 89416 54197 89423
rect 53960 89346 54007 89416
rect 55342 89347 55638 89772
rect 53908 89339 53960 89346
rect 53982 89340 54007 89346
rect 53908 89186 53982 89339
rect 55321 89197 55638 89347
rect 53787 89179 53908 89186
rect 53930 89179 53982 89186
rect 55282 89187 55321 89196
rect 55342 89187 55638 89197
rect 53787 89110 53930 89179
rect 55282 89120 55342 89187
rect 55201 89110 55282 89120
rect 55303 89110 55342 89120
rect 53787 88813 53908 89110
rect 55201 88961 55303 89110
rect 55011 88951 55201 88960
rect 55222 88951 55303 88961
rect 55011 88950 55222 88951
rect 55032 88813 55222 88950
rect 53140 88806 53787 88813
rect 53809 88806 53930 88813
rect 53140 88577 53809 88806
rect 55011 88587 55222 88813
rect 54002 88577 55011 88587
rect 55032 88577 55222 88587
rect 53140 86821 53787 88577
rect 53115 86814 53140 86821
rect 53162 86814 53809 86821
rect 53115 86745 53162 86814
rect 54023 86745 55032 88577
rect 53063 86738 53115 86745
rect 53137 86738 53162 86745
rect 53063 86585 53137 86738
rect 54002 86595 55032 86745
rect 52942 86578 53063 86585
rect 53085 86578 53137 86585
rect 53963 86585 54002 86595
rect 54023 86585 55032 86595
rect 52942 86509 53085 86578
rect 53963 86519 54023 86585
rect 53882 86509 53963 86519
rect 53984 86509 54023 86519
rect 52942 86211 53063 86509
rect 53882 86359 53984 86509
rect 53693 86349 53882 86359
rect 53903 86349 53984 86359
rect 53714 86211 53903 86349
rect 52599 86204 52942 86211
rect 52964 86204 53085 86211
rect 52599 85975 52964 86204
rect 53693 85985 53903 86211
rect 53157 85975 53693 85985
rect 53714 85975 53903 85985
rect 52599 85154 52942 85975
rect 52574 85147 52599 85154
rect 52621 85147 52964 85154
rect 52574 85077 52621 85147
rect 52596 85076 52621 85077
rect 52573 85074 52621 85076
rect 52596 85073 52621 85074
rect 52572 85071 52621 85073
rect 52571 85068 52595 85070
rect 52570 85065 52594 85067
rect 52569 85061 52593 85064
rect 52568 85058 52593 85061
rect 53178 85058 53714 85975
rect 52522 85037 52593 85058
rect 52522 85034 52592 85037
rect 52522 84911 52589 85034
rect 53157 84928 53714 85058
rect 53118 84918 53157 84928
rect 53178 84918 53714 84928
rect 52522 84863 52546 84911
rect 52522 84845 52577 84863
rect 53118 84852 53178 84918
rect 52522 84844 52593 84845
rect 52522 84843 52595 84844
rect 52522 84842 52597 84843
rect 53113 84842 53118 84851
rect 53139 84842 53178 84852
rect 52522 84837 52598 84842
rect 53109 84840 53118 84842
rect 52522 84821 52716 84837
rect 53109 84833 53114 84840
rect 53134 84831 53139 84842
rect 53106 84828 53107 84830
rect 52570 84820 52716 84821
rect 52571 84819 52716 84820
rect 52573 84818 52716 84819
rect 52574 84777 52716 84818
rect 53076 84822 53106 84828
rect 53129 84822 53134 84831
rect 53076 84821 53129 84822
rect 53076 84818 53106 84821
rect 53127 84818 53128 84820
rect 52574 84758 52707 84777
rect 52716 84758 52811 84777
rect 53076 84768 53127 84818
rect 52707 84738 52811 84758
rect 53054 84758 53076 84768
rect 53097 84758 53127 84768
rect 53054 84738 53097 84758
rect 52707 84737 52828 84738
rect 52707 84736 52830 84737
rect 53050 84736 53097 84738
rect 52707 84735 52832 84736
rect 52707 84734 52834 84735
rect 53049 84734 53097 84736
rect 52707 84733 52836 84734
rect 52707 84732 52838 84733
rect 53048 84732 53097 84734
rect 52707 84731 52840 84732
rect 52707 84730 52842 84731
rect 53047 84730 53097 84732
rect 52707 84729 52845 84730
rect 52707 84728 52848 84729
rect 53046 84728 53097 84730
rect 52707 84727 52850 84728
rect 52707 84726 52852 84727
rect 53045 84726 53097 84728
rect 52707 84725 52855 84726
rect 52707 84720 52856 84725
rect 52707 84715 52971 84720
rect 52802 84714 52971 84715
rect 52804 84713 52971 84714
rect 52806 84712 52971 84713
rect 52808 84711 52971 84712
rect 53044 84715 53097 84726
rect 53044 84714 53075 84715
rect 53044 84712 53074 84714
rect 53044 84711 53073 84712
rect 52810 84710 52971 84711
rect 52812 84709 52971 84710
rect 52815 84708 52971 84709
rect 52817 84707 52971 84708
rect 52819 84706 52971 84707
rect 52821 84705 52971 84706
rect 52824 84704 52971 84705
rect 52827 84703 52971 84704
rect 52829 84702 52971 84703
rect 52831 84701 52971 84702
rect 52832 84666 52971 84701
rect 53017 84710 53073 84711
rect 53017 84708 53072 84710
rect 53017 84706 53071 84708
rect 53017 84704 53070 84706
rect 53017 84702 53069 84704
rect 53017 84666 53068 84702
rect 52832 84642 53068 84666
rect 67802 82454 71518 82478
rect 67802 75866 67826 82454
rect 70827 82118 71518 82454
rect 70827 82102 71507 82118
rect 70827 82098 71518 82102
rect 71502 81678 71518 82098
rect 71502 81666 71942 81678
rect 71958 81666 72198 81678
rect 71502 81662 72198 81666
rect 71939 81318 72198 81662
rect 71939 81306 72179 81318
rect 72198 81305 72251 81318
rect 69134 81259 70346 81266
rect 69134 81242 70482 81259
rect 72178 81242 72251 81305
rect 69134 79558 69158 81242
rect 70322 81238 70335 81242
rect 70341 81238 70482 81242
rect 72198 81238 72251 81242
rect 70335 81219 70482 81238
rect 72178 81225 72231 81238
rect 72251 81226 72278 81238
rect 70335 81198 70476 81219
rect 70482 81198 70608 81219
rect 70476 81183 70608 81198
rect 72232 81198 72278 81226
rect 72232 81195 72259 81198
rect 72232 81186 72275 81195
rect 70476 81162 70602 81183
rect 70615 81162 70735 81181
rect 70602 81101 70735 81162
rect 70602 81082 70722 81101
rect 70735 81097 70741 81101
rect 70722 81078 70728 81082
rect 70741 81078 70855 81097
rect 70728 81021 70855 81078
rect 72255 81075 72275 81186
rect 72278 81078 72298 81198
rect 70728 81002 70842 81021
rect 70862 81002 70886 81014
rect 70842 80974 70886 81002
rect 72275 80999 72288 81075
rect 72298 81002 72311 81078
rect 70842 80962 70866 80974
rect 70886 80962 70958 80974
rect 70866 80854 70958 80962
rect 72288 80879 72308 80999
rect 72311 80879 72331 81002
rect 72288 80878 72331 80879
rect 72288 80876 72308 80878
rect 70866 80842 70938 80854
rect 70958 80842 70982 80854
rect 70938 80814 70982 80842
rect 70938 80802 70962 80814
rect 70962 80766 70980 80802
rect 70983 80776 71001 80812
rect 72308 80803 72321 80875
rect 72331 80803 72344 80878
rect 72308 80802 72344 80803
rect 72308 80800 72321 80802
rect 72344 80799 72371 80802
rect 71001 80766 71063 80776
rect 70980 80653 71063 80766
rect 70980 80643 71042 80653
rect 71063 80643 71101 80653
rect 72321 80643 72371 80799
rect 71042 80639 71080 80643
rect 72344 80639 72371 80643
rect 71042 80577 71101 80639
rect 72321 80638 72371 80639
rect 72321 80636 72348 80638
rect 71042 80567 71080 80577
rect 71101 80572 71103 80576
rect 71080 80566 71104 80567
rect 71080 80562 71082 80566
rect 72348 80564 72360 80635
rect 72371 80567 72383 80638
rect 71082 80358 71106 80562
rect 72360 80558 72362 80562
rect 72383 80558 72385 80567
rect 72360 80553 72385 80558
rect 72362 80547 72386 80552
rect 72363 80478 72375 80543
rect 72386 80478 72398 80547
rect 72363 80474 72398 80478
rect 72374 80404 72398 80474
rect 72363 80402 72398 80404
rect 71002 80352 71082 80358
rect 71002 80078 71105 80352
rect 72363 80311 72375 80402
rect 72363 80309 72364 80311
rect 72386 80309 72398 80402
rect 72362 80304 72386 80309
rect 72385 80301 72386 80304
rect 72361 80297 72385 80301
rect 72360 80294 72385 80297
rect 72360 80285 72362 80294
rect 72335 80282 72360 80284
rect 72383 80282 72385 80294
rect 72335 80081 72383 80282
rect 70802 80065 71002 80078
rect 71025 80072 71105 80078
rect 72325 80079 72335 80081
rect 72358 80079 72383 80081
rect 72325 80078 72358 80079
rect 70802 80002 71021 80065
rect 72325 80005 72335 80078
rect 70802 79798 71002 80002
rect 72305 79844 72325 80004
rect 72348 80002 72358 80078
rect 72300 79801 72305 79844
rect 72328 79842 72348 80002
rect 72295 79799 72300 79801
rect 72323 79799 72328 79842
rect 72295 79798 72323 79799
rect 70482 79780 70802 79798
rect 70821 79785 71021 79798
rect 70482 79762 70816 79780
rect 72295 79772 72300 79798
rect 72277 79765 72300 79772
rect 70482 79558 70802 79762
rect 72277 79732 72297 79765
rect 72318 79762 72323 79798
rect 72197 79722 72277 79732
rect 72298 79722 72318 79762
rect 72197 79572 72298 79722
rect 72195 79568 72197 79572
rect 72157 79558 72195 79568
rect 72218 79562 72298 79572
rect 72216 79558 72218 79562
rect 69134 79540 70816 79558
rect 69134 79534 70506 79540
rect 72157 79492 72216 79558
rect 72077 79482 72157 79492
rect 72178 79482 72216 79492
rect 72077 79332 72178 79482
rect 72017 79322 72077 79332
rect 72098 79322 72178 79332
rect 72017 79217 72098 79322
rect 71621 79212 72098 79217
rect 71621 79202 72021 79212
rect 72038 79202 72098 79212
rect 71621 78780 72038 79202
rect 71066 78777 72038 78780
rect 71066 78762 71626 78777
rect 71638 78762 72038 78777
rect 71066 78423 71638 78762
rect 70434 78420 71638 78423
rect 70434 78402 71074 78420
rect 71078 78402 71638 78420
rect 70434 78303 71078 78402
rect 70438 78282 71078 78303
rect 69158 78242 70438 78282
rect 69134 75866 69158 78242
rect 67802 75842 69158 75866
<< via4 >>
tri 55542 94217 55562 94278 se
rect 55562 94217 55638 94278
tri 55638 94217 55779 94278 sw
tri 55539 94208 55542 94217 se
rect 55542 94208 55779 94217
tri 55779 94208 55798 94217 sw
tri 55402 93785 55539 94208 se
rect 55539 93785 55798 94208
tri 55798 93785 56771 94208 sw
tri 55302 93478 55402 93785 se
rect 55402 93638 56771 93785
tri 56771 93638 57110 93785 sw
rect 55402 93512 57110 93638
tri 57110 93512 57399 93638 sw
rect 55402 93507 57399 93512
tri 57399 93507 57410 93512 sw
rect 55402 93478 57412 93507
tri 57412 93478 57478 93507 sw
tri 55227 93246 55302 93478 se
rect 55302 93402 57478 93478
rect 55302 93269 57411 93402
tri 57411 93271 57478 93402 nw
rect 55302 93246 57399 93269
tri 57399 93247 57411 93269 nw
tri 54175 90008 55227 93246 se
rect 55227 93245 57399 93246
rect 55227 93243 57398 93245
rect 55227 93242 57397 93243
rect 55227 93170 57361 93242
tri 57361 93170 57397 93242 nw
rect 55227 93010 57280 93170
tri 57280 93011 57361 93170 nw
rect 55227 90008 55638 93010
tri 53985 89423 54175 90008 se
rect 54175 89772 55638 90008
tri 55638 89772 57280 93010 nw
rect 54175 89423 55342 89772
tri 53960 89347 53985 89423 se
rect 53985 89347 55342 89423
tri 53908 89186 53960 89346 se
rect 53960 89186 55342 89347
tri 55342 89187 55638 89772 nw
tri 53787 88813 53908 89186 se
rect 53908 89110 55303 89186
tri 55303 89110 55342 89186 nw
rect 53908 88950 55222 89110
tri 55222 88951 55303 89110 nw
rect 53908 88813 55032 88950
tri 53140 86821 53787 88813 se
rect 53787 88577 55032 88813
tri 55032 88577 55222 88950 nw
rect 53787 86821 54023 88577
tri 53115 86745 53140 86821 se
rect 53140 86745 54023 86821
tri 53063 86585 53115 86745 se
rect 53115 86585 54023 86745
tri 54023 86585 55032 88577 nw
tri 52942 86211 53063 86585 se
rect 53063 86509 53984 86585
tri 53984 86509 54023 86585 nw
rect 53063 86349 53903 86509
tri 53903 86349 53984 86509 nw
rect 53063 86211 53714 86349
tri 52599 85154 52942 86211 se
rect 52942 85975 53714 86211
tri 53714 85975 53903 86349 nw
rect 52942 85154 53178 85975
tri 52574 85078 52599 85154 se
rect 52599 85078 53178 85154
tri 52573 85076 52574 85077 se
rect 52574 85076 53178 85078
tri 52572 85073 52573 85074 se
rect 52573 85073 53178 85076
tri 52571 85070 52572 85071 se
rect 52572 85070 53178 85073
tri 52570 85067 52571 85068 se
rect 52571 85067 53178 85070
tri 52569 85064 52570 85065 se
rect 52570 85064 53178 85067
rect 52569 85061 53178 85064
rect 52568 85058 53178 85061
tri 52522 84918 52567 85058 se
rect 52567 84918 53178 85058
tri 53178 84918 53714 85975 nw
rect 52522 84842 53139 84918
tri 53139 84842 53178 84918 nw
tri 52522 84821 52567 84842 ne
rect 52567 84831 53134 84842
tri 53134 84831 53139 84842 nw
rect 52567 84821 53129 84831
tri 53129 84822 53134 84831 nw
tri 52569 84820 52570 84821 ne
rect 52570 84820 53128 84821
tri 53128 84820 53129 84821 nw
rect 52571 84819 53127 84820
rect 52573 84818 53127 84819
tri 53127 84818 53128 84820 nw
tri 52574 84758 52707 84818 ne
rect 52707 84758 53097 84818
tri 53097 84758 53127 84818 nw
tri 52707 84715 52802 84758 ne
rect 52802 84714 53075 84758
tri 53075 84715 53097 84758 nw
rect 52804 84713 53074 84714
rect 52806 84712 53074 84713
rect 52808 84711 53073 84712
rect 52810 84710 53073 84711
rect 52812 84709 53072 84710
tri 52814 84708 52815 84709 ne
rect 52815 84708 53072 84709
tri 52816 84707 52817 84708 ne
rect 52817 84707 53071 84708
tri 52818 84706 52819 84707 ne
rect 52819 84706 53071 84707
rect 52821 84705 53070 84706
rect 52824 84704 53070 84705
tri 52826 84703 52827 84704 ne
rect 52827 84703 53069 84704
tri 52828 84702 52829 84703 ne
rect 52829 84702 53069 84703
rect 52831 84701 53068 84702
tri 52832 84642 52962 84701 ne
rect 52962 84642 53038 84701
tri 53038 84642 53068 84701 nw
rect 67802 82118 70838 82478
tri 70838 82118 71518 82478 sw
rect 67802 81678 71518 82118
tri 71518 81678 71958 82118 sw
rect 67802 81318 71958 81678
tri 71958 81318 72198 81678 sw
rect 67802 81242 72198 81318
rect 67802 79558 69158 81242
tri 70322 81238 70335 81242 ne
rect 70335 81238 72198 81242
tri 72198 81238 72251 81318 sw
tri 70335 81198 70476 81238 ne
rect 70476 81198 72251 81238
tri 72251 81198 72278 81238 sw
tri 70476 81162 70602 81198 ne
rect 70602 81162 72278 81198
tri 70602 81082 70722 81162 ne
rect 70722 81082 72278 81162
tri 70722 81078 70728 81082 ne
rect 70728 81078 72278 81082
tri 72278 81078 72298 81198 sw
tri 70728 81002 70842 81078 ne
rect 70842 81002 72298 81078
tri 72298 81002 72311 81078 sw
tri 70842 80962 70866 81002 ne
rect 70866 80962 72311 81002
tri 70866 80842 70938 80962 ne
rect 70938 80879 72311 80962
tri 72311 80879 72331 81002 sw
rect 70938 80842 72331 80879
tri 70938 80802 70962 80842 ne
rect 70962 80803 72331 80842
tri 72331 80803 72344 80878 sw
rect 70962 80802 72344 80803
tri 70962 80766 70980 80802 ne
rect 70980 80766 72344 80802
tri 70980 80643 71042 80766 ne
rect 71042 80643 72344 80766
tri 71042 80567 71080 80643 ne
rect 71080 80639 72344 80643
tri 72344 80639 72371 80802 sw
rect 71080 80567 72371 80639
tri 72371 80567 72383 80638 sw
rect 71080 80566 72383 80567
tri 71080 80562 71082 80566 ne
rect 71082 80558 72383 80566
tri 72383 80558 72385 80567 sw
rect 71082 80552 72385 80558
tri 72385 80552 72386 80553 sw
rect 71082 80478 72386 80552
tri 72386 80478 72398 80547 sw
rect 71082 80402 72398 80478
tri 71002 80078 71082 80358 se
rect 71082 80304 72386 80402
tri 72386 80309 72398 80402 nw
rect 71082 80294 72385 80304
tri 72385 80301 72386 80304 nw
rect 71082 80282 72383 80294
tri 72383 80282 72385 80294 nw
rect 71082 80078 72358 80282
tri 72358 80079 72383 80282 nw
tri 70802 79798 71002 80078 se
rect 71002 80002 72348 80078
tri 72348 80002 72358 80078 nw
rect 71002 79842 72328 80002
tri 72328 79842 72348 80002 nw
rect 71002 79798 72323 79842
tri 72323 79799 72328 79842 nw
tri 70482 79558 70802 79798 se
rect 70802 79762 72318 79798
tri 72318 79762 72323 79798 nw
rect 70802 79722 72298 79762
tri 72298 79722 72318 79762 nw
rect 70802 79562 72218 79722
tri 72218 79562 72298 79722 nw
rect 70802 79558 72216 79562
tri 72216 79558 72218 79562 nw
rect 67802 79482 72178 79558
tri 72178 79482 72216 79558 nw
rect 67802 79322 72098 79482
tri 72098 79322 72178 79482 nw
rect 67802 79202 72038 79322
tri 72038 79202 72098 79322 nw
rect 67802 78762 71638 79202
tri 71638 78762 72038 79202 nw
rect 67802 78402 71078 78762
tri 71078 78402 71638 78762 nw
rect 67802 78282 70438 78402
tri 70438 78282 71078 78402 nw
rect 67802 75842 69158 78282
tri 69158 78242 70438 78282 nw
<< end >>
