magic
tech sky130A
magscale 1 2
timestamp 1683806952
<< error_p >>
rect -147 890 -89 896
rect -29 890 29 896
rect 89 890 147 896
rect -147 856 -135 890
rect -29 856 -17 890
rect 89 856 101 890
rect -147 850 -89 856
rect -29 850 29 856
rect 89 850 147 856
rect -147 380 -89 386
rect -29 380 29 386
rect 89 380 147 386
rect -147 346 -135 380
rect -29 346 -17 380
rect 89 346 101 380
rect -147 340 -89 346
rect -29 340 29 346
rect 89 340 147 346
rect -147 272 -89 278
rect -29 272 29 278
rect 89 272 147 278
rect -147 238 -135 272
rect -29 238 -17 272
rect 89 238 101 272
rect -147 232 -89 238
rect -29 232 29 238
rect 89 232 147 238
rect -147 -238 -89 -232
rect -29 -238 29 -232
rect 89 -238 147 -232
rect -147 -272 -135 -238
rect -29 -272 -17 -238
rect 89 -272 101 -238
rect -147 -278 -89 -272
rect -29 -278 29 -272
rect 89 -278 147 -272
rect -147 -346 -89 -340
rect -29 -346 29 -340
rect 89 -346 147 -340
rect -147 -380 -135 -346
rect -29 -380 -17 -346
rect 89 -380 101 -346
rect -147 -386 -89 -380
rect -29 -386 29 -380
rect 89 -386 147 -380
rect -147 -856 -89 -850
rect -29 -856 29 -850
rect 89 -856 147 -850
rect -147 -890 -135 -856
rect -29 -890 -17 -856
rect 89 -890 101 -856
rect -147 -896 -89 -890
rect -29 -896 29 -890
rect 89 -896 147 -890
<< pwell >>
rect -344 -1028 344 1028
<< nmoslvt >>
rect -148 418 -88 818
rect -30 418 30 818
rect 88 418 148 818
rect -148 -200 -88 200
rect -30 -200 30 200
rect 88 -200 148 200
rect -148 -818 -88 -418
rect -30 -818 30 -418
rect 88 -818 148 -418
<< ndiff >>
rect -206 806 -148 818
rect -206 430 -194 806
rect -160 430 -148 806
rect -206 418 -148 430
rect -88 806 -30 818
rect -88 430 -76 806
rect -42 430 -30 806
rect -88 418 -30 430
rect 30 806 88 818
rect 30 430 42 806
rect 76 430 88 806
rect 30 418 88 430
rect 148 806 206 818
rect 148 430 160 806
rect 194 430 206 806
rect 148 418 206 430
rect -206 188 -148 200
rect -206 -188 -194 188
rect -160 -188 -148 188
rect -206 -200 -148 -188
rect -88 188 -30 200
rect -88 -188 -76 188
rect -42 -188 -30 188
rect -88 -200 -30 -188
rect 30 188 88 200
rect 30 -188 42 188
rect 76 -188 88 188
rect 30 -200 88 -188
rect 148 188 206 200
rect 148 -188 160 188
rect 194 -188 206 188
rect 148 -200 206 -188
rect -206 -430 -148 -418
rect -206 -806 -194 -430
rect -160 -806 -148 -430
rect -206 -818 -148 -806
rect -88 -430 -30 -418
rect -88 -806 -76 -430
rect -42 -806 -30 -430
rect -88 -818 -30 -806
rect 30 -430 88 -418
rect 30 -806 42 -430
rect 76 -806 88 -430
rect 30 -818 88 -806
rect 148 -430 206 -418
rect 148 -806 160 -430
rect 194 -806 206 -430
rect 148 -818 206 -806
<< ndiffc >>
rect -194 430 -160 806
rect -76 430 -42 806
rect 42 430 76 806
rect 160 430 194 806
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect -194 -806 -160 -430
rect -76 -806 -42 -430
rect 42 -806 76 -430
rect 160 -806 194 -430
<< psubdiff >>
rect -308 958 -212 992
rect 212 958 308 992
rect -308 896 -274 958
rect 274 896 308 958
rect -308 -958 -274 -896
rect 274 -958 308 -896
rect -308 -992 -212 -958
rect 212 -992 308 -958
<< psubdiffcont >>
rect -212 958 212 992
rect -308 -896 -274 896
rect 274 -896 308 896
rect -212 -992 212 -958
<< poly >>
rect -151 890 -85 906
rect -151 856 -135 890
rect -101 856 -85 890
rect -151 840 -85 856
rect -33 890 33 906
rect -33 856 -17 890
rect 17 856 33 890
rect -33 840 33 856
rect 85 890 151 906
rect 85 856 101 890
rect 135 856 151 890
rect 85 840 151 856
rect -148 818 -88 840
rect -30 818 30 840
rect 88 818 148 840
rect -148 396 -88 418
rect -30 396 30 418
rect 88 396 148 418
rect -151 380 -85 396
rect -151 346 -135 380
rect -101 346 -85 380
rect -151 330 -85 346
rect -33 380 33 396
rect -33 346 -17 380
rect 17 346 33 380
rect -33 330 33 346
rect 85 380 151 396
rect 85 346 101 380
rect 135 346 151 380
rect 85 330 151 346
rect -151 272 -85 288
rect -151 238 -135 272
rect -101 238 -85 272
rect -151 222 -85 238
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -33 222 33 238
rect 85 272 151 288
rect 85 238 101 272
rect 135 238 151 272
rect 85 222 151 238
rect -148 200 -88 222
rect -30 200 30 222
rect 88 200 148 222
rect -148 -222 -88 -200
rect -30 -222 30 -200
rect 88 -222 148 -200
rect -151 -238 -85 -222
rect -151 -272 -135 -238
rect -101 -272 -85 -238
rect -151 -288 -85 -272
rect -33 -238 33 -222
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 85 -238 151 -222
rect 85 -272 101 -238
rect 135 -272 151 -238
rect 85 -288 151 -272
rect -151 -346 -85 -330
rect -151 -380 -135 -346
rect -101 -380 -85 -346
rect -151 -396 -85 -380
rect -33 -346 33 -330
rect -33 -380 -17 -346
rect 17 -380 33 -346
rect -33 -396 33 -380
rect 85 -346 151 -330
rect 85 -380 101 -346
rect 135 -380 151 -346
rect 85 -396 151 -380
rect -148 -418 -88 -396
rect -30 -418 30 -396
rect 88 -418 148 -396
rect -148 -840 -88 -818
rect -30 -840 30 -818
rect 88 -840 148 -818
rect -151 -856 -85 -840
rect -151 -890 -135 -856
rect -101 -890 -85 -856
rect -151 -906 -85 -890
rect -33 -856 33 -840
rect -33 -890 -17 -856
rect 17 -890 33 -856
rect -33 -906 33 -890
rect 85 -856 151 -840
rect 85 -890 101 -856
rect 135 -890 151 -856
rect 85 -906 151 -890
<< polycont >>
rect -135 856 -101 890
rect -17 856 17 890
rect 101 856 135 890
rect -135 346 -101 380
rect -17 346 17 380
rect 101 346 135 380
rect -135 238 -101 272
rect -17 238 17 272
rect 101 238 135 272
rect -135 -272 -101 -238
rect -17 -272 17 -238
rect 101 -272 135 -238
rect -135 -380 -101 -346
rect -17 -380 17 -346
rect 101 -380 135 -346
rect -135 -890 -101 -856
rect -17 -890 17 -856
rect 101 -890 135 -856
<< locali >>
rect -308 958 -212 992
rect 212 958 308 992
rect -308 896 -274 958
rect 274 896 308 958
rect -151 856 -135 890
rect -101 856 -85 890
rect -33 856 -17 890
rect 17 856 33 890
rect 85 856 101 890
rect 135 856 151 890
rect -194 806 -160 822
rect -194 414 -160 430
rect -76 806 -42 822
rect -76 414 -42 430
rect 42 806 76 822
rect 42 414 76 430
rect 160 806 194 822
rect 160 414 194 430
rect -151 346 -135 380
rect -101 346 -85 380
rect -33 346 -17 380
rect 17 346 33 380
rect 85 346 101 380
rect 135 346 151 380
rect -151 238 -135 272
rect -101 238 -85 272
rect -33 238 -17 272
rect 17 238 33 272
rect 85 238 101 272
rect 135 238 151 272
rect -194 188 -160 204
rect -194 -204 -160 -188
rect -76 188 -42 204
rect -76 -204 -42 -188
rect 42 188 76 204
rect 42 -204 76 -188
rect 160 188 194 204
rect 160 -204 194 -188
rect -151 -272 -135 -238
rect -101 -272 -85 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 85 -272 101 -238
rect 135 -272 151 -238
rect -151 -380 -135 -346
rect -101 -380 -85 -346
rect -33 -380 -17 -346
rect 17 -380 33 -346
rect 85 -380 101 -346
rect 135 -380 151 -346
rect -194 -430 -160 -414
rect -194 -822 -160 -806
rect -76 -430 -42 -414
rect -76 -822 -42 -806
rect 42 -430 76 -414
rect 42 -822 76 -806
rect 160 -430 194 -414
rect 160 -822 194 -806
rect -151 -890 -135 -856
rect -101 -890 -85 -856
rect -33 -890 -17 -856
rect 17 -890 33 -856
rect 85 -890 101 -856
rect 135 -890 151 -856
rect -308 -958 -274 -896
rect 274 -958 308 -896
rect -308 -992 -212 -958
rect 212 -992 308 -958
<< viali >>
rect -135 856 -101 890
rect -17 856 17 890
rect 101 856 135 890
rect -194 430 -160 806
rect -76 430 -42 806
rect 42 430 76 806
rect 160 430 194 806
rect -135 346 -101 380
rect -17 346 17 380
rect 101 346 135 380
rect -135 238 -101 272
rect -17 238 17 272
rect 101 238 135 272
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect -135 -272 -101 -238
rect -17 -272 17 -238
rect 101 -272 135 -238
rect -135 -380 -101 -346
rect -17 -380 17 -346
rect 101 -380 135 -346
rect -194 -806 -160 -430
rect -76 -806 -42 -430
rect 42 -806 76 -430
rect 160 -806 194 -430
rect -135 -890 -101 -856
rect -17 -890 17 -856
rect 101 -890 135 -856
<< metal1 >>
rect -147 890 -89 896
rect -147 856 -135 890
rect -101 856 -89 890
rect -147 850 -89 856
rect -29 890 29 896
rect -29 856 -17 890
rect 17 856 29 890
rect -29 850 29 856
rect 89 890 147 896
rect 89 856 101 890
rect 135 856 147 890
rect 89 850 147 856
rect -200 806 -154 818
rect -200 430 -194 806
rect -160 430 -154 806
rect -200 418 -154 430
rect -82 806 -36 818
rect -82 430 -76 806
rect -42 430 -36 806
rect -82 418 -36 430
rect 36 806 82 818
rect 36 430 42 806
rect 76 430 82 806
rect 36 418 82 430
rect 154 806 200 818
rect 154 430 160 806
rect 194 430 200 806
rect 154 418 200 430
rect -147 380 -89 386
rect -147 346 -135 380
rect -101 346 -89 380
rect -147 340 -89 346
rect -29 380 29 386
rect -29 346 -17 380
rect 17 346 29 380
rect -29 340 29 346
rect 89 380 147 386
rect 89 346 101 380
rect 135 346 147 380
rect 89 340 147 346
rect -147 272 -89 278
rect -147 238 -135 272
rect -101 238 -89 272
rect -147 232 -89 238
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect 89 272 147 278
rect 89 238 101 272
rect 135 238 147 272
rect 89 232 147 238
rect -200 188 -154 200
rect -200 -188 -194 188
rect -160 -188 -154 188
rect -200 -200 -154 -188
rect -82 188 -36 200
rect -82 -188 -76 188
rect -42 -188 -36 188
rect -82 -200 -36 -188
rect 36 188 82 200
rect 36 -188 42 188
rect 76 -188 82 188
rect 36 -200 82 -188
rect 154 188 200 200
rect 154 -188 160 188
rect 194 -188 200 188
rect 154 -200 200 -188
rect -147 -238 -89 -232
rect -147 -272 -135 -238
rect -101 -272 -89 -238
rect -147 -278 -89 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 89 -238 147 -232
rect 89 -272 101 -238
rect 135 -272 147 -238
rect 89 -278 147 -272
rect -147 -346 -89 -340
rect -147 -380 -135 -346
rect -101 -380 -89 -346
rect -147 -386 -89 -380
rect -29 -346 29 -340
rect -29 -380 -17 -346
rect 17 -380 29 -346
rect -29 -386 29 -380
rect 89 -346 147 -340
rect 89 -380 101 -346
rect 135 -380 147 -346
rect 89 -386 147 -380
rect -200 -430 -154 -418
rect -200 -806 -194 -430
rect -160 -806 -154 -430
rect -200 -818 -154 -806
rect -82 -430 -36 -418
rect -82 -806 -76 -430
rect -42 -806 -36 -430
rect -82 -818 -36 -806
rect 36 -430 82 -418
rect 36 -806 42 -430
rect 76 -806 82 -430
rect 36 -818 82 -806
rect 154 -430 200 -418
rect 154 -806 160 -430
rect 194 -806 200 -430
rect 154 -818 200 -806
rect -147 -856 -89 -850
rect -147 -890 -135 -856
rect -101 -890 -89 -856
rect -147 -896 -89 -890
rect -29 -856 29 -850
rect -29 -890 -17 -856
rect 17 -890 29 -856
rect -29 -896 29 -890
rect 89 -856 147 -850
rect 89 -890 101 -856
rect 135 -890 147 -856
rect 89 -896 147 -890
<< properties >>
string FIXED_BBOX -291 -975 291 975
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.3 m 3 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
