magic
tech sky130A
magscale 1 2
timestamp 1683561438
<< nwell >>
rect -6173 963 -3907 1545
rect -3653 963 -1387 1545
rect -1133 963 1133 1545
rect 1387 963 3653 1545
rect 3907 963 6173 1545
rect -6173 127 -3907 709
rect -3653 127 -1387 709
rect -1133 127 1133 709
rect 1387 127 3653 709
rect 3907 127 6173 709
rect -6173 -709 -3907 -127
rect -3653 -709 -1387 -127
rect -1133 -709 1133 -127
rect 1387 -709 3653 -127
rect 3907 -709 6173 -127
rect -6173 -1545 -3907 -963
rect -3653 -1545 -1387 -963
rect -1133 -1545 1133 -963
rect 1387 -1545 3653 -963
rect 3907 -1545 6173 -963
<< pwell >>
rect -6283 1545 6283 1655
rect -6283 963 -6173 1545
rect -3907 963 -3653 1545
rect -1387 963 -1133 1545
rect 1133 963 1387 1545
rect 3653 963 3907 1545
rect 6173 963 6283 1545
rect -6283 709 6283 963
rect -6283 127 -6173 709
rect -3907 127 -3653 709
rect -1387 127 -1133 709
rect 1133 127 1387 709
rect 3653 127 3907 709
rect 6173 127 6283 709
rect -6283 -127 6283 127
rect -6283 -709 -6173 -127
rect -3907 -709 -3653 -127
rect -1387 -709 -1133 -127
rect 1133 -709 1387 -127
rect 3653 -709 3907 -127
rect 6173 -709 6283 -127
rect -6283 -963 6283 -709
rect -6283 -1545 -6173 -963
rect -3907 -1545 -3653 -963
rect -1387 -1545 -1133 -963
rect 1133 -1545 1387 -963
rect 3653 -1545 3907 -963
rect 6173 -1545 6283 -963
rect -6283 -1655 6283 -1545
<< varactor >>
rect -6040 1054 -4040 1454
rect -3520 1054 -1520 1454
rect -1000 1054 1000 1454
rect 1520 1054 3520 1454
rect 4040 1054 6040 1454
rect -6040 218 -4040 618
rect -3520 218 -1520 618
rect -1000 218 1000 618
rect 1520 218 3520 618
rect 4040 218 6040 618
rect -6040 -618 -4040 -218
rect -3520 -618 -1520 -218
rect -1000 -618 1000 -218
rect 1520 -618 3520 -218
rect 4040 -618 6040 -218
rect -6040 -1454 -4040 -1054
rect -3520 -1454 -1520 -1054
rect -1000 -1454 1000 -1054
rect 1520 -1454 3520 -1054
rect 4040 -1454 6040 -1054
<< psubdiff >>
rect -6247 1585 -6151 1619
rect 6151 1585 6247 1619
rect -6247 1523 -6213 1585
rect 6213 1523 6247 1585
rect -6247 -1585 -6213 -1523
rect 6213 -1585 6247 -1523
rect -6247 -1619 -6151 -1585
rect 6151 -1619 6247 -1585
<< nsubdiff >>
rect -6137 1430 -6040 1454
rect -6137 1078 -6125 1430
rect -6091 1078 -6040 1430
rect -6137 1054 -6040 1078
rect -4040 1430 -3943 1454
rect -4040 1078 -3989 1430
rect -3955 1078 -3943 1430
rect -4040 1054 -3943 1078
rect -3617 1430 -3520 1454
rect -3617 1078 -3605 1430
rect -3571 1078 -3520 1430
rect -3617 1054 -3520 1078
rect -1520 1430 -1423 1454
rect -1520 1078 -1469 1430
rect -1435 1078 -1423 1430
rect -1520 1054 -1423 1078
rect -1097 1430 -1000 1454
rect -1097 1078 -1085 1430
rect -1051 1078 -1000 1430
rect -1097 1054 -1000 1078
rect 1000 1430 1097 1454
rect 1000 1078 1051 1430
rect 1085 1078 1097 1430
rect 1000 1054 1097 1078
rect 1423 1430 1520 1454
rect 1423 1078 1435 1430
rect 1469 1078 1520 1430
rect 1423 1054 1520 1078
rect 3520 1430 3617 1454
rect 3520 1078 3571 1430
rect 3605 1078 3617 1430
rect 3520 1054 3617 1078
rect 3943 1430 4040 1454
rect 3943 1078 3955 1430
rect 3989 1078 4040 1430
rect 3943 1054 4040 1078
rect 6040 1430 6137 1454
rect 6040 1078 6091 1430
rect 6125 1078 6137 1430
rect 6040 1054 6137 1078
rect -6137 594 -6040 618
rect -6137 242 -6125 594
rect -6091 242 -6040 594
rect -6137 218 -6040 242
rect -4040 594 -3943 618
rect -4040 242 -3989 594
rect -3955 242 -3943 594
rect -4040 218 -3943 242
rect -3617 594 -3520 618
rect -3617 242 -3605 594
rect -3571 242 -3520 594
rect -3617 218 -3520 242
rect -1520 594 -1423 618
rect -1520 242 -1469 594
rect -1435 242 -1423 594
rect -1520 218 -1423 242
rect -1097 594 -1000 618
rect -1097 242 -1085 594
rect -1051 242 -1000 594
rect -1097 218 -1000 242
rect 1000 594 1097 618
rect 1000 242 1051 594
rect 1085 242 1097 594
rect 1000 218 1097 242
rect 1423 594 1520 618
rect 1423 242 1435 594
rect 1469 242 1520 594
rect 1423 218 1520 242
rect 3520 594 3617 618
rect 3520 242 3571 594
rect 3605 242 3617 594
rect 3520 218 3617 242
rect 3943 594 4040 618
rect 3943 242 3955 594
rect 3989 242 4040 594
rect 3943 218 4040 242
rect 6040 594 6137 618
rect 6040 242 6091 594
rect 6125 242 6137 594
rect 6040 218 6137 242
rect -6137 -242 -6040 -218
rect -6137 -594 -6125 -242
rect -6091 -594 -6040 -242
rect -6137 -618 -6040 -594
rect -4040 -242 -3943 -218
rect -4040 -594 -3989 -242
rect -3955 -594 -3943 -242
rect -4040 -618 -3943 -594
rect -3617 -242 -3520 -218
rect -3617 -594 -3605 -242
rect -3571 -594 -3520 -242
rect -3617 -618 -3520 -594
rect -1520 -242 -1423 -218
rect -1520 -594 -1469 -242
rect -1435 -594 -1423 -242
rect -1520 -618 -1423 -594
rect -1097 -242 -1000 -218
rect -1097 -594 -1085 -242
rect -1051 -594 -1000 -242
rect -1097 -618 -1000 -594
rect 1000 -242 1097 -218
rect 1000 -594 1051 -242
rect 1085 -594 1097 -242
rect 1000 -618 1097 -594
rect 1423 -242 1520 -218
rect 1423 -594 1435 -242
rect 1469 -594 1520 -242
rect 1423 -618 1520 -594
rect 3520 -242 3617 -218
rect 3520 -594 3571 -242
rect 3605 -594 3617 -242
rect 3520 -618 3617 -594
rect 3943 -242 4040 -218
rect 3943 -594 3955 -242
rect 3989 -594 4040 -242
rect 3943 -618 4040 -594
rect 6040 -242 6137 -218
rect 6040 -594 6091 -242
rect 6125 -594 6137 -242
rect 6040 -618 6137 -594
rect -6137 -1078 -6040 -1054
rect -6137 -1430 -6125 -1078
rect -6091 -1430 -6040 -1078
rect -6137 -1454 -6040 -1430
rect -4040 -1078 -3943 -1054
rect -4040 -1430 -3989 -1078
rect -3955 -1430 -3943 -1078
rect -4040 -1454 -3943 -1430
rect -3617 -1078 -3520 -1054
rect -3617 -1430 -3605 -1078
rect -3571 -1430 -3520 -1078
rect -3617 -1454 -3520 -1430
rect -1520 -1078 -1423 -1054
rect -1520 -1430 -1469 -1078
rect -1435 -1430 -1423 -1078
rect -1520 -1454 -1423 -1430
rect -1097 -1078 -1000 -1054
rect -1097 -1430 -1085 -1078
rect -1051 -1430 -1000 -1078
rect -1097 -1454 -1000 -1430
rect 1000 -1078 1097 -1054
rect 1000 -1430 1051 -1078
rect 1085 -1430 1097 -1078
rect 1000 -1454 1097 -1430
rect 1423 -1078 1520 -1054
rect 1423 -1430 1435 -1078
rect 1469 -1430 1520 -1078
rect 1423 -1454 1520 -1430
rect 3520 -1078 3617 -1054
rect 3520 -1430 3571 -1078
rect 3605 -1430 3617 -1078
rect 3520 -1454 3617 -1430
rect 3943 -1078 4040 -1054
rect 3943 -1430 3955 -1078
rect 3989 -1430 4040 -1078
rect 3943 -1454 4040 -1430
rect 6040 -1078 6137 -1054
rect 6040 -1430 6091 -1078
rect 6125 -1430 6137 -1078
rect 6040 -1454 6137 -1430
<< psubdiffcont >>
rect -6151 1585 6151 1619
rect -6247 -1523 -6213 1523
rect 6213 -1523 6247 1523
rect -6151 -1619 6151 -1585
<< nsubdiffcont >>
rect -6125 1078 -6091 1430
rect -3989 1078 -3955 1430
rect -3605 1078 -3571 1430
rect -1469 1078 -1435 1430
rect -1085 1078 -1051 1430
rect 1051 1078 1085 1430
rect 1435 1078 1469 1430
rect 3571 1078 3605 1430
rect 3955 1078 3989 1430
rect 6091 1078 6125 1430
rect -6125 242 -6091 594
rect -3989 242 -3955 594
rect -3605 242 -3571 594
rect -1469 242 -1435 594
rect -1085 242 -1051 594
rect 1051 242 1085 594
rect 1435 242 1469 594
rect 3571 242 3605 594
rect 3955 242 3989 594
rect 6091 242 6125 594
rect -6125 -594 -6091 -242
rect -3989 -594 -3955 -242
rect -3605 -594 -3571 -242
rect -1469 -594 -1435 -242
rect -1085 -594 -1051 -242
rect 1051 -594 1085 -242
rect 1435 -594 1469 -242
rect 3571 -594 3605 -242
rect 3955 -594 3989 -242
rect 6091 -594 6125 -242
rect -6125 -1430 -6091 -1078
rect -3989 -1430 -3955 -1078
rect -3605 -1430 -3571 -1078
rect -1469 -1430 -1435 -1078
rect -1085 -1430 -1051 -1078
rect 1051 -1430 1085 -1078
rect 1435 -1430 1469 -1078
rect 3571 -1430 3605 -1078
rect 3955 -1430 3989 -1078
rect 6091 -1430 6125 -1078
<< poly >>
rect -6040 1526 -4040 1542
rect -6040 1492 -6024 1526
rect -4056 1492 -4040 1526
rect -6040 1454 -4040 1492
rect -3520 1526 -1520 1542
rect -3520 1492 -3504 1526
rect -1536 1492 -1520 1526
rect -3520 1454 -1520 1492
rect -1000 1526 1000 1542
rect -1000 1492 -984 1526
rect 984 1492 1000 1526
rect -1000 1454 1000 1492
rect 1520 1526 3520 1542
rect 1520 1492 1536 1526
rect 3504 1492 3520 1526
rect 1520 1454 3520 1492
rect 4040 1526 6040 1542
rect 4040 1492 4056 1526
rect 6024 1492 6040 1526
rect 4040 1454 6040 1492
rect -6040 1016 -4040 1054
rect -6040 982 -6024 1016
rect -4056 982 -4040 1016
rect -6040 966 -4040 982
rect -3520 1016 -1520 1054
rect -3520 982 -3504 1016
rect -1536 982 -1520 1016
rect -3520 966 -1520 982
rect -1000 1016 1000 1054
rect -1000 982 -984 1016
rect 984 982 1000 1016
rect -1000 966 1000 982
rect 1520 1016 3520 1054
rect 1520 982 1536 1016
rect 3504 982 3520 1016
rect 1520 966 3520 982
rect 4040 1016 6040 1054
rect 4040 982 4056 1016
rect 6024 982 6040 1016
rect 4040 966 6040 982
rect -6040 690 -4040 706
rect -6040 656 -6024 690
rect -4056 656 -4040 690
rect -6040 618 -4040 656
rect -3520 690 -1520 706
rect -3520 656 -3504 690
rect -1536 656 -1520 690
rect -3520 618 -1520 656
rect -1000 690 1000 706
rect -1000 656 -984 690
rect 984 656 1000 690
rect -1000 618 1000 656
rect 1520 690 3520 706
rect 1520 656 1536 690
rect 3504 656 3520 690
rect 1520 618 3520 656
rect 4040 690 6040 706
rect 4040 656 4056 690
rect 6024 656 6040 690
rect 4040 618 6040 656
rect -6040 180 -4040 218
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -6040 130 -4040 146
rect -3520 180 -1520 218
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -3520 130 -1520 146
rect -1000 180 1000 218
rect -1000 146 -984 180
rect 984 146 1000 180
rect -1000 130 1000 146
rect 1520 180 3520 218
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 1520 130 3520 146
rect 4040 180 6040 218
rect 4040 146 4056 180
rect 6024 146 6040 180
rect 4040 130 6040 146
rect -6040 -146 -4040 -130
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -6040 -218 -4040 -180
rect -3520 -146 -1520 -130
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -3520 -218 -1520 -180
rect -1000 -146 1000 -130
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect -1000 -218 1000 -180
rect 1520 -146 3520 -130
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 1520 -218 3520 -180
rect 4040 -146 6040 -130
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect 4040 -218 6040 -180
rect -6040 -656 -4040 -618
rect -6040 -690 -6024 -656
rect -4056 -690 -4040 -656
rect -6040 -706 -4040 -690
rect -3520 -656 -1520 -618
rect -3520 -690 -3504 -656
rect -1536 -690 -1520 -656
rect -3520 -706 -1520 -690
rect -1000 -656 1000 -618
rect -1000 -690 -984 -656
rect 984 -690 1000 -656
rect -1000 -706 1000 -690
rect 1520 -656 3520 -618
rect 1520 -690 1536 -656
rect 3504 -690 3520 -656
rect 1520 -706 3520 -690
rect 4040 -656 6040 -618
rect 4040 -690 4056 -656
rect 6024 -690 6040 -656
rect 4040 -706 6040 -690
rect -6040 -982 -4040 -966
rect -6040 -1016 -6024 -982
rect -4056 -1016 -4040 -982
rect -6040 -1054 -4040 -1016
rect -3520 -982 -1520 -966
rect -3520 -1016 -3504 -982
rect -1536 -1016 -1520 -982
rect -3520 -1054 -1520 -1016
rect -1000 -982 1000 -966
rect -1000 -1016 -984 -982
rect 984 -1016 1000 -982
rect -1000 -1054 1000 -1016
rect 1520 -982 3520 -966
rect 1520 -1016 1536 -982
rect 3504 -1016 3520 -982
rect 1520 -1054 3520 -1016
rect 4040 -982 6040 -966
rect 4040 -1016 4056 -982
rect 6024 -1016 6040 -982
rect 4040 -1054 6040 -1016
rect -6040 -1492 -4040 -1454
rect -6040 -1526 -6024 -1492
rect -4056 -1526 -4040 -1492
rect -6040 -1542 -4040 -1526
rect -3520 -1492 -1520 -1454
rect -3520 -1526 -3504 -1492
rect -1536 -1526 -1520 -1492
rect -3520 -1542 -1520 -1526
rect -1000 -1492 1000 -1454
rect -1000 -1526 -984 -1492
rect 984 -1526 1000 -1492
rect -1000 -1542 1000 -1526
rect 1520 -1492 3520 -1454
rect 1520 -1526 1536 -1492
rect 3504 -1526 3520 -1492
rect 1520 -1542 3520 -1526
rect 4040 -1492 6040 -1454
rect 4040 -1526 4056 -1492
rect 6024 -1526 6040 -1492
rect 4040 -1542 6040 -1526
<< polycont >>
rect -6024 1492 -4056 1526
rect -3504 1492 -1536 1526
rect -984 1492 984 1526
rect 1536 1492 3504 1526
rect 4056 1492 6024 1526
rect -6024 982 -4056 1016
rect -3504 982 -1536 1016
rect -984 982 984 1016
rect 1536 982 3504 1016
rect 4056 982 6024 1016
rect -6024 656 -4056 690
rect -3504 656 -1536 690
rect -984 656 984 690
rect 1536 656 3504 690
rect 4056 656 6024 690
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6024 -690 -4056 -656
rect -3504 -690 -1536 -656
rect -984 -690 984 -656
rect 1536 -690 3504 -656
rect 4056 -690 6024 -656
rect -6024 -1016 -4056 -982
rect -3504 -1016 -1536 -982
rect -984 -1016 984 -982
rect 1536 -1016 3504 -982
rect 4056 -1016 6024 -982
rect -6024 -1526 -4056 -1492
rect -3504 -1526 -1536 -1492
rect -984 -1526 984 -1492
rect 1536 -1526 3504 -1492
rect 4056 -1526 6024 -1492
<< locali >>
rect -6247 1585 -6151 1619
rect 6151 1585 6247 1619
rect -6247 1523 -6213 1585
rect -6040 1492 -6024 1526
rect -4056 1492 -4040 1526
rect -3520 1492 -3504 1526
rect -1536 1492 -1520 1526
rect -1000 1492 -984 1526
rect 984 1492 1000 1526
rect 1520 1492 1536 1526
rect 3504 1492 3520 1526
rect 4040 1492 4056 1526
rect 6024 1492 6040 1526
rect 6213 1523 6247 1585
rect -6125 1430 -6091 1446
rect -6125 1062 -6091 1078
rect -3989 1430 -3955 1446
rect -3989 1062 -3955 1078
rect -3605 1430 -3571 1446
rect -3605 1062 -3571 1078
rect -1469 1430 -1435 1446
rect -1469 1062 -1435 1078
rect -1085 1430 -1051 1446
rect -1085 1062 -1051 1078
rect 1051 1430 1085 1446
rect 1051 1062 1085 1078
rect 1435 1430 1469 1446
rect 1435 1062 1469 1078
rect 3571 1430 3605 1446
rect 3571 1062 3605 1078
rect 3955 1430 3989 1446
rect 3955 1062 3989 1078
rect 6091 1430 6125 1446
rect 6091 1062 6125 1078
rect -6040 982 -6024 1016
rect -4056 982 -4040 1016
rect -3520 982 -3504 1016
rect -1536 982 -1520 1016
rect -1000 982 -984 1016
rect 984 982 1000 1016
rect 1520 982 1536 1016
rect 3504 982 3520 1016
rect 4040 982 4056 1016
rect 6024 982 6040 1016
rect -6040 656 -6024 690
rect -4056 656 -4040 690
rect -3520 656 -3504 690
rect -1536 656 -1520 690
rect -1000 656 -984 690
rect 984 656 1000 690
rect 1520 656 1536 690
rect 3504 656 3520 690
rect 4040 656 4056 690
rect 6024 656 6040 690
rect -6125 594 -6091 610
rect -6125 226 -6091 242
rect -3989 594 -3955 610
rect -3989 226 -3955 242
rect -3605 594 -3571 610
rect -3605 226 -3571 242
rect -1469 594 -1435 610
rect -1469 226 -1435 242
rect -1085 594 -1051 610
rect -1085 226 -1051 242
rect 1051 594 1085 610
rect 1051 226 1085 242
rect 1435 594 1469 610
rect 1435 226 1469 242
rect 3571 594 3605 610
rect 3571 226 3605 242
rect 3955 594 3989 610
rect 3955 226 3989 242
rect 6091 594 6125 610
rect 6091 226 6125 242
rect -6040 146 -6024 180
rect -4056 146 -4040 180
rect -3520 146 -3504 180
rect -1536 146 -1520 180
rect -1000 146 -984 180
rect 984 146 1000 180
rect 1520 146 1536 180
rect 3504 146 3520 180
rect 4040 146 4056 180
rect 6024 146 6040 180
rect -6040 -180 -6024 -146
rect -4056 -180 -4040 -146
rect -3520 -180 -3504 -146
rect -1536 -180 -1520 -146
rect -1000 -180 -984 -146
rect 984 -180 1000 -146
rect 1520 -180 1536 -146
rect 3504 -180 3520 -146
rect 4040 -180 4056 -146
rect 6024 -180 6040 -146
rect -6125 -242 -6091 -226
rect -6125 -610 -6091 -594
rect -3989 -242 -3955 -226
rect -3989 -610 -3955 -594
rect -3605 -242 -3571 -226
rect -3605 -610 -3571 -594
rect -1469 -242 -1435 -226
rect -1469 -610 -1435 -594
rect -1085 -242 -1051 -226
rect -1085 -610 -1051 -594
rect 1051 -242 1085 -226
rect 1051 -610 1085 -594
rect 1435 -242 1469 -226
rect 1435 -610 1469 -594
rect 3571 -242 3605 -226
rect 3571 -610 3605 -594
rect 3955 -242 3989 -226
rect 3955 -610 3989 -594
rect 6091 -242 6125 -226
rect 6091 -610 6125 -594
rect -6040 -690 -6024 -656
rect -4056 -690 -4040 -656
rect -3520 -690 -3504 -656
rect -1536 -690 -1520 -656
rect -1000 -690 -984 -656
rect 984 -690 1000 -656
rect 1520 -690 1536 -656
rect 3504 -690 3520 -656
rect 4040 -690 4056 -656
rect 6024 -690 6040 -656
rect -6040 -1016 -6024 -982
rect -4056 -1016 -4040 -982
rect -3520 -1016 -3504 -982
rect -1536 -1016 -1520 -982
rect -1000 -1016 -984 -982
rect 984 -1016 1000 -982
rect 1520 -1016 1536 -982
rect 3504 -1016 3520 -982
rect 4040 -1016 4056 -982
rect 6024 -1016 6040 -982
rect -6125 -1078 -6091 -1062
rect -6125 -1446 -6091 -1430
rect -3989 -1078 -3955 -1062
rect -3989 -1446 -3955 -1430
rect -3605 -1078 -3571 -1062
rect -3605 -1446 -3571 -1430
rect -1469 -1078 -1435 -1062
rect -1469 -1446 -1435 -1430
rect -1085 -1078 -1051 -1062
rect -1085 -1446 -1051 -1430
rect 1051 -1078 1085 -1062
rect 1051 -1446 1085 -1430
rect 1435 -1078 1469 -1062
rect 1435 -1446 1469 -1430
rect 3571 -1078 3605 -1062
rect 3571 -1446 3605 -1430
rect 3955 -1078 3989 -1062
rect 3955 -1446 3989 -1430
rect 6091 -1078 6125 -1062
rect 6091 -1446 6125 -1430
rect -6247 -1585 -6213 -1523
rect -6040 -1526 -6024 -1492
rect -4056 -1526 -4040 -1492
rect -3520 -1526 -3504 -1492
rect -1536 -1526 -1520 -1492
rect -1000 -1526 -984 -1492
rect 984 -1526 1000 -1492
rect 1520 -1526 1536 -1492
rect 3504 -1526 3520 -1492
rect 4040 -1526 4056 -1492
rect 6024 -1526 6040 -1492
rect 6213 -1585 6247 -1523
rect -6247 -1619 -6151 -1585
rect 6151 -1619 6247 -1585
<< viali >>
rect -6024 1492 -4056 1526
rect -3504 1492 -1536 1526
rect -984 1492 984 1526
rect 1536 1492 3504 1526
rect 4056 1492 6024 1526
rect -6125 1078 -6091 1430
rect -3989 1078 -3955 1430
rect -3605 1078 -3571 1430
rect -1469 1078 -1435 1430
rect -1085 1078 -1051 1430
rect 1051 1078 1085 1430
rect 1435 1078 1469 1430
rect 3571 1078 3605 1430
rect 3955 1078 3989 1430
rect 6091 1078 6125 1430
rect -6024 982 -4056 1016
rect -3504 982 -1536 1016
rect -984 982 984 1016
rect 1536 982 3504 1016
rect 4056 982 6024 1016
rect -6024 656 -4056 690
rect -3504 656 -1536 690
rect -984 656 984 690
rect 1536 656 3504 690
rect 4056 656 6024 690
rect -6125 242 -6091 594
rect -3989 242 -3955 594
rect -3605 242 -3571 594
rect -1469 242 -1435 594
rect -1085 242 -1051 594
rect 1051 242 1085 594
rect 1435 242 1469 594
rect 3571 242 3605 594
rect 3955 242 3989 594
rect 6091 242 6125 594
rect -6024 146 -4056 180
rect -3504 146 -1536 180
rect -984 146 984 180
rect 1536 146 3504 180
rect 4056 146 6024 180
rect -6024 -180 -4056 -146
rect -3504 -180 -1536 -146
rect -984 -180 984 -146
rect 1536 -180 3504 -146
rect 4056 -180 6024 -146
rect -6125 -594 -6091 -242
rect -3989 -594 -3955 -242
rect -3605 -594 -3571 -242
rect -1469 -594 -1435 -242
rect -1085 -594 -1051 -242
rect 1051 -594 1085 -242
rect 1435 -594 1469 -242
rect 3571 -594 3605 -242
rect 3955 -594 3989 -242
rect 6091 -594 6125 -242
rect -6024 -690 -4056 -656
rect -3504 -690 -1536 -656
rect -984 -690 984 -656
rect 1536 -690 3504 -656
rect 4056 -690 6024 -656
rect -6024 -1016 -4056 -982
rect -3504 -1016 -1536 -982
rect -984 -1016 984 -982
rect 1536 -1016 3504 -982
rect 4056 -1016 6024 -982
rect -6125 -1430 -6091 -1078
rect -3989 -1430 -3955 -1078
rect -3605 -1430 -3571 -1078
rect -1469 -1430 -1435 -1078
rect -1085 -1430 -1051 -1078
rect 1051 -1430 1085 -1078
rect 1435 -1430 1469 -1078
rect 3571 -1430 3605 -1078
rect 3955 -1430 3989 -1078
rect 6091 -1430 6125 -1078
rect -6024 -1526 -4056 -1492
rect -3504 -1526 -1536 -1492
rect -984 -1526 984 -1492
rect 1536 -1526 3504 -1492
rect 4056 -1526 6024 -1492
<< metal1 >>
rect -6036 1526 -4044 1532
rect -6036 1492 -6024 1526
rect -4056 1492 -4044 1526
rect -6036 1486 -4044 1492
rect -3516 1526 -1524 1532
rect -3516 1492 -3504 1526
rect -1536 1492 -1524 1526
rect -3516 1486 -1524 1492
rect -996 1526 996 1532
rect -996 1492 -984 1526
rect 984 1492 996 1526
rect -996 1486 996 1492
rect 1524 1526 3516 1532
rect 1524 1492 1536 1526
rect 3504 1492 3516 1526
rect 1524 1486 3516 1492
rect 4044 1526 6036 1532
rect 4044 1492 4056 1526
rect 6024 1492 6036 1526
rect 4044 1486 6036 1492
rect -6131 1430 -6085 1442
rect -3995 1430 -3949 1442
rect -6131 1078 -6125 1430
rect -6091 1078 -3989 1430
rect -3955 1078 -3949 1430
rect -6131 1066 -6085 1078
rect -3995 1066 -3949 1078
rect -3611 1430 -3565 1442
rect -1475 1430 -1429 1442
rect -3611 1078 -3605 1430
rect -3571 1078 -1469 1430
rect -1435 1078 -1429 1430
rect -3611 1066 -3565 1078
rect -1475 1066 -1429 1078
rect -1091 1430 -1045 1442
rect 1045 1430 1091 1442
rect -1091 1078 -1085 1430
rect -1051 1078 1051 1430
rect 1085 1078 1091 1430
rect -1091 1066 -1045 1078
rect 1045 1066 1091 1078
rect 1429 1430 1475 1442
rect 3565 1430 3611 1442
rect 1429 1078 1435 1430
rect 1469 1078 3571 1430
rect 3605 1078 3611 1430
rect 1429 1066 1475 1078
rect 3565 1066 3611 1078
rect 3949 1430 3995 1442
rect 6085 1430 6131 1442
rect 3949 1078 3955 1430
rect 3989 1078 6091 1430
rect 6125 1078 6131 1430
rect 3949 1066 3995 1078
rect 6085 1066 6131 1078
rect -6036 1016 -4044 1022
rect -6036 982 -6024 1016
rect -4056 982 -4044 1016
rect -6036 976 -4044 982
rect -3516 1016 -1524 1022
rect -3516 982 -3504 1016
rect -1536 982 -1524 1016
rect -3516 976 -1524 982
rect -996 1016 996 1022
rect -996 982 -984 1016
rect 984 982 996 1016
rect -996 976 996 982
rect 1524 1016 3516 1022
rect 1524 982 1536 1016
rect 3504 982 3516 1016
rect 1524 976 3516 982
rect 4044 1016 6036 1022
rect 4044 982 4056 1016
rect 6024 982 6036 1016
rect 4044 976 6036 982
rect -6036 690 -4044 696
rect -6036 656 -6024 690
rect -4056 656 -4044 690
rect -6036 650 -4044 656
rect -3516 690 -1524 696
rect -3516 656 -3504 690
rect -1536 656 -1524 690
rect -3516 650 -1524 656
rect -996 690 996 696
rect -996 656 -984 690
rect 984 656 996 690
rect -996 650 996 656
rect 1524 690 3516 696
rect 1524 656 1536 690
rect 3504 656 3516 690
rect 1524 650 3516 656
rect 4044 690 6036 696
rect 4044 656 4056 690
rect 6024 656 6036 690
rect 4044 650 6036 656
rect -6131 594 -6085 606
rect -3995 594 -3949 606
rect -6131 242 -6125 594
rect -6091 242 -3989 594
rect -3955 242 -3949 594
rect -6131 230 -6085 242
rect -3995 230 -3949 242
rect -3611 594 -3565 606
rect -1475 594 -1429 606
rect -3611 242 -3605 594
rect -3571 242 -1469 594
rect -1435 242 -1429 594
rect -3611 230 -3565 242
rect -1475 230 -1429 242
rect -1091 594 -1045 606
rect 1045 594 1091 606
rect -1091 242 -1085 594
rect -1051 242 1051 594
rect 1085 242 1091 594
rect -1091 230 -1045 242
rect 1045 230 1091 242
rect 1429 594 1475 606
rect 3565 594 3611 606
rect 1429 242 1435 594
rect 1469 242 3571 594
rect 3605 242 3611 594
rect 1429 230 1475 242
rect 3565 230 3611 242
rect 3949 594 3995 606
rect 6085 594 6131 606
rect 3949 242 3955 594
rect 3989 242 6091 594
rect 6125 242 6131 594
rect 3949 230 3995 242
rect 6085 230 6131 242
rect -6036 180 -4044 186
rect -6036 146 -6024 180
rect -4056 146 -4044 180
rect -6036 140 -4044 146
rect -3516 180 -1524 186
rect -3516 146 -3504 180
rect -1536 146 -1524 180
rect -3516 140 -1524 146
rect -996 180 996 186
rect -996 146 -984 180
rect 984 146 996 180
rect -996 140 996 146
rect 1524 180 3516 186
rect 1524 146 1536 180
rect 3504 146 3516 180
rect 1524 140 3516 146
rect 4044 180 6036 186
rect 4044 146 4056 180
rect 6024 146 6036 180
rect 4044 140 6036 146
rect -6036 -146 -4044 -140
rect -6036 -180 -6024 -146
rect -4056 -180 -4044 -146
rect -6036 -186 -4044 -180
rect -3516 -146 -1524 -140
rect -3516 -180 -3504 -146
rect -1536 -180 -1524 -146
rect -3516 -186 -1524 -180
rect -996 -146 996 -140
rect -996 -180 -984 -146
rect 984 -180 996 -146
rect -996 -186 996 -180
rect 1524 -146 3516 -140
rect 1524 -180 1536 -146
rect 3504 -180 3516 -146
rect 1524 -186 3516 -180
rect 4044 -146 6036 -140
rect 4044 -180 4056 -146
rect 6024 -180 6036 -146
rect 4044 -186 6036 -180
rect -6131 -242 -6085 -230
rect -3995 -242 -3949 -230
rect -6131 -594 -6125 -242
rect -6091 -594 -3989 -242
rect -3955 -594 -3949 -242
rect -6131 -606 -6085 -594
rect -3995 -606 -3949 -594
rect -3611 -242 -3565 -230
rect -1475 -242 -1429 -230
rect -3611 -594 -3605 -242
rect -3571 -594 -1469 -242
rect -1435 -594 -1429 -242
rect -3611 -606 -3565 -594
rect -1475 -606 -1429 -594
rect -1091 -242 -1045 -230
rect 1045 -242 1091 -230
rect -1091 -594 -1085 -242
rect -1051 -594 1051 -242
rect 1085 -594 1091 -242
rect -1091 -606 -1045 -594
rect 1045 -606 1091 -594
rect 1429 -242 1475 -230
rect 3565 -242 3611 -230
rect 1429 -594 1435 -242
rect 1469 -594 3571 -242
rect 3605 -594 3611 -242
rect 1429 -606 1475 -594
rect 3565 -606 3611 -594
rect 3949 -242 3995 -230
rect 6085 -242 6131 -230
rect 3949 -594 3955 -242
rect 3989 -594 6091 -242
rect 6125 -594 6131 -242
rect 3949 -606 3995 -594
rect 6085 -606 6131 -594
rect -6036 -656 -4044 -650
rect -6036 -690 -6024 -656
rect -4056 -690 -4044 -656
rect -6036 -696 -4044 -690
rect -3516 -656 -1524 -650
rect -3516 -690 -3504 -656
rect -1536 -690 -1524 -656
rect -3516 -696 -1524 -690
rect -996 -656 996 -650
rect -996 -690 -984 -656
rect 984 -690 996 -656
rect -996 -696 996 -690
rect 1524 -656 3516 -650
rect 1524 -690 1536 -656
rect 3504 -690 3516 -656
rect 1524 -696 3516 -690
rect 4044 -656 6036 -650
rect 4044 -690 4056 -656
rect 6024 -690 6036 -656
rect 4044 -696 6036 -690
rect -6036 -982 -4044 -976
rect -6036 -1016 -6024 -982
rect -4056 -1016 -4044 -982
rect -6036 -1022 -4044 -1016
rect -3516 -982 -1524 -976
rect -3516 -1016 -3504 -982
rect -1536 -1016 -1524 -982
rect -3516 -1022 -1524 -1016
rect -996 -982 996 -976
rect -996 -1016 -984 -982
rect 984 -1016 996 -982
rect -996 -1022 996 -1016
rect 1524 -982 3516 -976
rect 1524 -1016 1536 -982
rect 3504 -1016 3516 -982
rect 1524 -1022 3516 -1016
rect 4044 -982 6036 -976
rect 4044 -1016 4056 -982
rect 6024 -1016 6036 -982
rect 4044 -1022 6036 -1016
rect -6131 -1078 -6085 -1066
rect -3995 -1078 -3949 -1066
rect -6131 -1430 -6125 -1078
rect -6091 -1430 -3989 -1078
rect -3955 -1430 -3949 -1078
rect -6131 -1442 -6085 -1430
rect -3995 -1442 -3949 -1430
rect -3611 -1078 -3565 -1066
rect -1475 -1078 -1429 -1066
rect -3611 -1430 -3605 -1078
rect -3571 -1430 -1469 -1078
rect -1435 -1430 -1429 -1078
rect -3611 -1442 -3565 -1430
rect -1475 -1442 -1429 -1430
rect -1091 -1078 -1045 -1066
rect 1045 -1078 1091 -1066
rect -1091 -1430 -1085 -1078
rect -1051 -1430 1051 -1078
rect 1085 -1430 1091 -1078
rect -1091 -1442 -1045 -1430
rect 1045 -1442 1091 -1430
rect 1429 -1078 1475 -1066
rect 3565 -1078 3611 -1066
rect 1429 -1430 1435 -1078
rect 1469 -1430 3571 -1078
rect 3605 -1430 3611 -1078
rect 1429 -1442 1475 -1430
rect 3565 -1442 3611 -1430
rect 3949 -1078 3995 -1066
rect 6085 -1078 6131 -1066
rect 3949 -1430 3955 -1078
rect 3989 -1430 6091 -1078
rect 6125 -1430 6131 -1078
rect 3949 -1442 3995 -1430
rect 6085 -1442 6131 -1430
rect -6036 -1492 -4044 -1486
rect -6036 -1526 -6024 -1492
rect -4056 -1526 -4044 -1492
rect -6036 -1532 -4044 -1526
rect -3516 -1492 -1524 -1486
rect -3516 -1526 -3504 -1492
rect -1536 -1526 -1524 -1492
rect -3516 -1532 -1524 -1526
rect -996 -1492 996 -1486
rect -996 -1526 -984 -1492
rect 984 -1526 996 -1492
rect -996 -1532 996 -1526
rect 1524 -1492 3516 -1486
rect 1524 -1526 1536 -1492
rect 3504 -1526 3516 -1492
rect 1524 -1532 3516 -1526
rect 4044 -1492 6036 -1486
rect 4044 -1526 4056 -1492
rect 6024 -1526 6036 -1492
rect 4044 -1532 6036 -1526
<< properties >>
string FIXED_BBOX -6230 -1602 6230 1602
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 10 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
