magic
tech sky130A
magscale 1 2
timestamp 1683728594
<< nwell >>
rect 2300 800 4554 2274
<< pwell >>
rect -240 280 2264 2276
rect -20 -1820 2234 236
rect 2300 -760 4554 678
rect -2600 -4200 -1306 -2144
rect -800 -4200 494 -2144
rect 1000 -4200 2294 -2144
rect 2800 -4200 4094 -2144
rect 4800 -3520 7054 2244
rect -2600 -8200 -976 -4290
rect -800 -8200 824 -4290
rect 1000 -8200 2624 -4290
rect 2800 -8200 4424 -4290
<< pmos >>
rect 2500 1655 2530 2055
rect 2596 1655 2626 2055
rect 2692 1655 2722 2055
rect 2788 1655 2818 2055
rect 2884 1655 2914 2055
rect 2980 1655 3010 2055
rect 3076 1655 3106 2055
rect 3172 1655 3202 2055
rect 3268 1655 3298 2055
rect 3364 1655 3394 2055
rect 3460 1655 3490 2055
rect 3556 1655 3586 2055
rect 3652 1655 3682 2055
rect 3748 1655 3778 2055
rect 3844 1655 3874 2055
rect 3940 1655 3970 2055
rect 4036 1655 4066 2055
rect 4132 1655 4162 2055
rect 4228 1655 4258 2055
rect 4324 1655 4354 2055
rect 2500 1019 2530 1419
rect 2596 1019 2626 1419
rect 2692 1019 2722 1419
rect 2788 1019 2818 1419
rect 2884 1019 2914 1419
rect 2980 1019 3010 1419
rect 3076 1019 3106 1419
rect 3172 1019 3202 1419
rect 3268 1019 3298 1419
rect 3364 1019 3394 1419
rect 3460 1019 3490 1419
rect 3556 1019 3586 1419
rect 3652 1019 3682 1419
rect 3748 1019 3778 1419
rect 3844 1019 3874 1419
rect 3940 1019 3970 1419
rect 4036 1019 4066 1419
rect 4132 1019 4162 1419
rect 4228 1019 4258 1419
rect 4324 1019 4354 1419
<< nmoslvt >>
rect 180 -374 210 26
rect 276 -374 306 26
rect 372 -374 402 26
rect 468 -374 498 26
rect 564 -374 594 26
rect 660 -374 690 26
rect 756 -374 786 26
rect 852 -374 882 26
rect 948 -374 978 26
rect 1044 -374 1074 26
rect 1140 -374 1170 26
rect 1236 -374 1266 26
rect 1332 -374 1362 26
rect 1428 -374 1458 26
rect 1524 -374 1554 26
rect 1620 -374 1650 26
rect 1716 -374 1746 26
rect 1812 -374 1842 26
rect 1908 -374 1938 26
rect 2004 -374 2034 26
rect 180 -992 210 -592
rect 276 -992 306 -592
rect 372 -992 402 -592
rect 468 -992 498 -592
rect 564 -992 594 -592
rect 660 -992 690 -592
rect 756 -992 786 -592
rect 852 -992 882 -592
rect 948 -992 978 -592
rect 1044 -992 1074 -592
rect 1140 -992 1170 -592
rect 1236 -992 1266 -592
rect 1332 -992 1362 -592
rect 1428 -992 1458 -592
rect 1524 -992 1554 -592
rect 1620 -992 1650 -592
rect 1716 -992 1746 -592
rect 1812 -992 1842 -592
rect 1908 -992 1938 -592
rect 2004 -992 2034 -592
rect 180 -1610 210 -1210
rect 276 -1610 306 -1210
rect 372 -1610 402 -1210
rect 468 -1610 498 -1210
rect 564 -1610 594 -1210
rect 660 -1610 690 -1210
rect 756 -1610 786 -1210
rect 852 -1610 882 -1210
rect 948 -1610 978 -1210
rect 1044 -1610 1074 -1210
rect 1140 -1610 1170 -1210
rect 1236 -1610 1266 -1210
rect 1332 -1610 1362 -1210
rect 1428 -1610 1458 -1210
rect 1524 -1610 1554 -1210
rect 1620 -1610 1650 -1210
rect 1716 -1610 1746 -1210
rect 1812 -1610 1842 -1210
rect 1908 -1610 1938 -1210
rect 2004 -1610 2034 -1210
rect 2500 68 2530 468
rect 2596 68 2626 468
rect 2692 68 2722 468
rect 2788 68 2818 468
rect 2884 68 2914 468
rect 2980 68 3010 468
rect 3076 68 3106 468
rect 3172 68 3202 468
rect 3268 68 3298 468
rect 3364 68 3394 468
rect 3460 68 3490 468
rect 3556 68 3586 468
rect 3652 68 3682 468
rect 3748 68 3778 468
rect 3844 68 3874 468
rect 3940 68 3970 468
rect 4036 68 4066 468
rect 4132 68 4162 468
rect 4228 68 4258 468
rect 4324 68 4354 468
rect 2500 -550 2530 -150
rect 2596 -550 2626 -150
rect 2692 -550 2722 -150
rect 2788 -550 2818 -150
rect 2884 -550 2914 -150
rect 2980 -550 3010 -150
rect 3076 -550 3106 -150
rect 3172 -550 3202 -150
rect 3268 -550 3298 -150
rect 3364 -550 3394 -150
rect 3460 -550 3490 -150
rect 3556 -550 3586 -150
rect 3652 -550 3682 -150
rect 3748 -550 3778 -150
rect 3844 -550 3874 -150
rect 3940 -550 3970 -150
rect 4036 -550 4066 -150
rect 4132 -550 4162 -150
rect 4228 -550 4258 -150
rect 4324 -550 4354 -150
rect -2400 -2754 -2370 -2354
rect -2304 -2754 -2274 -2354
rect -2208 -2754 -2178 -2354
rect -2112 -2754 -2082 -2354
rect -2016 -2754 -1986 -2354
rect -1920 -2754 -1890 -2354
rect -1824 -2754 -1794 -2354
rect -1728 -2754 -1698 -2354
rect -1632 -2754 -1602 -2354
rect -1536 -2754 -1506 -2354
rect -2400 -3372 -2370 -2972
rect -2304 -3372 -2274 -2972
rect -2208 -3372 -2178 -2972
rect -2112 -3372 -2082 -2972
rect -2016 -3372 -1986 -2972
rect -1920 -3372 -1890 -2972
rect -1824 -3372 -1794 -2972
rect -1728 -3372 -1698 -2972
rect -1632 -3372 -1602 -2972
rect -1536 -3372 -1506 -2972
rect -2400 -3990 -2370 -3590
rect -2304 -3990 -2274 -3590
rect -2208 -3990 -2178 -3590
rect -2112 -3990 -2082 -3590
rect -2016 -3990 -1986 -3590
rect -1920 -3990 -1890 -3590
rect -1824 -3990 -1794 -3590
rect -1728 -3990 -1698 -3590
rect -1632 -3990 -1602 -3590
rect -1536 -3990 -1506 -3590
rect -600 -2754 -570 -2354
rect -504 -2754 -474 -2354
rect -408 -2754 -378 -2354
rect -312 -2754 -282 -2354
rect -216 -2754 -186 -2354
rect -120 -2754 -90 -2354
rect -24 -2754 6 -2354
rect 72 -2754 102 -2354
rect 168 -2754 198 -2354
rect 264 -2754 294 -2354
rect -600 -3372 -570 -2972
rect -504 -3372 -474 -2972
rect -408 -3372 -378 -2972
rect -312 -3372 -282 -2972
rect -216 -3372 -186 -2972
rect -120 -3372 -90 -2972
rect -24 -3372 6 -2972
rect 72 -3372 102 -2972
rect 168 -3372 198 -2972
rect 264 -3372 294 -2972
rect -600 -3990 -570 -3590
rect -504 -3990 -474 -3590
rect -408 -3990 -378 -3590
rect -312 -3990 -282 -3590
rect -216 -3990 -186 -3590
rect -120 -3990 -90 -3590
rect -24 -3990 6 -3590
rect 72 -3990 102 -3590
rect 168 -3990 198 -3590
rect 264 -3990 294 -3590
rect 1200 -2754 1230 -2354
rect 1296 -2754 1326 -2354
rect 1392 -2754 1422 -2354
rect 1488 -2754 1518 -2354
rect 1584 -2754 1614 -2354
rect 1680 -2754 1710 -2354
rect 1776 -2754 1806 -2354
rect 1872 -2754 1902 -2354
rect 1968 -2754 1998 -2354
rect 2064 -2754 2094 -2354
rect 1200 -3372 1230 -2972
rect 1296 -3372 1326 -2972
rect 1392 -3372 1422 -2972
rect 1488 -3372 1518 -2972
rect 1584 -3372 1614 -2972
rect 1680 -3372 1710 -2972
rect 1776 -3372 1806 -2972
rect 1872 -3372 1902 -2972
rect 1968 -3372 1998 -2972
rect 2064 -3372 2094 -2972
rect 1200 -3990 1230 -3590
rect 1296 -3990 1326 -3590
rect 1392 -3990 1422 -3590
rect 1488 -3990 1518 -3590
rect 1584 -3990 1614 -3590
rect 1680 -3990 1710 -3590
rect 1776 -3990 1806 -3590
rect 1872 -3990 1902 -3590
rect 1968 -3990 1998 -3590
rect 2064 -3990 2094 -3590
rect 3000 -2754 3030 -2354
rect 3096 -2754 3126 -2354
rect 3192 -2754 3222 -2354
rect 3288 -2754 3318 -2354
rect 3384 -2754 3414 -2354
rect 3480 -2754 3510 -2354
rect 3576 -2754 3606 -2354
rect 3672 -2754 3702 -2354
rect 3768 -2754 3798 -2354
rect 3864 -2754 3894 -2354
rect 3000 -3372 3030 -2972
rect 3096 -3372 3126 -2972
rect 3192 -3372 3222 -2972
rect 3288 -3372 3318 -2972
rect 3384 -3372 3414 -2972
rect 3480 -3372 3510 -2972
rect 3576 -3372 3606 -2972
rect 3672 -3372 3702 -2972
rect 3768 -3372 3798 -2972
rect 3864 -3372 3894 -2972
rect 3000 -3990 3030 -3590
rect 3096 -3990 3126 -3590
rect 3192 -3990 3222 -3590
rect 3288 -3990 3318 -3590
rect 3384 -3990 3414 -3590
rect 3480 -3990 3510 -3590
rect 3576 -3990 3606 -3590
rect 3672 -3990 3702 -3590
rect 3768 -3990 3798 -3590
rect 3864 -3990 3894 -3590
rect 5000 1634 5030 2034
rect 5096 1634 5126 2034
rect 5192 1634 5222 2034
rect 5288 1634 5318 2034
rect 5384 1634 5414 2034
rect 5480 1634 5510 2034
rect 5576 1634 5606 2034
rect 5672 1634 5702 2034
rect 5768 1634 5798 2034
rect 5864 1634 5894 2034
rect 5960 1634 5990 2034
rect 6056 1634 6086 2034
rect 6152 1634 6182 2034
rect 6248 1634 6278 2034
rect 6344 1634 6374 2034
rect 6440 1634 6470 2034
rect 6536 1634 6566 2034
rect 6632 1634 6662 2034
rect 6728 1634 6758 2034
rect 6824 1634 6854 2034
rect 5000 1016 5030 1416
rect 5096 1016 5126 1416
rect 5192 1016 5222 1416
rect 5288 1016 5318 1416
rect 5384 1016 5414 1416
rect 5480 1016 5510 1416
rect 5576 1016 5606 1416
rect 5672 1016 5702 1416
rect 5768 1016 5798 1416
rect 5864 1016 5894 1416
rect 5960 1016 5990 1416
rect 6056 1016 6086 1416
rect 6152 1016 6182 1416
rect 6248 1016 6278 1416
rect 6344 1016 6374 1416
rect 6440 1016 6470 1416
rect 6536 1016 6566 1416
rect 6632 1016 6662 1416
rect 6728 1016 6758 1416
rect 6824 1016 6854 1416
rect 5000 398 5030 798
rect 5096 398 5126 798
rect 5192 398 5222 798
rect 5288 398 5318 798
rect 5384 398 5414 798
rect 5480 398 5510 798
rect 5576 398 5606 798
rect 5672 398 5702 798
rect 5768 398 5798 798
rect 5864 398 5894 798
rect 5960 398 5990 798
rect 6056 398 6086 798
rect 6152 398 6182 798
rect 6248 398 6278 798
rect 6344 398 6374 798
rect 6440 398 6470 798
rect 6536 398 6566 798
rect 6632 398 6662 798
rect 6728 398 6758 798
rect 6824 398 6854 798
rect 5000 -220 5030 180
rect 5096 -220 5126 180
rect 5192 -220 5222 180
rect 5288 -220 5318 180
rect 5384 -220 5414 180
rect 5480 -220 5510 180
rect 5576 -220 5606 180
rect 5672 -220 5702 180
rect 5768 -220 5798 180
rect 5864 -220 5894 180
rect 5960 -220 5990 180
rect 6056 -220 6086 180
rect 6152 -220 6182 180
rect 6248 -220 6278 180
rect 6344 -220 6374 180
rect 6440 -220 6470 180
rect 6536 -220 6566 180
rect 6632 -220 6662 180
rect 6728 -220 6758 180
rect 6824 -220 6854 180
rect 5000 -838 5030 -438
rect 5096 -838 5126 -438
rect 5192 -838 5222 -438
rect 5288 -838 5318 -438
rect 5384 -838 5414 -438
rect 5480 -838 5510 -438
rect 5576 -838 5606 -438
rect 5672 -838 5702 -438
rect 5768 -838 5798 -438
rect 5864 -838 5894 -438
rect 5960 -838 5990 -438
rect 6056 -838 6086 -438
rect 6152 -838 6182 -438
rect 6248 -838 6278 -438
rect 6344 -838 6374 -438
rect 6440 -838 6470 -438
rect 6536 -838 6566 -438
rect 6632 -838 6662 -438
rect 6728 -838 6758 -438
rect 6824 -838 6854 -438
rect 5000 -1456 5030 -1056
rect 5096 -1456 5126 -1056
rect 5192 -1456 5222 -1056
rect 5288 -1456 5318 -1056
rect 5384 -1456 5414 -1056
rect 5480 -1456 5510 -1056
rect 5576 -1456 5606 -1056
rect 5672 -1456 5702 -1056
rect 5768 -1456 5798 -1056
rect 5864 -1456 5894 -1056
rect 5960 -1456 5990 -1056
rect 6056 -1456 6086 -1056
rect 6152 -1456 6182 -1056
rect 6248 -1456 6278 -1056
rect 6344 -1456 6374 -1056
rect 6440 -1456 6470 -1056
rect 6536 -1456 6566 -1056
rect 6632 -1456 6662 -1056
rect 6728 -1456 6758 -1056
rect 6824 -1456 6854 -1056
rect 5000 -2074 5030 -1674
rect 5096 -2074 5126 -1674
rect 5192 -2074 5222 -1674
rect 5288 -2074 5318 -1674
rect 5384 -2074 5414 -1674
rect 5480 -2074 5510 -1674
rect 5576 -2074 5606 -1674
rect 5672 -2074 5702 -1674
rect 5768 -2074 5798 -1674
rect 5864 -2074 5894 -1674
rect 5960 -2074 5990 -1674
rect 6056 -2074 6086 -1674
rect 6152 -2074 6182 -1674
rect 6248 -2074 6278 -1674
rect 6344 -2074 6374 -1674
rect 6440 -2074 6470 -1674
rect 6536 -2074 6566 -1674
rect 6632 -2074 6662 -1674
rect 6728 -2074 6758 -1674
rect 6824 -2074 6854 -1674
rect 5000 -2692 5030 -2292
rect 5096 -2692 5126 -2292
rect 5192 -2692 5222 -2292
rect 5288 -2692 5318 -2292
rect 5384 -2692 5414 -2292
rect 5480 -2692 5510 -2292
rect 5576 -2692 5606 -2292
rect 5672 -2692 5702 -2292
rect 5768 -2692 5798 -2292
rect 5864 -2692 5894 -2292
rect 5960 -2692 5990 -2292
rect 6056 -2692 6086 -2292
rect 6152 -2692 6182 -2292
rect 6248 -2692 6278 -2292
rect 6344 -2692 6374 -2292
rect 6440 -2692 6470 -2292
rect 6536 -2692 6566 -2292
rect 6632 -2692 6662 -2292
rect 6728 -2692 6758 -2292
rect 6824 -2692 6854 -2292
rect 5000 -3310 5030 -2910
rect 5096 -3310 5126 -2910
rect 5192 -3310 5222 -2910
rect 5288 -3310 5318 -2910
rect 5384 -3310 5414 -2910
rect 5480 -3310 5510 -2910
rect 5576 -3310 5606 -2910
rect 5672 -3310 5702 -2910
rect 5768 -3310 5798 -2910
rect 5864 -3310 5894 -2910
rect 5960 -3310 5990 -2910
rect 6056 -3310 6086 -2910
rect 6152 -3310 6182 -2910
rect 6248 -3310 6278 -2910
rect 6344 -3310 6374 -2910
rect 6440 -3310 6470 -2910
rect 6536 -3310 6566 -2910
rect 6632 -3310 6662 -2910
rect 6728 -3310 6758 -2910
rect 6824 -3310 6854 -2910
rect -2404 -4900 -2204 -4500
rect -2146 -4900 -1946 -4500
rect -1888 -4900 -1688 -4500
rect -1630 -4900 -1430 -4500
rect -1372 -4900 -1172 -4500
rect -2404 -5518 -2204 -5118
rect -2146 -5518 -1946 -5118
rect -1888 -5518 -1688 -5118
rect -1630 -5518 -1430 -5118
rect -1372 -5518 -1172 -5118
rect -2404 -6136 -2204 -5736
rect -2146 -6136 -1946 -5736
rect -1888 -6136 -1688 -5736
rect -1630 -6136 -1430 -5736
rect -1372 -6136 -1172 -5736
rect -2404 -6754 -2204 -6354
rect -2146 -6754 -1946 -6354
rect -1888 -6754 -1688 -6354
rect -1630 -6754 -1430 -6354
rect -1372 -6754 -1172 -6354
rect -2404 -7372 -2204 -6972
rect -2146 -7372 -1946 -6972
rect -1888 -7372 -1688 -6972
rect -1630 -7372 -1430 -6972
rect -1372 -7372 -1172 -6972
rect -2404 -7990 -2204 -7590
rect -2146 -7990 -1946 -7590
rect -1888 -7990 -1688 -7590
rect -1630 -7990 -1430 -7590
rect -1372 -7990 -1172 -7590
rect -604 -4900 -404 -4500
rect -346 -4900 -146 -4500
rect -88 -4900 112 -4500
rect 170 -4900 370 -4500
rect 428 -4900 628 -4500
rect -604 -5518 -404 -5118
rect -346 -5518 -146 -5118
rect -88 -5518 112 -5118
rect 170 -5518 370 -5118
rect 428 -5518 628 -5118
rect -604 -6136 -404 -5736
rect -346 -6136 -146 -5736
rect -88 -6136 112 -5736
rect 170 -6136 370 -5736
rect 428 -6136 628 -5736
rect -604 -6754 -404 -6354
rect -346 -6754 -146 -6354
rect -88 -6754 112 -6354
rect 170 -6754 370 -6354
rect 428 -6754 628 -6354
rect -604 -7372 -404 -6972
rect -346 -7372 -146 -6972
rect -88 -7372 112 -6972
rect 170 -7372 370 -6972
rect 428 -7372 628 -6972
rect -604 -7990 -404 -7590
rect -346 -7990 -146 -7590
rect -88 -7990 112 -7590
rect 170 -7990 370 -7590
rect 428 -7990 628 -7590
rect 1196 -4900 1396 -4500
rect 1454 -4900 1654 -4500
rect 1712 -4900 1912 -4500
rect 1970 -4900 2170 -4500
rect 2228 -4900 2428 -4500
rect 1196 -5518 1396 -5118
rect 1454 -5518 1654 -5118
rect 1712 -5518 1912 -5118
rect 1970 -5518 2170 -5118
rect 2228 -5518 2428 -5118
rect 1196 -6136 1396 -5736
rect 1454 -6136 1654 -5736
rect 1712 -6136 1912 -5736
rect 1970 -6136 2170 -5736
rect 2228 -6136 2428 -5736
rect 1196 -6754 1396 -6354
rect 1454 -6754 1654 -6354
rect 1712 -6754 1912 -6354
rect 1970 -6754 2170 -6354
rect 2228 -6754 2428 -6354
rect 1196 -7372 1396 -6972
rect 1454 -7372 1654 -6972
rect 1712 -7372 1912 -6972
rect 1970 -7372 2170 -6972
rect 2228 -7372 2428 -6972
rect 1196 -7990 1396 -7590
rect 1454 -7990 1654 -7590
rect 1712 -7990 1912 -7590
rect 1970 -7990 2170 -7590
rect 2228 -7990 2428 -7590
rect 2996 -4900 3196 -4500
rect 3254 -4900 3454 -4500
rect 3512 -4900 3712 -4500
rect 3770 -4900 3970 -4500
rect 4028 -4900 4228 -4500
rect 2996 -5518 3196 -5118
rect 3254 -5518 3454 -5118
rect 3512 -5518 3712 -5118
rect 3770 -5518 3970 -5118
rect 4028 -5518 4228 -5118
rect 2996 -6136 3196 -5736
rect 3254 -6136 3454 -5736
rect 3512 -6136 3712 -5736
rect 3770 -6136 3970 -5736
rect 4028 -6136 4228 -5736
rect 2996 -6754 3196 -6354
rect 3254 -6754 3454 -6354
rect 3512 -6754 3712 -6354
rect 3770 -6754 3970 -6354
rect 4028 -6754 4228 -6354
rect 2996 -7372 3196 -6972
rect 3254 -7372 3454 -6972
rect 3512 -7372 3712 -6972
rect 3770 -7372 3970 -6972
rect 4028 -7372 4228 -6972
rect 2996 -7990 3196 -7590
rect 3254 -7990 3454 -7590
rect 3512 -7990 3712 -7590
rect 3770 -7990 3970 -7590
rect 4028 -7990 4228 -7590
<< ndiff >>
rect 118 14 180 26
rect 118 -362 130 14
rect 164 -362 180 14
rect 118 -374 180 -362
rect 210 14 276 26
rect 210 -362 226 14
rect 260 -362 276 14
rect 210 -374 276 -362
rect 306 14 372 26
rect 306 -362 322 14
rect 356 -362 372 14
rect 306 -374 372 -362
rect 402 14 468 26
rect 402 -362 418 14
rect 452 -362 468 14
rect 402 -374 468 -362
rect 498 14 564 26
rect 498 -362 514 14
rect 548 -362 564 14
rect 498 -374 564 -362
rect 594 14 660 26
rect 594 -362 610 14
rect 644 -362 660 14
rect 594 -374 660 -362
rect 690 14 756 26
rect 690 -362 706 14
rect 740 -362 756 14
rect 690 -374 756 -362
rect 786 14 852 26
rect 786 -362 802 14
rect 836 -362 852 14
rect 786 -374 852 -362
rect 882 14 948 26
rect 882 -362 898 14
rect 932 -362 948 14
rect 882 -374 948 -362
rect 978 14 1044 26
rect 978 -362 994 14
rect 1028 -362 1044 14
rect 978 -374 1044 -362
rect 1074 14 1140 26
rect 1074 -362 1090 14
rect 1124 -362 1140 14
rect 1074 -374 1140 -362
rect 1170 14 1236 26
rect 1170 -362 1186 14
rect 1220 -362 1236 14
rect 1170 -374 1236 -362
rect 1266 14 1332 26
rect 1266 -362 1282 14
rect 1316 -362 1332 14
rect 1266 -374 1332 -362
rect 1362 14 1428 26
rect 1362 -362 1378 14
rect 1412 -362 1428 14
rect 1362 -374 1428 -362
rect 1458 14 1524 26
rect 1458 -362 1474 14
rect 1508 -362 1524 14
rect 1458 -374 1524 -362
rect 1554 14 1620 26
rect 1554 -362 1570 14
rect 1604 -362 1620 14
rect 1554 -374 1620 -362
rect 1650 14 1716 26
rect 1650 -362 1666 14
rect 1700 -362 1716 14
rect 1650 -374 1716 -362
rect 1746 14 1812 26
rect 1746 -362 1762 14
rect 1796 -362 1812 14
rect 1746 -374 1812 -362
rect 1842 14 1908 26
rect 1842 -362 1858 14
rect 1892 -362 1908 14
rect 1842 -374 1908 -362
rect 1938 14 2004 26
rect 1938 -362 1954 14
rect 1988 -362 2004 14
rect 1938 -374 2004 -362
rect 2034 14 2096 26
rect 2034 -362 2050 14
rect 2084 -362 2096 14
rect 2034 -374 2096 -362
rect 118 -604 180 -592
rect 118 -980 130 -604
rect 164 -980 180 -604
rect 118 -992 180 -980
rect 210 -604 276 -592
rect 210 -980 226 -604
rect 260 -980 276 -604
rect 210 -992 276 -980
rect 306 -604 372 -592
rect 306 -980 322 -604
rect 356 -980 372 -604
rect 306 -992 372 -980
rect 402 -604 468 -592
rect 402 -980 418 -604
rect 452 -980 468 -604
rect 402 -992 468 -980
rect 498 -604 564 -592
rect 498 -980 514 -604
rect 548 -980 564 -604
rect 498 -992 564 -980
rect 594 -604 660 -592
rect 594 -980 610 -604
rect 644 -980 660 -604
rect 594 -992 660 -980
rect 690 -604 756 -592
rect 690 -980 706 -604
rect 740 -980 756 -604
rect 690 -992 756 -980
rect 786 -604 852 -592
rect 786 -980 802 -604
rect 836 -980 852 -604
rect 786 -992 852 -980
rect 882 -604 948 -592
rect 882 -980 898 -604
rect 932 -980 948 -604
rect 882 -992 948 -980
rect 978 -604 1044 -592
rect 978 -980 994 -604
rect 1028 -980 1044 -604
rect 978 -992 1044 -980
rect 1074 -604 1140 -592
rect 1074 -980 1090 -604
rect 1124 -980 1140 -604
rect 1074 -992 1140 -980
rect 1170 -604 1236 -592
rect 1170 -980 1186 -604
rect 1220 -980 1236 -604
rect 1170 -992 1236 -980
rect 1266 -604 1332 -592
rect 1266 -980 1282 -604
rect 1316 -980 1332 -604
rect 1266 -992 1332 -980
rect 1362 -604 1428 -592
rect 1362 -980 1378 -604
rect 1412 -980 1428 -604
rect 1362 -992 1428 -980
rect 1458 -604 1524 -592
rect 1458 -980 1474 -604
rect 1508 -980 1524 -604
rect 1458 -992 1524 -980
rect 1554 -604 1620 -592
rect 1554 -980 1570 -604
rect 1604 -980 1620 -604
rect 1554 -992 1620 -980
rect 1650 -604 1716 -592
rect 1650 -980 1666 -604
rect 1700 -980 1716 -604
rect 1650 -992 1716 -980
rect 1746 -604 1812 -592
rect 1746 -980 1762 -604
rect 1796 -980 1812 -604
rect 1746 -992 1812 -980
rect 1842 -604 1908 -592
rect 1842 -980 1858 -604
rect 1892 -980 1908 -604
rect 1842 -992 1908 -980
rect 1938 -604 2004 -592
rect 1938 -980 1954 -604
rect 1988 -980 2004 -604
rect 1938 -992 2004 -980
rect 2034 -604 2096 -592
rect 2034 -980 2050 -604
rect 2084 -980 2096 -604
rect 2034 -992 2096 -980
rect 118 -1222 180 -1210
rect 118 -1598 130 -1222
rect 164 -1598 180 -1222
rect 118 -1610 180 -1598
rect 210 -1222 276 -1210
rect 210 -1598 226 -1222
rect 260 -1598 276 -1222
rect 210 -1610 276 -1598
rect 306 -1222 372 -1210
rect 306 -1598 322 -1222
rect 356 -1598 372 -1222
rect 306 -1610 372 -1598
rect 402 -1222 468 -1210
rect 402 -1598 418 -1222
rect 452 -1598 468 -1222
rect 402 -1610 468 -1598
rect 498 -1222 564 -1210
rect 498 -1598 514 -1222
rect 548 -1598 564 -1222
rect 498 -1610 564 -1598
rect 594 -1222 660 -1210
rect 594 -1598 610 -1222
rect 644 -1598 660 -1222
rect 594 -1610 660 -1598
rect 690 -1222 756 -1210
rect 690 -1598 706 -1222
rect 740 -1598 756 -1222
rect 690 -1610 756 -1598
rect 786 -1222 852 -1210
rect 786 -1598 802 -1222
rect 836 -1598 852 -1222
rect 786 -1610 852 -1598
rect 882 -1222 948 -1210
rect 882 -1598 898 -1222
rect 932 -1598 948 -1222
rect 882 -1610 948 -1598
rect 978 -1222 1044 -1210
rect 978 -1598 994 -1222
rect 1028 -1598 1044 -1222
rect 978 -1610 1044 -1598
rect 1074 -1222 1140 -1210
rect 1074 -1598 1090 -1222
rect 1124 -1598 1140 -1222
rect 1074 -1610 1140 -1598
rect 1170 -1222 1236 -1210
rect 1170 -1598 1186 -1222
rect 1220 -1598 1236 -1222
rect 1170 -1610 1236 -1598
rect 1266 -1222 1332 -1210
rect 1266 -1598 1282 -1222
rect 1316 -1598 1332 -1222
rect 1266 -1610 1332 -1598
rect 1362 -1222 1428 -1210
rect 1362 -1598 1378 -1222
rect 1412 -1598 1428 -1222
rect 1362 -1610 1428 -1598
rect 1458 -1222 1524 -1210
rect 1458 -1598 1474 -1222
rect 1508 -1598 1524 -1222
rect 1458 -1610 1524 -1598
rect 1554 -1222 1620 -1210
rect 1554 -1598 1570 -1222
rect 1604 -1598 1620 -1222
rect 1554 -1610 1620 -1598
rect 1650 -1222 1716 -1210
rect 1650 -1598 1666 -1222
rect 1700 -1598 1716 -1222
rect 1650 -1610 1716 -1598
rect 1746 -1222 1812 -1210
rect 1746 -1598 1762 -1222
rect 1796 -1598 1812 -1222
rect 1746 -1610 1812 -1598
rect 1842 -1222 1908 -1210
rect 1842 -1598 1858 -1222
rect 1892 -1598 1908 -1222
rect 1842 -1610 1908 -1598
rect 1938 -1222 2004 -1210
rect 1938 -1598 1954 -1222
rect 1988 -1598 2004 -1222
rect 1938 -1610 2004 -1598
rect 2034 -1222 2096 -1210
rect 2034 -1598 2050 -1222
rect 2084 -1598 2096 -1222
rect 2034 -1610 2096 -1598
rect 2438 456 2500 468
rect 2438 80 2450 456
rect 2484 80 2500 456
rect 2438 68 2500 80
rect 2530 456 2596 468
rect 2530 80 2546 456
rect 2580 80 2596 456
rect 2530 68 2596 80
rect 2626 456 2692 468
rect 2626 80 2642 456
rect 2676 80 2692 456
rect 2626 68 2692 80
rect 2722 456 2788 468
rect 2722 80 2738 456
rect 2772 80 2788 456
rect 2722 68 2788 80
rect 2818 456 2884 468
rect 2818 80 2834 456
rect 2868 80 2884 456
rect 2818 68 2884 80
rect 2914 456 2980 468
rect 2914 80 2930 456
rect 2964 80 2980 456
rect 2914 68 2980 80
rect 3010 456 3076 468
rect 3010 80 3026 456
rect 3060 80 3076 456
rect 3010 68 3076 80
rect 3106 456 3172 468
rect 3106 80 3122 456
rect 3156 80 3172 456
rect 3106 68 3172 80
rect 3202 456 3268 468
rect 3202 80 3218 456
rect 3252 80 3268 456
rect 3202 68 3268 80
rect 3298 456 3364 468
rect 3298 80 3314 456
rect 3348 80 3364 456
rect 3298 68 3364 80
rect 3394 456 3460 468
rect 3394 80 3410 456
rect 3444 80 3460 456
rect 3394 68 3460 80
rect 3490 456 3556 468
rect 3490 80 3506 456
rect 3540 80 3556 456
rect 3490 68 3556 80
rect 3586 456 3652 468
rect 3586 80 3602 456
rect 3636 80 3652 456
rect 3586 68 3652 80
rect 3682 456 3748 468
rect 3682 80 3698 456
rect 3732 80 3748 456
rect 3682 68 3748 80
rect 3778 456 3844 468
rect 3778 80 3794 456
rect 3828 80 3844 456
rect 3778 68 3844 80
rect 3874 456 3940 468
rect 3874 80 3890 456
rect 3924 80 3940 456
rect 3874 68 3940 80
rect 3970 456 4036 468
rect 3970 80 3986 456
rect 4020 80 4036 456
rect 3970 68 4036 80
rect 4066 456 4132 468
rect 4066 80 4082 456
rect 4116 80 4132 456
rect 4066 68 4132 80
rect 4162 456 4228 468
rect 4162 80 4178 456
rect 4212 80 4228 456
rect 4162 68 4228 80
rect 4258 456 4324 468
rect 4258 80 4274 456
rect 4308 80 4324 456
rect 4258 68 4324 80
rect 4354 456 4416 468
rect 4354 80 4370 456
rect 4404 80 4416 456
rect 4354 68 4416 80
rect 2438 -162 2500 -150
rect 2438 -538 2450 -162
rect 2484 -538 2500 -162
rect 2438 -550 2500 -538
rect 2530 -162 2596 -150
rect 2530 -538 2546 -162
rect 2580 -538 2596 -162
rect 2530 -550 2596 -538
rect 2626 -162 2692 -150
rect 2626 -538 2642 -162
rect 2676 -538 2692 -162
rect 2626 -550 2692 -538
rect 2722 -162 2788 -150
rect 2722 -538 2738 -162
rect 2772 -538 2788 -162
rect 2722 -550 2788 -538
rect 2818 -162 2884 -150
rect 2818 -538 2834 -162
rect 2868 -538 2884 -162
rect 2818 -550 2884 -538
rect 2914 -162 2980 -150
rect 2914 -538 2930 -162
rect 2964 -538 2980 -162
rect 2914 -550 2980 -538
rect 3010 -162 3076 -150
rect 3010 -538 3026 -162
rect 3060 -538 3076 -162
rect 3010 -550 3076 -538
rect 3106 -162 3172 -150
rect 3106 -538 3122 -162
rect 3156 -538 3172 -162
rect 3106 -550 3172 -538
rect 3202 -162 3268 -150
rect 3202 -538 3218 -162
rect 3252 -538 3268 -162
rect 3202 -550 3268 -538
rect 3298 -162 3364 -150
rect 3298 -538 3314 -162
rect 3348 -538 3364 -162
rect 3298 -550 3364 -538
rect 3394 -162 3460 -150
rect 3394 -538 3410 -162
rect 3444 -538 3460 -162
rect 3394 -550 3460 -538
rect 3490 -162 3556 -150
rect 3490 -538 3506 -162
rect 3540 -538 3556 -162
rect 3490 -550 3556 -538
rect 3586 -162 3652 -150
rect 3586 -538 3602 -162
rect 3636 -538 3652 -162
rect 3586 -550 3652 -538
rect 3682 -162 3748 -150
rect 3682 -538 3698 -162
rect 3732 -538 3748 -162
rect 3682 -550 3748 -538
rect 3778 -162 3844 -150
rect 3778 -538 3794 -162
rect 3828 -538 3844 -162
rect 3778 -550 3844 -538
rect 3874 -162 3940 -150
rect 3874 -538 3890 -162
rect 3924 -538 3940 -162
rect 3874 -550 3940 -538
rect 3970 -162 4036 -150
rect 3970 -538 3986 -162
rect 4020 -538 4036 -162
rect 3970 -550 4036 -538
rect 4066 -162 4132 -150
rect 4066 -538 4082 -162
rect 4116 -538 4132 -162
rect 4066 -550 4132 -538
rect 4162 -162 4228 -150
rect 4162 -538 4178 -162
rect 4212 -538 4228 -162
rect 4162 -550 4228 -538
rect 4258 -162 4324 -150
rect 4258 -538 4274 -162
rect 4308 -538 4324 -162
rect 4258 -550 4324 -538
rect 4354 -162 4416 -150
rect 4354 -538 4370 -162
rect 4404 -538 4416 -162
rect 4354 -550 4416 -538
rect -2462 -2366 -2400 -2354
rect -2462 -2742 -2450 -2366
rect -2416 -2742 -2400 -2366
rect -2462 -2754 -2400 -2742
rect -2370 -2366 -2304 -2354
rect -2370 -2742 -2354 -2366
rect -2320 -2742 -2304 -2366
rect -2370 -2754 -2304 -2742
rect -2274 -2366 -2208 -2354
rect -2274 -2742 -2258 -2366
rect -2224 -2742 -2208 -2366
rect -2274 -2754 -2208 -2742
rect -2178 -2366 -2112 -2354
rect -2178 -2742 -2162 -2366
rect -2128 -2742 -2112 -2366
rect -2178 -2754 -2112 -2742
rect -2082 -2366 -2016 -2354
rect -2082 -2742 -2066 -2366
rect -2032 -2742 -2016 -2366
rect -2082 -2754 -2016 -2742
rect -1986 -2366 -1920 -2354
rect -1986 -2742 -1970 -2366
rect -1936 -2742 -1920 -2366
rect -1986 -2754 -1920 -2742
rect -1890 -2366 -1824 -2354
rect -1890 -2742 -1874 -2366
rect -1840 -2742 -1824 -2366
rect -1890 -2754 -1824 -2742
rect -1794 -2366 -1728 -2354
rect -1794 -2742 -1778 -2366
rect -1744 -2742 -1728 -2366
rect -1794 -2754 -1728 -2742
rect -1698 -2366 -1632 -2354
rect -1698 -2742 -1682 -2366
rect -1648 -2742 -1632 -2366
rect -1698 -2754 -1632 -2742
rect -1602 -2366 -1536 -2354
rect -1602 -2742 -1586 -2366
rect -1552 -2742 -1536 -2366
rect -1602 -2754 -1536 -2742
rect -1506 -2366 -1444 -2354
rect -1506 -2742 -1490 -2366
rect -1456 -2742 -1444 -2366
rect -1506 -2754 -1444 -2742
rect -2462 -2984 -2400 -2972
rect -2462 -3360 -2450 -2984
rect -2416 -3360 -2400 -2984
rect -2462 -3372 -2400 -3360
rect -2370 -2984 -2304 -2972
rect -2370 -3360 -2354 -2984
rect -2320 -3360 -2304 -2984
rect -2370 -3372 -2304 -3360
rect -2274 -2984 -2208 -2972
rect -2274 -3360 -2258 -2984
rect -2224 -3360 -2208 -2984
rect -2274 -3372 -2208 -3360
rect -2178 -2984 -2112 -2972
rect -2178 -3360 -2162 -2984
rect -2128 -3360 -2112 -2984
rect -2178 -3372 -2112 -3360
rect -2082 -2984 -2016 -2972
rect -2082 -3360 -2066 -2984
rect -2032 -3360 -2016 -2984
rect -2082 -3372 -2016 -3360
rect -1986 -2984 -1920 -2972
rect -1986 -3360 -1970 -2984
rect -1936 -3360 -1920 -2984
rect -1986 -3372 -1920 -3360
rect -1890 -2984 -1824 -2972
rect -1890 -3360 -1874 -2984
rect -1840 -3360 -1824 -2984
rect -1890 -3372 -1824 -3360
rect -1794 -2984 -1728 -2972
rect -1794 -3360 -1778 -2984
rect -1744 -3360 -1728 -2984
rect -1794 -3372 -1728 -3360
rect -1698 -2984 -1632 -2972
rect -1698 -3360 -1682 -2984
rect -1648 -3360 -1632 -2984
rect -1698 -3372 -1632 -3360
rect -1602 -2984 -1536 -2972
rect -1602 -3360 -1586 -2984
rect -1552 -3360 -1536 -2984
rect -1602 -3372 -1536 -3360
rect -1506 -2984 -1444 -2972
rect -1506 -3360 -1490 -2984
rect -1456 -3360 -1444 -2984
rect -1506 -3372 -1444 -3360
rect -2462 -3602 -2400 -3590
rect -2462 -3978 -2450 -3602
rect -2416 -3978 -2400 -3602
rect -2462 -3990 -2400 -3978
rect -2370 -3602 -2304 -3590
rect -2370 -3978 -2354 -3602
rect -2320 -3978 -2304 -3602
rect -2370 -3990 -2304 -3978
rect -2274 -3602 -2208 -3590
rect -2274 -3978 -2258 -3602
rect -2224 -3978 -2208 -3602
rect -2274 -3990 -2208 -3978
rect -2178 -3602 -2112 -3590
rect -2178 -3978 -2162 -3602
rect -2128 -3978 -2112 -3602
rect -2178 -3990 -2112 -3978
rect -2082 -3602 -2016 -3590
rect -2082 -3978 -2066 -3602
rect -2032 -3978 -2016 -3602
rect -2082 -3990 -2016 -3978
rect -1986 -3602 -1920 -3590
rect -1986 -3978 -1970 -3602
rect -1936 -3978 -1920 -3602
rect -1986 -3990 -1920 -3978
rect -1890 -3602 -1824 -3590
rect -1890 -3978 -1874 -3602
rect -1840 -3978 -1824 -3602
rect -1890 -3990 -1824 -3978
rect -1794 -3602 -1728 -3590
rect -1794 -3978 -1778 -3602
rect -1744 -3978 -1728 -3602
rect -1794 -3990 -1728 -3978
rect -1698 -3602 -1632 -3590
rect -1698 -3978 -1682 -3602
rect -1648 -3978 -1632 -3602
rect -1698 -3990 -1632 -3978
rect -1602 -3602 -1536 -3590
rect -1602 -3978 -1586 -3602
rect -1552 -3978 -1536 -3602
rect -1602 -3990 -1536 -3978
rect -1506 -3602 -1444 -3590
rect -1506 -3978 -1490 -3602
rect -1456 -3978 -1444 -3602
rect -1506 -3990 -1444 -3978
rect -662 -2366 -600 -2354
rect -662 -2742 -650 -2366
rect -616 -2742 -600 -2366
rect -662 -2754 -600 -2742
rect -570 -2366 -504 -2354
rect -570 -2742 -554 -2366
rect -520 -2742 -504 -2366
rect -570 -2754 -504 -2742
rect -474 -2366 -408 -2354
rect -474 -2742 -458 -2366
rect -424 -2742 -408 -2366
rect -474 -2754 -408 -2742
rect -378 -2366 -312 -2354
rect -378 -2742 -362 -2366
rect -328 -2742 -312 -2366
rect -378 -2754 -312 -2742
rect -282 -2366 -216 -2354
rect -282 -2742 -266 -2366
rect -232 -2742 -216 -2366
rect -282 -2754 -216 -2742
rect -186 -2366 -120 -2354
rect -186 -2742 -170 -2366
rect -136 -2742 -120 -2366
rect -186 -2754 -120 -2742
rect -90 -2366 -24 -2354
rect -90 -2742 -74 -2366
rect -40 -2742 -24 -2366
rect -90 -2754 -24 -2742
rect 6 -2366 72 -2354
rect 6 -2742 22 -2366
rect 56 -2742 72 -2366
rect 6 -2754 72 -2742
rect 102 -2366 168 -2354
rect 102 -2742 118 -2366
rect 152 -2742 168 -2366
rect 102 -2754 168 -2742
rect 198 -2366 264 -2354
rect 198 -2742 214 -2366
rect 248 -2742 264 -2366
rect 198 -2754 264 -2742
rect 294 -2366 356 -2354
rect 294 -2742 310 -2366
rect 344 -2742 356 -2366
rect 294 -2754 356 -2742
rect -662 -2984 -600 -2972
rect -662 -3360 -650 -2984
rect -616 -3360 -600 -2984
rect -662 -3372 -600 -3360
rect -570 -2984 -504 -2972
rect -570 -3360 -554 -2984
rect -520 -3360 -504 -2984
rect -570 -3372 -504 -3360
rect -474 -2984 -408 -2972
rect -474 -3360 -458 -2984
rect -424 -3360 -408 -2984
rect -474 -3372 -408 -3360
rect -378 -2984 -312 -2972
rect -378 -3360 -362 -2984
rect -328 -3360 -312 -2984
rect -378 -3372 -312 -3360
rect -282 -2984 -216 -2972
rect -282 -3360 -266 -2984
rect -232 -3360 -216 -2984
rect -282 -3372 -216 -3360
rect -186 -2984 -120 -2972
rect -186 -3360 -170 -2984
rect -136 -3360 -120 -2984
rect -186 -3372 -120 -3360
rect -90 -2984 -24 -2972
rect -90 -3360 -74 -2984
rect -40 -3360 -24 -2984
rect -90 -3372 -24 -3360
rect 6 -2984 72 -2972
rect 6 -3360 22 -2984
rect 56 -3360 72 -2984
rect 6 -3372 72 -3360
rect 102 -2984 168 -2972
rect 102 -3360 118 -2984
rect 152 -3360 168 -2984
rect 102 -3372 168 -3360
rect 198 -2984 264 -2972
rect 198 -3360 214 -2984
rect 248 -3360 264 -2984
rect 198 -3372 264 -3360
rect 294 -2984 356 -2972
rect 294 -3360 310 -2984
rect 344 -3360 356 -2984
rect 294 -3372 356 -3360
rect -662 -3602 -600 -3590
rect -662 -3978 -650 -3602
rect -616 -3978 -600 -3602
rect -662 -3990 -600 -3978
rect -570 -3602 -504 -3590
rect -570 -3978 -554 -3602
rect -520 -3978 -504 -3602
rect -570 -3990 -504 -3978
rect -474 -3602 -408 -3590
rect -474 -3978 -458 -3602
rect -424 -3978 -408 -3602
rect -474 -3990 -408 -3978
rect -378 -3602 -312 -3590
rect -378 -3978 -362 -3602
rect -328 -3978 -312 -3602
rect -378 -3990 -312 -3978
rect -282 -3602 -216 -3590
rect -282 -3978 -266 -3602
rect -232 -3978 -216 -3602
rect -282 -3990 -216 -3978
rect -186 -3602 -120 -3590
rect -186 -3978 -170 -3602
rect -136 -3978 -120 -3602
rect -186 -3990 -120 -3978
rect -90 -3602 -24 -3590
rect -90 -3978 -74 -3602
rect -40 -3978 -24 -3602
rect -90 -3990 -24 -3978
rect 6 -3602 72 -3590
rect 6 -3978 22 -3602
rect 56 -3978 72 -3602
rect 6 -3990 72 -3978
rect 102 -3602 168 -3590
rect 102 -3978 118 -3602
rect 152 -3978 168 -3602
rect 102 -3990 168 -3978
rect 198 -3602 264 -3590
rect 198 -3978 214 -3602
rect 248 -3978 264 -3602
rect 198 -3990 264 -3978
rect 294 -3602 356 -3590
rect 294 -3978 310 -3602
rect 344 -3978 356 -3602
rect 294 -3990 356 -3978
rect 1138 -2366 1200 -2354
rect 1138 -2742 1150 -2366
rect 1184 -2742 1200 -2366
rect 1138 -2754 1200 -2742
rect 1230 -2366 1296 -2354
rect 1230 -2742 1246 -2366
rect 1280 -2742 1296 -2366
rect 1230 -2754 1296 -2742
rect 1326 -2366 1392 -2354
rect 1326 -2742 1342 -2366
rect 1376 -2742 1392 -2366
rect 1326 -2754 1392 -2742
rect 1422 -2366 1488 -2354
rect 1422 -2742 1438 -2366
rect 1472 -2742 1488 -2366
rect 1422 -2754 1488 -2742
rect 1518 -2366 1584 -2354
rect 1518 -2742 1534 -2366
rect 1568 -2742 1584 -2366
rect 1518 -2754 1584 -2742
rect 1614 -2366 1680 -2354
rect 1614 -2742 1630 -2366
rect 1664 -2742 1680 -2366
rect 1614 -2754 1680 -2742
rect 1710 -2366 1776 -2354
rect 1710 -2742 1726 -2366
rect 1760 -2742 1776 -2366
rect 1710 -2754 1776 -2742
rect 1806 -2366 1872 -2354
rect 1806 -2742 1822 -2366
rect 1856 -2742 1872 -2366
rect 1806 -2754 1872 -2742
rect 1902 -2366 1968 -2354
rect 1902 -2742 1918 -2366
rect 1952 -2742 1968 -2366
rect 1902 -2754 1968 -2742
rect 1998 -2366 2064 -2354
rect 1998 -2742 2014 -2366
rect 2048 -2742 2064 -2366
rect 1998 -2754 2064 -2742
rect 2094 -2366 2156 -2354
rect 2094 -2742 2110 -2366
rect 2144 -2742 2156 -2366
rect 2094 -2754 2156 -2742
rect 1138 -2984 1200 -2972
rect 1138 -3360 1150 -2984
rect 1184 -3360 1200 -2984
rect 1138 -3372 1200 -3360
rect 1230 -2984 1296 -2972
rect 1230 -3360 1246 -2984
rect 1280 -3360 1296 -2984
rect 1230 -3372 1296 -3360
rect 1326 -2984 1392 -2972
rect 1326 -3360 1342 -2984
rect 1376 -3360 1392 -2984
rect 1326 -3372 1392 -3360
rect 1422 -2984 1488 -2972
rect 1422 -3360 1438 -2984
rect 1472 -3360 1488 -2984
rect 1422 -3372 1488 -3360
rect 1518 -2984 1584 -2972
rect 1518 -3360 1534 -2984
rect 1568 -3360 1584 -2984
rect 1518 -3372 1584 -3360
rect 1614 -2984 1680 -2972
rect 1614 -3360 1630 -2984
rect 1664 -3360 1680 -2984
rect 1614 -3372 1680 -3360
rect 1710 -2984 1776 -2972
rect 1710 -3360 1726 -2984
rect 1760 -3360 1776 -2984
rect 1710 -3372 1776 -3360
rect 1806 -2984 1872 -2972
rect 1806 -3360 1822 -2984
rect 1856 -3360 1872 -2984
rect 1806 -3372 1872 -3360
rect 1902 -2984 1968 -2972
rect 1902 -3360 1918 -2984
rect 1952 -3360 1968 -2984
rect 1902 -3372 1968 -3360
rect 1998 -2984 2064 -2972
rect 1998 -3360 2014 -2984
rect 2048 -3360 2064 -2984
rect 1998 -3372 2064 -3360
rect 2094 -2984 2156 -2972
rect 2094 -3360 2110 -2984
rect 2144 -3360 2156 -2984
rect 2094 -3372 2156 -3360
rect 1138 -3602 1200 -3590
rect 1138 -3978 1150 -3602
rect 1184 -3978 1200 -3602
rect 1138 -3990 1200 -3978
rect 1230 -3602 1296 -3590
rect 1230 -3978 1246 -3602
rect 1280 -3978 1296 -3602
rect 1230 -3990 1296 -3978
rect 1326 -3602 1392 -3590
rect 1326 -3978 1342 -3602
rect 1376 -3978 1392 -3602
rect 1326 -3990 1392 -3978
rect 1422 -3602 1488 -3590
rect 1422 -3978 1438 -3602
rect 1472 -3978 1488 -3602
rect 1422 -3990 1488 -3978
rect 1518 -3602 1584 -3590
rect 1518 -3978 1534 -3602
rect 1568 -3978 1584 -3602
rect 1518 -3990 1584 -3978
rect 1614 -3602 1680 -3590
rect 1614 -3978 1630 -3602
rect 1664 -3978 1680 -3602
rect 1614 -3990 1680 -3978
rect 1710 -3602 1776 -3590
rect 1710 -3978 1726 -3602
rect 1760 -3978 1776 -3602
rect 1710 -3990 1776 -3978
rect 1806 -3602 1872 -3590
rect 1806 -3978 1822 -3602
rect 1856 -3978 1872 -3602
rect 1806 -3990 1872 -3978
rect 1902 -3602 1968 -3590
rect 1902 -3978 1918 -3602
rect 1952 -3978 1968 -3602
rect 1902 -3990 1968 -3978
rect 1998 -3602 2064 -3590
rect 1998 -3978 2014 -3602
rect 2048 -3978 2064 -3602
rect 1998 -3990 2064 -3978
rect 2094 -3602 2156 -3590
rect 2094 -3978 2110 -3602
rect 2144 -3978 2156 -3602
rect 2094 -3990 2156 -3978
rect 2938 -2366 3000 -2354
rect 2938 -2742 2950 -2366
rect 2984 -2742 3000 -2366
rect 2938 -2754 3000 -2742
rect 3030 -2366 3096 -2354
rect 3030 -2742 3046 -2366
rect 3080 -2742 3096 -2366
rect 3030 -2754 3096 -2742
rect 3126 -2366 3192 -2354
rect 3126 -2742 3142 -2366
rect 3176 -2742 3192 -2366
rect 3126 -2754 3192 -2742
rect 3222 -2366 3288 -2354
rect 3222 -2742 3238 -2366
rect 3272 -2742 3288 -2366
rect 3222 -2754 3288 -2742
rect 3318 -2366 3384 -2354
rect 3318 -2742 3334 -2366
rect 3368 -2742 3384 -2366
rect 3318 -2754 3384 -2742
rect 3414 -2366 3480 -2354
rect 3414 -2742 3430 -2366
rect 3464 -2742 3480 -2366
rect 3414 -2754 3480 -2742
rect 3510 -2366 3576 -2354
rect 3510 -2742 3526 -2366
rect 3560 -2742 3576 -2366
rect 3510 -2754 3576 -2742
rect 3606 -2366 3672 -2354
rect 3606 -2742 3622 -2366
rect 3656 -2742 3672 -2366
rect 3606 -2754 3672 -2742
rect 3702 -2366 3768 -2354
rect 3702 -2742 3718 -2366
rect 3752 -2742 3768 -2366
rect 3702 -2754 3768 -2742
rect 3798 -2366 3864 -2354
rect 3798 -2742 3814 -2366
rect 3848 -2742 3864 -2366
rect 3798 -2754 3864 -2742
rect 3894 -2366 3956 -2354
rect 3894 -2742 3910 -2366
rect 3944 -2742 3956 -2366
rect 3894 -2754 3956 -2742
rect 2938 -2984 3000 -2972
rect 2938 -3360 2950 -2984
rect 2984 -3360 3000 -2984
rect 2938 -3372 3000 -3360
rect 3030 -2984 3096 -2972
rect 3030 -3360 3046 -2984
rect 3080 -3360 3096 -2984
rect 3030 -3372 3096 -3360
rect 3126 -2984 3192 -2972
rect 3126 -3360 3142 -2984
rect 3176 -3360 3192 -2984
rect 3126 -3372 3192 -3360
rect 3222 -2984 3288 -2972
rect 3222 -3360 3238 -2984
rect 3272 -3360 3288 -2984
rect 3222 -3372 3288 -3360
rect 3318 -2984 3384 -2972
rect 3318 -3360 3334 -2984
rect 3368 -3360 3384 -2984
rect 3318 -3372 3384 -3360
rect 3414 -2984 3480 -2972
rect 3414 -3360 3430 -2984
rect 3464 -3360 3480 -2984
rect 3414 -3372 3480 -3360
rect 3510 -2984 3576 -2972
rect 3510 -3360 3526 -2984
rect 3560 -3360 3576 -2984
rect 3510 -3372 3576 -3360
rect 3606 -2984 3672 -2972
rect 3606 -3360 3622 -2984
rect 3656 -3360 3672 -2984
rect 3606 -3372 3672 -3360
rect 3702 -2984 3768 -2972
rect 3702 -3360 3718 -2984
rect 3752 -3360 3768 -2984
rect 3702 -3372 3768 -3360
rect 3798 -2984 3864 -2972
rect 3798 -3360 3814 -2984
rect 3848 -3360 3864 -2984
rect 3798 -3372 3864 -3360
rect 3894 -2984 3956 -2972
rect 3894 -3360 3910 -2984
rect 3944 -3360 3956 -2984
rect 3894 -3372 3956 -3360
rect 2938 -3602 3000 -3590
rect 2938 -3978 2950 -3602
rect 2984 -3978 3000 -3602
rect 2938 -3990 3000 -3978
rect 3030 -3602 3096 -3590
rect 3030 -3978 3046 -3602
rect 3080 -3978 3096 -3602
rect 3030 -3990 3096 -3978
rect 3126 -3602 3192 -3590
rect 3126 -3978 3142 -3602
rect 3176 -3978 3192 -3602
rect 3126 -3990 3192 -3978
rect 3222 -3602 3288 -3590
rect 3222 -3978 3238 -3602
rect 3272 -3978 3288 -3602
rect 3222 -3990 3288 -3978
rect 3318 -3602 3384 -3590
rect 3318 -3978 3334 -3602
rect 3368 -3978 3384 -3602
rect 3318 -3990 3384 -3978
rect 3414 -3602 3480 -3590
rect 3414 -3978 3430 -3602
rect 3464 -3978 3480 -3602
rect 3414 -3990 3480 -3978
rect 3510 -3602 3576 -3590
rect 3510 -3978 3526 -3602
rect 3560 -3978 3576 -3602
rect 3510 -3990 3576 -3978
rect 3606 -3602 3672 -3590
rect 3606 -3978 3622 -3602
rect 3656 -3978 3672 -3602
rect 3606 -3990 3672 -3978
rect 3702 -3602 3768 -3590
rect 3702 -3978 3718 -3602
rect 3752 -3978 3768 -3602
rect 3702 -3990 3768 -3978
rect 3798 -3602 3864 -3590
rect 3798 -3978 3814 -3602
rect 3848 -3978 3864 -3602
rect 3798 -3990 3864 -3978
rect 3894 -3602 3956 -3590
rect 3894 -3978 3910 -3602
rect 3944 -3978 3956 -3602
rect 3894 -3990 3956 -3978
rect 4938 2022 5000 2034
rect 4938 1646 4950 2022
rect 4984 1646 5000 2022
rect 4938 1634 5000 1646
rect 5030 2022 5096 2034
rect 5030 1646 5046 2022
rect 5080 1646 5096 2022
rect 5030 1634 5096 1646
rect 5126 2022 5192 2034
rect 5126 1646 5142 2022
rect 5176 1646 5192 2022
rect 5126 1634 5192 1646
rect 5222 2022 5288 2034
rect 5222 1646 5238 2022
rect 5272 1646 5288 2022
rect 5222 1634 5288 1646
rect 5318 2022 5384 2034
rect 5318 1646 5334 2022
rect 5368 1646 5384 2022
rect 5318 1634 5384 1646
rect 5414 2022 5480 2034
rect 5414 1646 5430 2022
rect 5464 1646 5480 2022
rect 5414 1634 5480 1646
rect 5510 2022 5576 2034
rect 5510 1646 5526 2022
rect 5560 1646 5576 2022
rect 5510 1634 5576 1646
rect 5606 2022 5672 2034
rect 5606 1646 5622 2022
rect 5656 1646 5672 2022
rect 5606 1634 5672 1646
rect 5702 2022 5768 2034
rect 5702 1646 5718 2022
rect 5752 1646 5768 2022
rect 5702 1634 5768 1646
rect 5798 2022 5864 2034
rect 5798 1646 5814 2022
rect 5848 1646 5864 2022
rect 5798 1634 5864 1646
rect 5894 2022 5960 2034
rect 5894 1646 5910 2022
rect 5944 1646 5960 2022
rect 5894 1634 5960 1646
rect 5990 2022 6056 2034
rect 5990 1646 6006 2022
rect 6040 1646 6056 2022
rect 5990 1634 6056 1646
rect 6086 2022 6152 2034
rect 6086 1646 6102 2022
rect 6136 1646 6152 2022
rect 6086 1634 6152 1646
rect 6182 2022 6248 2034
rect 6182 1646 6198 2022
rect 6232 1646 6248 2022
rect 6182 1634 6248 1646
rect 6278 2022 6344 2034
rect 6278 1646 6294 2022
rect 6328 1646 6344 2022
rect 6278 1634 6344 1646
rect 6374 2022 6440 2034
rect 6374 1646 6390 2022
rect 6424 1646 6440 2022
rect 6374 1634 6440 1646
rect 6470 2022 6536 2034
rect 6470 1646 6486 2022
rect 6520 1646 6536 2022
rect 6470 1634 6536 1646
rect 6566 2022 6632 2034
rect 6566 1646 6582 2022
rect 6616 1646 6632 2022
rect 6566 1634 6632 1646
rect 6662 2022 6728 2034
rect 6662 1646 6678 2022
rect 6712 1646 6728 2022
rect 6662 1634 6728 1646
rect 6758 2022 6824 2034
rect 6758 1646 6774 2022
rect 6808 1646 6824 2022
rect 6758 1634 6824 1646
rect 6854 2022 6916 2034
rect 6854 1646 6870 2022
rect 6904 1646 6916 2022
rect 6854 1634 6916 1646
rect 4938 1404 5000 1416
rect 4938 1028 4950 1404
rect 4984 1028 5000 1404
rect 4938 1016 5000 1028
rect 5030 1404 5096 1416
rect 5030 1028 5046 1404
rect 5080 1028 5096 1404
rect 5030 1016 5096 1028
rect 5126 1404 5192 1416
rect 5126 1028 5142 1404
rect 5176 1028 5192 1404
rect 5126 1016 5192 1028
rect 5222 1404 5288 1416
rect 5222 1028 5238 1404
rect 5272 1028 5288 1404
rect 5222 1016 5288 1028
rect 5318 1404 5384 1416
rect 5318 1028 5334 1404
rect 5368 1028 5384 1404
rect 5318 1016 5384 1028
rect 5414 1404 5480 1416
rect 5414 1028 5430 1404
rect 5464 1028 5480 1404
rect 5414 1016 5480 1028
rect 5510 1404 5576 1416
rect 5510 1028 5526 1404
rect 5560 1028 5576 1404
rect 5510 1016 5576 1028
rect 5606 1404 5672 1416
rect 5606 1028 5622 1404
rect 5656 1028 5672 1404
rect 5606 1016 5672 1028
rect 5702 1404 5768 1416
rect 5702 1028 5718 1404
rect 5752 1028 5768 1404
rect 5702 1016 5768 1028
rect 5798 1404 5864 1416
rect 5798 1028 5814 1404
rect 5848 1028 5864 1404
rect 5798 1016 5864 1028
rect 5894 1404 5960 1416
rect 5894 1028 5910 1404
rect 5944 1028 5960 1404
rect 5894 1016 5960 1028
rect 5990 1404 6056 1416
rect 5990 1028 6006 1404
rect 6040 1028 6056 1404
rect 5990 1016 6056 1028
rect 6086 1404 6152 1416
rect 6086 1028 6102 1404
rect 6136 1028 6152 1404
rect 6086 1016 6152 1028
rect 6182 1404 6248 1416
rect 6182 1028 6198 1404
rect 6232 1028 6248 1404
rect 6182 1016 6248 1028
rect 6278 1404 6344 1416
rect 6278 1028 6294 1404
rect 6328 1028 6344 1404
rect 6278 1016 6344 1028
rect 6374 1404 6440 1416
rect 6374 1028 6390 1404
rect 6424 1028 6440 1404
rect 6374 1016 6440 1028
rect 6470 1404 6536 1416
rect 6470 1028 6486 1404
rect 6520 1028 6536 1404
rect 6470 1016 6536 1028
rect 6566 1404 6632 1416
rect 6566 1028 6582 1404
rect 6616 1028 6632 1404
rect 6566 1016 6632 1028
rect 6662 1404 6728 1416
rect 6662 1028 6678 1404
rect 6712 1028 6728 1404
rect 6662 1016 6728 1028
rect 6758 1404 6824 1416
rect 6758 1028 6774 1404
rect 6808 1028 6824 1404
rect 6758 1016 6824 1028
rect 6854 1404 6916 1416
rect 6854 1028 6870 1404
rect 6904 1028 6916 1404
rect 6854 1016 6916 1028
rect 4938 786 5000 798
rect 4938 410 4950 786
rect 4984 410 5000 786
rect 4938 398 5000 410
rect 5030 786 5096 798
rect 5030 410 5046 786
rect 5080 410 5096 786
rect 5030 398 5096 410
rect 5126 786 5192 798
rect 5126 410 5142 786
rect 5176 410 5192 786
rect 5126 398 5192 410
rect 5222 786 5288 798
rect 5222 410 5238 786
rect 5272 410 5288 786
rect 5222 398 5288 410
rect 5318 786 5384 798
rect 5318 410 5334 786
rect 5368 410 5384 786
rect 5318 398 5384 410
rect 5414 786 5480 798
rect 5414 410 5430 786
rect 5464 410 5480 786
rect 5414 398 5480 410
rect 5510 786 5576 798
rect 5510 410 5526 786
rect 5560 410 5576 786
rect 5510 398 5576 410
rect 5606 786 5672 798
rect 5606 410 5622 786
rect 5656 410 5672 786
rect 5606 398 5672 410
rect 5702 786 5768 798
rect 5702 410 5718 786
rect 5752 410 5768 786
rect 5702 398 5768 410
rect 5798 786 5864 798
rect 5798 410 5814 786
rect 5848 410 5864 786
rect 5798 398 5864 410
rect 5894 786 5960 798
rect 5894 410 5910 786
rect 5944 410 5960 786
rect 5894 398 5960 410
rect 5990 786 6056 798
rect 5990 410 6006 786
rect 6040 410 6056 786
rect 5990 398 6056 410
rect 6086 786 6152 798
rect 6086 410 6102 786
rect 6136 410 6152 786
rect 6086 398 6152 410
rect 6182 786 6248 798
rect 6182 410 6198 786
rect 6232 410 6248 786
rect 6182 398 6248 410
rect 6278 786 6344 798
rect 6278 410 6294 786
rect 6328 410 6344 786
rect 6278 398 6344 410
rect 6374 786 6440 798
rect 6374 410 6390 786
rect 6424 410 6440 786
rect 6374 398 6440 410
rect 6470 786 6536 798
rect 6470 410 6486 786
rect 6520 410 6536 786
rect 6470 398 6536 410
rect 6566 786 6632 798
rect 6566 410 6582 786
rect 6616 410 6632 786
rect 6566 398 6632 410
rect 6662 786 6728 798
rect 6662 410 6678 786
rect 6712 410 6728 786
rect 6662 398 6728 410
rect 6758 786 6824 798
rect 6758 410 6774 786
rect 6808 410 6824 786
rect 6758 398 6824 410
rect 6854 786 6916 798
rect 6854 410 6870 786
rect 6904 410 6916 786
rect 6854 398 6916 410
rect 4938 168 5000 180
rect 4938 -208 4950 168
rect 4984 -208 5000 168
rect 4938 -220 5000 -208
rect 5030 168 5096 180
rect 5030 -208 5046 168
rect 5080 -208 5096 168
rect 5030 -220 5096 -208
rect 5126 168 5192 180
rect 5126 -208 5142 168
rect 5176 -208 5192 168
rect 5126 -220 5192 -208
rect 5222 168 5288 180
rect 5222 -208 5238 168
rect 5272 -208 5288 168
rect 5222 -220 5288 -208
rect 5318 168 5384 180
rect 5318 -208 5334 168
rect 5368 -208 5384 168
rect 5318 -220 5384 -208
rect 5414 168 5480 180
rect 5414 -208 5430 168
rect 5464 -208 5480 168
rect 5414 -220 5480 -208
rect 5510 168 5576 180
rect 5510 -208 5526 168
rect 5560 -208 5576 168
rect 5510 -220 5576 -208
rect 5606 168 5672 180
rect 5606 -208 5622 168
rect 5656 -208 5672 168
rect 5606 -220 5672 -208
rect 5702 168 5768 180
rect 5702 -208 5718 168
rect 5752 -208 5768 168
rect 5702 -220 5768 -208
rect 5798 168 5864 180
rect 5798 -208 5814 168
rect 5848 -208 5864 168
rect 5798 -220 5864 -208
rect 5894 168 5960 180
rect 5894 -208 5910 168
rect 5944 -208 5960 168
rect 5894 -220 5960 -208
rect 5990 168 6056 180
rect 5990 -208 6006 168
rect 6040 -208 6056 168
rect 5990 -220 6056 -208
rect 6086 168 6152 180
rect 6086 -208 6102 168
rect 6136 -208 6152 168
rect 6086 -220 6152 -208
rect 6182 168 6248 180
rect 6182 -208 6198 168
rect 6232 -208 6248 168
rect 6182 -220 6248 -208
rect 6278 168 6344 180
rect 6278 -208 6294 168
rect 6328 -208 6344 168
rect 6278 -220 6344 -208
rect 6374 168 6440 180
rect 6374 -208 6390 168
rect 6424 -208 6440 168
rect 6374 -220 6440 -208
rect 6470 168 6536 180
rect 6470 -208 6486 168
rect 6520 -208 6536 168
rect 6470 -220 6536 -208
rect 6566 168 6632 180
rect 6566 -208 6582 168
rect 6616 -208 6632 168
rect 6566 -220 6632 -208
rect 6662 168 6728 180
rect 6662 -208 6678 168
rect 6712 -208 6728 168
rect 6662 -220 6728 -208
rect 6758 168 6824 180
rect 6758 -208 6774 168
rect 6808 -208 6824 168
rect 6758 -220 6824 -208
rect 6854 168 6916 180
rect 6854 -208 6870 168
rect 6904 -208 6916 168
rect 6854 -220 6916 -208
rect 4938 -450 5000 -438
rect 4938 -826 4950 -450
rect 4984 -826 5000 -450
rect 4938 -838 5000 -826
rect 5030 -450 5096 -438
rect 5030 -826 5046 -450
rect 5080 -826 5096 -450
rect 5030 -838 5096 -826
rect 5126 -450 5192 -438
rect 5126 -826 5142 -450
rect 5176 -826 5192 -450
rect 5126 -838 5192 -826
rect 5222 -450 5288 -438
rect 5222 -826 5238 -450
rect 5272 -826 5288 -450
rect 5222 -838 5288 -826
rect 5318 -450 5384 -438
rect 5318 -826 5334 -450
rect 5368 -826 5384 -450
rect 5318 -838 5384 -826
rect 5414 -450 5480 -438
rect 5414 -826 5430 -450
rect 5464 -826 5480 -450
rect 5414 -838 5480 -826
rect 5510 -450 5576 -438
rect 5510 -826 5526 -450
rect 5560 -826 5576 -450
rect 5510 -838 5576 -826
rect 5606 -450 5672 -438
rect 5606 -826 5622 -450
rect 5656 -826 5672 -450
rect 5606 -838 5672 -826
rect 5702 -450 5768 -438
rect 5702 -826 5718 -450
rect 5752 -826 5768 -450
rect 5702 -838 5768 -826
rect 5798 -450 5864 -438
rect 5798 -826 5814 -450
rect 5848 -826 5864 -450
rect 5798 -838 5864 -826
rect 5894 -450 5960 -438
rect 5894 -826 5910 -450
rect 5944 -826 5960 -450
rect 5894 -838 5960 -826
rect 5990 -450 6056 -438
rect 5990 -826 6006 -450
rect 6040 -826 6056 -450
rect 5990 -838 6056 -826
rect 6086 -450 6152 -438
rect 6086 -826 6102 -450
rect 6136 -826 6152 -450
rect 6086 -838 6152 -826
rect 6182 -450 6248 -438
rect 6182 -826 6198 -450
rect 6232 -826 6248 -450
rect 6182 -838 6248 -826
rect 6278 -450 6344 -438
rect 6278 -826 6294 -450
rect 6328 -826 6344 -450
rect 6278 -838 6344 -826
rect 6374 -450 6440 -438
rect 6374 -826 6390 -450
rect 6424 -826 6440 -450
rect 6374 -838 6440 -826
rect 6470 -450 6536 -438
rect 6470 -826 6486 -450
rect 6520 -826 6536 -450
rect 6470 -838 6536 -826
rect 6566 -450 6632 -438
rect 6566 -826 6582 -450
rect 6616 -826 6632 -450
rect 6566 -838 6632 -826
rect 6662 -450 6728 -438
rect 6662 -826 6678 -450
rect 6712 -826 6728 -450
rect 6662 -838 6728 -826
rect 6758 -450 6824 -438
rect 6758 -826 6774 -450
rect 6808 -826 6824 -450
rect 6758 -838 6824 -826
rect 6854 -450 6916 -438
rect 6854 -826 6870 -450
rect 6904 -826 6916 -450
rect 6854 -838 6916 -826
rect 4938 -1068 5000 -1056
rect 4938 -1444 4950 -1068
rect 4984 -1444 5000 -1068
rect 4938 -1456 5000 -1444
rect 5030 -1068 5096 -1056
rect 5030 -1444 5046 -1068
rect 5080 -1444 5096 -1068
rect 5030 -1456 5096 -1444
rect 5126 -1068 5192 -1056
rect 5126 -1444 5142 -1068
rect 5176 -1444 5192 -1068
rect 5126 -1456 5192 -1444
rect 5222 -1068 5288 -1056
rect 5222 -1444 5238 -1068
rect 5272 -1444 5288 -1068
rect 5222 -1456 5288 -1444
rect 5318 -1068 5384 -1056
rect 5318 -1444 5334 -1068
rect 5368 -1444 5384 -1068
rect 5318 -1456 5384 -1444
rect 5414 -1068 5480 -1056
rect 5414 -1444 5430 -1068
rect 5464 -1444 5480 -1068
rect 5414 -1456 5480 -1444
rect 5510 -1068 5576 -1056
rect 5510 -1444 5526 -1068
rect 5560 -1444 5576 -1068
rect 5510 -1456 5576 -1444
rect 5606 -1068 5672 -1056
rect 5606 -1444 5622 -1068
rect 5656 -1444 5672 -1068
rect 5606 -1456 5672 -1444
rect 5702 -1068 5768 -1056
rect 5702 -1444 5718 -1068
rect 5752 -1444 5768 -1068
rect 5702 -1456 5768 -1444
rect 5798 -1068 5864 -1056
rect 5798 -1444 5814 -1068
rect 5848 -1444 5864 -1068
rect 5798 -1456 5864 -1444
rect 5894 -1068 5960 -1056
rect 5894 -1444 5910 -1068
rect 5944 -1444 5960 -1068
rect 5894 -1456 5960 -1444
rect 5990 -1068 6056 -1056
rect 5990 -1444 6006 -1068
rect 6040 -1444 6056 -1068
rect 5990 -1456 6056 -1444
rect 6086 -1068 6152 -1056
rect 6086 -1444 6102 -1068
rect 6136 -1444 6152 -1068
rect 6086 -1456 6152 -1444
rect 6182 -1068 6248 -1056
rect 6182 -1444 6198 -1068
rect 6232 -1444 6248 -1068
rect 6182 -1456 6248 -1444
rect 6278 -1068 6344 -1056
rect 6278 -1444 6294 -1068
rect 6328 -1444 6344 -1068
rect 6278 -1456 6344 -1444
rect 6374 -1068 6440 -1056
rect 6374 -1444 6390 -1068
rect 6424 -1444 6440 -1068
rect 6374 -1456 6440 -1444
rect 6470 -1068 6536 -1056
rect 6470 -1444 6486 -1068
rect 6520 -1444 6536 -1068
rect 6470 -1456 6536 -1444
rect 6566 -1068 6632 -1056
rect 6566 -1444 6582 -1068
rect 6616 -1444 6632 -1068
rect 6566 -1456 6632 -1444
rect 6662 -1068 6728 -1056
rect 6662 -1444 6678 -1068
rect 6712 -1444 6728 -1068
rect 6662 -1456 6728 -1444
rect 6758 -1068 6824 -1056
rect 6758 -1444 6774 -1068
rect 6808 -1444 6824 -1068
rect 6758 -1456 6824 -1444
rect 6854 -1068 6916 -1056
rect 6854 -1444 6870 -1068
rect 6904 -1444 6916 -1068
rect 6854 -1456 6916 -1444
rect 4938 -1686 5000 -1674
rect 4938 -2062 4950 -1686
rect 4984 -2062 5000 -1686
rect 4938 -2074 5000 -2062
rect 5030 -1686 5096 -1674
rect 5030 -2062 5046 -1686
rect 5080 -2062 5096 -1686
rect 5030 -2074 5096 -2062
rect 5126 -1686 5192 -1674
rect 5126 -2062 5142 -1686
rect 5176 -2062 5192 -1686
rect 5126 -2074 5192 -2062
rect 5222 -1686 5288 -1674
rect 5222 -2062 5238 -1686
rect 5272 -2062 5288 -1686
rect 5222 -2074 5288 -2062
rect 5318 -1686 5384 -1674
rect 5318 -2062 5334 -1686
rect 5368 -2062 5384 -1686
rect 5318 -2074 5384 -2062
rect 5414 -1686 5480 -1674
rect 5414 -2062 5430 -1686
rect 5464 -2062 5480 -1686
rect 5414 -2074 5480 -2062
rect 5510 -1686 5576 -1674
rect 5510 -2062 5526 -1686
rect 5560 -2062 5576 -1686
rect 5510 -2074 5576 -2062
rect 5606 -1686 5672 -1674
rect 5606 -2062 5622 -1686
rect 5656 -2062 5672 -1686
rect 5606 -2074 5672 -2062
rect 5702 -1686 5768 -1674
rect 5702 -2062 5718 -1686
rect 5752 -2062 5768 -1686
rect 5702 -2074 5768 -2062
rect 5798 -1686 5864 -1674
rect 5798 -2062 5814 -1686
rect 5848 -2062 5864 -1686
rect 5798 -2074 5864 -2062
rect 5894 -1686 5960 -1674
rect 5894 -2062 5910 -1686
rect 5944 -2062 5960 -1686
rect 5894 -2074 5960 -2062
rect 5990 -1686 6056 -1674
rect 5990 -2062 6006 -1686
rect 6040 -2062 6056 -1686
rect 5990 -2074 6056 -2062
rect 6086 -1686 6152 -1674
rect 6086 -2062 6102 -1686
rect 6136 -2062 6152 -1686
rect 6086 -2074 6152 -2062
rect 6182 -1686 6248 -1674
rect 6182 -2062 6198 -1686
rect 6232 -2062 6248 -1686
rect 6182 -2074 6248 -2062
rect 6278 -1686 6344 -1674
rect 6278 -2062 6294 -1686
rect 6328 -2062 6344 -1686
rect 6278 -2074 6344 -2062
rect 6374 -1686 6440 -1674
rect 6374 -2062 6390 -1686
rect 6424 -2062 6440 -1686
rect 6374 -2074 6440 -2062
rect 6470 -1686 6536 -1674
rect 6470 -2062 6486 -1686
rect 6520 -2062 6536 -1686
rect 6470 -2074 6536 -2062
rect 6566 -1686 6632 -1674
rect 6566 -2062 6582 -1686
rect 6616 -2062 6632 -1686
rect 6566 -2074 6632 -2062
rect 6662 -1686 6728 -1674
rect 6662 -2062 6678 -1686
rect 6712 -2062 6728 -1686
rect 6662 -2074 6728 -2062
rect 6758 -1686 6824 -1674
rect 6758 -2062 6774 -1686
rect 6808 -2062 6824 -1686
rect 6758 -2074 6824 -2062
rect 6854 -1686 6916 -1674
rect 6854 -2062 6870 -1686
rect 6904 -2062 6916 -1686
rect 6854 -2074 6916 -2062
rect 4938 -2304 5000 -2292
rect 4938 -2680 4950 -2304
rect 4984 -2680 5000 -2304
rect 4938 -2692 5000 -2680
rect 5030 -2304 5096 -2292
rect 5030 -2680 5046 -2304
rect 5080 -2680 5096 -2304
rect 5030 -2692 5096 -2680
rect 5126 -2304 5192 -2292
rect 5126 -2680 5142 -2304
rect 5176 -2680 5192 -2304
rect 5126 -2692 5192 -2680
rect 5222 -2304 5288 -2292
rect 5222 -2680 5238 -2304
rect 5272 -2680 5288 -2304
rect 5222 -2692 5288 -2680
rect 5318 -2304 5384 -2292
rect 5318 -2680 5334 -2304
rect 5368 -2680 5384 -2304
rect 5318 -2692 5384 -2680
rect 5414 -2304 5480 -2292
rect 5414 -2680 5430 -2304
rect 5464 -2680 5480 -2304
rect 5414 -2692 5480 -2680
rect 5510 -2304 5576 -2292
rect 5510 -2680 5526 -2304
rect 5560 -2680 5576 -2304
rect 5510 -2692 5576 -2680
rect 5606 -2304 5672 -2292
rect 5606 -2680 5622 -2304
rect 5656 -2680 5672 -2304
rect 5606 -2692 5672 -2680
rect 5702 -2304 5768 -2292
rect 5702 -2680 5718 -2304
rect 5752 -2680 5768 -2304
rect 5702 -2692 5768 -2680
rect 5798 -2304 5864 -2292
rect 5798 -2680 5814 -2304
rect 5848 -2680 5864 -2304
rect 5798 -2692 5864 -2680
rect 5894 -2304 5960 -2292
rect 5894 -2680 5910 -2304
rect 5944 -2680 5960 -2304
rect 5894 -2692 5960 -2680
rect 5990 -2304 6056 -2292
rect 5990 -2680 6006 -2304
rect 6040 -2680 6056 -2304
rect 5990 -2692 6056 -2680
rect 6086 -2304 6152 -2292
rect 6086 -2680 6102 -2304
rect 6136 -2680 6152 -2304
rect 6086 -2692 6152 -2680
rect 6182 -2304 6248 -2292
rect 6182 -2680 6198 -2304
rect 6232 -2680 6248 -2304
rect 6182 -2692 6248 -2680
rect 6278 -2304 6344 -2292
rect 6278 -2680 6294 -2304
rect 6328 -2680 6344 -2304
rect 6278 -2692 6344 -2680
rect 6374 -2304 6440 -2292
rect 6374 -2680 6390 -2304
rect 6424 -2680 6440 -2304
rect 6374 -2692 6440 -2680
rect 6470 -2304 6536 -2292
rect 6470 -2680 6486 -2304
rect 6520 -2680 6536 -2304
rect 6470 -2692 6536 -2680
rect 6566 -2304 6632 -2292
rect 6566 -2680 6582 -2304
rect 6616 -2680 6632 -2304
rect 6566 -2692 6632 -2680
rect 6662 -2304 6728 -2292
rect 6662 -2680 6678 -2304
rect 6712 -2680 6728 -2304
rect 6662 -2692 6728 -2680
rect 6758 -2304 6824 -2292
rect 6758 -2680 6774 -2304
rect 6808 -2680 6824 -2304
rect 6758 -2692 6824 -2680
rect 6854 -2304 6916 -2292
rect 6854 -2680 6870 -2304
rect 6904 -2680 6916 -2304
rect 6854 -2692 6916 -2680
rect 4938 -2922 5000 -2910
rect 4938 -3298 4950 -2922
rect 4984 -3298 5000 -2922
rect 4938 -3310 5000 -3298
rect 5030 -2922 5096 -2910
rect 5030 -3298 5046 -2922
rect 5080 -3298 5096 -2922
rect 5030 -3310 5096 -3298
rect 5126 -2922 5192 -2910
rect 5126 -3298 5142 -2922
rect 5176 -3298 5192 -2922
rect 5126 -3310 5192 -3298
rect 5222 -2922 5288 -2910
rect 5222 -3298 5238 -2922
rect 5272 -3298 5288 -2922
rect 5222 -3310 5288 -3298
rect 5318 -2922 5384 -2910
rect 5318 -3298 5334 -2922
rect 5368 -3298 5384 -2922
rect 5318 -3310 5384 -3298
rect 5414 -2922 5480 -2910
rect 5414 -3298 5430 -2922
rect 5464 -3298 5480 -2922
rect 5414 -3310 5480 -3298
rect 5510 -2922 5576 -2910
rect 5510 -3298 5526 -2922
rect 5560 -3298 5576 -2922
rect 5510 -3310 5576 -3298
rect 5606 -2922 5672 -2910
rect 5606 -3298 5622 -2922
rect 5656 -3298 5672 -2922
rect 5606 -3310 5672 -3298
rect 5702 -2922 5768 -2910
rect 5702 -3298 5718 -2922
rect 5752 -3298 5768 -2922
rect 5702 -3310 5768 -3298
rect 5798 -2922 5864 -2910
rect 5798 -3298 5814 -2922
rect 5848 -3298 5864 -2922
rect 5798 -3310 5864 -3298
rect 5894 -2922 5960 -2910
rect 5894 -3298 5910 -2922
rect 5944 -3298 5960 -2922
rect 5894 -3310 5960 -3298
rect 5990 -2922 6056 -2910
rect 5990 -3298 6006 -2922
rect 6040 -3298 6056 -2922
rect 5990 -3310 6056 -3298
rect 6086 -2922 6152 -2910
rect 6086 -3298 6102 -2922
rect 6136 -3298 6152 -2922
rect 6086 -3310 6152 -3298
rect 6182 -2922 6248 -2910
rect 6182 -3298 6198 -2922
rect 6232 -3298 6248 -2922
rect 6182 -3310 6248 -3298
rect 6278 -2922 6344 -2910
rect 6278 -3298 6294 -2922
rect 6328 -3298 6344 -2922
rect 6278 -3310 6344 -3298
rect 6374 -2922 6440 -2910
rect 6374 -3298 6390 -2922
rect 6424 -3298 6440 -2922
rect 6374 -3310 6440 -3298
rect 6470 -2922 6536 -2910
rect 6470 -3298 6486 -2922
rect 6520 -3298 6536 -2922
rect 6470 -3310 6536 -3298
rect 6566 -2922 6632 -2910
rect 6566 -3298 6582 -2922
rect 6616 -3298 6632 -2922
rect 6566 -3310 6632 -3298
rect 6662 -2922 6728 -2910
rect 6662 -3298 6678 -2922
rect 6712 -3298 6728 -2922
rect 6662 -3310 6728 -3298
rect 6758 -2922 6824 -2910
rect 6758 -3298 6774 -2922
rect 6808 -3298 6824 -2922
rect 6758 -3310 6824 -3298
rect 6854 -2922 6916 -2910
rect 6854 -3298 6870 -2922
rect 6904 -3298 6916 -2922
rect 6854 -3310 6916 -3298
rect -2462 -4512 -2404 -4500
rect -2462 -4888 -2450 -4512
rect -2416 -4888 -2404 -4512
rect -2462 -4900 -2404 -4888
rect -2204 -4512 -2146 -4500
rect -2204 -4888 -2192 -4512
rect -2158 -4888 -2146 -4512
rect -2204 -4900 -2146 -4888
rect -1946 -4512 -1888 -4500
rect -1946 -4888 -1934 -4512
rect -1900 -4888 -1888 -4512
rect -1946 -4900 -1888 -4888
rect -1688 -4512 -1630 -4500
rect -1688 -4888 -1676 -4512
rect -1642 -4888 -1630 -4512
rect -1688 -4900 -1630 -4888
rect -1430 -4512 -1372 -4500
rect -1430 -4888 -1418 -4512
rect -1384 -4888 -1372 -4512
rect -1430 -4900 -1372 -4888
rect -1172 -4512 -1114 -4500
rect -1172 -4888 -1160 -4512
rect -1126 -4888 -1114 -4512
rect -1172 -4900 -1114 -4888
rect -2462 -5130 -2404 -5118
rect -2462 -5506 -2450 -5130
rect -2416 -5506 -2404 -5130
rect -2462 -5518 -2404 -5506
rect -2204 -5130 -2146 -5118
rect -2204 -5506 -2192 -5130
rect -2158 -5506 -2146 -5130
rect -2204 -5518 -2146 -5506
rect -1946 -5130 -1888 -5118
rect -1946 -5506 -1934 -5130
rect -1900 -5506 -1888 -5130
rect -1946 -5518 -1888 -5506
rect -1688 -5130 -1630 -5118
rect -1688 -5506 -1676 -5130
rect -1642 -5506 -1630 -5130
rect -1688 -5518 -1630 -5506
rect -1430 -5130 -1372 -5118
rect -1430 -5506 -1418 -5130
rect -1384 -5506 -1372 -5130
rect -1430 -5518 -1372 -5506
rect -1172 -5130 -1114 -5118
rect -1172 -5506 -1160 -5130
rect -1126 -5506 -1114 -5130
rect -1172 -5518 -1114 -5506
rect -2462 -5748 -2404 -5736
rect -2462 -6124 -2450 -5748
rect -2416 -6124 -2404 -5748
rect -2462 -6136 -2404 -6124
rect -2204 -5748 -2146 -5736
rect -2204 -6124 -2192 -5748
rect -2158 -6124 -2146 -5748
rect -2204 -6136 -2146 -6124
rect -1946 -5748 -1888 -5736
rect -1946 -6124 -1934 -5748
rect -1900 -6124 -1888 -5748
rect -1946 -6136 -1888 -6124
rect -1688 -5748 -1630 -5736
rect -1688 -6124 -1676 -5748
rect -1642 -6124 -1630 -5748
rect -1688 -6136 -1630 -6124
rect -1430 -5748 -1372 -5736
rect -1430 -6124 -1418 -5748
rect -1384 -6124 -1372 -5748
rect -1430 -6136 -1372 -6124
rect -1172 -5748 -1114 -5736
rect -1172 -6124 -1160 -5748
rect -1126 -6124 -1114 -5748
rect -1172 -6136 -1114 -6124
rect -2462 -6366 -2404 -6354
rect -2462 -6742 -2450 -6366
rect -2416 -6742 -2404 -6366
rect -2462 -6754 -2404 -6742
rect -2204 -6366 -2146 -6354
rect -2204 -6742 -2192 -6366
rect -2158 -6742 -2146 -6366
rect -2204 -6754 -2146 -6742
rect -1946 -6366 -1888 -6354
rect -1946 -6742 -1934 -6366
rect -1900 -6742 -1888 -6366
rect -1946 -6754 -1888 -6742
rect -1688 -6366 -1630 -6354
rect -1688 -6742 -1676 -6366
rect -1642 -6742 -1630 -6366
rect -1688 -6754 -1630 -6742
rect -1430 -6366 -1372 -6354
rect -1430 -6742 -1418 -6366
rect -1384 -6742 -1372 -6366
rect -1430 -6754 -1372 -6742
rect -1172 -6366 -1114 -6354
rect -1172 -6742 -1160 -6366
rect -1126 -6742 -1114 -6366
rect -1172 -6754 -1114 -6742
rect -2462 -6984 -2404 -6972
rect -2462 -7360 -2450 -6984
rect -2416 -7360 -2404 -6984
rect -2462 -7372 -2404 -7360
rect -2204 -6984 -2146 -6972
rect -2204 -7360 -2192 -6984
rect -2158 -7360 -2146 -6984
rect -2204 -7372 -2146 -7360
rect -1946 -6984 -1888 -6972
rect -1946 -7360 -1934 -6984
rect -1900 -7360 -1888 -6984
rect -1946 -7372 -1888 -7360
rect -1688 -6984 -1630 -6972
rect -1688 -7360 -1676 -6984
rect -1642 -7360 -1630 -6984
rect -1688 -7372 -1630 -7360
rect -1430 -6984 -1372 -6972
rect -1430 -7360 -1418 -6984
rect -1384 -7360 -1372 -6984
rect -1430 -7372 -1372 -7360
rect -1172 -6984 -1114 -6972
rect -1172 -7360 -1160 -6984
rect -1126 -7360 -1114 -6984
rect -1172 -7372 -1114 -7360
rect -2462 -7602 -2404 -7590
rect -2462 -7978 -2450 -7602
rect -2416 -7978 -2404 -7602
rect -2462 -7990 -2404 -7978
rect -2204 -7602 -2146 -7590
rect -2204 -7978 -2192 -7602
rect -2158 -7978 -2146 -7602
rect -2204 -7990 -2146 -7978
rect -1946 -7602 -1888 -7590
rect -1946 -7978 -1934 -7602
rect -1900 -7978 -1888 -7602
rect -1946 -7990 -1888 -7978
rect -1688 -7602 -1630 -7590
rect -1688 -7978 -1676 -7602
rect -1642 -7978 -1630 -7602
rect -1688 -7990 -1630 -7978
rect -1430 -7602 -1372 -7590
rect -1430 -7978 -1418 -7602
rect -1384 -7978 -1372 -7602
rect -1430 -7990 -1372 -7978
rect -1172 -7602 -1114 -7590
rect -1172 -7978 -1160 -7602
rect -1126 -7978 -1114 -7602
rect -1172 -7990 -1114 -7978
rect -662 -4512 -604 -4500
rect -662 -4888 -650 -4512
rect -616 -4888 -604 -4512
rect -662 -4900 -604 -4888
rect -404 -4512 -346 -4500
rect -404 -4888 -392 -4512
rect -358 -4888 -346 -4512
rect -404 -4900 -346 -4888
rect -146 -4512 -88 -4500
rect -146 -4888 -134 -4512
rect -100 -4888 -88 -4512
rect -146 -4900 -88 -4888
rect 112 -4512 170 -4500
rect 112 -4888 124 -4512
rect 158 -4888 170 -4512
rect 112 -4900 170 -4888
rect 370 -4512 428 -4500
rect 370 -4888 382 -4512
rect 416 -4888 428 -4512
rect 370 -4900 428 -4888
rect 628 -4512 686 -4500
rect 628 -4888 640 -4512
rect 674 -4888 686 -4512
rect 628 -4900 686 -4888
rect -662 -5130 -604 -5118
rect -662 -5506 -650 -5130
rect -616 -5506 -604 -5130
rect -662 -5518 -604 -5506
rect -404 -5130 -346 -5118
rect -404 -5506 -392 -5130
rect -358 -5506 -346 -5130
rect -404 -5518 -346 -5506
rect -146 -5130 -88 -5118
rect -146 -5506 -134 -5130
rect -100 -5506 -88 -5130
rect -146 -5518 -88 -5506
rect 112 -5130 170 -5118
rect 112 -5506 124 -5130
rect 158 -5506 170 -5130
rect 112 -5518 170 -5506
rect 370 -5130 428 -5118
rect 370 -5506 382 -5130
rect 416 -5506 428 -5130
rect 370 -5518 428 -5506
rect 628 -5130 686 -5118
rect 628 -5506 640 -5130
rect 674 -5506 686 -5130
rect 628 -5518 686 -5506
rect -662 -5748 -604 -5736
rect -662 -6124 -650 -5748
rect -616 -6124 -604 -5748
rect -662 -6136 -604 -6124
rect -404 -5748 -346 -5736
rect -404 -6124 -392 -5748
rect -358 -6124 -346 -5748
rect -404 -6136 -346 -6124
rect -146 -5748 -88 -5736
rect -146 -6124 -134 -5748
rect -100 -6124 -88 -5748
rect -146 -6136 -88 -6124
rect 112 -5748 170 -5736
rect 112 -6124 124 -5748
rect 158 -6124 170 -5748
rect 112 -6136 170 -6124
rect 370 -5748 428 -5736
rect 370 -6124 382 -5748
rect 416 -6124 428 -5748
rect 370 -6136 428 -6124
rect 628 -5748 686 -5736
rect 628 -6124 640 -5748
rect 674 -6124 686 -5748
rect 628 -6136 686 -6124
rect -662 -6366 -604 -6354
rect -662 -6742 -650 -6366
rect -616 -6742 -604 -6366
rect -662 -6754 -604 -6742
rect -404 -6366 -346 -6354
rect -404 -6742 -392 -6366
rect -358 -6742 -346 -6366
rect -404 -6754 -346 -6742
rect -146 -6366 -88 -6354
rect -146 -6742 -134 -6366
rect -100 -6742 -88 -6366
rect -146 -6754 -88 -6742
rect 112 -6366 170 -6354
rect 112 -6742 124 -6366
rect 158 -6742 170 -6366
rect 112 -6754 170 -6742
rect 370 -6366 428 -6354
rect 370 -6742 382 -6366
rect 416 -6742 428 -6366
rect 370 -6754 428 -6742
rect 628 -6366 686 -6354
rect 628 -6742 640 -6366
rect 674 -6742 686 -6366
rect 628 -6754 686 -6742
rect -662 -6984 -604 -6972
rect -662 -7360 -650 -6984
rect -616 -7360 -604 -6984
rect -662 -7372 -604 -7360
rect -404 -6984 -346 -6972
rect -404 -7360 -392 -6984
rect -358 -7360 -346 -6984
rect -404 -7372 -346 -7360
rect -146 -6984 -88 -6972
rect -146 -7360 -134 -6984
rect -100 -7360 -88 -6984
rect -146 -7372 -88 -7360
rect 112 -6984 170 -6972
rect 112 -7360 124 -6984
rect 158 -7360 170 -6984
rect 112 -7372 170 -7360
rect 370 -6984 428 -6972
rect 370 -7360 382 -6984
rect 416 -7360 428 -6984
rect 370 -7372 428 -7360
rect 628 -6984 686 -6972
rect 628 -7360 640 -6984
rect 674 -7360 686 -6984
rect 628 -7372 686 -7360
rect -662 -7602 -604 -7590
rect -662 -7978 -650 -7602
rect -616 -7978 -604 -7602
rect -662 -7990 -604 -7978
rect -404 -7602 -346 -7590
rect -404 -7978 -392 -7602
rect -358 -7978 -346 -7602
rect -404 -7990 -346 -7978
rect -146 -7602 -88 -7590
rect -146 -7978 -134 -7602
rect -100 -7978 -88 -7602
rect -146 -7990 -88 -7978
rect 112 -7602 170 -7590
rect 112 -7978 124 -7602
rect 158 -7978 170 -7602
rect 112 -7990 170 -7978
rect 370 -7602 428 -7590
rect 370 -7978 382 -7602
rect 416 -7978 428 -7602
rect 370 -7990 428 -7978
rect 628 -7602 686 -7590
rect 628 -7978 640 -7602
rect 674 -7978 686 -7602
rect 628 -7990 686 -7978
rect 1138 -4512 1196 -4500
rect 1138 -4888 1150 -4512
rect 1184 -4888 1196 -4512
rect 1138 -4900 1196 -4888
rect 1396 -4512 1454 -4500
rect 1396 -4888 1408 -4512
rect 1442 -4888 1454 -4512
rect 1396 -4900 1454 -4888
rect 1654 -4512 1712 -4500
rect 1654 -4888 1666 -4512
rect 1700 -4888 1712 -4512
rect 1654 -4900 1712 -4888
rect 1912 -4512 1970 -4500
rect 1912 -4888 1924 -4512
rect 1958 -4888 1970 -4512
rect 1912 -4900 1970 -4888
rect 2170 -4512 2228 -4500
rect 2170 -4888 2182 -4512
rect 2216 -4888 2228 -4512
rect 2170 -4900 2228 -4888
rect 2428 -4512 2486 -4500
rect 2428 -4888 2440 -4512
rect 2474 -4888 2486 -4512
rect 2428 -4900 2486 -4888
rect 1138 -5130 1196 -5118
rect 1138 -5506 1150 -5130
rect 1184 -5506 1196 -5130
rect 1138 -5518 1196 -5506
rect 1396 -5130 1454 -5118
rect 1396 -5506 1408 -5130
rect 1442 -5506 1454 -5130
rect 1396 -5518 1454 -5506
rect 1654 -5130 1712 -5118
rect 1654 -5506 1666 -5130
rect 1700 -5506 1712 -5130
rect 1654 -5518 1712 -5506
rect 1912 -5130 1970 -5118
rect 1912 -5506 1924 -5130
rect 1958 -5506 1970 -5130
rect 1912 -5518 1970 -5506
rect 2170 -5130 2228 -5118
rect 2170 -5506 2182 -5130
rect 2216 -5506 2228 -5130
rect 2170 -5518 2228 -5506
rect 2428 -5130 2486 -5118
rect 2428 -5506 2440 -5130
rect 2474 -5506 2486 -5130
rect 2428 -5518 2486 -5506
rect 1138 -5748 1196 -5736
rect 1138 -6124 1150 -5748
rect 1184 -6124 1196 -5748
rect 1138 -6136 1196 -6124
rect 1396 -5748 1454 -5736
rect 1396 -6124 1408 -5748
rect 1442 -6124 1454 -5748
rect 1396 -6136 1454 -6124
rect 1654 -5748 1712 -5736
rect 1654 -6124 1666 -5748
rect 1700 -6124 1712 -5748
rect 1654 -6136 1712 -6124
rect 1912 -5748 1970 -5736
rect 1912 -6124 1924 -5748
rect 1958 -6124 1970 -5748
rect 1912 -6136 1970 -6124
rect 2170 -5748 2228 -5736
rect 2170 -6124 2182 -5748
rect 2216 -6124 2228 -5748
rect 2170 -6136 2228 -6124
rect 2428 -5748 2486 -5736
rect 2428 -6124 2440 -5748
rect 2474 -6124 2486 -5748
rect 2428 -6136 2486 -6124
rect 1138 -6366 1196 -6354
rect 1138 -6742 1150 -6366
rect 1184 -6742 1196 -6366
rect 1138 -6754 1196 -6742
rect 1396 -6366 1454 -6354
rect 1396 -6742 1408 -6366
rect 1442 -6742 1454 -6366
rect 1396 -6754 1454 -6742
rect 1654 -6366 1712 -6354
rect 1654 -6742 1666 -6366
rect 1700 -6742 1712 -6366
rect 1654 -6754 1712 -6742
rect 1912 -6366 1970 -6354
rect 1912 -6742 1924 -6366
rect 1958 -6742 1970 -6366
rect 1912 -6754 1970 -6742
rect 2170 -6366 2228 -6354
rect 2170 -6742 2182 -6366
rect 2216 -6742 2228 -6366
rect 2170 -6754 2228 -6742
rect 2428 -6366 2486 -6354
rect 2428 -6742 2440 -6366
rect 2474 -6742 2486 -6366
rect 2428 -6754 2486 -6742
rect 1138 -6984 1196 -6972
rect 1138 -7360 1150 -6984
rect 1184 -7360 1196 -6984
rect 1138 -7372 1196 -7360
rect 1396 -6984 1454 -6972
rect 1396 -7360 1408 -6984
rect 1442 -7360 1454 -6984
rect 1396 -7372 1454 -7360
rect 1654 -6984 1712 -6972
rect 1654 -7360 1666 -6984
rect 1700 -7360 1712 -6984
rect 1654 -7372 1712 -7360
rect 1912 -6984 1970 -6972
rect 1912 -7360 1924 -6984
rect 1958 -7360 1970 -6984
rect 1912 -7372 1970 -7360
rect 2170 -6984 2228 -6972
rect 2170 -7360 2182 -6984
rect 2216 -7360 2228 -6984
rect 2170 -7372 2228 -7360
rect 2428 -6984 2486 -6972
rect 2428 -7360 2440 -6984
rect 2474 -7360 2486 -6984
rect 2428 -7372 2486 -7360
rect 1138 -7602 1196 -7590
rect 1138 -7978 1150 -7602
rect 1184 -7978 1196 -7602
rect 1138 -7990 1196 -7978
rect 1396 -7602 1454 -7590
rect 1396 -7978 1408 -7602
rect 1442 -7978 1454 -7602
rect 1396 -7990 1454 -7978
rect 1654 -7602 1712 -7590
rect 1654 -7978 1666 -7602
rect 1700 -7978 1712 -7602
rect 1654 -7990 1712 -7978
rect 1912 -7602 1970 -7590
rect 1912 -7978 1924 -7602
rect 1958 -7978 1970 -7602
rect 1912 -7990 1970 -7978
rect 2170 -7602 2228 -7590
rect 2170 -7978 2182 -7602
rect 2216 -7978 2228 -7602
rect 2170 -7990 2228 -7978
rect 2428 -7602 2486 -7590
rect 2428 -7978 2440 -7602
rect 2474 -7978 2486 -7602
rect 2428 -7990 2486 -7978
rect 2938 -4512 2996 -4500
rect 2938 -4888 2950 -4512
rect 2984 -4888 2996 -4512
rect 2938 -4900 2996 -4888
rect 3196 -4512 3254 -4500
rect 3196 -4888 3208 -4512
rect 3242 -4888 3254 -4512
rect 3196 -4900 3254 -4888
rect 3454 -4512 3512 -4500
rect 3454 -4888 3466 -4512
rect 3500 -4888 3512 -4512
rect 3454 -4900 3512 -4888
rect 3712 -4512 3770 -4500
rect 3712 -4888 3724 -4512
rect 3758 -4888 3770 -4512
rect 3712 -4900 3770 -4888
rect 3970 -4512 4028 -4500
rect 3970 -4888 3982 -4512
rect 4016 -4888 4028 -4512
rect 3970 -4900 4028 -4888
rect 4228 -4512 4286 -4500
rect 4228 -4888 4240 -4512
rect 4274 -4888 4286 -4512
rect 4228 -4900 4286 -4888
rect 2938 -5130 2996 -5118
rect 2938 -5506 2950 -5130
rect 2984 -5506 2996 -5130
rect 2938 -5518 2996 -5506
rect 3196 -5130 3254 -5118
rect 3196 -5506 3208 -5130
rect 3242 -5506 3254 -5130
rect 3196 -5518 3254 -5506
rect 3454 -5130 3512 -5118
rect 3454 -5506 3466 -5130
rect 3500 -5506 3512 -5130
rect 3454 -5518 3512 -5506
rect 3712 -5130 3770 -5118
rect 3712 -5506 3724 -5130
rect 3758 -5506 3770 -5130
rect 3712 -5518 3770 -5506
rect 3970 -5130 4028 -5118
rect 3970 -5506 3982 -5130
rect 4016 -5506 4028 -5130
rect 3970 -5518 4028 -5506
rect 4228 -5130 4286 -5118
rect 4228 -5506 4240 -5130
rect 4274 -5506 4286 -5130
rect 4228 -5518 4286 -5506
rect 2938 -5748 2996 -5736
rect 2938 -6124 2950 -5748
rect 2984 -6124 2996 -5748
rect 2938 -6136 2996 -6124
rect 3196 -5748 3254 -5736
rect 3196 -6124 3208 -5748
rect 3242 -6124 3254 -5748
rect 3196 -6136 3254 -6124
rect 3454 -5748 3512 -5736
rect 3454 -6124 3466 -5748
rect 3500 -6124 3512 -5748
rect 3454 -6136 3512 -6124
rect 3712 -5748 3770 -5736
rect 3712 -6124 3724 -5748
rect 3758 -6124 3770 -5748
rect 3712 -6136 3770 -6124
rect 3970 -5748 4028 -5736
rect 3970 -6124 3982 -5748
rect 4016 -6124 4028 -5748
rect 3970 -6136 4028 -6124
rect 4228 -5748 4286 -5736
rect 4228 -6124 4240 -5748
rect 4274 -6124 4286 -5748
rect 4228 -6136 4286 -6124
rect 2938 -6366 2996 -6354
rect 2938 -6742 2950 -6366
rect 2984 -6742 2996 -6366
rect 2938 -6754 2996 -6742
rect 3196 -6366 3254 -6354
rect 3196 -6742 3208 -6366
rect 3242 -6742 3254 -6366
rect 3196 -6754 3254 -6742
rect 3454 -6366 3512 -6354
rect 3454 -6742 3466 -6366
rect 3500 -6742 3512 -6366
rect 3454 -6754 3512 -6742
rect 3712 -6366 3770 -6354
rect 3712 -6742 3724 -6366
rect 3758 -6742 3770 -6366
rect 3712 -6754 3770 -6742
rect 3970 -6366 4028 -6354
rect 3970 -6742 3982 -6366
rect 4016 -6742 4028 -6366
rect 3970 -6754 4028 -6742
rect 4228 -6366 4286 -6354
rect 4228 -6742 4240 -6366
rect 4274 -6742 4286 -6366
rect 4228 -6754 4286 -6742
rect 2938 -6984 2996 -6972
rect 2938 -7360 2950 -6984
rect 2984 -7360 2996 -6984
rect 2938 -7372 2996 -7360
rect 3196 -6984 3254 -6972
rect 3196 -7360 3208 -6984
rect 3242 -7360 3254 -6984
rect 3196 -7372 3254 -7360
rect 3454 -6984 3512 -6972
rect 3454 -7360 3466 -6984
rect 3500 -7360 3512 -6984
rect 3454 -7372 3512 -7360
rect 3712 -6984 3770 -6972
rect 3712 -7360 3724 -6984
rect 3758 -7360 3770 -6984
rect 3712 -7372 3770 -7360
rect 3970 -6984 4028 -6972
rect 3970 -7360 3982 -6984
rect 4016 -7360 4028 -6984
rect 3970 -7372 4028 -7360
rect 4228 -6984 4286 -6972
rect 4228 -7360 4240 -6984
rect 4274 -7360 4286 -6984
rect 4228 -7372 4286 -7360
rect 2938 -7602 2996 -7590
rect 2938 -7978 2950 -7602
rect 2984 -7978 2996 -7602
rect 2938 -7990 2996 -7978
rect 3196 -7602 3254 -7590
rect 3196 -7978 3208 -7602
rect 3242 -7978 3254 -7602
rect 3196 -7990 3254 -7978
rect 3454 -7602 3512 -7590
rect 3454 -7978 3466 -7602
rect 3500 -7978 3512 -7602
rect 3454 -7990 3512 -7978
rect 3712 -7602 3770 -7590
rect 3712 -7978 3724 -7602
rect 3758 -7978 3770 -7602
rect 3712 -7990 3770 -7978
rect 3970 -7602 4028 -7590
rect 3970 -7978 3982 -7602
rect 4016 -7978 4028 -7602
rect 3970 -7990 4028 -7978
rect 4228 -7602 4286 -7590
rect 4228 -7978 4240 -7602
rect 4274 -7978 4286 -7602
rect 4228 -7990 4286 -7978
<< pdiff >>
rect 2438 2043 2500 2055
rect 2438 1667 2450 2043
rect 2484 1667 2500 2043
rect 2438 1655 2500 1667
rect 2530 2043 2596 2055
rect 2530 1667 2546 2043
rect 2580 1667 2596 2043
rect 2530 1655 2596 1667
rect 2626 2043 2692 2055
rect 2626 1667 2642 2043
rect 2676 1667 2692 2043
rect 2626 1655 2692 1667
rect 2722 2043 2788 2055
rect 2722 1667 2738 2043
rect 2772 1667 2788 2043
rect 2722 1655 2788 1667
rect 2818 2043 2884 2055
rect 2818 1667 2834 2043
rect 2868 1667 2884 2043
rect 2818 1655 2884 1667
rect 2914 2043 2980 2055
rect 2914 1667 2930 2043
rect 2964 1667 2980 2043
rect 2914 1655 2980 1667
rect 3010 2043 3076 2055
rect 3010 1667 3026 2043
rect 3060 1667 3076 2043
rect 3010 1655 3076 1667
rect 3106 2043 3172 2055
rect 3106 1667 3122 2043
rect 3156 1667 3172 2043
rect 3106 1655 3172 1667
rect 3202 2043 3268 2055
rect 3202 1667 3218 2043
rect 3252 1667 3268 2043
rect 3202 1655 3268 1667
rect 3298 2043 3364 2055
rect 3298 1667 3314 2043
rect 3348 1667 3364 2043
rect 3298 1655 3364 1667
rect 3394 2043 3460 2055
rect 3394 1667 3410 2043
rect 3444 1667 3460 2043
rect 3394 1655 3460 1667
rect 3490 2043 3556 2055
rect 3490 1667 3506 2043
rect 3540 1667 3556 2043
rect 3490 1655 3556 1667
rect 3586 2043 3652 2055
rect 3586 1667 3602 2043
rect 3636 1667 3652 2043
rect 3586 1655 3652 1667
rect 3682 2043 3748 2055
rect 3682 1667 3698 2043
rect 3732 1667 3748 2043
rect 3682 1655 3748 1667
rect 3778 2043 3844 2055
rect 3778 1667 3794 2043
rect 3828 1667 3844 2043
rect 3778 1655 3844 1667
rect 3874 2043 3940 2055
rect 3874 1667 3890 2043
rect 3924 1667 3940 2043
rect 3874 1655 3940 1667
rect 3970 2043 4036 2055
rect 3970 1667 3986 2043
rect 4020 1667 4036 2043
rect 3970 1655 4036 1667
rect 4066 2043 4132 2055
rect 4066 1667 4082 2043
rect 4116 1667 4132 2043
rect 4066 1655 4132 1667
rect 4162 2043 4228 2055
rect 4162 1667 4178 2043
rect 4212 1667 4228 2043
rect 4162 1655 4228 1667
rect 4258 2043 4324 2055
rect 4258 1667 4274 2043
rect 4308 1667 4324 2043
rect 4258 1655 4324 1667
rect 4354 2043 4416 2055
rect 4354 1667 4370 2043
rect 4404 1667 4416 2043
rect 4354 1655 4416 1667
rect 2438 1407 2500 1419
rect 2438 1031 2450 1407
rect 2484 1031 2500 1407
rect 2438 1019 2500 1031
rect 2530 1407 2596 1419
rect 2530 1031 2546 1407
rect 2580 1031 2596 1407
rect 2530 1019 2596 1031
rect 2626 1407 2692 1419
rect 2626 1031 2642 1407
rect 2676 1031 2692 1407
rect 2626 1019 2692 1031
rect 2722 1407 2788 1419
rect 2722 1031 2738 1407
rect 2772 1031 2788 1407
rect 2722 1019 2788 1031
rect 2818 1407 2884 1419
rect 2818 1031 2834 1407
rect 2868 1031 2884 1407
rect 2818 1019 2884 1031
rect 2914 1407 2980 1419
rect 2914 1031 2930 1407
rect 2964 1031 2980 1407
rect 2914 1019 2980 1031
rect 3010 1407 3076 1419
rect 3010 1031 3026 1407
rect 3060 1031 3076 1407
rect 3010 1019 3076 1031
rect 3106 1407 3172 1419
rect 3106 1031 3122 1407
rect 3156 1031 3172 1407
rect 3106 1019 3172 1031
rect 3202 1407 3268 1419
rect 3202 1031 3218 1407
rect 3252 1031 3268 1407
rect 3202 1019 3268 1031
rect 3298 1407 3364 1419
rect 3298 1031 3314 1407
rect 3348 1031 3364 1407
rect 3298 1019 3364 1031
rect 3394 1407 3460 1419
rect 3394 1031 3410 1407
rect 3444 1031 3460 1407
rect 3394 1019 3460 1031
rect 3490 1407 3556 1419
rect 3490 1031 3506 1407
rect 3540 1031 3556 1407
rect 3490 1019 3556 1031
rect 3586 1407 3652 1419
rect 3586 1031 3602 1407
rect 3636 1031 3652 1407
rect 3586 1019 3652 1031
rect 3682 1407 3748 1419
rect 3682 1031 3698 1407
rect 3732 1031 3748 1407
rect 3682 1019 3748 1031
rect 3778 1407 3844 1419
rect 3778 1031 3794 1407
rect 3828 1031 3844 1407
rect 3778 1019 3844 1031
rect 3874 1407 3940 1419
rect 3874 1031 3890 1407
rect 3924 1031 3940 1407
rect 3874 1019 3940 1031
rect 3970 1407 4036 1419
rect 3970 1031 3986 1407
rect 4020 1031 4036 1407
rect 3970 1019 4036 1031
rect 4066 1407 4132 1419
rect 4066 1031 4082 1407
rect 4116 1031 4132 1407
rect 4066 1019 4132 1031
rect 4162 1407 4228 1419
rect 4162 1031 4178 1407
rect 4212 1031 4228 1407
rect 4162 1019 4228 1031
rect 4258 1407 4324 1419
rect 4258 1031 4274 1407
rect 4308 1031 4324 1407
rect 4258 1019 4324 1031
rect 4354 1407 4416 1419
rect 4354 1031 4370 1407
rect 4404 1031 4416 1407
rect 4354 1019 4416 1031
<< ndiffc >>
rect 130 -362 164 14
rect 226 -362 260 14
rect 322 -362 356 14
rect 418 -362 452 14
rect 514 -362 548 14
rect 610 -362 644 14
rect 706 -362 740 14
rect 802 -362 836 14
rect 898 -362 932 14
rect 994 -362 1028 14
rect 1090 -362 1124 14
rect 1186 -362 1220 14
rect 1282 -362 1316 14
rect 1378 -362 1412 14
rect 1474 -362 1508 14
rect 1570 -362 1604 14
rect 1666 -362 1700 14
rect 1762 -362 1796 14
rect 1858 -362 1892 14
rect 1954 -362 1988 14
rect 2050 -362 2084 14
rect 130 -980 164 -604
rect 226 -980 260 -604
rect 322 -980 356 -604
rect 418 -980 452 -604
rect 514 -980 548 -604
rect 610 -980 644 -604
rect 706 -980 740 -604
rect 802 -980 836 -604
rect 898 -980 932 -604
rect 994 -980 1028 -604
rect 1090 -980 1124 -604
rect 1186 -980 1220 -604
rect 1282 -980 1316 -604
rect 1378 -980 1412 -604
rect 1474 -980 1508 -604
rect 1570 -980 1604 -604
rect 1666 -980 1700 -604
rect 1762 -980 1796 -604
rect 1858 -980 1892 -604
rect 1954 -980 1988 -604
rect 2050 -980 2084 -604
rect 130 -1598 164 -1222
rect 226 -1598 260 -1222
rect 322 -1598 356 -1222
rect 418 -1598 452 -1222
rect 514 -1598 548 -1222
rect 610 -1598 644 -1222
rect 706 -1598 740 -1222
rect 802 -1598 836 -1222
rect 898 -1598 932 -1222
rect 994 -1598 1028 -1222
rect 1090 -1598 1124 -1222
rect 1186 -1598 1220 -1222
rect 1282 -1598 1316 -1222
rect 1378 -1598 1412 -1222
rect 1474 -1598 1508 -1222
rect 1570 -1598 1604 -1222
rect 1666 -1598 1700 -1222
rect 1762 -1598 1796 -1222
rect 1858 -1598 1892 -1222
rect 1954 -1598 1988 -1222
rect 2050 -1598 2084 -1222
rect 2450 80 2484 456
rect 2546 80 2580 456
rect 2642 80 2676 456
rect 2738 80 2772 456
rect 2834 80 2868 456
rect 2930 80 2964 456
rect 3026 80 3060 456
rect 3122 80 3156 456
rect 3218 80 3252 456
rect 3314 80 3348 456
rect 3410 80 3444 456
rect 3506 80 3540 456
rect 3602 80 3636 456
rect 3698 80 3732 456
rect 3794 80 3828 456
rect 3890 80 3924 456
rect 3986 80 4020 456
rect 4082 80 4116 456
rect 4178 80 4212 456
rect 4274 80 4308 456
rect 4370 80 4404 456
rect 2450 -538 2484 -162
rect 2546 -538 2580 -162
rect 2642 -538 2676 -162
rect 2738 -538 2772 -162
rect 2834 -538 2868 -162
rect 2930 -538 2964 -162
rect 3026 -538 3060 -162
rect 3122 -538 3156 -162
rect 3218 -538 3252 -162
rect 3314 -538 3348 -162
rect 3410 -538 3444 -162
rect 3506 -538 3540 -162
rect 3602 -538 3636 -162
rect 3698 -538 3732 -162
rect 3794 -538 3828 -162
rect 3890 -538 3924 -162
rect 3986 -538 4020 -162
rect 4082 -538 4116 -162
rect 4178 -538 4212 -162
rect 4274 -538 4308 -162
rect 4370 -538 4404 -162
rect -2450 -2742 -2416 -2366
rect -2354 -2742 -2320 -2366
rect -2258 -2742 -2224 -2366
rect -2162 -2742 -2128 -2366
rect -2066 -2742 -2032 -2366
rect -1970 -2742 -1936 -2366
rect -1874 -2742 -1840 -2366
rect -1778 -2742 -1744 -2366
rect -1682 -2742 -1648 -2366
rect -1586 -2742 -1552 -2366
rect -1490 -2742 -1456 -2366
rect -2450 -3360 -2416 -2984
rect -2354 -3360 -2320 -2984
rect -2258 -3360 -2224 -2984
rect -2162 -3360 -2128 -2984
rect -2066 -3360 -2032 -2984
rect -1970 -3360 -1936 -2984
rect -1874 -3360 -1840 -2984
rect -1778 -3360 -1744 -2984
rect -1682 -3360 -1648 -2984
rect -1586 -3360 -1552 -2984
rect -1490 -3360 -1456 -2984
rect -2450 -3978 -2416 -3602
rect -2354 -3978 -2320 -3602
rect -2258 -3978 -2224 -3602
rect -2162 -3978 -2128 -3602
rect -2066 -3978 -2032 -3602
rect -1970 -3978 -1936 -3602
rect -1874 -3978 -1840 -3602
rect -1778 -3978 -1744 -3602
rect -1682 -3978 -1648 -3602
rect -1586 -3978 -1552 -3602
rect -1490 -3978 -1456 -3602
rect -650 -2742 -616 -2366
rect -554 -2742 -520 -2366
rect -458 -2742 -424 -2366
rect -362 -2742 -328 -2366
rect -266 -2742 -232 -2366
rect -170 -2742 -136 -2366
rect -74 -2742 -40 -2366
rect 22 -2742 56 -2366
rect 118 -2742 152 -2366
rect 214 -2742 248 -2366
rect 310 -2742 344 -2366
rect -650 -3360 -616 -2984
rect -554 -3360 -520 -2984
rect -458 -3360 -424 -2984
rect -362 -3360 -328 -2984
rect -266 -3360 -232 -2984
rect -170 -3360 -136 -2984
rect -74 -3360 -40 -2984
rect 22 -3360 56 -2984
rect 118 -3360 152 -2984
rect 214 -3360 248 -2984
rect 310 -3360 344 -2984
rect -650 -3978 -616 -3602
rect -554 -3978 -520 -3602
rect -458 -3978 -424 -3602
rect -362 -3978 -328 -3602
rect -266 -3978 -232 -3602
rect -170 -3978 -136 -3602
rect -74 -3978 -40 -3602
rect 22 -3978 56 -3602
rect 118 -3978 152 -3602
rect 214 -3978 248 -3602
rect 310 -3978 344 -3602
rect 1150 -2742 1184 -2366
rect 1246 -2742 1280 -2366
rect 1342 -2742 1376 -2366
rect 1438 -2742 1472 -2366
rect 1534 -2742 1568 -2366
rect 1630 -2742 1664 -2366
rect 1726 -2742 1760 -2366
rect 1822 -2742 1856 -2366
rect 1918 -2742 1952 -2366
rect 2014 -2742 2048 -2366
rect 2110 -2742 2144 -2366
rect 1150 -3360 1184 -2984
rect 1246 -3360 1280 -2984
rect 1342 -3360 1376 -2984
rect 1438 -3360 1472 -2984
rect 1534 -3360 1568 -2984
rect 1630 -3360 1664 -2984
rect 1726 -3360 1760 -2984
rect 1822 -3360 1856 -2984
rect 1918 -3360 1952 -2984
rect 2014 -3360 2048 -2984
rect 2110 -3360 2144 -2984
rect 1150 -3978 1184 -3602
rect 1246 -3978 1280 -3602
rect 1342 -3978 1376 -3602
rect 1438 -3978 1472 -3602
rect 1534 -3978 1568 -3602
rect 1630 -3978 1664 -3602
rect 1726 -3978 1760 -3602
rect 1822 -3978 1856 -3602
rect 1918 -3978 1952 -3602
rect 2014 -3978 2048 -3602
rect 2110 -3978 2144 -3602
rect 2950 -2742 2984 -2366
rect 3046 -2742 3080 -2366
rect 3142 -2742 3176 -2366
rect 3238 -2742 3272 -2366
rect 3334 -2742 3368 -2366
rect 3430 -2742 3464 -2366
rect 3526 -2742 3560 -2366
rect 3622 -2742 3656 -2366
rect 3718 -2742 3752 -2366
rect 3814 -2742 3848 -2366
rect 3910 -2742 3944 -2366
rect 2950 -3360 2984 -2984
rect 3046 -3360 3080 -2984
rect 3142 -3360 3176 -2984
rect 3238 -3360 3272 -2984
rect 3334 -3360 3368 -2984
rect 3430 -3360 3464 -2984
rect 3526 -3360 3560 -2984
rect 3622 -3360 3656 -2984
rect 3718 -3360 3752 -2984
rect 3814 -3360 3848 -2984
rect 3910 -3360 3944 -2984
rect 2950 -3978 2984 -3602
rect 3046 -3978 3080 -3602
rect 3142 -3978 3176 -3602
rect 3238 -3978 3272 -3602
rect 3334 -3978 3368 -3602
rect 3430 -3978 3464 -3602
rect 3526 -3978 3560 -3602
rect 3622 -3978 3656 -3602
rect 3718 -3978 3752 -3602
rect 3814 -3978 3848 -3602
rect 3910 -3978 3944 -3602
rect 4950 1646 4984 2022
rect 5046 1646 5080 2022
rect 5142 1646 5176 2022
rect 5238 1646 5272 2022
rect 5334 1646 5368 2022
rect 5430 1646 5464 2022
rect 5526 1646 5560 2022
rect 5622 1646 5656 2022
rect 5718 1646 5752 2022
rect 5814 1646 5848 2022
rect 5910 1646 5944 2022
rect 6006 1646 6040 2022
rect 6102 1646 6136 2022
rect 6198 1646 6232 2022
rect 6294 1646 6328 2022
rect 6390 1646 6424 2022
rect 6486 1646 6520 2022
rect 6582 1646 6616 2022
rect 6678 1646 6712 2022
rect 6774 1646 6808 2022
rect 6870 1646 6904 2022
rect 4950 1028 4984 1404
rect 5046 1028 5080 1404
rect 5142 1028 5176 1404
rect 5238 1028 5272 1404
rect 5334 1028 5368 1404
rect 5430 1028 5464 1404
rect 5526 1028 5560 1404
rect 5622 1028 5656 1404
rect 5718 1028 5752 1404
rect 5814 1028 5848 1404
rect 5910 1028 5944 1404
rect 6006 1028 6040 1404
rect 6102 1028 6136 1404
rect 6198 1028 6232 1404
rect 6294 1028 6328 1404
rect 6390 1028 6424 1404
rect 6486 1028 6520 1404
rect 6582 1028 6616 1404
rect 6678 1028 6712 1404
rect 6774 1028 6808 1404
rect 6870 1028 6904 1404
rect 4950 410 4984 786
rect 5046 410 5080 786
rect 5142 410 5176 786
rect 5238 410 5272 786
rect 5334 410 5368 786
rect 5430 410 5464 786
rect 5526 410 5560 786
rect 5622 410 5656 786
rect 5718 410 5752 786
rect 5814 410 5848 786
rect 5910 410 5944 786
rect 6006 410 6040 786
rect 6102 410 6136 786
rect 6198 410 6232 786
rect 6294 410 6328 786
rect 6390 410 6424 786
rect 6486 410 6520 786
rect 6582 410 6616 786
rect 6678 410 6712 786
rect 6774 410 6808 786
rect 6870 410 6904 786
rect 4950 -208 4984 168
rect 5046 -208 5080 168
rect 5142 -208 5176 168
rect 5238 -208 5272 168
rect 5334 -208 5368 168
rect 5430 -208 5464 168
rect 5526 -208 5560 168
rect 5622 -208 5656 168
rect 5718 -208 5752 168
rect 5814 -208 5848 168
rect 5910 -208 5944 168
rect 6006 -208 6040 168
rect 6102 -208 6136 168
rect 6198 -208 6232 168
rect 6294 -208 6328 168
rect 6390 -208 6424 168
rect 6486 -208 6520 168
rect 6582 -208 6616 168
rect 6678 -208 6712 168
rect 6774 -208 6808 168
rect 6870 -208 6904 168
rect 4950 -826 4984 -450
rect 5046 -826 5080 -450
rect 5142 -826 5176 -450
rect 5238 -826 5272 -450
rect 5334 -826 5368 -450
rect 5430 -826 5464 -450
rect 5526 -826 5560 -450
rect 5622 -826 5656 -450
rect 5718 -826 5752 -450
rect 5814 -826 5848 -450
rect 5910 -826 5944 -450
rect 6006 -826 6040 -450
rect 6102 -826 6136 -450
rect 6198 -826 6232 -450
rect 6294 -826 6328 -450
rect 6390 -826 6424 -450
rect 6486 -826 6520 -450
rect 6582 -826 6616 -450
rect 6678 -826 6712 -450
rect 6774 -826 6808 -450
rect 6870 -826 6904 -450
rect 4950 -1444 4984 -1068
rect 5046 -1444 5080 -1068
rect 5142 -1444 5176 -1068
rect 5238 -1444 5272 -1068
rect 5334 -1444 5368 -1068
rect 5430 -1444 5464 -1068
rect 5526 -1444 5560 -1068
rect 5622 -1444 5656 -1068
rect 5718 -1444 5752 -1068
rect 5814 -1444 5848 -1068
rect 5910 -1444 5944 -1068
rect 6006 -1444 6040 -1068
rect 6102 -1444 6136 -1068
rect 6198 -1444 6232 -1068
rect 6294 -1444 6328 -1068
rect 6390 -1444 6424 -1068
rect 6486 -1444 6520 -1068
rect 6582 -1444 6616 -1068
rect 6678 -1444 6712 -1068
rect 6774 -1444 6808 -1068
rect 6870 -1444 6904 -1068
rect 4950 -2062 4984 -1686
rect 5046 -2062 5080 -1686
rect 5142 -2062 5176 -1686
rect 5238 -2062 5272 -1686
rect 5334 -2062 5368 -1686
rect 5430 -2062 5464 -1686
rect 5526 -2062 5560 -1686
rect 5622 -2062 5656 -1686
rect 5718 -2062 5752 -1686
rect 5814 -2062 5848 -1686
rect 5910 -2062 5944 -1686
rect 6006 -2062 6040 -1686
rect 6102 -2062 6136 -1686
rect 6198 -2062 6232 -1686
rect 6294 -2062 6328 -1686
rect 6390 -2062 6424 -1686
rect 6486 -2062 6520 -1686
rect 6582 -2062 6616 -1686
rect 6678 -2062 6712 -1686
rect 6774 -2062 6808 -1686
rect 6870 -2062 6904 -1686
rect 4950 -2680 4984 -2304
rect 5046 -2680 5080 -2304
rect 5142 -2680 5176 -2304
rect 5238 -2680 5272 -2304
rect 5334 -2680 5368 -2304
rect 5430 -2680 5464 -2304
rect 5526 -2680 5560 -2304
rect 5622 -2680 5656 -2304
rect 5718 -2680 5752 -2304
rect 5814 -2680 5848 -2304
rect 5910 -2680 5944 -2304
rect 6006 -2680 6040 -2304
rect 6102 -2680 6136 -2304
rect 6198 -2680 6232 -2304
rect 6294 -2680 6328 -2304
rect 6390 -2680 6424 -2304
rect 6486 -2680 6520 -2304
rect 6582 -2680 6616 -2304
rect 6678 -2680 6712 -2304
rect 6774 -2680 6808 -2304
rect 6870 -2680 6904 -2304
rect 4950 -3298 4984 -2922
rect 5046 -3298 5080 -2922
rect 5142 -3298 5176 -2922
rect 5238 -3298 5272 -2922
rect 5334 -3298 5368 -2922
rect 5430 -3298 5464 -2922
rect 5526 -3298 5560 -2922
rect 5622 -3298 5656 -2922
rect 5718 -3298 5752 -2922
rect 5814 -3298 5848 -2922
rect 5910 -3298 5944 -2922
rect 6006 -3298 6040 -2922
rect 6102 -3298 6136 -2922
rect 6198 -3298 6232 -2922
rect 6294 -3298 6328 -2922
rect 6390 -3298 6424 -2922
rect 6486 -3298 6520 -2922
rect 6582 -3298 6616 -2922
rect 6678 -3298 6712 -2922
rect 6774 -3298 6808 -2922
rect 6870 -3298 6904 -2922
rect -2450 -4888 -2416 -4512
rect -2192 -4888 -2158 -4512
rect -1934 -4888 -1900 -4512
rect -1676 -4888 -1642 -4512
rect -1418 -4888 -1384 -4512
rect -1160 -4888 -1126 -4512
rect -2450 -5506 -2416 -5130
rect -2192 -5506 -2158 -5130
rect -1934 -5506 -1900 -5130
rect -1676 -5506 -1642 -5130
rect -1418 -5506 -1384 -5130
rect -1160 -5506 -1126 -5130
rect -2450 -6124 -2416 -5748
rect -2192 -6124 -2158 -5748
rect -1934 -6124 -1900 -5748
rect -1676 -6124 -1642 -5748
rect -1418 -6124 -1384 -5748
rect -1160 -6124 -1126 -5748
rect -2450 -6742 -2416 -6366
rect -2192 -6742 -2158 -6366
rect -1934 -6742 -1900 -6366
rect -1676 -6742 -1642 -6366
rect -1418 -6742 -1384 -6366
rect -1160 -6742 -1126 -6366
rect -2450 -7360 -2416 -6984
rect -2192 -7360 -2158 -6984
rect -1934 -7360 -1900 -6984
rect -1676 -7360 -1642 -6984
rect -1418 -7360 -1384 -6984
rect -1160 -7360 -1126 -6984
rect -2450 -7978 -2416 -7602
rect -2192 -7978 -2158 -7602
rect -1934 -7978 -1900 -7602
rect -1676 -7978 -1642 -7602
rect -1418 -7978 -1384 -7602
rect -1160 -7978 -1126 -7602
rect -650 -4888 -616 -4512
rect -392 -4888 -358 -4512
rect -134 -4888 -100 -4512
rect 124 -4888 158 -4512
rect 382 -4888 416 -4512
rect 640 -4888 674 -4512
rect -650 -5506 -616 -5130
rect -392 -5506 -358 -5130
rect -134 -5506 -100 -5130
rect 124 -5506 158 -5130
rect 382 -5506 416 -5130
rect 640 -5506 674 -5130
rect -650 -6124 -616 -5748
rect -392 -6124 -358 -5748
rect -134 -6124 -100 -5748
rect 124 -6124 158 -5748
rect 382 -6124 416 -5748
rect 640 -6124 674 -5748
rect -650 -6742 -616 -6366
rect -392 -6742 -358 -6366
rect -134 -6742 -100 -6366
rect 124 -6742 158 -6366
rect 382 -6742 416 -6366
rect 640 -6742 674 -6366
rect -650 -7360 -616 -6984
rect -392 -7360 -358 -6984
rect -134 -7360 -100 -6984
rect 124 -7360 158 -6984
rect 382 -7360 416 -6984
rect 640 -7360 674 -6984
rect -650 -7978 -616 -7602
rect -392 -7978 -358 -7602
rect -134 -7978 -100 -7602
rect 124 -7978 158 -7602
rect 382 -7978 416 -7602
rect 640 -7978 674 -7602
rect 1150 -4888 1184 -4512
rect 1408 -4888 1442 -4512
rect 1666 -4888 1700 -4512
rect 1924 -4888 1958 -4512
rect 2182 -4888 2216 -4512
rect 2440 -4888 2474 -4512
rect 1150 -5506 1184 -5130
rect 1408 -5506 1442 -5130
rect 1666 -5506 1700 -5130
rect 1924 -5506 1958 -5130
rect 2182 -5506 2216 -5130
rect 2440 -5506 2474 -5130
rect 1150 -6124 1184 -5748
rect 1408 -6124 1442 -5748
rect 1666 -6124 1700 -5748
rect 1924 -6124 1958 -5748
rect 2182 -6124 2216 -5748
rect 2440 -6124 2474 -5748
rect 1150 -6742 1184 -6366
rect 1408 -6742 1442 -6366
rect 1666 -6742 1700 -6366
rect 1924 -6742 1958 -6366
rect 2182 -6742 2216 -6366
rect 2440 -6742 2474 -6366
rect 1150 -7360 1184 -6984
rect 1408 -7360 1442 -6984
rect 1666 -7360 1700 -6984
rect 1924 -7360 1958 -6984
rect 2182 -7360 2216 -6984
rect 2440 -7360 2474 -6984
rect 1150 -7978 1184 -7602
rect 1408 -7978 1442 -7602
rect 1666 -7978 1700 -7602
rect 1924 -7978 1958 -7602
rect 2182 -7978 2216 -7602
rect 2440 -7978 2474 -7602
rect 2950 -4888 2984 -4512
rect 3208 -4888 3242 -4512
rect 3466 -4888 3500 -4512
rect 3724 -4888 3758 -4512
rect 3982 -4888 4016 -4512
rect 4240 -4888 4274 -4512
rect 2950 -5506 2984 -5130
rect 3208 -5506 3242 -5130
rect 3466 -5506 3500 -5130
rect 3724 -5506 3758 -5130
rect 3982 -5506 4016 -5130
rect 4240 -5506 4274 -5130
rect 2950 -6124 2984 -5748
rect 3208 -6124 3242 -5748
rect 3466 -6124 3500 -5748
rect 3724 -6124 3758 -5748
rect 3982 -6124 4016 -5748
rect 4240 -6124 4274 -5748
rect 2950 -6742 2984 -6366
rect 3208 -6742 3242 -6366
rect 3466 -6742 3500 -6366
rect 3724 -6742 3758 -6366
rect 3982 -6742 4016 -6366
rect 4240 -6742 4274 -6366
rect 2950 -7360 2984 -6984
rect 3208 -7360 3242 -6984
rect 3466 -7360 3500 -6984
rect 3724 -7360 3758 -6984
rect 3982 -7360 4016 -6984
rect 4240 -7360 4274 -6984
rect 2950 -7978 2984 -7602
rect 3208 -7978 3242 -7602
rect 3466 -7978 3500 -7602
rect 3724 -7978 3758 -7602
rect 3982 -7978 4016 -7602
rect 4240 -7978 4274 -7602
<< pdiffc >>
rect 2450 1667 2484 2043
rect 2546 1667 2580 2043
rect 2642 1667 2676 2043
rect 2738 1667 2772 2043
rect 2834 1667 2868 2043
rect 2930 1667 2964 2043
rect 3026 1667 3060 2043
rect 3122 1667 3156 2043
rect 3218 1667 3252 2043
rect 3314 1667 3348 2043
rect 3410 1667 3444 2043
rect 3506 1667 3540 2043
rect 3602 1667 3636 2043
rect 3698 1667 3732 2043
rect 3794 1667 3828 2043
rect 3890 1667 3924 2043
rect 3986 1667 4020 2043
rect 4082 1667 4116 2043
rect 4178 1667 4212 2043
rect 4274 1667 4308 2043
rect 4370 1667 4404 2043
rect 2450 1031 2484 1407
rect 2546 1031 2580 1407
rect 2642 1031 2676 1407
rect 2738 1031 2772 1407
rect 2834 1031 2868 1407
rect 2930 1031 2964 1407
rect 3026 1031 3060 1407
rect 3122 1031 3156 1407
rect 3218 1031 3252 1407
rect 3314 1031 3348 1407
rect 3410 1031 3444 1407
rect 3506 1031 3540 1407
rect 3602 1031 3636 1407
rect 3698 1031 3732 1407
rect 3794 1031 3828 1407
rect 3890 1031 3924 1407
rect 3986 1031 4020 1407
rect 4082 1031 4116 1407
rect 4178 1031 4212 1407
rect 4274 1031 4308 1407
rect 4370 1031 4404 1407
<< psubdiff >>
rect -204 2206 -108 2240
rect 2132 2206 2228 2240
rect -204 2144 -170 2206
rect 2194 2144 2228 2206
rect -204 350 -170 412
rect 4836 2174 4932 2208
rect 6922 2174 7018 2208
rect 4836 2112 4870 2174
rect 2194 350 2228 412
rect -204 316 -108 350
rect 2132 316 2228 350
rect 2336 608 2432 642
rect 4422 608 4518 642
rect 2336 546 2370 608
rect 16 166 112 200
rect 2102 166 2198 200
rect 16 104 50 166
rect 2164 104 2198 166
rect 16 -1750 50 -1688
rect 4484 546 4518 608
rect 2336 -690 2370 -628
rect 4484 -690 4518 -628
rect 2336 -724 2432 -690
rect 4422 -724 4518 -690
rect 2164 -1750 2198 -1688
rect 16 -1784 112 -1750
rect 2102 -1784 2198 -1750
rect -2564 -2214 -2468 -2180
rect -1438 -2214 -1342 -2180
rect -2564 -2276 -2530 -2214
rect -1376 -2276 -1342 -2214
rect -2564 -4130 -2530 -4068
rect -1376 -4130 -1342 -4068
rect -2564 -4164 -2468 -4130
rect -1438 -4164 -1342 -4130
rect -764 -2214 -668 -2180
rect 362 -2214 458 -2180
rect -764 -2276 -730 -2214
rect 424 -2276 458 -2214
rect -764 -4130 -730 -4068
rect 424 -4130 458 -4068
rect -764 -4164 -668 -4130
rect 362 -4164 458 -4130
rect 1036 -2214 1132 -2180
rect 2162 -2214 2258 -2180
rect 1036 -2276 1070 -2214
rect 2224 -2276 2258 -2214
rect 1036 -4130 1070 -4068
rect 2224 -4130 2258 -4068
rect 1036 -4164 1132 -4130
rect 2162 -4164 2258 -4130
rect 2836 -2214 2932 -2180
rect 3962 -2214 4058 -2180
rect 2836 -2276 2870 -2214
rect 4024 -2276 4058 -2214
rect 2836 -4130 2870 -4068
rect 6984 2112 7018 2174
rect 4836 -3450 4870 -3388
rect 6984 -3450 7018 -3388
rect 4836 -3484 4932 -3450
rect 6922 -3484 7018 -3450
rect 4024 -4130 4058 -4068
rect 2836 -4164 2932 -4130
rect 3962 -4164 4058 -4130
rect -2564 -4360 -2468 -4326
rect -1108 -4360 -1012 -4326
rect -2564 -4422 -2530 -4360
rect -1046 -4422 -1012 -4360
rect -2564 -8130 -2530 -8068
rect -1046 -8130 -1012 -8068
rect -2564 -8164 -2468 -8130
rect -1108 -8164 -1012 -8130
rect -764 -4360 -668 -4326
rect 692 -4360 788 -4326
rect -764 -4422 -730 -4360
rect 754 -4422 788 -4360
rect -764 -8130 -730 -8068
rect 754 -8130 788 -8068
rect -764 -8164 -668 -8130
rect 692 -8164 788 -8130
rect 1036 -4360 1132 -4326
rect 2492 -4360 2588 -4326
rect 1036 -4422 1070 -4360
rect 2554 -4422 2588 -4360
rect 1036 -8130 1070 -8068
rect 2554 -8130 2588 -8068
rect 1036 -8164 1132 -8130
rect 2492 -8164 2588 -8130
rect 2836 -4360 2932 -4326
rect 4292 -4360 4388 -4326
rect 2836 -4422 2870 -4360
rect 4354 -4422 4388 -4360
rect 2836 -8130 2870 -8068
rect 4354 -8130 4388 -8068
rect 2836 -8164 2932 -8130
rect 4292 -8164 4388 -8130
rect -5468 -9416 -5444 -8610
rect -4636 -9416 -4612 -8610
<< nsubdiff >>
rect 2336 2204 2432 2238
rect 4422 2204 4518 2238
rect 2336 2142 2370 2204
rect 4484 2142 4518 2204
rect 2336 870 2370 932
rect 4484 870 4518 932
rect 2336 836 2432 870
rect 4422 836 4518 870
<< psubdiffcont >>
rect -108 2206 2132 2240
rect -204 412 -170 2144
rect 2194 412 2228 2144
rect 4932 2174 6922 2208
rect -108 316 2132 350
rect 2432 608 4422 642
rect 112 166 2102 200
rect 16 -1688 50 104
rect 2164 -1688 2198 104
rect 2336 -628 2370 546
rect 4484 -628 4518 546
rect 2432 -724 4422 -690
rect 112 -1784 2102 -1750
rect -2468 -2214 -1438 -2180
rect -2564 -4068 -2530 -2276
rect -1376 -4068 -1342 -2276
rect -2468 -4164 -1438 -4130
rect -668 -2214 362 -2180
rect -764 -4068 -730 -2276
rect 424 -4068 458 -2276
rect -668 -4164 362 -4130
rect 1132 -2214 2162 -2180
rect 1036 -4068 1070 -2276
rect 2224 -4068 2258 -2276
rect 1132 -4164 2162 -4130
rect 2932 -2214 3962 -2180
rect 2836 -4068 2870 -2276
rect 4024 -4068 4058 -2276
rect 4836 -3388 4870 2112
rect 6984 -3388 7018 2112
rect 4932 -3484 6922 -3450
rect 2932 -4164 3962 -4130
rect -2468 -4360 -1108 -4326
rect -2564 -8068 -2530 -4422
rect -1046 -8068 -1012 -4422
rect -2468 -8164 -1108 -8130
rect -668 -4360 692 -4326
rect -764 -8068 -730 -4422
rect 754 -8068 788 -4422
rect -668 -8164 692 -8130
rect 1132 -4360 2492 -4326
rect 1036 -8068 1070 -4422
rect 2554 -8068 2588 -4422
rect 1132 -8164 2492 -8130
rect 2932 -4360 4292 -4326
rect 2836 -8068 2870 -4422
rect 4354 -8068 4388 -4422
rect 2932 -8164 4292 -8130
rect -5444 -9416 -4636 -8610
<< nsubdiffcont >>
rect 2432 2204 4422 2238
rect 2336 932 2370 2142
rect 4484 932 4518 2142
rect 2432 836 4422 870
<< poly >>
rect 2482 2136 2548 2152
rect 2482 2102 2498 2136
rect 2532 2102 2548 2136
rect 2482 2086 2548 2102
rect 2674 2136 2740 2152
rect 2674 2102 2690 2136
rect 2724 2102 2740 2136
rect 2674 2086 2740 2102
rect 2866 2136 2932 2152
rect 2866 2102 2882 2136
rect 2916 2102 2932 2136
rect 2866 2086 2932 2102
rect 3058 2136 3124 2152
rect 3058 2102 3074 2136
rect 3108 2102 3124 2136
rect 3058 2086 3124 2102
rect 3250 2136 3316 2152
rect 3250 2102 3266 2136
rect 3300 2102 3316 2136
rect 3250 2086 3316 2102
rect 3442 2136 3508 2152
rect 3442 2102 3458 2136
rect 3492 2102 3508 2136
rect 3442 2086 3508 2102
rect 3634 2136 3700 2152
rect 3634 2102 3650 2136
rect 3684 2102 3700 2136
rect 3634 2086 3700 2102
rect 3826 2136 3892 2152
rect 3826 2102 3842 2136
rect 3876 2102 3892 2136
rect 3826 2086 3892 2102
rect 4018 2136 4084 2152
rect 4018 2102 4034 2136
rect 4068 2102 4084 2136
rect 4018 2086 4084 2102
rect 4210 2136 4276 2152
rect 4210 2102 4226 2136
rect 4260 2102 4276 2136
rect 4210 2086 4276 2102
rect 2500 2055 2530 2086
rect 2596 2055 2626 2081
rect 2692 2055 2722 2086
rect 2788 2055 2818 2081
rect 2884 2055 2914 2086
rect 2980 2055 3010 2081
rect 3076 2055 3106 2086
rect 3172 2055 3202 2081
rect 3268 2055 3298 2086
rect 3364 2055 3394 2081
rect 3460 2055 3490 2086
rect 3556 2055 3586 2081
rect 3652 2055 3682 2086
rect 3748 2055 3778 2081
rect 3844 2055 3874 2086
rect 3940 2055 3970 2081
rect 4036 2055 4066 2086
rect 4132 2055 4162 2081
rect 4228 2055 4258 2086
rect 4324 2055 4354 2081
rect 2500 1629 2530 1655
rect 2596 1624 2626 1655
rect 2692 1629 2722 1655
rect 2788 1624 2818 1655
rect 2884 1629 2914 1655
rect 2980 1624 3010 1655
rect 3076 1629 3106 1655
rect 3172 1624 3202 1655
rect 3268 1629 3298 1655
rect 3364 1624 3394 1655
rect 3460 1629 3490 1655
rect 3556 1624 3586 1655
rect 3652 1629 3682 1655
rect 3748 1624 3778 1655
rect 3844 1629 3874 1655
rect 3940 1624 3970 1655
rect 4036 1629 4066 1655
rect 4132 1624 4162 1655
rect 4228 1629 4258 1655
rect 4324 1624 4354 1655
rect 2578 1608 2644 1624
rect 2578 1574 2594 1608
rect 2628 1574 2644 1608
rect 2578 1558 2644 1574
rect 2770 1608 2836 1624
rect 2770 1574 2786 1608
rect 2820 1574 2836 1608
rect 2770 1558 2836 1574
rect 2962 1608 3028 1624
rect 2962 1574 2978 1608
rect 3012 1574 3028 1608
rect 2962 1558 3028 1574
rect 3154 1608 3220 1624
rect 3154 1574 3170 1608
rect 3204 1574 3220 1608
rect 3154 1558 3220 1574
rect 3346 1608 3412 1624
rect 3346 1574 3362 1608
rect 3396 1574 3412 1608
rect 3346 1558 3412 1574
rect 3538 1608 3604 1624
rect 3538 1574 3554 1608
rect 3588 1574 3604 1608
rect 3538 1558 3604 1574
rect 3730 1608 3796 1624
rect 3730 1574 3746 1608
rect 3780 1574 3796 1608
rect 3730 1558 3796 1574
rect 3922 1608 3988 1624
rect 3922 1574 3938 1608
rect 3972 1574 3988 1608
rect 3922 1558 3988 1574
rect 4114 1608 4180 1624
rect 4114 1574 4130 1608
rect 4164 1574 4180 1608
rect 4114 1558 4180 1574
rect 4306 1608 4372 1624
rect 4306 1574 4322 1608
rect 4356 1574 4372 1608
rect 4306 1558 4372 1574
rect 2578 1500 2644 1516
rect 2578 1466 2594 1500
rect 2628 1466 2644 1500
rect 2578 1450 2644 1466
rect 2770 1500 2836 1516
rect 2770 1466 2786 1500
rect 2820 1466 2836 1500
rect 2770 1450 2836 1466
rect 2962 1500 3028 1516
rect 2962 1466 2978 1500
rect 3012 1466 3028 1500
rect 2962 1450 3028 1466
rect 3154 1500 3220 1516
rect 3154 1466 3170 1500
rect 3204 1466 3220 1500
rect 3154 1450 3220 1466
rect 3346 1500 3412 1516
rect 3346 1466 3362 1500
rect 3396 1466 3412 1500
rect 3346 1450 3412 1466
rect 3538 1500 3604 1516
rect 3538 1466 3554 1500
rect 3588 1466 3604 1500
rect 3538 1450 3604 1466
rect 3730 1500 3796 1516
rect 3730 1466 3746 1500
rect 3780 1466 3796 1500
rect 3730 1450 3796 1466
rect 3922 1500 3988 1516
rect 3922 1466 3938 1500
rect 3972 1466 3988 1500
rect 3922 1450 3988 1466
rect 4114 1500 4180 1516
rect 4114 1466 4130 1500
rect 4164 1466 4180 1500
rect 4114 1450 4180 1466
rect 4306 1500 4372 1516
rect 4306 1466 4322 1500
rect 4356 1466 4372 1500
rect 4306 1450 4372 1466
rect 2500 1419 2530 1445
rect 2596 1419 2626 1450
rect 2692 1419 2722 1445
rect 2788 1419 2818 1450
rect 2884 1419 2914 1445
rect 2980 1419 3010 1450
rect 3076 1419 3106 1445
rect 3172 1419 3202 1450
rect 3268 1419 3298 1445
rect 3364 1419 3394 1450
rect 3460 1419 3490 1445
rect 3556 1419 3586 1450
rect 3652 1419 3682 1445
rect 3748 1419 3778 1450
rect 3844 1419 3874 1445
rect 3940 1419 3970 1450
rect 4036 1419 4066 1445
rect 4132 1419 4162 1450
rect 4228 1419 4258 1445
rect 4324 1419 4354 1450
rect 2500 988 2530 1019
rect 2596 993 2626 1019
rect 2692 988 2722 1019
rect 2788 993 2818 1019
rect 2884 988 2914 1019
rect 2980 993 3010 1019
rect 3076 988 3106 1019
rect 3172 993 3202 1019
rect 3268 988 3298 1019
rect 3364 993 3394 1019
rect 3460 988 3490 1019
rect 3556 993 3586 1019
rect 3652 988 3682 1019
rect 3748 993 3778 1019
rect 3844 988 3874 1019
rect 3940 993 3970 1019
rect 4036 988 4066 1019
rect 4132 993 4162 1019
rect 4228 988 4258 1019
rect 4324 993 4354 1019
rect 2482 972 2548 988
rect 2482 938 2498 972
rect 2532 938 2548 972
rect 2482 922 2548 938
rect 2674 972 2740 988
rect 2674 938 2690 972
rect 2724 938 2740 972
rect 2674 922 2740 938
rect 2866 972 2932 988
rect 2866 938 2882 972
rect 2916 938 2932 972
rect 2866 922 2932 938
rect 3058 972 3124 988
rect 3058 938 3074 972
rect 3108 938 3124 972
rect 3058 922 3124 938
rect 3250 972 3316 988
rect 3250 938 3266 972
rect 3300 938 3316 972
rect 3250 922 3316 938
rect 3442 972 3508 988
rect 3442 938 3458 972
rect 3492 938 3508 972
rect 3442 922 3508 938
rect 3634 972 3700 988
rect 3634 938 3650 972
rect 3684 938 3700 972
rect 3634 922 3700 938
rect 3826 972 3892 988
rect 3826 938 3842 972
rect 3876 938 3892 972
rect 3826 922 3892 938
rect 4018 972 4084 988
rect 4018 938 4034 972
rect 4068 938 4084 972
rect 4018 922 4084 938
rect 4210 972 4276 988
rect 4210 938 4226 972
rect 4260 938 4276 972
rect 4210 922 4276 938
rect 258 98 324 114
rect 258 64 274 98
rect 308 64 324 98
rect 180 26 210 52
rect 258 48 324 64
rect 450 98 516 114
rect 450 64 466 98
rect 500 64 516 98
rect 276 26 306 48
rect 372 26 402 52
rect 450 48 516 64
rect 642 98 708 114
rect 642 64 658 98
rect 692 64 708 98
rect 468 26 498 48
rect 564 26 594 52
rect 642 48 708 64
rect 834 98 900 114
rect 834 64 850 98
rect 884 64 900 98
rect 660 26 690 48
rect 756 26 786 52
rect 834 48 900 64
rect 1026 98 1092 114
rect 1026 64 1042 98
rect 1076 64 1092 98
rect 852 26 882 48
rect 948 26 978 52
rect 1026 48 1092 64
rect 1218 98 1284 114
rect 1218 64 1234 98
rect 1268 64 1284 98
rect 1044 26 1074 48
rect 1140 26 1170 52
rect 1218 48 1284 64
rect 1410 98 1476 114
rect 1410 64 1426 98
rect 1460 64 1476 98
rect 1236 26 1266 48
rect 1332 26 1362 52
rect 1410 48 1476 64
rect 1602 98 1668 114
rect 1602 64 1618 98
rect 1652 64 1668 98
rect 1428 26 1458 48
rect 1524 26 1554 52
rect 1602 48 1668 64
rect 1794 98 1860 114
rect 1794 64 1810 98
rect 1844 64 1860 98
rect 1620 26 1650 48
rect 1716 26 1746 52
rect 1794 48 1860 64
rect 1986 98 2052 114
rect 1986 64 2002 98
rect 2036 64 2052 98
rect 1812 26 1842 48
rect 1908 26 1938 52
rect 1986 48 2052 64
rect 2004 26 2034 48
rect 180 -396 210 -374
rect 162 -412 228 -396
rect 276 -400 306 -374
rect 372 -396 402 -374
rect 162 -446 178 -412
rect 212 -446 228 -412
rect 162 -462 228 -446
rect 354 -412 420 -396
rect 468 -400 498 -374
rect 564 -396 594 -374
rect 354 -446 370 -412
rect 404 -446 420 -412
rect 354 -462 420 -446
rect 546 -412 612 -396
rect 660 -400 690 -374
rect 756 -396 786 -374
rect 546 -446 562 -412
rect 596 -446 612 -412
rect 546 -462 612 -446
rect 738 -412 804 -396
rect 852 -400 882 -374
rect 948 -396 978 -374
rect 738 -446 754 -412
rect 788 -446 804 -412
rect 738 -462 804 -446
rect 930 -412 996 -396
rect 1044 -400 1074 -374
rect 1140 -396 1170 -374
rect 930 -446 946 -412
rect 980 -446 996 -412
rect 930 -462 996 -446
rect 1122 -412 1188 -396
rect 1236 -400 1266 -374
rect 1332 -396 1362 -374
rect 1122 -446 1138 -412
rect 1172 -446 1188 -412
rect 1122 -462 1188 -446
rect 1314 -412 1380 -396
rect 1428 -400 1458 -374
rect 1524 -396 1554 -374
rect 1314 -446 1330 -412
rect 1364 -446 1380 -412
rect 1314 -462 1380 -446
rect 1506 -412 1572 -396
rect 1620 -400 1650 -374
rect 1716 -396 1746 -374
rect 1506 -446 1522 -412
rect 1556 -446 1572 -412
rect 1506 -462 1572 -446
rect 1698 -412 1764 -396
rect 1812 -400 1842 -374
rect 1908 -396 1938 -374
rect 1698 -446 1714 -412
rect 1748 -446 1764 -412
rect 1698 -462 1764 -446
rect 1890 -412 1956 -396
rect 2004 -400 2034 -374
rect 1890 -446 1906 -412
rect 1940 -446 1956 -412
rect 1890 -462 1956 -446
rect 162 -520 228 -504
rect 162 -554 178 -520
rect 212 -554 228 -520
rect 162 -570 228 -554
rect 354 -520 420 -504
rect 354 -554 370 -520
rect 404 -554 420 -520
rect 180 -592 210 -570
rect 276 -592 306 -566
rect 354 -570 420 -554
rect 546 -520 612 -504
rect 546 -554 562 -520
rect 596 -554 612 -520
rect 372 -592 402 -570
rect 468 -592 498 -566
rect 546 -570 612 -554
rect 738 -520 804 -504
rect 738 -554 754 -520
rect 788 -554 804 -520
rect 564 -592 594 -570
rect 660 -592 690 -566
rect 738 -570 804 -554
rect 930 -520 996 -504
rect 930 -554 946 -520
rect 980 -554 996 -520
rect 756 -592 786 -570
rect 852 -592 882 -566
rect 930 -570 996 -554
rect 1122 -520 1188 -504
rect 1122 -554 1138 -520
rect 1172 -554 1188 -520
rect 948 -592 978 -570
rect 1044 -592 1074 -566
rect 1122 -570 1188 -554
rect 1314 -520 1380 -504
rect 1314 -554 1330 -520
rect 1364 -554 1380 -520
rect 1140 -592 1170 -570
rect 1236 -592 1266 -566
rect 1314 -570 1380 -554
rect 1506 -520 1572 -504
rect 1506 -554 1522 -520
rect 1556 -554 1572 -520
rect 1332 -592 1362 -570
rect 1428 -592 1458 -566
rect 1506 -570 1572 -554
rect 1698 -520 1764 -504
rect 1698 -554 1714 -520
rect 1748 -554 1764 -520
rect 1524 -592 1554 -570
rect 1620 -592 1650 -566
rect 1698 -570 1764 -554
rect 1890 -520 1956 -504
rect 1890 -554 1906 -520
rect 1940 -554 1956 -520
rect 1716 -592 1746 -570
rect 1812 -592 1842 -566
rect 1890 -570 1956 -554
rect 1908 -592 1938 -570
rect 2004 -592 2034 -566
rect 180 -1018 210 -992
rect 276 -1014 306 -992
rect 258 -1030 324 -1014
rect 372 -1018 402 -992
rect 468 -1014 498 -992
rect 258 -1064 274 -1030
rect 308 -1064 324 -1030
rect 258 -1080 324 -1064
rect 450 -1030 516 -1014
rect 564 -1018 594 -992
rect 660 -1014 690 -992
rect 450 -1064 466 -1030
rect 500 -1064 516 -1030
rect 450 -1080 516 -1064
rect 642 -1030 708 -1014
rect 756 -1018 786 -992
rect 852 -1014 882 -992
rect 642 -1064 658 -1030
rect 692 -1064 708 -1030
rect 642 -1080 708 -1064
rect 834 -1030 900 -1014
rect 948 -1018 978 -992
rect 1044 -1014 1074 -992
rect 834 -1064 850 -1030
rect 884 -1064 900 -1030
rect 834 -1080 900 -1064
rect 1026 -1030 1092 -1014
rect 1140 -1018 1170 -992
rect 1236 -1014 1266 -992
rect 1026 -1064 1042 -1030
rect 1076 -1064 1092 -1030
rect 1026 -1080 1092 -1064
rect 1218 -1030 1284 -1014
rect 1332 -1018 1362 -992
rect 1428 -1014 1458 -992
rect 1218 -1064 1234 -1030
rect 1268 -1064 1284 -1030
rect 1218 -1080 1284 -1064
rect 1410 -1030 1476 -1014
rect 1524 -1018 1554 -992
rect 1620 -1014 1650 -992
rect 1410 -1064 1426 -1030
rect 1460 -1064 1476 -1030
rect 1410 -1080 1476 -1064
rect 1602 -1030 1668 -1014
rect 1716 -1018 1746 -992
rect 1812 -1014 1842 -992
rect 1602 -1064 1618 -1030
rect 1652 -1064 1668 -1030
rect 1602 -1080 1668 -1064
rect 1794 -1030 1860 -1014
rect 1908 -1018 1938 -992
rect 2004 -1014 2034 -992
rect 1794 -1064 1810 -1030
rect 1844 -1064 1860 -1030
rect 1794 -1080 1860 -1064
rect 1986 -1030 2052 -1014
rect 1986 -1064 2002 -1030
rect 2036 -1064 2052 -1030
rect 1986 -1080 2052 -1064
rect 258 -1138 324 -1122
rect 258 -1172 274 -1138
rect 308 -1172 324 -1138
rect 180 -1210 210 -1184
rect 258 -1188 324 -1172
rect 450 -1138 516 -1122
rect 450 -1172 466 -1138
rect 500 -1172 516 -1138
rect 276 -1210 306 -1188
rect 372 -1210 402 -1184
rect 450 -1188 516 -1172
rect 642 -1138 708 -1122
rect 642 -1172 658 -1138
rect 692 -1172 708 -1138
rect 468 -1210 498 -1188
rect 564 -1210 594 -1184
rect 642 -1188 708 -1172
rect 834 -1138 900 -1122
rect 834 -1172 850 -1138
rect 884 -1172 900 -1138
rect 660 -1210 690 -1188
rect 756 -1210 786 -1184
rect 834 -1188 900 -1172
rect 1026 -1138 1092 -1122
rect 1026 -1172 1042 -1138
rect 1076 -1172 1092 -1138
rect 852 -1210 882 -1188
rect 948 -1210 978 -1184
rect 1026 -1188 1092 -1172
rect 1218 -1138 1284 -1122
rect 1218 -1172 1234 -1138
rect 1268 -1172 1284 -1138
rect 1044 -1210 1074 -1188
rect 1140 -1210 1170 -1184
rect 1218 -1188 1284 -1172
rect 1410 -1138 1476 -1122
rect 1410 -1172 1426 -1138
rect 1460 -1172 1476 -1138
rect 1236 -1210 1266 -1188
rect 1332 -1210 1362 -1184
rect 1410 -1188 1476 -1172
rect 1602 -1138 1668 -1122
rect 1602 -1172 1618 -1138
rect 1652 -1172 1668 -1138
rect 1428 -1210 1458 -1188
rect 1524 -1210 1554 -1184
rect 1602 -1188 1668 -1172
rect 1794 -1138 1860 -1122
rect 1794 -1172 1810 -1138
rect 1844 -1172 1860 -1138
rect 1620 -1210 1650 -1188
rect 1716 -1210 1746 -1184
rect 1794 -1188 1860 -1172
rect 1986 -1138 2052 -1122
rect 1986 -1172 2002 -1138
rect 2036 -1172 2052 -1138
rect 1812 -1210 1842 -1188
rect 1908 -1210 1938 -1184
rect 1986 -1188 2052 -1172
rect 2004 -1210 2034 -1188
rect 180 -1632 210 -1610
rect 162 -1648 228 -1632
rect 276 -1636 306 -1610
rect 372 -1632 402 -1610
rect 162 -1682 178 -1648
rect 212 -1682 228 -1648
rect 162 -1698 228 -1682
rect 354 -1648 420 -1632
rect 468 -1636 498 -1610
rect 564 -1632 594 -1610
rect 354 -1682 370 -1648
rect 404 -1682 420 -1648
rect 354 -1698 420 -1682
rect 546 -1648 612 -1632
rect 660 -1636 690 -1610
rect 756 -1632 786 -1610
rect 546 -1682 562 -1648
rect 596 -1682 612 -1648
rect 546 -1698 612 -1682
rect 738 -1648 804 -1632
rect 852 -1636 882 -1610
rect 948 -1632 978 -1610
rect 738 -1682 754 -1648
rect 788 -1682 804 -1648
rect 738 -1698 804 -1682
rect 930 -1648 996 -1632
rect 1044 -1636 1074 -1610
rect 1140 -1632 1170 -1610
rect 930 -1682 946 -1648
rect 980 -1682 996 -1648
rect 930 -1698 996 -1682
rect 1122 -1648 1188 -1632
rect 1236 -1636 1266 -1610
rect 1332 -1632 1362 -1610
rect 1122 -1682 1138 -1648
rect 1172 -1682 1188 -1648
rect 1122 -1698 1188 -1682
rect 1314 -1648 1380 -1632
rect 1428 -1636 1458 -1610
rect 1524 -1632 1554 -1610
rect 1314 -1682 1330 -1648
rect 1364 -1682 1380 -1648
rect 1314 -1698 1380 -1682
rect 1506 -1648 1572 -1632
rect 1620 -1636 1650 -1610
rect 1716 -1632 1746 -1610
rect 1506 -1682 1522 -1648
rect 1556 -1682 1572 -1648
rect 1506 -1698 1572 -1682
rect 1698 -1648 1764 -1632
rect 1812 -1636 1842 -1610
rect 1908 -1632 1938 -1610
rect 1698 -1682 1714 -1648
rect 1748 -1682 1764 -1648
rect 1698 -1698 1764 -1682
rect 1890 -1648 1956 -1632
rect 2004 -1636 2034 -1610
rect 1890 -1682 1906 -1648
rect 1940 -1682 1956 -1648
rect 1890 -1698 1956 -1682
rect 2482 540 2548 556
rect 2482 506 2498 540
rect 2532 506 2548 540
rect 2482 490 2548 506
rect 2674 540 2740 556
rect 2674 506 2690 540
rect 2724 506 2740 540
rect 2500 468 2530 490
rect 2596 468 2626 494
rect 2674 490 2740 506
rect 2866 540 2932 556
rect 2866 506 2882 540
rect 2916 506 2932 540
rect 2692 468 2722 490
rect 2788 468 2818 494
rect 2866 490 2932 506
rect 3058 540 3124 556
rect 3058 506 3074 540
rect 3108 506 3124 540
rect 2884 468 2914 490
rect 2980 468 3010 494
rect 3058 490 3124 506
rect 3250 540 3316 556
rect 3250 506 3266 540
rect 3300 506 3316 540
rect 3076 468 3106 490
rect 3172 468 3202 494
rect 3250 490 3316 506
rect 3442 540 3508 556
rect 3442 506 3458 540
rect 3492 506 3508 540
rect 3268 468 3298 490
rect 3364 468 3394 494
rect 3442 490 3508 506
rect 3634 540 3700 556
rect 3634 506 3650 540
rect 3684 506 3700 540
rect 3460 468 3490 490
rect 3556 468 3586 494
rect 3634 490 3700 506
rect 3826 540 3892 556
rect 3826 506 3842 540
rect 3876 506 3892 540
rect 3652 468 3682 490
rect 3748 468 3778 494
rect 3826 490 3892 506
rect 4018 540 4084 556
rect 4018 506 4034 540
rect 4068 506 4084 540
rect 3844 468 3874 490
rect 3940 468 3970 494
rect 4018 490 4084 506
rect 4210 540 4276 556
rect 4210 506 4226 540
rect 4260 506 4276 540
rect 4036 468 4066 490
rect 4132 468 4162 494
rect 4210 490 4276 506
rect 4228 468 4258 490
rect 4324 468 4354 494
rect 2500 42 2530 68
rect 2596 46 2626 68
rect 2578 30 2644 46
rect 2692 42 2722 68
rect 2788 46 2818 68
rect 2578 -4 2594 30
rect 2628 -4 2644 30
rect 2578 -20 2644 -4
rect 2770 30 2836 46
rect 2884 42 2914 68
rect 2980 46 3010 68
rect 2770 -4 2786 30
rect 2820 -4 2836 30
rect 2770 -20 2836 -4
rect 2962 30 3028 46
rect 3076 42 3106 68
rect 3172 46 3202 68
rect 2962 -4 2978 30
rect 3012 -4 3028 30
rect 2962 -20 3028 -4
rect 3154 30 3220 46
rect 3268 42 3298 68
rect 3364 46 3394 68
rect 3154 -4 3170 30
rect 3204 -4 3220 30
rect 3154 -20 3220 -4
rect 3346 30 3412 46
rect 3460 42 3490 68
rect 3556 46 3586 68
rect 3346 -4 3362 30
rect 3396 -4 3412 30
rect 3346 -20 3412 -4
rect 3538 30 3604 46
rect 3652 42 3682 68
rect 3748 46 3778 68
rect 3538 -4 3554 30
rect 3588 -4 3604 30
rect 3538 -20 3604 -4
rect 3730 30 3796 46
rect 3844 42 3874 68
rect 3940 46 3970 68
rect 3730 -4 3746 30
rect 3780 -4 3796 30
rect 3730 -20 3796 -4
rect 3922 30 3988 46
rect 4036 42 4066 68
rect 4132 46 4162 68
rect 3922 -4 3938 30
rect 3972 -4 3988 30
rect 3922 -20 3988 -4
rect 4114 30 4180 46
rect 4228 42 4258 68
rect 4324 46 4354 68
rect 4114 -4 4130 30
rect 4164 -4 4180 30
rect 4114 -20 4180 -4
rect 4306 30 4372 46
rect 4306 -4 4322 30
rect 4356 -4 4372 30
rect 4306 -20 4372 -4
rect 2578 -78 2644 -62
rect 2578 -112 2594 -78
rect 2628 -112 2644 -78
rect 2500 -150 2530 -124
rect 2578 -128 2644 -112
rect 2770 -78 2836 -62
rect 2770 -112 2786 -78
rect 2820 -112 2836 -78
rect 2596 -150 2626 -128
rect 2692 -150 2722 -124
rect 2770 -128 2836 -112
rect 2962 -78 3028 -62
rect 2962 -112 2978 -78
rect 3012 -112 3028 -78
rect 2788 -150 2818 -128
rect 2884 -150 2914 -124
rect 2962 -128 3028 -112
rect 3154 -78 3220 -62
rect 3154 -112 3170 -78
rect 3204 -112 3220 -78
rect 2980 -150 3010 -128
rect 3076 -150 3106 -124
rect 3154 -128 3220 -112
rect 3346 -78 3412 -62
rect 3346 -112 3362 -78
rect 3396 -112 3412 -78
rect 3172 -150 3202 -128
rect 3268 -150 3298 -124
rect 3346 -128 3412 -112
rect 3538 -78 3604 -62
rect 3538 -112 3554 -78
rect 3588 -112 3604 -78
rect 3364 -150 3394 -128
rect 3460 -150 3490 -124
rect 3538 -128 3604 -112
rect 3730 -78 3796 -62
rect 3730 -112 3746 -78
rect 3780 -112 3796 -78
rect 3556 -150 3586 -128
rect 3652 -150 3682 -124
rect 3730 -128 3796 -112
rect 3922 -78 3988 -62
rect 3922 -112 3938 -78
rect 3972 -112 3988 -78
rect 3748 -150 3778 -128
rect 3844 -150 3874 -124
rect 3922 -128 3988 -112
rect 4114 -78 4180 -62
rect 4114 -112 4130 -78
rect 4164 -112 4180 -78
rect 3940 -150 3970 -128
rect 4036 -150 4066 -124
rect 4114 -128 4180 -112
rect 4306 -78 4372 -62
rect 4306 -112 4322 -78
rect 4356 -112 4372 -78
rect 4132 -150 4162 -128
rect 4228 -150 4258 -124
rect 4306 -128 4372 -112
rect 4324 -150 4354 -128
rect 2500 -572 2530 -550
rect 2482 -588 2548 -572
rect 2596 -576 2626 -550
rect 2692 -572 2722 -550
rect 2482 -622 2498 -588
rect 2532 -622 2548 -588
rect 2482 -638 2548 -622
rect 2674 -588 2740 -572
rect 2788 -576 2818 -550
rect 2884 -572 2914 -550
rect 2674 -622 2690 -588
rect 2724 -622 2740 -588
rect 2674 -638 2740 -622
rect 2866 -588 2932 -572
rect 2980 -576 3010 -550
rect 3076 -572 3106 -550
rect 2866 -622 2882 -588
rect 2916 -622 2932 -588
rect 2866 -638 2932 -622
rect 3058 -588 3124 -572
rect 3172 -576 3202 -550
rect 3268 -572 3298 -550
rect 3058 -622 3074 -588
rect 3108 -622 3124 -588
rect 3058 -638 3124 -622
rect 3250 -588 3316 -572
rect 3364 -576 3394 -550
rect 3460 -572 3490 -550
rect 3250 -622 3266 -588
rect 3300 -622 3316 -588
rect 3250 -638 3316 -622
rect 3442 -588 3508 -572
rect 3556 -576 3586 -550
rect 3652 -572 3682 -550
rect 3442 -622 3458 -588
rect 3492 -622 3508 -588
rect 3442 -638 3508 -622
rect 3634 -588 3700 -572
rect 3748 -576 3778 -550
rect 3844 -572 3874 -550
rect 3634 -622 3650 -588
rect 3684 -622 3700 -588
rect 3634 -638 3700 -622
rect 3826 -588 3892 -572
rect 3940 -576 3970 -550
rect 4036 -572 4066 -550
rect 3826 -622 3842 -588
rect 3876 -622 3892 -588
rect 3826 -638 3892 -622
rect 4018 -588 4084 -572
rect 4132 -576 4162 -550
rect 4228 -572 4258 -550
rect 4018 -622 4034 -588
rect 4068 -622 4084 -588
rect 4018 -638 4084 -622
rect 4210 -588 4276 -572
rect 4324 -576 4354 -550
rect 4210 -622 4226 -588
rect 4260 -622 4276 -588
rect 4210 -638 4276 -622
rect -2322 -2282 -2256 -2266
rect -2322 -2316 -2306 -2282
rect -2272 -2316 -2256 -2282
rect -2400 -2354 -2370 -2328
rect -2322 -2332 -2256 -2316
rect -2130 -2282 -2064 -2266
rect -2130 -2316 -2114 -2282
rect -2080 -2316 -2064 -2282
rect -2304 -2354 -2274 -2332
rect -2208 -2354 -2178 -2328
rect -2130 -2332 -2064 -2316
rect -1938 -2282 -1872 -2266
rect -1938 -2316 -1922 -2282
rect -1888 -2316 -1872 -2282
rect -2112 -2354 -2082 -2332
rect -2016 -2354 -1986 -2328
rect -1938 -2332 -1872 -2316
rect -1746 -2282 -1680 -2266
rect -1746 -2316 -1730 -2282
rect -1696 -2316 -1680 -2282
rect -1920 -2354 -1890 -2332
rect -1824 -2354 -1794 -2328
rect -1746 -2332 -1680 -2316
rect -1554 -2282 -1488 -2266
rect -1554 -2316 -1538 -2282
rect -1504 -2316 -1488 -2282
rect -1728 -2354 -1698 -2332
rect -1632 -2354 -1602 -2328
rect -1554 -2332 -1488 -2316
rect -1536 -2354 -1506 -2332
rect -2400 -2776 -2370 -2754
rect -2418 -2792 -2352 -2776
rect -2304 -2780 -2274 -2754
rect -2208 -2776 -2178 -2754
rect -2418 -2826 -2402 -2792
rect -2368 -2826 -2352 -2792
rect -2418 -2842 -2352 -2826
rect -2226 -2792 -2160 -2776
rect -2112 -2780 -2082 -2754
rect -2016 -2776 -1986 -2754
rect -2226 -2826 -2210 -2792
rect -2176 -2826 -2160 -2792
rect -2226 -2842 -2160 -2826
rect -2034 -2792 -1968 -2776
rect -1920 -2780 -1890 -2754
rect -1824 -2776 -1794 -2754
rect -2034 -2826 -2018 -2792
rect -1984 -2826 -1968 -2792
rect -2034 -2842 -1968 -2826
rect -1842 -2792 -1776 -2776
rect -1728 -2780 -1698 -2754
rect -1632 -2776 -1602 -2754
rect -1842 -2826 -1826 -2792
rect -1792 -2826 -1776 -2792
rect -1842 -2842 -1776 -2826
rect -1650 -2792 -1584 -2776
rect -1536 -2780 -1506 -2754
rect -1650 -2826 -1634 -2792
rect -1600 -2826 -1584 -2792
rect -1650 -2842 -1584 -2826
rect -2418 -2900 -2352 -2884
rect -2418 -2934 -2402 -2900
rect -2368 -2934 -2352 -2900
rect -2418 -2950 -2352 -2934
rect -2226 -2900 -2160 -2884
rect -2226 -2934 -2210 -2900
rect -2176 -2934 -2160 -2900
rect -2400 -2972 -2370 -2950
rect -2304 -2972 -2274 -2946
rect -2226 -2950 -2160 -2934
rect -2034 -2900 -1968 -2884
rect -2034 -2934 -2018 -2900
rect -1984 -2934 -1968 -2900
rect -2208 -2972 -2178 -2950
rect -2112 -2972 -2082 -2946
rect -2034 -2950 -1968 -2934
rect -1842 -2900 -1776 -2884
rect -1842 -2934 -1826 -2900
rect -1792 -2934 -1776 -2900
rect -2016 -2972 -1986 -2950
rect -1920 -2972 -1890 -2946
rect -1842 -2950 -1776 -2934
rect -1650 -2900 -1584 -2884
rect -1650 -2934 -1634 -2900
rect -1600 -2934 -1584 -2900
rect -1824 -2972 -1794 -2950
rect -1728 -2972 -1698 -2946
rect -1650 -2950 -1584 -2934
rect -1632 -2972 -1602 -2950
rect -1536 -2972 -1506 -2946
rect -2400 -3398 -2370 -3372
rect -2304 -3394 -2274 -3372
rect -2322 -3410 -2256 -3394
rect -2208 -3398 -2178 -3372
rect -2112 -3394 -2082 -3372
rect -2322 -3444 -2306 -3410
rect -2272 -3444 -2256 -3410
rect -2322 -3460 -2256 -3444
rect -2130 -3410 -2064 -3394
rect -2016 -3398 -1986 -3372
rect -1920 -3394 -1890 -3372
rect -2130 -3444 -2114 -3410
rect -2080 -3444 -2064 -3410
rect -2130 -3460 -2064 -3444
rect -1938 -3410 -1872 -3394
rect -1824 -3398 -1794 -3372
rect -1728 -3394 -1698 -3372
rect -1938 -3444 -1922 -3410
rect -1888 -3444 -1872 -3410
rect -1938 -3460 -1872 -3444
rect -1746 -3410 -1680 -3394
rect -1632 -3398 -1602 -3372
rect -1536 -3394 -1506 -3372
rect -1746 -3444 -1730 -3410
rect -1696 -3444 -1680 -3410
rect -1746 -3460 -1680 -3444
rect -1554 -3410 -1488 -3394
rect -1554 -3444 -1538 -3410
rect -1504 -3444 -1488 -3410
rect -1554 -3460 -1488 -3444
rect -2322 -3518 -2256 -3502
rect -2322 -3552 -2306 -3518
rect -2272 -3552 -2256 -3518
rect -2400 -3590 -2370 -3564
rect -2322 -3568 -2256 -3552
rect -2130 -3518 -2064 -3502
rect -2130 -3552 -2114 -3518
rect -2080 -3552 -2064 -3518
rect -2304 -3590 -2274 -3568
rect -2208 -3590 -2178 -3564
rect -2130 -3568 -2064 -3552
rect -1938 -3518 -1872 -3502
rect -1938 -3552 -1922 -3518
rect -1888 -3552 -1872 -3518
rect -2112 -3590 -2082 -3568
rect -2016 -3590 -1986 -3564
rect -1938 -3568 -1872 -3552
rect -1746 -3518 -1680 -3502
rect -1746 -3552 -1730 -3518
rect -1696 -3552 -1680 -3518
rect -1920 -3590 -1890 -3568
rect -1824 -3590 -1794 -3564
rect -1746 -3568 -1680 -3552
rect -1554 -3518 -1488 -3502
rect -1554 -3552 -1538 -3518
rect -1504 -3552 -1488 -3518
rect -1728 -3590 -1698 -3568
rect -1632 -3590 -1602 -3564
rect -1554 -3568 -1488 -3552
rect -1536 -3590 -1506 -3568
rect -2400 -4012 -2370 -3990
rect -2418 -4028 -2352 -4012
rect -2304 -4016 -2274 -3990
rect -2208 -4012 -2178 -3990
rect -2418 -4062 -2402 -4028
rect -2368 -4062 -2352 -4028
rect -2418 -4078 -2352 -4062
rect -2226 -4028 -2160 -4012
rect -2112 -4016 -2082 -3990
rect -2016 -4012 -1986 -3990
rect -2226 -4062 -2210 -4028
rect -2176 -4062 -2160 -4028
rect -2226 -4078 -2160 -4062
rect -2034 -4028 -1968 -4012
rect -1920 -4016 -1890 -3990
rect -1824 -4012 -1794 -3990
rect -2034 -4062 -2018 -4028
rect -1984 -4062 -1968 -4028
rect -2034 -4078 -1968 -4062
rect -1842 -4028 -1776 -4012
rect -1728 -4016 -1698 -3990
rect -1632 -4012 -1602 -3990
rect -1842 -4062 -1826 -4028
rect -1792 -4062 -1776 -4028
rect -1842 -4078 -1776 -4062
rect -1650 -4028 -1584 -4012
rect -1536 -4016 -1506 -3990
rect -1650 -4062 -1634 -4028
rect -1600 -4062 -1584 -4028
rect -1650 -4078 -1584 -4062
rect -522 -2282 -456 -2266
rect -522 -2316 -506 -2282
rect -472 -2316 -456 -2282
rect -600 -2354 -570 -2328
rect -522 -2332 -456 -2316
rect -330 -2282 -264 -2266
rect -330 -2316 -314 -2282
rect -280 -2316 -264 -2282
rect -504 -2354 -474 -2332
rect -408 -2354 -378 -2328
rect -330 -2332 -264 -2316
rect -138 -2282 -72 -2266
rect -138 -2316 -122 -2282
rect -88 -2316 -72 -2282
rect -312 -2354 -282 -2332
rect -216 -2354 -186 -2328
rect -138 -2332 -72 -2316
rect 54 -2282 120 -2266
rect 54 -2316 70 -2282
rect 104 -2316 120 -2282
rect -120 -2354 -90 -2332
rect -24 -2354 6 -2328
rect 54 -2332 120 -2316
rect 246 -2282 312 -2266
rect 246 -2316 262 -2282
rect 296 -2316 312 -2282
rect 72 -2354 102 -2332
rect 168 -2354 198 -2328
rect 246 -2332 312 -2316
rect 264 -2354 294 -2332
rect -600 -2776 -570 -2754
rect -618 -2792 -552 -2776
rect -504 -2780 -474 -2754
rect -408 -2776 -378 -2754
rect -618 -2826 -602 -2792
rect -568 -2826 -552 -2792
rect -618 -2842 -552 -2826
rect -426 -2792 -360 -2776
rect -312 -2780 -282 -2754
rect -216 -2776 -186 -2754
rect -426 -2826 -410 -2792
rect -376 -2826 -360 -2792
rect -426 -2842 -360 -2826
rect -234 -2792 -168 -2776
rect -120 -2780 -90 -2754
rect -24 -2776 6 -2754
rect -234 -2826 -218 -2792
rect -184 -2826 -168 -2792
rect -234 -2842 -168 -2826
rect -42 -2792 24 -2776
rect 72 -2780 102 -2754
rect 168 -2776 198 -2754
rect -42 -2826 -26 -2792
rect 8 -2826 24 -2792
rect -42 -2842 24 -2826
rect 150 -2792 216 -2776
rect 264 -2780 294 -2754
rect 150 -2826 166 -2792
rect 200 -2826 216 -2792
rect 150 -2842 216 -2826
rect -618 -2900 -552 -2884
rect -618 -2934 -602 -2900
rect -568 -2934 -552 -2900
rect -618 -2950 -552 -2934
rect -426 -2900 -360 -2884
rect -426 -2934 -410 -2900
rect -376 -2934 -360 -2900
rect -600 -2972 -570 -2950
rect -504 -2972 -474 -2946
rect -426 -2950 -360 -2934
rect -234 -2900 -168 -2884
rect -234 -2934 -218 -2900
rect -184 -2934 -168 -2900
rect -408 -2972 -378 -2950
rect -312 -2972 -282 -2946
rect -234 -2950 -168 -2934
rect -42 -2900 24 -2884
rect -42 -2934 -26 -2900
rect 8 -2934 24 -2900
rect -216 -2972 -186 -2950
rect -120 -2972 -90 -2946
rect -42 -2950 24 -2934
rect 150 -2900 216 -2884
rect 150 -2934 166 -2900
rect 200 -2934 216 -2900
rect -24 -2972 6 -2950
rect 72 -2972 102 -2946
rect 150 -2950 216 -2934
rect 168 -2972 198 -2950
rect 264 -2972 294 -2946
rect -600 -3398 -570 -3372
rect -504 -3394 -474 -3372
rect -522 -3410 -456 -3394
rect -408 -3398 -378 -3372
rect -312 -3394 -282 -3372
rect -522 -3444 -506 -3410
rect -472 -3444 -456 -3410
rect -522 -3460 -456 -3444
rect -330 -3410 -264 -3394
rect -216 -3398 -186 -3372
rect -120 -3394 -90 -3372
rect -330 -3444 -314 -3410
rect -280 -3444 -264 -3410
rect -330 -3460 -264 -3444
rect -138 -3410 -72 -3394
rect -24 -3398 6 -3372
rect 72 -3394 102 -3372
rect -138 -3444 -122 -3410
rect -88 -3444 -72 -3410
rect -138 -3460 -72 -3444
rect 54 -3410 120 -3394
rect 168 -3398 198 -3372
rect 264 -3394 294 -3372
rect 54 -3444 70 -3410
rect 104 -3444 120 -3410
rect 54 -3460 120 -3444
rect 246 -3410 312 -3394
rect 246 -3444 262 -3410
rect 296 -3444 312 -3410
rect 246 -3460 312 -3444
rect -522 -3518 -456 -3502
rect -522 -3552 -506 -3518
rect -472 -3552 -456 -3518
rect -600 -3590 -570 -3564
rect -522 -3568 -456 -3552
rect -330 -3518 -264 -3502
rect -330 -3552 -314 -3518
rect -280 -3552 -264 -3518
rect -504 -3590 -474 -3568
rect -408 -3590 -378 -3564
rect -330 -3568 -264 -3552
rect -138 -3518 -72 -3502
rect -138 -3552 -122 -3518
rect -88 -3552 -72 -3518
rect -312 -3590 -282 -3568
rect -216 -3590 -186 -3564
rect -138 -3568 -72 -3552
rect 54 -3518 120 -3502
rect 54 -3552 70 -3518
rect 104 -3552 120 -3518
rect -120 -3590 -90 -3568
rect -24 -3590 6 -3564
rect 54 -3568 120 -3552
rect 246 -3518 312 -3502
rect 246 -3552 262 -3518
rect 296 -3552 312 -3518
rect 72 -3590 102 -3568
rect 168 -3590 198 -3564
rect 246 -3568 312 -3552
rect 264 -3590 294 -3568
rect -600 -4012 -570 -3990
rect -618 -4028 -552 -4012
rect -504 -4016 -474 -3990
rect -408 -4012 -378 -3990
rect -618 -4062 -602 -4028
rect -568 -4062 -552 -4028
rect -618 -4078 -552 -4062
rect -426 -4028 -360 -4012
rect -312 -4016 -282 -3990
rect -216 -4012 -186 -3990
rect -426 -4062 -410 -4028
rect -376 -4062 -360 -4028
rect -426 -4078 -360 -4062
rect -234 -4028 -168 -4012
rect -120 -4016 -90 -3990
rect -24 -4012 6 -3990
rect -234 -4062 -218 -4028
rect -184 -4062 -168 -4028
rect -234 -4078 -168 -4062
rect -42 -4028 24 -4012
rect 72 -4016 102 -3990
rect 168 -4012 198 -3990
rect -42 -4062 -26 -4028
rect 8 -4062 24 -4028
rect -42 -4078 24 -4062
rect 150 -4028 216 -4012
rect 264 -4016 294 -3990
rect 150 -4062 166 -4028
rect 200 -4062 216 -4028
rect 150 -4078 216 -4062
rect 1278 -2282 1344 -2266
rect 1278 -2316 1294 -2282
rect 1328 -2316 1344 -2282
rect 1200 -2354 1230 -2328
rect 1278 -2332 1344 -2316
rect 1470 -2282 1536 -2266
rect 1470 -2316 1486 -2282
rect 1520 -2316 1536 -2282
rect 1296 -2354 1326 -2332
rect 1392 -2354 1422 -2328
rect 1470 -2332 1536 -2316
rect 1662 -2282 1728 -2266
rect 1662 -2316 1678 -2282
rect 1712 -2316 1728 -2282
rect 1488 -2354 1518 -2332
rect 1584 -2354 1614 -2328
rect 1662 -2332 1728 -2316
rect 1854 -2282 1920 -2266
rect 1854 -2316 1870 -2282
rect 1904 -2316 1920 -2282
rect 1680 -2354 1710 -2332
rect 1776 -2354 1806 -2328
rect 1854 -2332 1920 -2316
rect 2046 -2282 2112 -2266
rect 2046 -2316 2062 -2282
rect 2096 -2316 2112 -2282
rect 1872 -2354 1902 -2332
rect 1968 -2354 1998 -2328
rect 2046 -2332 2112 -2316
rect 2064 -2354 2094 -2332
rect 1200 -2776 1230 -2754
rect 1182 -2792 1248 -2776
rect 1296 -2780 1326 -2754
rect 1392 -2776 1422 -2754
rect 1182 -2826 1198 -2792
rect 1232 -2826 1248 -2792
rect 1182 -2842 1248 -2826
rect 1374 -2792 1440 -2776
rect 1488 -2780 1518 -2754
rect 1584 -2776 1614 -2754
rect 1374 -2826 1390 -2792
rect 1424 -2826 1440 -2792
rect 1374 -2842 1440 -2826
rect 1566 -2792 1632 -2776
rect 1680 -2780 1710 -2754
rect 1776 -2776 1806 -2754
rect 1566 -2826 1582 -2792
rect 1616 -2826 1632 -2792
rect 1566 -2842 1632 -2826
rect 1758 -2792 1824 -2776
rect 1872 -2780 1902 -2754
rect 1968 -2776 1998 -2754
rect 1758 -2826 1774 -2792
rect 1808 -2826 1824 -2792
rect 1758 -2842 1824 -2826
rect 1950 -2792 2016 -2776
rect 2064 -2780 2094 -2754
rect 1950 -2826 1966 -2792
rect 2000 -2826 2016 -2792
rect 1950 -2842 2016 -2826
rect 1182 -2900 1248 -2884
rect 1182 -2934 1198 -2900
rect 1232 -2934 1248 -2900
rect 1182 -2950 1248 -2934
rect 1374 -2900 1440 -2884
rect 1374 -2934 1390 -2900
rect 1424 -2934 1440 -2900
rect 1200 -2972 1230 -2950
rect 1296 -2972 1326 -2946
rect 1374 -2950 1440 -2934
rect 1566 -2900 1632 -2884
rect 1566 -2934 1582 -2900
rect 1616 -2934 1632 -2900
rect 1392 -2972 1422 -2950
rect 1488 -2972 1518 -2946
rect 1566 -2950 1632 -2934
rect 1758 -2900 1824 -2884
rect 1758 -2934 1774 -2900
rect 1808 -2934 1824 -2900
rect 1584 -2972 1614 -2950
rect 1680 -2972 1710 -2946
rect 1758 -2950 1824 -2934
rect 1950 -2900 2016 -2884
rect 1950 -2934 1966 -2900
rect 2000 -2934 2016 -2900
rect 1776 -2972 1806 -2950
rect 1872 -2972 1902 -2946
rect 1950 -2950 2016 -2934
rect 1968 -2972 1998 -2950
rect 2064 -2972 2094 -2946
rect 1200 -3398 1230 -3372
rect 1296 -3394 1326 -3372
rect 1278 -3410 1344 -3394
rect 1392 -3398 1422 -3372
rect 1488 -3394 1518 -3372
rect 1278 -3444 1294 -3410
rect 1328 -3444 1344 -3410
rect 1278 -3460 1344 -3444
rect 1470 -3410 1536 -3394
rect 1584 -3398 1614 -3372
rect 1680 -3394 1710 -3372
rect 1470 -3444 1486 -3410
rect 1520 -3444 1536 -3410
rect 1470 -3460 1536 -3444
rect 1662 -3410 1728 -3394
rect 1776 -3398 1806 -3372
rect 1872 -3394 1902 -3372
rect 1662 -3444 1678 -3410
rect 1712 -3444 1728 -3410
rect 1662 -3460 1728 -3444
rect 1854 -3410 1920 -3394
rect 1968 -3398 1998 -3372
rect 2064 -3394 2094 -3372
rect 1854 -3444 1870 -3410
rect 1904 -3444 1920 -3410
rect 1854 -3460 1920 -3444
rect 2046 -3410 2112 -3394
rect 2046 -3444 2062 -3410
rect 2096 -3444 2112 -3410
rect 2046 -3460 2112 -3444
rect 1278 -3518 1344 -3502
rect 1278 -3552 1294 -3518
rect 1328 -3552 1344 -3518
rect 1200 -3590 1230 -3564
rect 1278 -3568 1344 -3552
rect 1470 -3518 1536 -3502
rect 1470 -3552 1486 -3518
rect 1520 -3552 1536 -3518
rect 1296 -3590 1326 -3568
rect 1392 -3590 1422 -3564
rect 1470 -3568 1536 -3552
rect 1662 -3518 1728 -3502
rect 1662 -3552 1678 -3518
rect 1712 -3552 1728 -3518
rect 1488 -3590 1518 -3568
rect 1584 -3590 1614 -3564
rect 1662 -3568 1728 -3552
rect 1854 -3518 1920 -3502
rect 1854 -3552 1870 -3518
rect 1904 -3552 1920 -3518
rect 1680 -3590 1710 -3568
rect 1776 -3590 1806 -3564
rect 1854 -3568 1920 -3552
rect 2046 -3518 2112 -3502
rect 2046 -3552 2062 -3518
rect 2096 -3552 2112 -3518
rect 1872 -3590 1902 -3568
rect 1968 -3590 1998 -3564
rect 2046 -3568 2112 -3552
rect 2064 -3590 2094 -3568
rect 1200 -4012 1230 -3990
rect 1182 -4028 1248 -4012
rect 1296 -4016 1326 -3990
rect 1392 -4012 1422 -3990
rect 1182 -4062 1198 -4028
rect 1232 -4062 1248 -4028
rect 1182 -4078 1248 -4062
rect 1374 -4028 1440 -4012
rect 1488 -4016 1518 -3990
rect 1584 -4012 1614 -3990
rect 1374 -4062 1390 -4028
rect 1424 -4062 1440 -4028
rect 1374 -4078 1440 -4062
rect 1566 -4028 1632 -4012
rect 1680 -4016 1710 -3990
rect 1776 -4012 1806 -3990
rect 1566 -4062 1582 -4028
rect 1616 -4062 1632 -4028
rect 1566 -4078 1632 -4062
rect 1758 -4028 1824 -4012
rect 1872 -4016 1902 -3990
rect 1968 -4012 1998 -3990
rect 1758 -4062 1774 -4028
rect 1808 -4062 1824 -4028
rect 1758 -4078 1824 -4062
rect 1950 -4028 2016 -4012
rect 2064 -4016 2094 -3990
rect 1950 -4062 1966 -4028
rect 2000 -4062 2016 -4028
rect 1950 -4078 2016 -4062
rect 3078 -2282 3144 -2266
rect 3078 -2316 3094 -2282
rect 3128 -2316 3144 -2282
rect 3000 -2354 3030 -2328
rect 3078 -2332 3144 -2316
rect 3270 -2282 3336 -2266
rect 3270 -2316 3286 -2282
rect 3320 -2316 3336 -2282
rect 3096 -2354 3126 -2332
rect 3192 -2354 3222 -2328
rect 3270 -2332 3336 -2316
rect 3462 -2282 3528 -2266
rect 3462 -2316 3478 -2282
rect 3512 -2316 3528 -2282
rect 3288 -2354 3318 -2332
rect 3384 -2354 3414 -2328
rect 3462 -2332 3528 -2316
rect 3654 -2282 3720 -2266
rect 3654 -2316 3670 -2282
rect 3704 -2316 3720 -2282
rect 3480 -2354 3510 -2332
rect 3576 -2354 3606 -2328
rect 3654 -2332 3720 -2316
rect 3846 -2282 3912 -2266
rect 3846 -2316 3862 -2282
rect 3896 -2316 3912 -2282
rect 3672 -2354 3702 -2332
rect 3768 -2354 3798 -2328
rect 3846 -2332 3912 -2316
rect 3864 -2354 3894 -2332
rect 3000 -2776 3030 -2754
rect 2982 -2792 3048 -2776
rect 3096 -2780 3126 -2754
rect 3192 -2776 3222 -2754
rect 2982 -2826 2998 -2792
rect 3032 -2826 3048 -2792
rect 2982 -2842 3048 -2826
rect 3174 -2792 3240 -2776
rect 3288 -2780 3318 -2754
rect 3384 -2776 3414 -2754
rect 3174 -2826 3190 -2792
rect 3224 -2826 3240 -2792
rect 3174 -2842 3240 -2826
rect 3366 -2792 3432 -2776
rect 3480 -2780 3510 -2754
rect 3576 -2776 3606 -2754
rect 3366 -2826 3382 -2792
rect 3416 -2826 3432 -2792
rect 3366 -2842 3432 -2826
rect 3558 -2792 3624 -2776
rect 3672 -2780 3702 -2754
rect 3768 -2776 3798 -2754
rect 3558 -2826 3574 -2792
rect 3608 -2826 3624 -2792
rect 3558 -2842 3624 -2826
rect 3750 -2792 3816 -2776
rect 3864 -2780 3894 -2754
rect 3750 -2826 3766 -2792
rect 3800 -2826 3816 -2792
rect 3750 -2842 3816 -2826
rect 2982 -2900 3048 -2884
rect 2982 -2934 2998 -2900
rect 3032 -2934 3048 -2900
rect 2982 -2950 3048 -2934
rect 3174 -2900 3240 -2884
rect 3174 -2934 3190 -2900
rect 3224 -2934 3240 -2900
rect 3000 -2972 3030 -2950
rect 3096 -2972 3126 -2946
rect 3174 -2950 3240 -2934
rect 3366 -2900 3432 -2884
rect 3366 -2934 3382 -2900
rect 3416 -2934 3432 -2900
rect 3192 -2972 3222 -2950
rect 3288 -2972 3318 -2946
rect 3366 -2950 3432 -2934
rect 3558 -2900 3624 -2884
rect 3558 -2934 3574 -2900
rect 3608 -2934 3624 -2900
rect 3384 -2972 3414 -2950
rect 3480 -2972 3510 -2946
rect 3558 -2950 3624 -2934
rect 3750 -2900 3816 -2884
rect 3750 -2934 3766 -2900
rect 3800 -2934 3816 -2900
rect 3576 -2972 3606 -2950
rect 3672 -2972 3702 -2946
rect 3750 -2950 3816 -2934
rect 3768 -2972 3798 -2950
rect 3864 -2972 3894 -2946
rect 3000 -3398 3030 -3372
rect 3096 -3394 3126 -3372
rect 3078 -3410 3144 -3394
rect 3192 -3398 3222 -3372
rect 3288 -3394 3318 -3372
rect 3078 -3444 3094 -3410
rect 3128 -3444 3144 -3410
rect 3078 -3460 3144 -3444
rect 3270 -3410 3336 -3394
rect 3384 -3398 3414 -3372
rect 3480 -3394 3510 -3372
rect 3270 -3444 3286 -3410
rect 3320 -3444 3336 -3410
rect 3270 -3460 3336 -3444
rect 3462 -3410 3528 -3394
rect 3576 -3398 3606 -3372
rect 3672 -3394 3702 -3372
rect 3462 -3444 3478 -3410
rect 3512 -3444 3528 -3410
rect 3462 -3460 3528 -3444
rect 3654 -3410 3720 -3394
rect 3768 -3398 3798 -3372
rect 3864 -3394 3894 -3372
rect 3654 -3444 3670 -3410
rect 3704 -3444 3720 -3410
rect 3654 -3460 3720 -3444
rect 3846 -3410 3912 -3394
rect 3846 -3444 3862 -3410
rect 3896 -3444 3912 -3410
rect 3846 -3460 3912 -3444
rect 3078 -3518 3144 -3502
rect 3078 -3552 3094 -3518
rect 3128 -3552 3144 -3518
rect 3000 -3590 3030 -3564
rect 3078 -3568 3144 -3552
rect 3270 -3518 3336 -3502
rect 3270 -3552 3286 -3518
rect 3320 -3552 3336 -3518
rect 3096 -3590 3126 -3568
rect 3192 -3590 3222 -3564
rect 3270 -3568 3336 -3552
rect 3462 -3518 3528 -3502
rect 3462 -3552 3478 -3518
rect 3512 -3552 3528 -3518
rect 3288 -3590 3318 -3568
rect 3384 -3590 3414 -3564
rect 3462 -3568 3528 -3552
rect 3654 -3518 3720 -3502
rect 3654 -3552 3670 -3518
rect 3704 -3552 3720 -3518
rect 3480 -3590 3510 -3568
rect 3576 -3590 3606 -3564
rect 3654 -3568 3720 -3552
rect 3846 -3518 3912 -3502
rect 3846 -3552 3862 -3518
rect 3896 -3552 3912 -3518
rect 3672 -3590 3702 -3568
rect 3768 -3590 3798 -3564
rect 3846 -3568 3912 -3552
rect 3864 -3590 3894 -3568
rect 3000 -4012 3030 -3990
rect 2982 -4028 3048 -4012
rect 3096 -4016 3126 -3990
rect 3192 -4012 3222 -3990
rect 2982 -4062 2998 -4028
rect 3032 -4062 3048 -4028
rect 2982 -4078 3048 -4062
rect 3174 -4028 3240 -4012
rect 3288 -4016 3318 -3990
rect 3384 -4012 3414 -3990
rect 3174 -4062 3190 -4028
rect 3224 -4062 3240 -4028
rect 3174 -4078 3240 -4062
rect 3366 -4028 3432 -4012
rect 3480 -4016 3510 -3990
rect 3576 -4012 3606 -3990
rect 3366 -4062 3382 -4028
rect 3416 -4062 3432 -4028
rect 3366 -4078 3432 -4062
rect 3558 -4028 3624 -4012
rect 3672 -4016 3702 -3990
rect 3768 -4012 3798 -3990
rect 3558 -4062 3574 -4028
rect 3608 -4062 3624 -4028
rect 3558 -4078 3624 -4062
rect 3750 -4028 3816 -4012
rect 3864 -4016 3894 -3990
rect 3750 -4062 3766 -4028
rect 3800 -4062 3816 -4028
rect 3750 -4078 3816 -4062
rect 5078 2106 5144 2122
rect 5078 2072 5094 2106
rect 5128 2072 5144 2106
rect 5000 2034 5030 2060
rect 5078 2056 5144 2072
rect 5270 2106 5336 2122
rect 5270 2072 5286 2106
rect 5320 2072 5336 2106
rect 5096 2034 5126 2056
rect 5192 2034 5222 2060
rect 5270 2056 5336 2072
rect 5462 2106 5528 2122
rect 5462 2072 5478 2106
rect 5512 2072 5528 2106
rect 5288 2034 5318 2056
rect 5384 2034 5414 2060
rect 5462 2056 5528 2072
rect 5654 2106 5720 2122
rect 5654 2072 5670 2106
rect 5704 2072 5720 2106
rect 5480 2034 5510 2056
rect 5576 2034 5606 2060
rect 5654 2056 5720 2072
rect 5846 2106 5912 2122
rect 5846 2072 5862 2106
rect 5896 2072 5912 2106
rect 5672 2034 5702 2056
rect 5768 2034 5798 2060
rect 5846 2056 5912 2072
rect 6038 2106 6104 2122
rect 6038 2072 6054 2106
rect 6088 2072 6104 2106
rect 5864 2034 5894 2056
rect 5960 2034 5990 2060
rect 6038 2056 6104 2072
rect 6230 2106 6296 2122
rect 6230 2072 6246 2106
rect 6280 2072 6296 2106
rect 6056 2034 6086 2056
rect 6152 2034 6182 2060
rect 6230 2056 6296 2072
rect 6422 2106 6488 2122
rect 6422 2072 6438 2106
rect 6472 2072 6488 2106
rect 6248 2034 6278 2056
rect 6344 2034 6374 2060
rect 6422 2056 6488 2072
rect 6614 2106 6680 2122
rect 6614 2072 6630 2106
rect 6664 2072 6680 2106
rect 6440 2034 6470 2056
rect 6536 2034 6566 2060
rect 6614 2056 6680 2072
rect 6806 2106 6872 2122
rect 6806 2072 6822 2106
rect 6856 2072 6872 2106
rect 6632 2034 6662 2056
rect 6728 2034 6758 2060
rect 6806 2056 6872 2072
rect 6824 2034 6854 2056
rect 5000 1612 5030 1634
rect 4982 1596 5048 1612
rect 5096 1608 5126 1634
rect 5192 1612 5222 1634
rect 4982 1562 4998 1596
rect 5032 1562 5048 1596
rect 4982 1546 5048 1562
rect 5174 1596 5240 1612
rect 5288 1608 5318 1634
rect 5384 1612 5414 1634
rect 5174 1562 5190 1596
rect 5224 1562 5240 1596
rect 5174 1546 5240 1562
rect 5366 1596 5432 1612
rect 5480 1608 5510 1634
rect 5576 1612 5606 1634
rect 5366 1562 5382 1596
rect 5416 1562 5432 1596
rect 5366 1546 5432 1562
rect 5558 1596 5624 1612
rect 5672 1608 5702 1634
rect 5768 1612 5798 1634
rect 5558 1562 5574 1596
rect 5608 1562 5624 1596
rect 5558 1546 5624 1562
rect 5750 1596 5816 1612
rect 5864 1608 5894 1634
rect 5960 1612 5990 1634
rect 5750 1562 5766 1596
rect 5800 1562 5816 1596
rect 5750 1546 5816 1562
rect 5942 1596 6008 1612
rect 6056 1608 6086 1634
rect 6152 1612 6182 1634
rect 5942 1562 5958 1596
rect 5992 1562 6008 1596
rect 5942 1546 6008 1562
rect 6134 1596 6200 1612
rect 6248 1608 6278 1634
rect 6344 1612 6374 1634
rect 6134 1562 6150 1596
rect 6184 1562 6200 1596
rect 6134 1546 6200 1562
rect 6326 1596 6392 1612
rect 6440 1608 6470 1634
rect 6536 1612 6566 1634
rect 6326 1562 6342 1596
rect 6376 1562 6392 1596
rect 6326 1546 6392 1562
rect 6518 1596 6584 1612
rect 6632 1608 6662 1634
rect 6728 1612 6758 1634
rect 6518 1562 6534 1596
rect 6568 1562 6584 1596
rect 6518 1546 6584 1562
rect 6710 1596 6776 1612
rect 6824 1608 6854 1634
rect 6710 1562 6726 1596
rect 6760 1562 6776 1596
rect 6710 1546 6776 1562
rect 4982 1488 5048 1504
rect 4982 1454 4998 1488
rect 5032 1454 5048 1488
rect 4982 1438 5048 1454
rect 5174 1488 5240 1504
rect 5174 1454 5190 1488
rect 5224 1454 5240 1488
rect 5000 1416 5030 1438
rect 5096 1416 5126 1442
rect 5174 1438 5240 1454
rect 5366 1488 5432 1504
rect 5366 1454 5382 1488
rect 5416 1454 5432 1488
rect 5192 1416 5222 1438
rect 5288 1416 5318 1442
rect 5366 1438 5432 1454
rect 5558 1488 5624 1504
rect 5558 1454 5574 1488
rect 5608 1454 5624 1488
rect 5384 1416 5414 1438
rect 5480 1416 5510 1442
rect 5558 1438 5624 1454
rect 5750 1488 5816 1504
rect 5750 1454 5766 1488
rect 5800 1454 5816 1488
rect 5576 1416 5606 1438
rect 5672 1416 5702 1442
rect 5750 1438 5816 1454
rect 5942 1488 6008 1504
rect 5942 1454 5958 1488
rect 5992 1454 6008 1488
rect 5768 1416 5798 1438
rect 5864 1416 5894 1442
rect 5942 1438 6008 1454
rect 6134 1488 6200 1504
rect 6134 1454 6150 1488
rect 6184 1454 6200 1488
rect 5960 1416 5990 1438
rect 6056 1416 6086 1442
rect 6134 1438 6200 1454
rect 6326 1488 6392 1504
rect 6326 1454 6342 1488
rect 6376 1454 6392 1488
rect 6152 1416 6182 1438
rect 6248 1416 6278 1442
rect 6326 1438 6392 1454
rect 6518 1488 6584 1504
rect 6518 1454 6534 1488
rect 6568 1454 6584 1488
rect 6344 1416 6374 1438
rect 6440 1416 6470 1442
rect 6518 1438 6584 1454
rect 6710 1488 6776 1504
rect 6710 1454 6726 1488
rect 6760 1454 6776 1488
rect 6536 1416 6566 1438
rect 6632 1416 6662 1442
rect 6710 1438 6776 1454
rect 6728 1416 6758 1438
rect 6824 1416 6854 1442
rect 5000 990 5030 1016
rect 5096 994 5126 1016
rect 5078 978 5144 994
rect 5192 990 5222 1016
rect 5288 994 5318 1016
rect 5078 944 5094 978
rect 5128 944 5144 978
rect 5078 928 5144 944
rect 5270 978 5336 994
rect 5384 990 5414 1016
rect 5480 994 5510 1016
rect 5270 944 5286 978
rect 5320 944 5336 978
rect 5270 928 5336 944
rect 5462 978 5528 994
rect 5576 990 5606 1016
rect 5672 994 5702 1016
rect 5462 944 5478 978
rect 5512 944 5528 978
rect 5462 928 5528 944
rect 5654 978 5720 994
rect 5768 990 5798 1016
rect 5864 994 5894 1016
rect 5654 944 5670 978
rect 5704 944 5720 978
rect 5654 928 5720 944
rect 5846 978 5912 994
rect 5960 990 5990 1016
rect 6056 994 6086 1016
rect 5846 944 5862 978
rect 5896 944 5912 978
rect 5846 928 5912 944
rect 6038 978 6104 994
rect 6152 990 6182 1016
rect 6248 994 6278 1016
rect 6038 944 6054 978
rect 6088 944 6104 978
rect 6038 928 6104 944
rect 6230 978 6296 994
rect 6344 990 6374 1016
rect 6440 994 6470 1016
rect 6230 944 6246 978
rect 6280 944 6296 978
rect 6230 928 6296 944
rect 6422 978 6488 994
rect 6536 990 6566 1016
rect 6632 994 6662 1016
rect 6422 944 6438 978
rect 6472 944 6488 978
rect 6422 928 6488 944
rect 6614 978 6680 994
rect 6728 990 6758 1016
rect 6824 994 6854 1016
rect 6614 944 6630 978
rect 6664 944 6680 978
rect 6614 928 6680 944
rect 6806 978 6872 994
rect 6806 944 6822 978
rect 6856 944 6872 978
rect 6806 928 6872 944
rect 5078 870 5144 886
rect 5078 836 5094 870
rect 5128 836 5144 870
rect 5000 798 5030 824
rect 5078 820 5144 836
rect 5270 870 5336 886
rect 5270 836 5286 870
rect 5320 836 5336 870
rect 5096 798 5126 820
rect 5192 798 5222 824
rect 5270 820 5336 836
rect 5462 870 5528 886
rect 5462 836 5478 870
rect 5512 836 5528 870
rect 5288 798 5318 820
rect 5384 798 5414 824
rect 5462 820 5528 836
rect 5654 870 5720 886
rect 5654 836 5670 870
rect 5704 836 5720 870
rect 5480 798 5510 820
rect 5576 798 5606 824
rect 5654 820 5720 836
rect 5846 870 5912 886
rect 5846 836 5862 870
rect 5896 836 5912 870
rect 5672 798 5702 820
rect 5768 798 5798 824
rect 5846 820 5912 836
rect 6038 870 6104 886
rect 6038 836 6054 870
rect 6088 836 6104 870
rect 5864 798 5894 820
rect 5960 798 5990 824
rect 6038 820 6104 836
rect 6230 870 6296 886
rect 6230 836 6246 870
rect 6280 836 6296 870
rect 6056 798 6086 820
rect 6152 798 6182 824
rect 6230 820 6296 836
rect 6422 870 6488 886
rect 6422 836 6438 870
rect 6472 836 6488 870
rect 6248 798 6278 820
rect 6344 798 6374 824
rect 6422 820 6488 836
rect 6614 870 6680 886
rect 6614 836 6630 870
rect 6664 836 6680 870
rect 6440 798 6470 820
rect 6536 798 6566 824
rect 6614 820 6680 836
rect 6806 870 6872 886
rect 6806 836 6822 870
rect 6856 836 6872 870
rect 6632 798 6662 820
rect 6728 798 6758 824
rect 6806 820 6872 836
rect 6824 798 6854 820
rect 5000 376 5030 398
rect 4982 360 5048 376
rect 5096 372 5126 398
rect 5192 376 5222 398
rect 4982 326 4998 360
rect 5032 326 5048 360
rect 4982 310 5048 326
rect 5174 360 5240 376
rect 5288 372 5318 398
rect 5384 376 5414 398
rect 5174 326 5190 360
rect 5224 326 5240 360
rect 5174 310 5240 326
rect 5366 360 5432 376
rect 5480 372 5510 398
rect 5576 376 5606 398
rect 5366 326 5382 360
rect 5416 326 5432 360
rect 5366 310 5432 326
rect 5558 360 5624 376
rect 5672 372 5702 398
rect 5768 376 5798 398
rect 5558 326 5574 360
rect 5608 326 5624 360
rect 5558 310 5624 326
rect 5750 360 5816 376
rect 5864 372 5894 398
rect 5960 376 5990 398
rect 5750 326 5766 360
rect 5800 326 5816 360
rect 5750 310 5816 326
rect 5942 360 6008 376
rect 6056 372 6086 398
rect 6152 376 6182 398
rect 5942 326 5958 360
rect 5992 326 6008 360
rect 5942 310 6008 326
rect 6134 360 6200 376
rect 6248 372 6278 398
rect 6344 376 6374 398
rect 6134 326 6150 360
rect 6184 326 6200 360
rect 6134 310 6200 326
rect 6326 360 6392 376
rect 6440 372 6470 398
rect 6536 376 6566 398
rect 6326 326 6342 360
rect 6376 326 6392 360
rect 6326 310 6392 326
rect 6518 360 6584 376
rect 6632 372 6662 398
rect 6728 376 6758 398
rect 6518 326 6534 360
rect 6568 326 6584 360
rect 6518 310 6584 326
rect 6710 360 6776 376
rect 6824 372 6854 398
rect 6710 326 6726 360
rect 6760 326 6776 360
rect 6710 310 6776 326
rect 4982 252 5048 268
rect 4982 218 4998 252
rect 5032 218 5048 252
rect 4982 202 5048 218
rect 5174 252 5240 268
rect 5174 218 5190 252
rect 5224 218 5240 252
rect 5000 180 5030 202
rect 5096 180 5126 206
rect 5174 202 5240 218
rect 5366 252 5432 268
rect 5366 218 5382 252
rect 5416 218 5432 252
rect 5192 180 5222 202
rect 5288 180 5318 206
rect 5366 202 5432 218
rect 5558 252 5624 268
rect 5558 218 5574 252
rect 5608 218 5624 252
rect 5384 180 5414 202
rect 5480 180 5510 206
rect 5558 202 5624 218
rect 5750 252 5816 268
rect 5750 218 5766 252
rect 5800 218 5816 252
rect 5576 180 5606 202
rect 5672 180 5702 206
rect 5750 202 5816 218
rect 5942 252 6008 268
rect 5942 218 5958 252
rect 5992 218 6008 252
rect 5768 180 5798 202
rect 5864 180 5894 206
rect 5942 202 6008 218
rect 6134 252 6200 268
rect 6134 218 6150 252
rect 6184 218 6200 252
rect 5960 180 5990 202
rect 6056 180 6086 206
rect 6134 202 6200 218
rect 6326 252 6392 268
rect 6326 218 6342 252
rect 6376 218 6392 252
rect 6152 180 6182 202
rect 6248 180 6278 206
rect 6326 202 6392 218
rect 6518 252 6584 268
rect 6518 218 6534 252
rect 6568 218 6584 252
rect 6344 180 6374 202
rect 6440 180 6470 206
rect 6518 202 6584 218
rect 6710 252 6776 268
rect 6710 218 6726 252
rect 6760 218 6776 252
rect 6536 180 6566 202
rect 6632 180 6662 206
rect 6710 202 6776 218
rect 6728 180 6758 202
rect 6824 180 6854 206
rect 5000 -246 5030 -220
rect 5096 -242 5126 -220
rect 5078 -258 5144 -242
rect 5192 -246 5222 -220
rect 5288 -242 5318 -220
rect 5078 -292 5094 -258
rect 5128 -292 5144 -258
rect 5078 -308 5144 -292
rect 5270 -258 5336 -242
rect 5384 -246 5414 -220
rect 5480 -242 5510 -220
rect 5270 -292 5286 -258
rect 5320 -292 5336 -258
rect 5270 -308 5336 -292
rect 5462 -258 5528 -242
rect 5576 -246 5606 -220
rect 5672 -242 5702 -220
rect 5462 -292 5478 -258
rect 5512 -292 5528 -258
rect 5462 -308 5528 -292
rect 5654 -258 5720 -242
rect 5768 -246 5798 -220
rect 5864 -242 5894 -220
rect 5654 -292 5670 -258
rect 5704 -292 5720 -258
rect 5654 -308 5720 -292
rect 5846 -258 5912 -242
rect 5960 -246 5990 -220
rect 6056 -242 6086 -220
rect 5846 -292 5862 -258
rect 5896 -292 5912 -258
rect 5846 -308 5912 -292
rect 6038 -258 6104 -242
rect 6152 -246 6182 -220
rect 6248 -242 6278 -220
rect 6038 -292 6054 -258
rect 6088 -292 6104 -258
rect 6038 -308 6104 -292
rect 6230 -258 6296 -242
rect 6344 -246 6374 -220
rect 6440 -242 6470 -220
rect 6230 -292 6246 -258
rect 6280 -292 6296 -258
rect 6230 -308 6296 -292
rect 6422 -258 6488 -242
rect 6536 -246 6566 -220
rect 6632 -242 6662 -220
rect 6422 -292 6438 -258
rect 6472 -292 6488 -258
rect 6422 -308 6488 -292
rect 6614 -258 6680 -242
rect 6728 -246 6758 -220
rect 6824 -242 6854 -220
rect 6614 -292 6630 -258
rect 6664 -292 6680 -258
rect 6614 -308 6680 -292
rect 6806 -258 6872 -242
rect 6806 -292 6822 -258
rect 6856 -292 6872 -258
rect 6806 -308 6872 -292
rect 5078 -366 5144 -350
rect 5078 -400 5094 -366
rect 5128 -400 5144 -366
rect 5000 -438 5030 -412
rect 5078 -416 5144 -400
rect 5270 -366 5336 -350
rect 5270 -400 5286 -366
rect 5320 -400 5336 -366
rect 5096 -438 5126 -416
rect 5192 -438 5222 -412
rect 5270 -416 5336 -400
rect 5462 -366 5528 -350
rect 5462 -400 5478 -366
rect 5512 -400 5528 -366
rect 5288 -438 5318 -416
rect 5384 -438 5414 -412
rect 5462 -416 5528 -400
rect 5654 -366 5720 -350
rect 5654 -400 5670 -366
rect 5704 -400 5720 -366
rect 5480 -438 5510 -416
rect 5576 -438 5606 -412
rect 5654 -416 5720 -400
rect 5846 -366 5912 -350
rect 5846 -400 5862 -366
rect 5896 -400 5912 -366
rect 5672 -438 5702 -416
rect 5768 -438 5798 -412
rect 5846 -416 5912 -400
rect 6038 -366 6104 -350
rect 6038 -400 6054 -366
rect 6088 -400 6104 -366
rect 5864 -438 5894 -416
rect 5960 -438 5990 -412
rect 6038 -416 6104 -400
rect 6230 -366 6296 -350
rect 6230 -400 6246 -366
rect 6280 -400 6296 -366
rect 6056 -438 6086 -416
rect 6152 -438 6182 -412
rect 6230 -416 6296 -400
rect 6422 -366 6488 -350
rect 6422 -400 6438 -366
rect 6472 -400 6488 -366
rect 6248 -438 6278 -416
rect 6344 -438 6374 -412
rect 6422 -416 6488 -400
rect 6614 -366 6680 -350
rect 6614 -400 6630 -366
rect 6664 -400 6680 -366
rect 6440 -438 6470 -416
rect 6536 -438 6566 -412
rect 6614 -416 6680 -400
rect 6806 -366 6872 -350
rect 6806 -400 6822 -366
rect 6856 -400 6872 -366
rect 6632 -438 6662 -416
rect 6728 -438 6758 -412
rect 6806 -416 6872 -400
rect 6824 -438 6854 -416
rect 5000 -860 5030 -838
rect 4982 -876 5048 -860
rect 5096 -864 5126 -838
rect 5192 -860 5222 -838
rect 4982 -910 4998 -876
rect 5032 -910 5048 -876
rect 4982 -926 5048 -910
rect 5174 -876 5240 -860
rect 5288 -864 5318 -838
rect 5384 -860 5414 -838
rect 5174 -910 5190 -876
rect 5224 -910 5240 -876
rect 5174 -926 5240 -910
rect 5366 -876 5432 -860
rect 5480 -864 5510 -838
rect 5576 -860 5606 -838
rect 5366 -910 5382 -876
rect 5416 -910 5432 -876
rect 5366 -926 5432 -910
rect 5558 -876 5624 -860
rect 5672 -864 5702 -838
rect 5768 -860 5798 -838
rect 5558 -910 5574 -876
rect 5608 -910 5624 -876
rect 5558 -926 5624 -910
rect 5750 -876 5816 -860
rect 5864 -864 5894 -838
rect 5960 -860 5990 -838
rect 5750 -910 5766 -876
rect 5800 -910 5816 -876
rect 5750 -926 5816 -910
rect 5942 -876 6008 -860
rect 6056 -864 6086 -838
rect 6152 -860 6182 -838
rect 5942 -910 5958 -876
rect 5992 -910 6008 -876
rect 5942 -926 6008 -910
rect 6134 -876 6200 -860
rect 6248 -864 6278 -838
rect 6344 -860 6374 -838
rect 6134 -910 6150 -876
rect 6184 -910 6200 -876
rect 6134 -926 6200 -910
rect 6326 -876 6392 -860
rect 6440 -864 6470 -838
rect 6536 -860 6566 -838
rect 6326 -910 6342 -876
rect 6376 -910 6392 -876
rect 6326 -926 6392 -910
rect 6518 -876 6584 -860
rect 6632 -864 6662 -838
rect 6728 -860 6758 -838
rect 6518 -910 6534 -876
rect 6568 -910 6584 -876
rect 6518 -926 6584 -910
rect 6710 -876 6776 -860
rect 6824 -864 6854 -838
rect 6710 -910 6726 -876
rect 6760 -910 6776 -876
rect 6710 -926 6776 -910
rect 4982 -984 5048 -968
rect 4982 -1018 4998 -984
rect 5032 -1018 5048 -984
rect 4982 -1034 5048 -1018
rect 5174 -984 5240 -968
rect 5174 -1018 5190 -984
rect 5224 -1018 5240 -984
rect 5000 -1056 5030 -1034
rect 5096 -1056 5126 -1030
rect 5174 -1034 5240 -1018
rect 5366 -984 5432 -968
rect 5366 -1018 5382 -984
rect 5416 -1018 5432 -984
rect 5192 -1056 5222 -1034
rect 5288 -1056 5318 -1030
rect 5366 -1034 5432 -1018
rect 5558 -984 5624 -968
rect 5558 -1018 5574 -984
rect 5608 -1018 5624 -984
rect 5384 -1056 5414 -1034
rect 5480 -1056 5510 -1030
rect 5558 -1034 5624 -1018
rect 5750 -984 5816 -968
rect 5750 -1018 5766 -984
rect 5800 -1018 5816 -984
rect 5576 -1056 5606 -1034
rect 5672 -1056 5702 -1030
rect 5750 -1034 5816 -1018
rect 5942 -984 6008 -968
rect 5942 -1018 5958 -984
rect 5992 -1018 6008 -984
rect 5768 -1056 5798 -1034
rect 5864 -1056 5894 -1030
rect 5942 -1034 6008 -1018
rect 6134 -984 6200 -968
rect 6134 -1018 6150 -984
rect 6184 -1018 6200 -984
rect 5960 -1056 5990 -1034
rect 6056 -1056 6086 -1030
rect 6134 -1034 6200 -1018
rect 6326 -984 6392 -968
rect 6326 -1018 6342 -984
rect 6376 -1018 6392 -984
rect 6152 -1056 6182 -1034
rect 6248 -1056 6278 -1030
rect 6326 -1034 6392 -1018
rect 6518 -984 6584 -968
rect 6518 -1018 6534 -984
rect 6568 -1018 6584 -984
rect 6344 -1056 6374 -1034
rect 6440 -1056 6470 -1030
rect 6518 -1034 6584 -1018
rect 6710 -984 6776 -968
rect 6710 -1018 6726 -984
rect 6760 -1018 6776 -984
rect 6536 -1056 6566 -1034
rect 6632 -1056 6662 -1030
rect 6710 -1034 6776 -1018
rect 6728 -1056 6758 -1034
rect 6824 -1056 6854 -1030
rect 5000 -1482 5030 -1456
rect 5096 -1478 5126 -1456
rect 5078 -1494 5144 -1478
rect 5192 -1482 5222 -1456
rect 5288 -1478 5318 -1456
rect 5078 -1528 5094 -1494
rect 5128 -1528 5144 -1494
rect 5078 -1544 5144 -1528
rect 5270 -1494 5336 -1478
rect 5384 -1482 5414 -1456
rect 5480 -1478 5510 -1456
rect 5270 -1528 5286 -1494
rect 5320 -1528 5336 -1494
rect 5270 -1544 5336 -1528
rect 5462 -1494 5528 -1478
rect 5576 -1482 5606 -1456
rect 5672 -1478 5702 -1456
rect 5462 -1528 5478 -1494
rect 5512 -1528 5528 -1494
rect 5462 -1544 5528 -1528
rect 5654 -1494 5720 -1478
rect 5768 -1482 5798 -1456
rect 5864 -1478 5894 -1456
rect 5654 -1528 5670 -1494
rect 5704 -1528 5720 -1494
rect 5654 -1544 5720 -1528
rect 5846 -1494 5912 -1478
rect 5960 -1482 5990 -1456
rect 6056 -1478 6086 -1456
rect 5846 -1528 5862 -1494
rect 5896 -1528 5912 -1494
rect 5846 -1544 5912 -1528
rect 6038 -1494 6104 -1478
rect 6152 -1482 6182 -1456
rect 6248 -1478 6278 -1456
rect 6038 -1528 6054 -1494
rect 6088 -1528 6104 -1494
rect 6038 -1544 6104 -1528
rect 6230 -1494 6296 -1478
rect 6344 -1482 6374 -1456
rect 6440 -1478 6470 -1456
rect 6230 -1528 6246 -1494
rect 6280 -1528 6296 -1494
rect 6230 -1544 6296 -1528
rect 6422 -1494 6488 -1478
rect 6536 -1482 6566 -1456
rect 6632 -1478 6662 -1456
rect 6422 -1528 6438 -1494
rect 6472 -1528 6488 -1494
rect 6422 -1544 6488 -1528
rect 6614 -1494 6680 -1478
rect 6728 -1482 6758 -1456
rect 6824 -1478 6854 -1456
rect 6614 -1528 6630 -1494
rect 6664 -1528 6680 -1494
rect 6614 -1544 6680 -1528
rect 6806 -1494 6872 -1478
rect 6806 -1528 6822 -1494
rect 6856 -1528 6872 -1494
rect 6806 -1544 6872 -1528
rect 5078 -1602 5144 -1586
rect 5078 -1636 5094 -1602
rect 5128 -1636 5144 -1602
rect 5000 -1674 5030 -1648
rect 5078 -1652 5144 -1636
rect 5270 -1602 5336 -1586
rect 5270 -1636 5286 -1602
rect 5320 -1636 5336 -1602
rect 5096 -1674 5126 -1652
rect 5192 -1674 5222 -1648
rect 5270 -1652 5336 -1636
rect 5462 -1602 5528 -1586
rect 5462 -1636 5478 -1602
rect 5512 -1636 5528 -1602
rect 5288 -1674 5318 -1652
rect 5384 -1674 5414 -1648
rect 5462 -1652 5528 -1636
rect 5654 -1602 5720 -1586
rect 5654 -1636 5670 -1602
rect 5704 -1636 5720 -1602
rect 5480 -1674 5510 -1652
rect 5576 -1674 5606 -1648
rect 5654 -1652 5720 -1636
rect 5846 -1602 5912 -1586
rect 5846 -1636 5862 -1602
rect 5896 -1636 5912 -1602
rect 5672 -1674 5702 -1652
rect 5768 -1674 5798 -1648
rect 5846 -1652 5912 -1636
rect 6038 -1602 6104 -1586
rect 6038 -1636 6054 -1602
rect 6088 -1636 6104 -1602
rect 5864 -1674 5894 -1652
rect 5960 -1674 5990 -1648
rect 6038 -1652 6104 -1636
rect 6230 -1602 6296 -1586
rect 6230 -1636 6246 -1602
rect 6280 -1636 6296 -1602
rect 6056 -1674 6086 -1652
rect 6152 -1674 6182 -1648
rect 6230 -1652 6296 -1636
rect 6422 -1602 6488 -1586
rect 6422 -1636 6438 -1602
rect 6472 -1636 6488 -1602
rect 6248 -1674 6278 -1652
rect 6344 -1674 6374 -1648
rect 6422 -1652 6488 -1636
rect 6614 -1602 6680 -1586
rect 6614 -1636 6630 -1602
rect 6664 -1636 6680 -1602
rect 6440 -1674 6470 -1652
rect 6536 -1674 6566 -1648
rect 6614 -1652 6680 -1636
rect 6806 -1602 6872 -1586
rect 6806 -1636 6822 -1602
rect 6856 -1636 6872 -1602
rect 6632 -1674 6662 -1652
rect 6728 -1674 6758 -1648
rect 6806 -1652 6872 -1636
rect 6824 -1674 6854 -1652
rect 5000 -2096 5030 -2074
rect 4982 -2112 5048 -2096
rect 5096 -2100 5126 -2074
rect 5192 -2096 5222 -2074
rect 4982 -2146 4998 -2112
rect 5032 -2146 5048 -2112
rect 4982 -2162 5048 -2146
rect 5174 -2112 5240 -2096
rect 5288 -2100 5318 -2074
rect 5384 -2096 5414 -2074
rect 5174 -2146 5190 -2112
rect 5224 -2146 5240 -2112
rect 5174 -2162 5240 -2146
rect 5366 -2112 5432 -2096
rect 5480 -2100 5510 -2074
rect 5576 -2096 5606 -2074
rect 5366 -2146 5382 -2112
rect 5416 -2146 5432 -2112
rect 5366 -2162 5432 -2146
rect 5558 -2112 5624 -2096
rect 5672 -2100 5702 -2074
rect 5768 -2096 5798 -2074
rect 5558 -2146 5574 -2112
rect 5608 -2146 5624 -2112
rect 5558 -2162 5624 -2146
rect 5750 -2112 5816 -2096
rect 5864 -2100 5894 -2074
rect 5960 -2096 5990 -2074
rect 5750 -2146 5766 -2112
rect 5800 -2146 5816 -2112
rect 5750 -2162 5816 -2146
rect 5942 -2112 6008 -2096
rect 6056 -2100 6086 -2074
rect 6152 -2096 6182 -2074
rect 5942 -2146 5958 -2112
rect 5992 -2146 6008 -2112
rect 5942 -2162 6008 -2146
rect 6134 -2112 6200 -2096
rect 6248 -2100 6278 -2074
rect 6344 -2096 6374 -2074
rect 6134 -2146 6150 -2112
rect 6184 -2146 6200 -2112
rect 6134 -2162 6200 -2146
rect 6326 -2112 6392 -2096
rect 6440 -2100 6470 -2074
rect 6536 -2096 6566 -2074
rect 6326 -2146 6342 -2112
rect 6376 -2146 6392 -2112
rect 6326 -2162 6392 -2146
rect 6518 -2112 6584 -2096
rect 6632 -2100 6662 -2074
rect 6728 -2096 6758 -2074
rect 6518 -2146 6534 -2112
rect 6568 -2146 6584 -2112
rect 6518 -2162 6584 -2146
rect 6710 -2112 6776 -2096
rect 6824 -2100 6854 -2074
rect 6710 -2146 6726 -2112
rect 6760 -2146 6776 -2112
rect 6710 -2162 6776 -2146
rect 4982 -2220 5048 -2204
rect 4982 -2254 4998 -2220
rect 5032 -2254 5048 -2220
rect 4982 -2270 5048 -2254
rect 5174 -2220 5240 -2204
rect 5174 -2254 5190 -2220
rect 5224 -2254 5240 -2220
rect 5000 -2292 5030 -2270
rect 5096 -2292 5126 -2266
rect 5174 -2270 5240 -2254
rect 5366 -2220 5432 -2204
rect 5366 -2254 5382 -2220
rect 5416 -2254 5432 -2220
rect 5192 -2292 5222 -2270
rect 5288 -2292 5318 -2266
rect 5366 -2270 5432 -2254
rect 5558 -2220 5624 -2204
rect 5558 -2254 5574 -2220
rect 5608 -2254 5624 -2220
rect 5384 -2292 5414 -2270
rect 5480 -2292 5510 -2266
rect 5558 -2270 5624 -2254
rect 5750 -2220 5816 -2204
rect 5750 -2254 5766 -2220
rect 5800 -2254 5816 -2220
rect 5576 -2292 5606 -2270
rect 5672 -2292 5702 -2266
rect 5750 -2270 5816 -2254
rect 5942 -2220 6008 -2204
rect 5942 -2254 5958 -2220
rect 5992 -2254 6008 -2220
rect 5768 -2292 5798 -2270
rect 5864 -2292 5894 -2266
rect 5942 -2270 6008 -2254
rect 6134 -2220 6200 -2204
rect 6134 -2254 6150 -2220
rect 6184 -2254 6200 -2220
rect 5960 -2292 5990 -2270
rect 6056 -2292 6086 -2266
rect 6134 -2270 6200 -2254
rect 6326 -2220 6392 -2204
rect 6326 -2254 6342 -2220
rect 6376 -2254 6392 -2220
rect 6152 -2292 6182 -2270
rect 6248 -2292 6278 -2266
rect 6326 -2270 6392 -2254
rect 6518 -2220 6584 -2204
rect 6518 -2254 6534 -2220
rect 6568 -2254 6584 -2220
rect 6344 -2292 6374 -2270
rect 6440 -2292 6470 -2266
rect 6518 -2270 6584 -2254
rect 6710 -2220 6776 -2204
rect 6710 -2254 6726 -2220
rect 6760 -2254 6776 -2220
rect 6536 -2292 6566 -2270
rect 6632 -2292 6662 -2266
rect 6710 -2270 6776 -2254
rect 6728 -2292 6758 -2270
rect 6824 -2292 6854 -2266
rect 5000 -2718 5030 -2692
rect 5096 -2714 5126 -2692
rect 5078 -2730 5144 -2714
rect 5192 -2718 5222 -2692
rect 5288 -2714 5318 -2692
rect 5078 -2764 5094 -2730
rect 5128 -2764 5144 -2730
rect 5078 -2780 5144 -2764
rect 5270 -2730 5336 -2714
rect 5384 -2718 5414 -2692
rect 5480 -2714 5510 -2692
rect 5270 -2764 5286 -2730
rect 5320 -2764 5336 -2730
rect 5270 -2780 5336 -2764
rect 5462 -2730 5528 -2714
rect 5576 -2718 5606 -2692
rect 5672 -2714 5702 -2692
rect 5462 -2764 5478 -2730
rect 5512 -2764 5528 -2730
rect 5462 -2780 5528 -2764
rect 5654 -2730 5720 -2714
rect 5768 -2718 5798 -2692
rect 5864 -2714 5894 -2692
rect 5654 -2764 5670 -2730
rect 5704 -2764 5720 -2730
rect 5654 -2780 5720 -2764
rect 5846 -2730 5912 -2714
rect 5960 -2718 5990 -2692
rect 6056 -2714 6086 -2692
rect 5846 -2764 5862 -2730
rect 5896 -2764 5912 -2730
rect 5846 -2780 5912 -2764
rect 6038 -2730 6104 -2714
rect 6152 -2718 6182 -2692
rect 6248 -2714 6278 -2692
rect 6038 -2764 6054 -2730
rect 6088 -2764 6104 -2730
rect 6038 -2780 6104 -2764
rect 6230 -2730 6296 -2714
rect 6344 -2718 6374 -2692
rect 6440 -2714 6470 -2692
rect 6230 -2764 6246 -2730
rect 6280 -2764 6296 -2730
rect 6230 -2780 6296 -2764
rect 6422 -2730 6488 -2714
rect 6536 -2718 6566 -2692
rect 6632 -2714 6662 -2692
rect 6422 -2764 6438 -2730
rect 6472 -2764 6488 -2730
rect 6422 -2780 6488 -2764
rect 6614 -2730 6680 -2714
rect 6728 -2718 6758 -2692
rect 6824 -2714 6854 -2692
rect 6614 -2764 6630 -2730
rect 6664 -2764 6680 -2730
rect 6614 -2780 6680 -2764
rect 6806 -2730 6872 -2714
rect 6806 -2764 6822 -2730
rect 6856 -2764 6872 -2730
rect 6806 -2780 6872 -2764
rect 5078 -2838 5144 -2822
rect 5078 -2872 5094 -2838
rect 5128 -2872 5144 -2838
rect 5000 -2910 5030 -2884
rect 5078 -2888 5144 -2872
rect 5270 -2838 5336 -2822
rect 5270 -2872 5286 -2838
rect 5320 -2872 5336 -2838
rect 5096 -2910 5126 -2888
rect 5192 -2910 5222 -2884
rect 5270 -2888 5336 -2872
rect 5462 -2838 5528 -2822
rect 5462 -2872 5478 -2838
rect 5512 -2872 5528 -2838
rect 5288 -2910 5318 -2888
rect 5384 -2910 5414 -2884
rect 5462 -2888 5528 -2872
rect 5654 -2838 5720 -2822
rect 5654 -2872 5670 -2838
rect 5704 -2872 5720 -2838
rect 5480 -2910 5510 -2888
rect 5576 -2910 5606 -2884
rect 5654 -2888 5720 -2872
rect 5846 -2838 5912 -2822
rect 5846 -2872 5862 -2838
rect 5896 -2872 5912 -2838
rect 5672 -2910 5702 -2888
rect 5768 -2910 5798 -2884
rect 5846 -2888 5912 -2872
rect 6038 -2838 6104 -2822
rect 6038 -2872 6054 -2838
rect 6088 -2872 6104 -2838
rect 5864 -2910 5894 -2888
rect 5960 -2910 5990 -2884
rect 6038 -2888 6104 -2872
rect 6230 -2838 6296 -2822
rect 6230 -2872 6246 -2838
rect 6280 -2872 6296 -2838
rect 6056 -2910 6086 -2888
rect 6152 -2910 6182 -2884
rect 6230 -2888 6296 -2872
rect 6422 -2838 6488 -2822
rect 6422 -2872 6438 -2838
rect 6472 -2872 6488 -2838
rect 6248 -2910 6278 -2888
rect 6344 -2910 6374 -2884
rect 6422 -2888 6488 -2872
rect 6614 -2838 6680 -2822
rect 6614 -2872 6630 -2838
rect 6664 -2872 6680 -2838
rect 6440 -2910 6470 -2888
rect 6536 -2910 6566 -2884
rect 6614 -2888 6680 -2872
rect 6806 -2838 6872 -2822
rect 6806 -2872 6822 -2838
rect 6856 -2872 6872 -2838
rect 6632 -2910 6662 -2888
rect 6728 -2910 6758 -2884
rect 6806 -2888 6872 -2872
rect 6824 -2910 6854 -2888
rect 5000 -3332 5030 -3310
rect 4982 -3348 5048 -3332
rect 5096 -3336 5126 -3310
rect 5192 -3332 5222 -3310
rect 4982 -3382 4998 -3348
rect 5032 -3382 5048 -3348
rect 4982 -3398 5048 -3382
rect 5174 -3348 5240 -3332
rect 5288 -3336 5318 -3310
rect 5384 -3332 5414 -3310
rect 5174 -3382 5190 -3348
rect 5224 -3382 5240 -3348
rect 5174 -3398 5240 -3382
rect 5366 -3348 5432 -3332
rect 5480 -3336 5510 -3310
rect 5576 -3332 5606 -3310
rect 5366 -3382 5382 -3348
rect 5416 -3382 5432 -3348
rect 5366 -3398 5432 -3382
rect 5558 -3348 5624 -3332
rect 5672 -3336 5702 -3310
rect 5768 -3332 5798 -3310
rect 5558 -3382 5574 -3348
rect 5608 -3382 5624 -3348
rect 5558 -3398 5624 -3382
rect 5750 -3348 5816 -3332
rect 5864 -3336 5894 -3310
rect 5960 -3332 5990 -3310
rect 5750 -3382 5766 -3348
rect 5800 -3382 5816 -3348
rect 5750 -3398 5816 -3382
rect 5942 -3348 6008 -3332
rect 6056 -3336 6086 -3310
rect 6152 -3332 6182 -3310
rect 5942 -3382 5958 -3348
rect 5992 -3382 6008 -3348
rect 5942 -3398 6008 -3382
rect 6134 -3348 6200 -3332
rect 6248 -3336 6278 -3310
rect 6344 -3332 6374 -3310
rect 6134 -3382 6150 -3348
rect 6184 -3382 6200 -3348
rect 6134 -3398 6200 -3382
rect 6326 -3348 6392 -3332
rect 6440 -3336 6470 -3310
rect 6536 -3332 6566 -3310
rect 6326 -3382 6342 -3348
rect 6376 -3382 6392 -3348
rect 6326 -3398 6392 -3382
rect 6518 -3348 6584 -3332
rect 6632 -3336 6662 -3310
rect 6728 -3332 6758 -3310
rect 6518 -3382 6534 -3348
rect 6568 -3382 6584 -3348
rect 6518 -3398 6584 -3382
rect 6710 -3348 6776 -3332
rect 6824 -3336 6854 -3310
rect 6710 -3382 6726 -3348
rect 6760 -3382 6776 -3348
rect 6710 -3398 6776 -3382
rect -2404 -4428 -2204 -4412
rect -2404 -4462 -2388 -4428
rect -2220 -4462 -2204 -4428
rect -2404 -4500 -2204 -4462
rect -2146 -4428 -1946 -4412
rect -2146 -4462 -2130 -4428
rect -1962 -4462 -1946 -4428
rect -2146 -4500 -1946 -4462
rect -1888 -4428 -1688 -4412
rect -1888 -4462 -1872 -4428
rect -1704 -4462 -1688 -4428
rect -1888 -4500 -1688 -4462
rect -1630 -4428 -1430 -4412
rect -1630 -4462 -1614 -4428
rect -1446 -4462 -1430 -4428
rect -1630 -4500 -1430 -4462
rect -1372 -4428 -1172 -4412
rect -1372 -4462 -1356 -4428
rect -1188 -4462 -1172 -4428
rect -1372 -4500 -1172 -4462
rect -2404 -4938 -2204 -4900
rect -2404 -4972 -2388 -4938
rect -2220 -4972 -2204 -4938
rect -2404 -4988 -2204 -4972
rect -2146 -4938 -1946 -4900
rect -2146 -4972 -2130 -4938
rect -1962 -4972 -1946 -4938
rect -2146 -4988 -1946 -4972
rect -1888 -4938 -1688 -4900
rect -1888 -4972 -1872 -4938
rect -1704 -4972 -1688 -4938
rect -1888 -4988 -1688 -4972
rect -1630 -4938 -1430 -4900
rect -1630 -4972 -1614 -4938
rect -1446 -4972 -1430 -4938
rect -1630 -4988 -1430 -4972
rect -1372 -4938 -1172 -4900
rect -1372 -4972 -1356 -4938
rect -1188 -4972 -1172 -4938
rect -1372 -4988 -1172 -4972
rect -2404 -5046 -2204 -5030
rect -2404 -5080 -2388 -5046
rect -2220 -5080 -2204 -5046
rect -2404 -5118 -2204 -5080
rect -2146 -5046 -1946 -5030
rect -2146 -5080 -2130 -5046
rect -1962 -5080 -1946 -5046
rect -2146 -5118 -1946 -5080
rect -1888 -5046 -1688 -5030
rect -1888 -5080 -1872 -5046
rect -1704 -5080 -1688 -5046
rect -1888 -5118 -1688 -5080
rect -1630 -5046 -1430 -5030
rect -1630 -5080 -1614 -5046
rect -1446 -5080 -1430 -5046
rect -1630 -5118 -1430 -5080
rect -1372 -5046 -1172 -5030
rect -1372 -5080 -1356 -5046
rect -1188 -5080 -1172 -5046
rect -1372 -5118 -1172 -5080
rect -2404 -5556 -2204 -5518
rect -2404 -5590 -2388 -5556
rect -2220 -5590 -2204 -5556
rect -2404 -5606 -2204 -5590
rect -2146 -5556 -1946 -5518
rect -2146 -5590 -2130 -5556
rect -1962 -5590 -1946 -5556
rect -2146 -5606 -1946 -5590
rect -1888 -5556 -1688 -5518
rect -1888 -5590 -1872 -5556
rect -1704 -5590 -1688 -5556
rect -1888 -5606 -1688 -5590
rect -1630 -5556 -1430 -5518
rect -1630 -5590 -1614 -5556
rect -1446 -5590 -1430 -5556
rect -1630 -5606 -1430 -5590
rect -1372 -5556 -1172 -5518
rect -1372 -5590 -1356 -5556
rect -1188 -5590 -1172 -5556
rect -1372 -5606 -1172 -5590
rect -2404 -5664 -2204 -5648
rect -2404 -5698 -2388 -5664
rect -2220 -5698 -2204 -5664
rect -2404 -5736 -2204 -5698
rect -2146 -5664 -1946 -5648
rect -2146 -5698 -2130 -5664
rect -1962 -5698 -1946 -5664
rect -2146 -5736 -1946 -5698
rect -1888 -5664 -1688 -5648
rect -1888 -5698 -1872 -5664
rect -1704 -5698 -1688 -5664
rect -1888 -5736 -1688 -5698
rect -1630 -5664 -1430 -5648
rect -1630 -5698 -1614 -5664
rect -1446 -5698 -1430 -5664
rect -1630 -5736 -1430 -5698
rect -1372 -5664 -1172 -5648
rect -1372 -5698 -1356 -5664
rect -1188 -5698 -1172 -5664
rect -1372 -5736 -1172 -5698
rect -2404 -6174 -2204 -6136
rect -2404 -6208 -2388 -6174
rect -2220 -6208 -2204 -6174
rect -2404 -6224 -2204 -6208
rect -2146 -6174 -1946 -6136
rect -2146 -6208 -2130 -6174
rect -1962 -6208 -1946 -6174
rect -2146 -6224 -1946 -6208
rect -1888 -6174 -1688 -6136
rect -1888 -6208 -1872 -6174
rect -1704 -6208 -1688 -6174
rect -1888 -6224 -1688 -6208
rect -1630 -6174 -1430 -6136
rect -1630 -6208 -1614 -6174
rect -1446 -6208 -1430 -6174
rect -1630 -6224 -1430 -6208
rect -1372 -6174 -1172 -6136
rect -1372 -6208 -1356 -6174
rect -1188 -6208 -1172 -6174
rect -1372 -6224 -1172 -6208
rect -2404 -6282 -2204 -6266
rect -2404 -6316 -2388 -6282
rect -2220 -6316 -2204 -6282
rect -2404 -6354 -2204 -6316
rect -2146 -6282 -1946 -6266
rect -2146 -6316 -2130 -6282
rect -1962 -6316 -1946 -6282
rect -2146 -6354 -1946 -6316
rect -1888 -6282 -1688 -6266
rect -1888 -6316 -1872 -6282
rect -1704 -6316 -1688 -6282
rect -1888 -6354 -1688 -6316
rect -1630 -6282 -1430 -6266
rect -1630 -6316 -1614 -6282
rect -1446 -6316 -1430 -6282
rect -1630 -6354 -1430 -6316
rect -1372 -6282 -1172 -6266
rect -1372 -6316 -1356 -6282
rect -1188 -6316 -1172 -6282
rect -1372 -6354 -1172 -6316
rect -2404 -6792 -2204 -6754
rect -2404 -6826 -2388 -6792
rect -2220 -6826 -2204 -6792
rect -2404 -6842 -2204 -6826
rect -2146 -6792 -1946 -6754
rect -2146 -6826 -2130 -6792
rect -1962 -6826 -1946 -6792
rect -2146 -6842 -1946 -6826
rect -1888 -6792 -1688 -6754
rect -1888 -6826 -1872 -6792
rect -1704 -6826 -1688 -6792
rect -1888 -6842 -1688 -6826
rect -1630 -6792 -1430 -6754
rect -1630 -6826 -1614 -6792
rect -1446 -6826 -1430 -6792
rect -1630 -6842 -1430 -6826
rect -1372 -6792 -1172 -6754
rect -1372 -6826 -1356 -6792
rect -1188 -6826 -1172 -6792
rect -1372 -6842 -1172 -6826
rect -2404 -6900 -2204 -6884
rect -2404 -6934 -2388 -6900
rect -2220 -6934 -2204 -6900
rect -2404 -6972 -2204 -6934
rect -2146 -6900 -1946 -6884
rect -2146 -6934 -2130 -6900
rect -1962 -6934 -1946 -6900
rect -2146 -6972 -1946 -6934
rect -1888 -6900 -1688 -6884
rect -1888 -6934 -1872 -6900
rect -1704 -6934 -1688 -6900
rect -1888 -6972 -1688 -6934
rect -1630 -6900 -1430 -6884
rect -1630 -6934 -1614 -6900
rect -1446 -6934 -1430 -6900
rect -1630 -6972 -1430 -6934
rect -1372 -6900 -1172 -6884
rect -1372 -6934 -1356 -6900
rect -1188 -6934 -1172 -6900
rect -1372 -6972 -1172 -6934
rect -2404 -7410 -2204 -7372
rect -2404 -7444 -2388 -7410
rect -2220 -7444 -2204 -7410
rect -2404 -7460 -2204 -7444
rect -2146 -7410 -1946 -7372
rect -2146 -7444 -2130 -7410
rect -1962 -7444 -1946 -7410
rect -2146 -7460 -1946 -7444
rect -1888 -7410 -1688 -7372
rect -1888 -7444 -1872 -7410
rect -1704 -7444 -1688 -7410
rect -1888 -7460 -1688 -7444
rect -1630 -7410 -1430 -7372
rect -1630 -7444 -1614 -7410
rect -1446 -7444 -1430 -7410
rect -1630 -7460 -1430 -7444
rect -1372 -7410 -1172 -7372
rect -1372 -7444 -1356 -7410
rect -1188 -7444 -1172 -7410
rect -1372 -7460 -1172 -7444
rect -2404 -7518 -2204 -7502
rect -2404 -7552 -2388 -7518
rect -2220 -7552 -2204 -7518
rect -2404 -7590 -2204 -7552
rect -2146 -7518 -1946 -7502
rect -2146 -7552 -2130 -7518
rect -1962 -7552 -1946 -7518
rect -2146 -7590 -1946 -7552
rect -1888 -7518 -1688 -7502
rect -1888 -7552 -1872 -7518
rect -1704 -7552 -1688 -7518
rect -1888 -7590 -1688 -7552
rect -1630 -7518 -1430 -7502
rect -1630 -7552 -1614 -7518
rect -1446 -7552 -1430 -7518
rect -1630 -7590 -1430 -7552
rect -1372 -7518 -1172 -7502
rect -1372 -7552 -1356 -7518
rect -1188 -7552 -1172 -7518
rect -1372 -7590 -1172 -7552
rect -2404 -8028 -2204 -7990
rect -2404 -8062 -2388 -8028
rect -2220 -8062 -2204 -8028
rect -2404 -8078 -2204 -8062
rect -2146 -8028 -1946 -7990
rect -2146 -8062 -2130 -8028
rect -1962 -8062 -1946 -8028
rect -2146 -8078 -1946 -8062
rect -1888 -8028 -1688 -7990
rect -1888 -8062 -1872 -8028
rect -1704 -8062 -1688 -8028
rect -1888 -8078 -1688 -8062
rect -1630 -8028 -1430 -7990
rect -1630 -8062 -1614 -8028
rect -1446 -8062 -1430 -8028
rect -1630 -8078 -1430 -8062
rect -1372 -8028 -1172 -7990
rect -1372 -8062 -1356 -8028
rect -1188 -8062 -1172 -8028
rect -1372 -8078 -1172 -8062
rect -604 -4428 -404 -4412
rect -604 -4462 -588 -4428
rect -420 -4462 -404 -4428
rect -604 -4500 -404 -4462
rect -346 -4428 -146 -4412
rect -346 -4462 -330 -4428
rect -162 -4462 -146 -4428
rect -346 -4500 -146 -4462
rect -88 -4428 112 -4412
rect -88 -4462 -72 -4428
rect 96 -4462 112 -4428
rect -88 -4500 112 -4462
rect 170 -4428 370 -4412
rect 170 -4462 186 -4428
rect 354 -4462 370 -4428
rect 170 -4500 370 -4462
rect 428 -4428 628 -4412
rect 428 -4462 444 -4428
rect 612 -4462 628 -4428
rect 428 -4500 628 -4462
rect -604 -4938 -404 -4900
rect -604 -4972 -588 -4938
rect -420 -4972 -404 -4938
rect -604 -4988 -404 -4972
rect -346 -4938 -146 -4900
rect -346 -4972 -330 -4938
rect -162 -4972 -146 -4938
rect -346 -4988 -146 -4972
rect -88 -4938 112 -4900
rect -88 -4972 -72 -4938
rect 96 -4972 112 -4938
rect -88 -4988 112 -4972
rect 170 -4938 370 -4900
rect 170 -4972 186 -4938
rect 354 -4972 370 -4938
rect 170 -4988 370 -4972
rect 428 -4938 628 -4900
rect 428 -4972 444 -4938
rect 612 -4972 628 -4938
rect 428 -4988 628 -4972
rect -604 -5046 -404 -5030
rect -604 -5080 -588 -5046
rect -420 -5080 -404 -5046
rect -604 -5118 -404 -5080
rect -346 -5046 -146 -5030
rect -346 -5080 -330 -5046
rect -162 -5080 -146 -5046
rect -346 -5118 -146 -5080
rect -88 -5046 112 -5030
rect -88 -5080 -72 -5046
rect 96 -5080 112 -5046
rect -88 -5118 112 -5080
rect 170 -5046 370 -5030
rect 170 -5080 186 -5046
rect 354 -5080 370 -5046
rect 170 -5118 370 -5080
rect 428 -5046 628 -5030
rect 428 -5080 444 -5046
rect 612 -5080 628 -5046
rect 428 -5118 628 -5080
rect -604 -5556 -404 -5518
rect -604 -5590 -588 -5556
rect -420 -5590 -404 -5556
rect -604 -5606 -404 -5590
rect -346 -5556 -146 -5518
rect -346 -5590 -330 -5556
rect -162 -5590 -146 -5556
rect -346 -5606 -146 -5590
rect -88 -5556 112 -5518
rect -88 -5590 -72 -5556
rect 96 -5590 112 -5556
rect -88 -5606 112 -5590
rect 170 -5556 370 -5518
rect 170 -5590 186 -5556
rect 354 -5590 370 -5556
rect 170 -5606 370 -5590
rect 428 -5556 628 -5518
rect 428 -5590 444 -5556
rect 612 -5590 628 -5556
rect 428 -5606 628 -5590
rect -604 -5664 -404 -5648
rect -604 -5698 -588 -5664
rect -420 -5698 -404 -5664
rect -604 -5736 -404 -5698
rect -346 -5664 -146 -5648
rect -346 -5698 -330 -5664
rect -162 -5698 -146 -5664
rect -346 -5736 -146 -5698
rect -88 -5664 112 -5648
rect -88 -5698 -72 -5664
rect 96 -5698 112 -5664
rect -88 -5736 112 -5698
rect 170 -5664 370 -5648
rect 170 -5698 186 -5664
rect 354 -5698 370 -5664
rect 170 -5736 370 -5698
rect 428 -5664 628 -5648
rect 428 -5698 444 -5664
rect 612 -5698 628 -5664
rect 428 -5736 628 -5698
rect -604 -6174 -404 -6136
rect -604 -6208 -588 -6174
rect -420 -6208 -404 -6174
rect -604 -6224 -404 -6208
rect -346 -6174 -146 -6136
rect -346 -6208 -330 -6174
rect -162 -6208 -146 -6174
rect -346 -6224 -146 -6208
rect -88 -6174 112 -6136
rect -88 -6208 -72 -6174
rect 96 -6208 112 -6174
rect -88 -6224 112 -6208
rect 170 -6174 370 -6136
rect 170 -6208 186 -6174
rect 354 -6208 370 -6174
rect 170 -6224 370 -6208
rect 428 -6174 628 -6136
rect 428 -6208 444 -6174
rect 612 -6208 628 -6174
rect 428 -6224 628 -6208
rect -604 -6282 -404 -6266
rect -604 -6316 -588 -6282
rect -420 -6316 -404 -6282
rect -604 -6354 -404 -6316
rect -346 -6282 -146 -6266
rect -346 -6316 -330 -6282
rect -162 -6316 -146 -6282
rect -346 -6354 -146 -6316
rect -88 -6282 112 -6266
rect -88 -6316 -72 -6282
rect 96 -6316 112 -6282
rect -88 -6354 112 -6316
rect 170 -6282 370 -6266
rect 170 -6316 186 -6282
rect 354 -6316 370 -6282
rect 170 -6354 370 -6316
rect 428 -6282 628 -6266
rect 428 -6316 444 -6282
rect 612 -6316 628 -6282
rect 428 -6354 628 -6316
rect -604 -6792 -404 -6754
rect -604 -6826 -588 -6792
rect -420 -6826 -404 -6792
rect -604 -6842 -404 -6826
rect -346 -6792 -146 -6754
rect -346 -6826 -330 -6792
rect -162 -6826 -146 -6792
rect -346 -6842 -146 -6826
rect -88 -6792 112 -6754
rect -88 -6826 -72 -6792
rect 96 -6826 112 -6792
rect -88 -6842 112 -6826
rect 170 -6792 370 -6754
rect 170 -6826 186 -6792
rect 354 -6826 370 -6792
rect 170 -6842 370 -6826
rect 428 -6792 628 -6754
rect 428 -6826 444 -6792
rect 612 -6826 628 -6792
rect 428 -6842 628 -6826
rect -604 -6900 -404 -6884
rect -604 -6934 -588 -6900
rect -420 -6934 -404 -6900
rect -604 -6972 -404 -6934
rect -346 -6900 -146 -6884
rect -346 -6934 -330 -6900
rect -162 -6934 -146 -6900
rect -346 -6972 -146 -6934
rect -88 -6900 112 -6884
rect -88 -6934 -72 -6900
rect 96 -6934 112 -6900
rect -88 -6972 112 -6934
rect 170 -6900 370 -6884
rect 170 -6934 186 -6900
rect 354 -6934 370 -6900
rect 170 -6972 370 -6934
rect 428 -6900 628 -6884
rect 428 -6934 444 -6900
rect 612 -6934 628 -6900
rect 428 -6972 628 -6934
rect -604 -7410 -404 -7372
rect -604 -7444 -588 -7410
rect -420 -7444 -404 -7410
rect -604 -7460 -404 -7444
rect -346 -7410 -146 -7372
rect -346 -7444 -330 -7410
rect -162 -7444 -146 -7410
rect -346 -7460 -146 -7444
rect -88 -7410 112 -7372
rect -88 -7444 -72 -7410
rect 96 -7444 112 -7410
rect -88 -7460 112 -7444
rect 170 -7410 370 -7372
rect 170 -7444 186 -7410
rect 354 -7444 370 -7410
rect 170 -7460 370 -7444
rect 428 -7410 628 -7372
rect 428 -7444 444 -7410
rect 612 -7444 628 -7410
rect 428 -7460 628 -7444
rect -604 -7518 -404 -7502
rect -604 -7552 -588 -7518
rect -420 -7552 -404 -7518
rect -604 -7590 -404 -7552
rect -346 -7518 -146 -7502
rect -346 -7552 -330 -7518
rect -162 -7552 -146 -7518
rect -346 -7590 -146 -7552
rect -88 -7518 112 -7502
rect -88 -7552 -72 -7518
rect 96 -7552 112 -7518
rect -88 -7590 112 -7552
rect 170 -7518 370 -7502
rect 170 -7552 186 -7518
rect 354 -7552 370 -7518
rect 170 -7590 370 -7552
rect 428 -7518 628 -7502
rect 428 -7552 444 -7518
rect 612 -7552 628 -7518
rect 428 -7590 628 -7552
rect -604 -8028 -404 -7990
rect -604 -8062 -588 -8028
rect -420 -8062 -404 -8028
rect -604 -8078 -404 -8062
rect -346 -8028 -146 -7990
rect -346 -8062 -330 -8028
rect -162 -8062 -146 -8028
rect -346 -8078 -146 -8062
rect -88 -8028 112 -7990
rect -88 -8062 -72 -8028
rect 96 -8062 112 -8028
rect -88 -8078 112 -8062
rect 170 -8028 370 -7990
rect 170 -8062 186 -8028
rect 354 -8062 370 -8028
rect 170 -8078 370 -8062
rect 428 -8028 628 -7990
rect 428 -8062 444 -8028
rect 612 -8062 628 -8028
rect 428 -8078 628 -8062
rect 1196 -4428 1396 -4412
rect 1196 -4462 1212 -4428
rect 1380 -4462 1396 -4428
rect 1196 -4500 1396 -4462
rect 1454 -4428 1654 -4412
rect 1454 -4462 1470 -4428
rect 1638 -4462 1654 -4428
rect 1454 -4500 1654 -4462
rect 1712 -4428 1912 -4412
rect 1712 -4462 1728 -4428
rect 1896 -4462 1912 -4428
rect 1712 -4500 1912 -4462
rect 1970 -4428 2170 -4412
rect 1970 -4462 1986 -4428
rect 2154 -4462 2170 -4428
rect 1970 -4500 2170 -4462
rect 2228 -4428 2428 -4412
rect 2228 -4462 2244 -4428
rect 2412 -4462 2428 -4428
rect 2228 -4500 2428 -4462
rect 1196 -4938 1396 -4900
rect 1196 -4972 1212 -4938
rect 1380 -4972 1396 -4938
rect 1196 -4988 1396 -4972
rect 1454 -4938 1654 -4900
rect 1454 -4972 1470 -4938
rect 1638 -4972 1654 -4938
rect 1454 -4988 1654 -4972
rect 1712 -4938 1912 -4900
rect 1712 -4972 1728 -4938
rect 1896 -4972 1912 -4938
rect 1712 -4988 1912 -4972
rect 1970 -4938 2170 -4900
rect 1970 -4972 1986 -4938
rect 2154 -4972 2170 -4938
rect 1970 -4988 2170 -4972
rect 2228 -4938 2428 -4900
rect 2228 -4972 2244 -4938
rect 2412 -4972 2428 -4938
rect 2228 -4988 2428 -4972
rect 1196 -5046 1396 -5030
rect 1196 -5080 1212 -5046
rect 1380 -5080 1396 -5046
rect 1196 -5118 1396 -5080
rect 1454 -5046 1654 -5030
rect 1454 -5080 1470 -5046
rect 1638 -5080 1654 -5046
rect 1454 -5118 1654 -5080
rect 1712 -5046 1912 -5030
rect 1712 -5080 1728 -5046
rect 1896 -5080 1912 -5046
rect 1712 -5118 1912 -5080
rect 1970 -5046 2170 -5030
rect 1970 -5080 1986 -5046
rect 2154 -5080 2170 -5046
rect 1970 -5118 2170 -5080
rect 2228 -5046 2428 -5030
rect 2228 -5080 2244 -5046
rect 2412 -5080 2428 -5046
rect 2228 -5118 2428 -5080
rect 1196 -5556 1396 -5518
rect 1196 -5590 1212 -5556
rect 1380 -5590 1396 -5556
rect 1196 -5606 1396 -5590
rect 1454 -5556 1654 -5518
rect 1454 -5590 1470 -5556
rect 1638 -5590 1654 -5556
rect 1454 -5606 1654 -5590
rect 1712 -5556 1912 -5518
rect 1712 -5590 1728 -5556
rect 1896 -5590 1912 -5556
rect 1712 -5606 1912 -5590
rect 1970 -5556 2170 -5518
rect 1970 -5590 1986 -5556
rect 2154 -5590 2170 -5556
rect 1970 -5606 2170 -5590
rect 2228 -5556 2428 -5518
rect 2228 -5590 2244 -5556
rect 2412 -5590 2428 -5556
rect 2228 -5606 2428 -5590
rect 1196 -5664 1396 -5648
rect 1196 -5698 1212 -5664
rect 1380 -5698 1396 -5664
rect 1196 -5736 1396 -5698
rect 1454 -5664 1654 -5648
rect 1454 -5698 1470 -5664
rect 1638 -5698 1654 -5664
rect 1454 -5736 1654 -5698
rect 1712 -5664 1912 -5648
rect 1712 -5698 1728 -5664
rect 1896 -5698 1912 -5664
rect 1712 -5736 1912 -5698
rect 1970 -5664 2170 -5648
rect 1970 -5698 1986 -5664
rect 2154 -5698 2170 -5664
rect 1970 -5736 2170 -5698
rect 2228 -5664 2428 -5648
rect 2228 -5698 2244 -5664
rect 2412 -5698 2428 -5664
rect 2228 -5736 2428 -5698
rect 1196 -6174 1396 -6136
rect 1196 -6208 1212 -6174
rect 1380 -6208 1396 -6174
rect 1196 -6224 1396 -6208
rect 1454 -6174 1654 -6136
rect 1454 -6208 1470 -6174
rect 1638 -6208 1654 -6174
rect 1454 -6224 1654 -6208
rect 1712 -6174 1912 -6136
rect 1712 -6208 1728 -6174
rect 1896 -6208 1912 -6174
rect 1712 -6224 1912 -6208
rect 1970 -6174 2170 -6136
rect 1970 -6208 1986 -6174
rect 2154 -6208 2170 -6174
rect 1970 -6224 2170 -6208
rect 2228 -6174 2428 -6136
rect 2228 -6208 2244 -6174
rect 2412 -6208 2428 -6174
rect 2228 -6224 2428 -6208
rect 1196 -6282 1396 -6266
rect 1196 -6316 1212 -6282
rect 1380 -6316 1396 -6282
rect 1196 -6354 1396 -6316
rect 1454 -6282 1654 -6266
rect 1454 -6316 1470 -6282
rect 1638 -6316 1654 -6282
rect 1454 -6354 1654 -6316
rect 1712 -6282 1912 -6266
rect 1712 -6316 1728 -6282
rect 1896 -6316 1912 -6282
rect 1712 -6354 1912 -6316
rect 1970 -6282 2170 -6266
rect 1970 -6316 1986 -6282
rect 2154 -6316 2170 -6282
rect 1970 -6354 2170 -6316
rect 2228 -6282 2428 -6266
rect 2228 -6316 2244 -6282
rect 2412 -6316 2428 -6282
rect 2228 -6354 2428 -6316
rect 1196 -6792 1396 -6754
rect 1196 -6826 1212 -6792
rect 1380 -6826 1396 -6792
rect 1196 -6842 1396 -6826
rect 1454 -6792 1654 -6754
rect 1454 -6826 1470 -6792
rect 1638 -6826 1654 -6792
rect 1454 -6842 1654 -6826
rect 1712 -6792 1912 -6754
rect 1712 -6826 1728 -6792
rect 1896 -6826 1912 -6792
rect 1712 -6842 1912 -6826
rect 1970 -6792 2170 -6754
rect 1970 -6826 1986 -6792
rect 2154 -6826 2170 -6792
rect 1970 -6842 2170 -6826
rect 2228 -6792 2428 -6754
rect 2228 -6826 2244 -6792
rect 2412 -6826 2428 -6792
rect 2228 -6842 2428 -6826
rect 1196 -6900 1396 -6884
rect 1196 -6934 1212 -6900
rect 1380 -6934 1396 -6900
rect 1196 -6972 1396 -6934
rect 1454 -6900 1654 -6884
rect 1454 -6934 1470 -6900
rect 1638 -6934 1654 -6900
rect 1454 -6972 1654 -6934
rect 1712 -6900 1912 -6884
rect 1712 -6934 1728 -6900
rect 1896 -6934 1912 -6900
rect 1712 -6972 1912 -6934
rect 1970 -6900 2170 -6884
rect 1970 -6934 1986 -6900
rect 2154 -6934 2170 -6900
rect 1970 -6972 2170 -6934
rect 2228 -6900 2428 -6884
rect 2228 -6934 2244 -6900
rect 2412 -6934 2428 -6900
rect 2228 -6972 2428 -6934
rect 1196 -7410 1396 -7372
rect 1196 -7444 1212 -7410
rect 1380 -7444 1396 -7410
rect 1196 -7460 1396 -7444
rect 1454 -7410 1654 -7372
rect 1454 -7444 1470 -7410
rect 1638 -7444 1654 -7410
rect 1454 -7460 1654 -7444
rect 1712 -7410 1912 -7372
rect 1712 -7444 1728 -7410
rect 1896 -7444 1912 -7410
rect 1712 -7460 1912 -7444
rect 1970 -7410 2170 -7372
rect 1970 -7444 1986 -7410
rect 2154 -7444 2170 -7410
rect 1970 -7460 2170 -7444
rect 2228 -7410 2428 -7372
rect 2228 -7444 2244 -7410
rect 2412 -7444 2428 -7410
rect 2228 -7460 2428 -7444
rect 1196 -7518 1396 -7502
rect 1196 -7552 1212 -7518
rect 1380 -7552 1396 -7518
rect 1196 -7590 1396 -7552
rect 1454 -7518 1654 -7502
rect 1454 -7552 1470 -7518
rect 1638 -7552 1654 -7518
rect 1454 -7590 1654 -7552
rect 1712 -7518 1912 -7502
rect 1712 -7552 1728 -7518
rect 1896 -7552 1912 -7518
rect 1712 -7590 1912 -7552
rect 1970 -7518 2170 -7502
rect 1970 -7552 1986 -7518
rect 2154 -7552 2170 -7518
rect 1970 -7590 2170 -7552
rect 2228 -7518 2428 -7502
rect 2228 -7552 2244 -7518
rect 2412 -7552 2428 -7518
rect 2228 -7590 2428 -7552
rect 1196 -8028 1396 -7990
rect 1196 -8062 1212 -8028
rect 1380 -8062 1396 -8028
rect 1196 -8078 1396 -8062
rect 1454 -8028 1654 -7990
rect 1454 -8062 1470 -8028
rect 1638 -8062 1654 -8028
rect 1454 -8078 1654 -8062
rect 1712 -8028 1912 -7990
rect 1712 -8062 1728 -8028
rect 1896 -8062 1912 -8028
rect 1712 -8078 1912 -8062
rect 1970 -8028 2170 -7990
rect 1970 -8062 1986 -8028
rect 2154 -8062 2170 -8028
rect 1970 -8078 2170 -8062
rect 2228 -8028 2428 -7990
rect 2228 -8062 2244 -8028
rect 2412 -8062 2428 -8028
rect 2228 -8078 2428 -8062
rect 2996 -4428 3196 -4412
rect 2996 -4462 3012 -4428
rect 3180 -4462 3196 -4428
rect 2996 -4500 3196 -4462
rect 3254 -4428 3454 -4412
rect 3254 -4462 3270 -4428
rect 3438 -4462 3454 -4428
rect 3254 -4500 3454 -4462
rect 3512 -4428 3712 -4412
rect 3512 -4462 3528 -4428
rect 3696 -4462 3712 -4428
rect 3512 -4500 3712 -4462
rect 3770 -4428 3970 -4412
rect 3770 -4462 3786 -4428
rect 3954 -4462 3970 -4428
rect 3770 -4500 3970 -4462
rect 4028 -4428 4228 -4412
rect 4028 -4462 4044 -4428
rect 4212 -4462 4228 -4428
rect 4028 -4500 4228 -4462
rect 2996 -4938 3196 -4900
rect 2996 -4972 3012 -4938
rect 3180 -4972 3196 -4938
rect 2996 -4988 3196 -4972
rect 3254 -4938 3454 -4900
rect 3254 -4972 3270 -4938
rect 3438 -4972 3454 -4938
rect 3254 -4988 3454 -4972
rect 3512 -4938 3712 -4900
rect 3512 -4972 3528 -4938
rect 3696 -4972 3712 -4938
rect 3512 -4988 3712 -4972
rect 3770 -4938 3970 -4900
rect 3770 -4972 3786 -4938
rect 3954 -4972 3970 -4938
rect 3770 -4988 3970 -4972
rect 4028 -4938 4228 -4900
rect 4028 -4972 4044 -4938
rect 4212 -4972 4228 -4938
rect 4028 -4988 4228 -4972
rect 2996 -5046 3196 -5030
rect 2996 -5080 3012 -5046
rect 3180 -5080 3196 -5046
rect 2996 -5118 3196 -5080
rect 3254 -5046 3454 -5030
rect 3254 -5080 3270 -5046
rect 3438 -5080 3454 -5046
rect 3254 -5118 3454 -5080
rect 3512 -5046 3712 -5030
rect 3512 -5080 3528 -5046
rect 3696 -5080 3712 -5046
rect 3512 -5118 3712 -5080
rect 3770 -5046 3970 -5030
rect 3770 -5080 3786 -5046
rect 3954 -5080 3970 -5046
rect 3770 -5118 3970 -5080
rect 4028 -5046 4228 -5030
rect 4028 -5080 4044 -5046
rect 4212 -5080 4228 -5046
rect 4028 -5118 4228 -5080
rect 2996 -5556 3196 -5518
rect 2996 -5590 3012 -5556
rect 3180 -5590 3196 -5556
rect 2996 -5606 3196 -5590
rect 3254 -5556 3454 -5518
rect 3254 -5590 3270 -5556
rect 3438 -5590 3454 -5556
rect 3254 -5606 3454 -5590
rect 3512 -5556 3712 -5518
rect 3512 -5590 3528 -5556
rect 3696 -5590 3712 -5556
rect 3512 -5606 3712 -5590
rect 3770 -5556 3970 -5518
rect 3770 -5590 3786 -5556
rect 3954 -5590 3970 -5556
rect 3770 -5606 3970 -5590
rect 4028 -5556 4228 -5518
rect 4028 -5590 4044 -5556
rect 4212 -5590 4228 -5556
rect 4028 -5606 4228 -5590
rect 2996 -5664 3196 -5648
rect 2996 -5698 3012 -5664
rect 3180 -5698 3196 -5664
rect 2996 -5736 3196 -5698
rect 3254 -5664 3454 -5648
rect 3254 -5698 3270 -5664
rect 3438 -5698 3454 -5664
rect 3254 -5736 3454 -5698
rect 3512 -5664 3712 -5648
rect 3512 -5698 3528 -5664
rect 3696 -5698 3712 -5664
rect 3512 -5736 3712 -5698
rect 3770 -5664 3970 -5648
rect 3770 -5698 3786 -5664
rect 3954 -5698 3970 -5664
rect 3770 -5736 3970 -5698
rect 4028 -5664 4228 -5648
rect 4028 -5698 4044 -5664
rect 4212 -5698 4228 -5664
rect 4028 -5736 4228 -5698
rect 2996 -6174 3196 -6136
rect 2996 -6208 3012 -6174
rect 3180 -6208 3196 -6174
rect 2996 -6224 3196 -6208
rect 3254 -6174 3454 -6136
rect 3254 -6208 3270 -6174
rect 3438 -6208 3454 -6174
rect 3254 -6224 3454 -6208
rect 3512 -6174 3712 -6136
rect 3512 -6208 3528 -6174
rect 3696 -6208 3712 -6174
rect 3512 -6224 3712 -6208
rect 3770 -6174 3970 -6136
rect 3770 -6208 3786 -6174
rect 3954 -6208 3970 -6174
rect 3770 -6224 3970 -6208
rect 4028 -6174 4228 -6136
rect 4028 -6208 4044 -6174
rect 4212 -6208 4228 -6174
rect 4028 -6224 4228 -6208
rect 2996 -6282 3196 -6266
rect 2996 -6316 3012 -6282
rect 3180 -6316 3196 -6282
rect 2996 -6354 3196 -6316
rect 3254 -6282 3454 -6266
rect 3254 -6316 3270 -6282
rect 3438 -6316 3454 -6282
rect 3254 -6354 3454 -6316
rect 3512 -6282 3712 -6266
rect 3512 -6316 3528 -6282
rect 3696 -6316 3712 -6282
rect 3512 -6354 3712 -6316
rect 3770 -6282 3970 -6266
rect 3770 -6316 3786 -6282
rect 3954 -6316 3970 -6282
rect 3770 -6354 3970 -6316
rect 4028 -6282 4228 -6266
rect 4028 -6316 4044 -6282
rect 4212 -6316 4228 -6282
rect 4028 -6354 4228 -6316
rect 2996 -6792 3196 -6754
rect 2996 -6826 3012 -6792
rect 3180 -6826 3196 -6792
rect 2996 -6842 3196 -6826
rect 3254 -6792 3454 -6754
rect 3254 -6826 3270 -6792
rect 3438 -6826 3454 -6792
rect 3254 -6842 3454 -6826
rect 3512 -6792 3712 -6754
rect 3512 -6826 3528 -6792
rect 3696 -6826 3712 -6792
rect 3512 -6842 3712 -6826
rect 3770 -6792 3970 -6754
rect 3770 -6826 3786 -6792
rect 3954 -6826 3970 -6792
rect 3770 -6842 3970 -6826
rect 4028 -6792 4228 -6754
rect 4028 -6826 4044 -6792
rect 4212 -6826 4228 -6792
rect 4028 -6842 4228 -6826
rect 2996 -6900 3196 -6884
rect 2996 -6934 3012 -6900
rect 3180 -6934 3196 -6900
rect 2996 -6972 3196 -6934
rect 3254 -6900 3454 -6884
rect 3254 -6934 3270 -6900
rect 3438 -6934 3454 -6900
rect 3254 -6972 3454 -6934
rect 3512 -6900 3712 -6884
rect 3512 -6934 3528 -6900
rect 3696 -6934 3712 -6900
rect 3512 -6972 3712 -6934
rect 3770 -6900 3970 -6884
rect 3770 -6934 3786 -6900
rect 3954 -6934 3970 -6900
rect 3770 -6972 3970 -6934
rect 4028 -6900 4228 -6884
rect 4028 -6934 4044 -6900
rect 4212 -6934 4228 -6900
rect 4028 -6972 4228 -6934
rect 2996 -7410 3196 -7372
rect 2996 -7444 3012 -7410
rect 3180 -7444 3196 -7410
rect 2996 -7460 3196 -7444
rect 3254 -7410 3454 -7372
rect 3254 -7444 3270 -7410
rect 3438 -7444 3454 -7410
rect 3254 -7460 3454 -7444
rect 3512 -7410 3712 -7372
rect 3512 -7444 3528 -7410
rect 3696 -7444 3712 -7410
rect 3512 -7460 3712 -7444
rect 3770 -7410 3970 -7372
rect 3770 -7444 3786 -7410
rect 3954 -7444 3970 -7410
rect 3770 -7460 3970 -7444
rect 4028 -7410 4228 -7372
rect 4028 -7444 4044 -7410
rect 4212 -7444 4228 -7410
rect 4028 -7460 4228 -7444
rect 2996 -7518 3196 -7502
rect 2996 -7552 3012 -7518
rect 3180 -7552 3196 -7518
rect 2996 -7590 3196 -7552
rect 3254 -7518 3454 -7502
rect 3254 -7552 3270 -7518
rect 3438 -7552 3454 -7518
rect 3254 -7590 3454 -7552
rect 3512 -7518 3712 -7502
rect 3512 -7552 3528 -7518
rect 3696 -7552 3712 -7518
rect 3512 -7590 3712 -7552
rect 3770 -7518 3970 -7502
rect 3770 -7552 3786 -7518
rect 3954 -7552 3970 -7518
rect 3770 -7590 3970 -7552
rect 4028 -7518 4228 -7502
rect 4028 -7552 4044 -7518
rect 4212 -7552 4228 -7518
rect 4028 -7590 4228 -7552
rect 2996 -8028 3196 -7990
rect 2996 -8062 3012 -8028
rect 3180 -8062 3196 -8028
rect 2996 -8078 3196 -8062
rect 3254 -8028 3454 -7990
rect 3254 -8062 3270 -8028
rect 3438 -8062 3454 -8028
rect 3254 -8078 3454 -8062
rect 3512 -8028 3712 -7990
rect 3512 -8062 3528 -8028
rect 3696 -8062 3712 -8028
rect 3512 -8078 3712 -8062
rect 3770 -8028 3970 -7990
rect 3770 -8062 3786 -8028
rect 3954 -8062 3970 -8028
rect 3770 -8078 3970 -8062
rect 4028 -8028 4228 -7990
rect 4028 -8062 4044 -8028
rect 4212 -8062 4228 -8028
rect 4028 -8078 4228 -8062
<< polycont >>
rect 2498 2102 2532 2136
rect 2690 2102 2724 2136
rect 2882 2102 2916 2136
rect 3074 2102 3108 2136
rect 3266 2102 3300 2136
rect 3458 2102 3492 2136
rect 3650 2102 3684 2136
rect 3842 2102 3876 2136
rect 4034 2102 4068 2136
rect 4226 2102 4260 2136
rect 2594 1574 2628 1608
rect 2786 1574 2820 1608
rect 2978 1574 3012 1608
rect 3170 1574 3204 1608
rect 3362 1574 3396 1608
rect 3554 1574 3588 1608
rect 3746 1574 3780 1608
rect 3938 1574 3972 1608
rect 4130 1574 4164 1608
rect 4322 1574 4356 1608
rect 2594 1466 2628 1500
rect 2786 1466 2820 1500
rect 2978 1466 3012 1500
rect 3170 1466 3204 1500
rect 3362 1466 3396 1500
rect 3554 1466 3588 1500
rect 3746 1466 3780 1500
rect 3938 1466 3972 1500
rect 4130 1466 4164 1500
rect 4322 1466 4356 1500
rect 2498 938 2532 972
rect 2690 938 2724 972
rect 2882 938 2916 972
rect 3074 938 3108 972
rect 3266 938 3300 972
rect 3458 938 3492 972
rect 3650 938 3684 972
rect 3842 938 3876 972
rect 4034 938 4068 972
rect 4226 938 4260 972
rect 274 64 308 98
rect 466 64 500 98
rect 658 64 692 98
rect 850 64 884 98
rect 1042 64 1076 98
rect 1234 64 1268 98
rect 1426 64 1460 98
rect 1618 64 1652 98
rect 1810 64 1844 98
rect 2002 64 2036 98
rect 178 -446 212 -412
rect 370 -446 404 -412
rect 562 -446 596 -412
rect 754 -446 788 -412
rect 946 -446 980 -412
rect 1138 -446 1172 -412
rect 1330 -446 1364 -412
rect 1522 -446 1556 -412
rect 1714 -446 1748 -412
rect 1906 -446 1940 -412
rect 178 -554 212 -520
rect 370 -554 404 -520
rect 562 -554 596 -520
rect 754 -554 788 -520
rect 946 -554 980 -520
rect 1138 -554 1172 -520
rect 1330 -554 1364 -520
rect 1522 -554 1556 -520
rect 1714 -554 1748 -520
rect 1906 -554 1940 -520
rect 274 -1064 308 -1030
rect 466 -1064 500 -1030
rect 658 -1064 692 -1030
rect 850 -1064 884 -1030
rect 1042 -1064 1076 -1030
rect 1234 -1064 1268 -1030
rect 1426 -1064 1460 -1030
rect 1618 -1064 1652 -1030
rect 1810 -1064 1844 -1030
rect 2002 -1064 2036 -1030
rect 274 -1172 308 -1138
rect 466 -1172 500 -1138
rect 658 -1172 692 -1138
rect 850 -1172 884 -1138
rect 1042 -1172 1076 -1138
rect 1234 -1172 1268 -1138
rect 1426 -1172 1460 -1138
rect 1618 -1172 1652 -1138
rect 1810 -1172 1844 -1138
rect 2002 -1172 2036 -1138
rect 178 -1682 212 -1648
rect 370 -1682 404 -1648
rect 562 -1682 596 -1648
rect 754 -1682 788 -1648
rect 946 -1682 980 -1648
rect 1138 -1682 1172 -1648
rect 1330 -1682 1364 -1648
rect 1522 -1682 1556 -1648
rect 1714 -1682 1748 -1648
rect 1906 -1682 1940 -1648
rect 2498 506 2532 540
rect 2690 506 2724 540
rect 2882 506 2916 540
rect 3074 506 3108 540
rect 3266 506 3300 540
rect 3458 506 3492 540
rect 3650 506 3684 540
rect 3842 506 3876 540
rect 4034 506 4068 540
rect 4226 506 4260 540
rect 2594 -4 2628 30
rect 2786 -4 2820 30
rect 2978 -4 3012 30
rect 3170 -4 3204 30
rect 3362 -4 3396 30
rect 3554 -4 3588 30
rect 3746 -4 3780 30
rect 3938 -4 3972 30
rect 4130 -4 4164 30
rect 4322 -4 4356 30
rect 2594 -112 2628 -78
rect 2786 -112 2820 -78
rect 2978 -112 3012 -78
rect 3170 -112 3204 -78
rect 3362 -112 3396 -78
rect 3554 -112 3588 -78
rect 3746 -112 3780 -78
rect 3938 -112 3972 -78
rect 4130 -112 4164 -78
rect 4322 -112 4356 -78
rect 2498 -622 2532 -588
rect 2690 -622 2724 -588
rect 2882 -622 2916 -588
rect 3074 -622 3108 -588
rect 3266 -622 3300 -588
rect 3458 -622 3492 -588
rect 3650 -622 3684 -588
rect 3842 -622 3876 -588
rect 4034 -622 4068 -588
rect 4226 -622 4260 -588
rect -2306 -2316 -2272 -2282
rect -2114 -2316 -2080 -2282
rect -1922 -2316 -1888 -2282
rect -1730 -2316 -1696 -2282
rect -1538 -2316 -1504 -2282
rect -2402 -2826 -2368 -2792
rect -2210 -2826 -2176 -2792
rect -2018 -2826 -1984 -2792
rect -1826 -2826 -1792 -2792
rect -1634 -2826 -1600 -2792
rect -2402 -2934 -2368 -2900
rect -2210 -2934 -2176 -2900
rect -2018 -2934 -1984 -2900
rect -1826 -2934 -1792 -2900
rect -1634 -2934 -1600 -2900
rect -2306 -3444 -2272 -3410
rect -2114 -3444 -2080 -3410
rect -1922 -3444 -1888 -3410
rect -1730 -3444 -1696 -3410
rect -1538 -3444 -1504 -3410
rect -2306 -3552 -2272 -3518
rect -2114 -3552 -2080 -3518
rect -1922 -3552 -1888 -3518
rect -1730 -3552 -1696 -3518
rect -1538 -3552 -1504 -3518
rect -2402 -4062 -2368 -4028
rect -2210 -4062 -2176 -4028
rect -2018 -4062 -1984 -4028
rect -1826 -4062 -1792 -4028
rect -1634 -4062 -1600 -4028
rect -506 -2316 -472 -2282
rect -314 -2316 -280 -2282
rect -122 -2316 -88 -2282
rect 70 -2316 104 -2282
rect 262 -2316 296 -2282
rect -602 -2826 -568 -2792
rect -410 -2826 -376 -2792
rect -218 -2826 -184 -2792
rect -26 -2826 8 -2792
rect 166 -2826 200 -2792
rect -602 -2934 -568 -2900
rect -410 -2934 -376 -2900
rect -218 -2934 -184 -2900
rect -26 -2934 8 -2900
rect 166 -2934 200 -2900
rect -506 -3444 -472 -3410
rect -314 -3444 -280 -3410
rect -122 -3444 -88 -3410
rect 70 -3444 104 -3410
rect 262 -3444 296 -3410
rect -506 -3552 -472 -3518
rect -314 -3552 -280 -3518
rect -122 -3552 -88 -3518
rect 70 -3552 104 -3518
rect 262 -3552 296 -3518
rect -602 -4062 -568 -4028
rect -410 -4062 -376 -4028
rect -218 -4062 -184 -4028
rect -26 -4062 8 -4028
rect 166 -4062 200 -4028
rect 1294 -2316 1328 -2282
rect 1486 -2316 1520 -2282
rect 1678 -2316 1712 -2282
rect 1870 -2316 1904 -2282
rect 2062 -2316 2096 -2282
rect 1198 -2826 1232 -2792
rect 1390 -2826 1424 -2792
rect 1582 -2826 1616 -2792
rect 1774 -2826 1808 -2792
rect 1966 -2826 2000 -2792
rect 1198 -2934 1232 -2900
rect 1390 -2934 1424 -2900
rect 1582 -2934 1616 -2900
rect 1774 -2934 1808 -2900
rect 1966 -2934 2000 -2900
rect 1294 -3444 1328 -3410
rect 1486 -3444 1520 -3410
rect 1678 -3444 1712 -3410
rect 1870 -3444 1904 -3410
rect 2062 -3444 2096 -3410
rect 1294 -3552 1328 -3518
rect 1486 -3552 1520 -3518
rect 1678 -3552 1712 -3518
rect 1870 -3552 1904 -3518
rect 2062 -3552 2096 -3518
rect 1198 -4062 1232 -4028
rect 1390 -4062 1424 -4028
rect 1582 -4062 1616 -4028
rect 1774 -4062 1808 -4028
rect 1966 -4062 2000 -4028
rect 3094 -2316 3128 -2282
rect 3286 -2316 3320 -2282
rect 3478 -2316 3512 -2282
rect 3670 -2316 3704 -2282
rect 3862 -2316 3896 -2282
rect 2998 -2826 3032 -2792
rect 3190 -2826 3224 -2792
rect 3382 -2826 3416 -2792
rect 3574 -2826 3608 -2792
rect 3766 -2826 3800 -2792
rect 2998 -2934 3032 -2900
rect 3190 -2934 3224 -2900
rect 3382 -2934 3416 -2900
rect 3574 -2934 3608 -2900
rect 3766 -2934 3800 -2900
rect 3094 -3444 3128 -3410
rect 3286 -3444 3320 -3410
rect 3478 -3444 3512 -3410
rect 3670 -3444 3704 -3410
rect 3862 -3444 3896 -3410
rect 3094 -3552 3128 -3518
rect 3286 -3552 3320 -3518
rect 3478 -3552 3512 -3518
rect 3670 -3552 3704 -3518
rect 3862 -3552 3896 -3518
rect 2998 -4062 3032 -4028
rect 3190 -4062 3224 -4028
rect 3382 -4062 3416 -4028
rect 3574 -4062 3608 -4028
rect 3766 -4062 3800 -4028
rect 5094 2072 5128 2106
rect 5286 2072 5320 2106
rect 5478 2072 5512 2106
rect 5670 2072 5704 2106
rect 5862 2072 5896 2106
rect 6054 2072 6088 2106
rect 6246 2072 6280 2106
rect 6438 2072 6472 2106
rect 6630 2072 6664 2106
rect 6822 2072 6856 2106
rect 4998 1562 5032 1596
rect 5190 1562 5224 1596
rect 5382 1562 5416 1596
rect 5574 1562 5608 1596
rect 5766 1562 5800 1596
rect 5958 1562 5992 1596
rect 6150 1562 6184 1596
rect 6342 1562 6376 1596
rect 6534 1562 6568 1596
rect 6726 1562 6760 1596
rect 4998 1454 5032 1488
rect 5190 1454 5224 1488
rect 5382 1454 5416 1488
rect 5574 1454 5608 1488
rect 5766 1454 5800 1488
rect 5958 1454 5992 1488
rect 6150 1454 6184 1488
rect 6342 1454 6376 1488
rect 6534 1454 6568 1488
rect 6726 1454 6760 1488
rect 5094 944 5128 978
rect 5286 944 5320 978
rect 5478 944 5512 978
rect 5670 944 5704 978
rect 5862 944 5896 978
rect 6054 944 6088 978
rect 6246 944 6280 978
rect 6438 944 6472 978
rect 6630 944 6664 978
rect 6822 944 6856 978
rect 5094 836 5128 870
rect 5286 836 5320 870
rect 5478 836 5512 870
rect 5670 836 5704 870
rect 5862 836 5896 870
rect 6054 836 6088 870
rect 6246 836 6280 870
rect 6438 836 6472 870
rect 6630 836 6664 870
rect 6822 836 6856 870
rect 4998 326 5032 360
rect 5190 326 5224 360
rect 5382 326 5416 360
rect 5574 326 5608 360
rect 5766 326 5800 360
rect 5958 326 5992 360
rect 6150 326 6184 360
rect 6342 326 6376 360
rect 6534 326 6568 360
rect 6726 326 6760 360
rect 4998 218 5032 252
rect 5190 218 5224 252
rect 5382 218 5416 252
rect 5574 218 5608 252
rect 5766 218 5800 252
rect 5958 218 5992 252
rect 6150 218 6184 252
rect 6342 218 6376 252
rect 6534 218 6568 252
rect 6726 218 6760 252
rect 5094 -292 5128 -258
rect 5286 -292 5320 -258
rect 5478 -292 5512 -258
rect 5670 -292 5704 -258
rect 5862 -292 5896 -258
rect 6054 -292 6088 -258
rect 6246 -292 6280 -258
rect 6438 -292 6472 -258
rect 6630 -292 6664 -258
rect 6822 -292 6856 -258
rect 5094 -400 5128 -366
rect 5286 -400 5320 -366
rect 5478 -400 5512 -366
rect 5670 -400 5704 -366
rect 5862 -400 5896 -366
rect 6054 -400 6088 -366
rect 6246 -400 6280 -366
rect 6438 -400 6472 -366
rect 6630 -400 6664 -366
rect 6822 -400 6856 -366
rect 4998 -910 5032 -876
rect 5190 -910 5224 -876
rect 5382 -910 5416 -876
rect 5574 -910 5608 -876
rect 5766 -910 5800 -876
rect 5958 -910 5992 -876
rect 6150 -910 6184 -876
rect 6342 -910 6376 -876
rect 6534 -910 6568 -876
rect 6726 -910 6760 -876
rect 4998 -1018 5032 -984
rect 5190 -1018 5224 -984
rect 5382 -1018 5416 -984
rect 5574 -1018 5608 -984
rect 5766 -1018 5800 -984
rect 5958 -1018 5992 -984
rect 6150 -1018 6184 -984
rect 6342 -1018 6376 -984
rect 6534 -1018 6568 -984
rect 6726 -1018 6760 -984
rect 5094 -1528 5128 -1494
rect 5286 -1528 5320 -1494
rect 5478 -1528 5512 -1494
rect 5670 -1528 5704 -1494
rect 5862 -1528 5896 -1494
rect 6054 -1528 6088 -1494
rect 6246 -1528 6280 -1494
rect 6438 -1528 6472 -1494
rect 6630 -1528 6664 -1494
rect 6822 -1528 6856 -1494
rect 5094 -1636 5128 -1602
rect 5286 -1636 5320 -1602
rect 5478 -1636 5512 -1602
rect 5670 -1636 5704 -1602
rect 5862 -1636 5896 -1602
rect 6054 -1636 6088 -1602
rect 6246 -1636 6280 -1602
rect 6438 -1636 6472 -1602
rect 6630 -1636 6664 -1602
rect 6822 -1636 6856 -1602
rect 4998 -2146 5032 -2112
rect 5190 -2146 5224 -2112
rect 5382 -2146 5416 -2112
rect 5574 -2146 5608 -2112
rect 5766 -2146 5800 -2112
rect 5958 -2146 5992 -2112
rect 6150 -2146 6184 -2112
rect 6342 -2146 6376 -2112
rect 6534 -2146 6568 -2112
rect 6726 -2146 6760 -2112
rect 4998 -2254 5032 -2220
rect 5190 -2254 5224 -2220
rect 5382 -2254 5416 -2220
rect 5574 -2254 5608 -2220
rect 5766 -2254 5800 -2220
rect 5958 -2254 5992 -2220
rect 6150 -2254 6184 -2220
rect 6342 -2254 6376 -2220
rect 6534 -2254 6568 -2220
rect 6726 -2254 6760 -2220
rect 5094 -2764 5128 -2730
rect 5286 -2764 5320 -2730
rect 5478 -2764 5512 -2730
rect 5670 -2764 5704 -2730
rect 5862 -2764 5896 -2730
rect 6054 -2764 6088 -2730
rect 6246 -2764 6280 -2730
rect 6438 -2764 6472 -2730
rect 6630 -2764 6664 -2730
rect 6822 -2764 6856 -2730
rect 5094 -2872 5128 -2838
rect 5286 -2872 5320 -2838
rect 5478 -2872 5512 -2838
rect 5670 -2872 5704 -2838
rect 5862 -2872 5896 -2838
rect 6054 -2872 6088 -2838
rect 6246 -2872 6280 -2838
rect 6438 -2872 6472 -2838
rect 6630 -2872 6664 -2838
rect 6822 -2872 6856 -2838
rect 4998 -3382 5032 -3348
rect 5190 -3382 5224 -3348
rect 5382 -3382 5416 -3348
rect 5574 -3382 5608 -3348
rect 5766 -3382 5800 -3348
rect 5958 -3382 5992 -3348
rect 6150 -3382 6184 -3348
rect 6342 -3382 6376 -3348
rect 6534 -3382 6568 -3348
rect 6726 -3382 6760 -3348
rect -2388 -4462 -2220 -4428
rect -2130 -4462 -1962 -4428
rect -1872 -4462 -1704 -4428
rect -1614 -4462 -1446 -4428
rect -1356 -4462 -1188 -4428
rect -2388 -4972 -2220 -4938
rect -2130 -4972 -1962 -4938
rect -1872 -4972 -1704 -4938
rect -1614 -4972 -1446 -4938
rect -1356 -4972 -1188 -4938
rect -2388 -5080 -2220 -5046
rect -2130 -5080 -1962 -5046
rect -1872 -5080 -1704 -5046
rect -1614 -5080 -1446 -5046
rect -1356 -5080 -1188 -5046
rect -2388 -5590 -2220 -5556
rect -2130 -5590 -1962 -5556
rect -1872 -5590 -1704 -5556
rect -1614 -5590 -1446 -5556
rect -1356 -5590 -1188 -5556
rect -2388 -5698 -2220 -5664
rect -2130 -5698 -1962 -5664
rect -1872 -5698 -1704 -5664
rect -1614 -5698 -1446 -5664
rect -1356 -5698 -1188 -5664
rect -2388 -6208 -2220 -6174
rect -2130 -6208 -1962 -6174
rect -1872 -6208 -1704 -6174
rect -1614 -6208 -1446 -6174
rect -1356 -6208 -1188 -6174
rect -2388 -6316 -2220 -6282
rect -2130 -6316 -1962 -6282
rect -1872 -6316 -1704 -6282
rect -1614 -6316 -1446 -6282
rect -1356 -6316 -1188 -6282
rect -2388 -6826 -2220 -6792
rect -2130 -6826 -1962 -6792
rect -1872 -6826 -1704 -6792
rect -1614 -6826 -1446 -6792
rect -1356 -6826 -1188 -6792
rect -2388 -6934 -2220 -6900
rect -2130 -6934 -1962 -6900
rect -1872 -6934 -1704 -6900
rect -1614 -6934 -1446 -6900
rect -1356 -6934 -1188 -6900
rect -2388 -7444 -2220 -7410
rect -2130 -7444 -1962 -7410
rect -1872 -7444 -1704 -7410
rect -1614 -7444 -1446 -7410
rect -1356 -7444 -1188 -7410
rect -2388 -7552 -2220 -7518
rect -2130 -7552 -1962 -7518
rect -1872 -7552 -1704 -7518
rect -1614 -7552 -1446 -7518
rect -1356 -7552 -1188 -7518
rect -2388 -8062 -2220 -8028
rect -2130 -8062 -1962 -8028
rect -1872 -8062 -1704 -8028
rect -1614 -8062 -1446 -8028
rect -1356 -8062 -1188 -8028
rect -588 -4462 -420 -4428
rect -330 -4462 -162 -4428
rect -72 -4462 96 -4428
rect 186 -4462 354 -4428
rect 444 -4462 612 -4428
rect -588 -4972 -420 -4938
rect -330 -4972 -162 -4938
rect -72 -4972 96 -4938
rect 186 -4972 354 -4938
rect 444 -4972 612 -4938
rect -588 -5080 -420 -5046
rect -330 -5080 -162 -5046
rect -72 -5080 96 -5046
rect 186 -5080 354 -5046
rect 444 -5080 612 -5046
rect -588 -5590 -420 -5556
rect -330 -5590 -162 -5556
rect -72 -5590 96 -5556
rect 186 -5590 354 -5556
rect 444 -5590 612 -5556
rect -588 -5698 -420 -5664
rect -330 -5698 -162 -5664
rect -72 -5698 96 -5664
rect 186 -5698 354 -5664
rect 444 -5698 612 -5664
rect -588 -6208 -420 -6174
rect -330 -6208 -162 -6174
rect -72 -6208 96 -6174
rect 186 -6208 354 -6174
rect 444 -6208 612 -6174
rect -588 -6316 -420 -6282
rect -330 -6316 -162 -6282
rect -72 -6316 96 -6282
rect 186 -6316 354 -6282
rect 444 -6316 612 -6282
rect -588 -6826 -420 -6792
rect -330 -6826 -162 -6792
rect -72 -6826 96 -6792
rect 186 -6826 354 -6792
rect 444 -6826 612 -6792
rect -588 -6934 -420 -6900
rect -330 -6934 -162 -6900
rect -72 -6934 96 -6900
rect 186 -6934 354 -6900
rect 444 -6934 612 -6900
rect -588 -7444 -420 -7410
rect -330 -7444 -162 -7410
rect -72 -7444 96 -7410
rect 186 -7444 354 -7410
rect 444 -7444 612 -7410
rect -588 -7552 -420 -7518
rect -330 -7552 -162 -7518
rect -72 -7552 96 -7518
rect 186 -7552 354 -7518
rect 444 -7552 612 -7518
rect -588 -8062 -420 -8028
rect -330 -8062 -162 -8028
rect -72 -8062 96 -8028
rect 186 -8062 354 -8028
rect 444 -8062 612 -8028
rect 1212 -4462 1380 -4428
rect 1470 -4462 1638 -4428
rect 1728 -4462 1896 -4428
rect 1986 -4462 2154 -4428
rect 2244 -4462 2412 -4428
rect 1212 -4972 1380 -4938
rect 1470 -4972 1638 -4938
rect 1728 -4972 1896 -4938
rect 1986 -4972 2154 -4938
rect 2244 -4972 2412 -4938
rect 1212 -5080 1380 -5046
rect 1470 -5080 1638 -5046
rect 1728 -5080 1896 -5046
rect 1986 -5080 2154 -5046
rect 2244 -5080 2412 -5046
rect 1212 -5590 1380 -5556
rect 1470 -5590 1638 -5556
rect 1728 -5590 1896 -5556
rect 1986 -5590 2154 -5556
rect 2244 -5590 2412 -5556
rect 1212 -5698 1380 -5664
rect 1470 -5698 1638 -5664
rect 1728 -5698 1896 -5664
rect 1986 -5698 2154 -5664
rect 2244 -5698 2412 -5664
rect 1212 -6208 1380 -6174
rect 1470 -6208 1638 -6174
rect 1728 -6208 1896 -6174
rect 1986 -6208 2154 -6174
rect 2244 -6208 2412 -6174
rect 1212 -6316 1380 -6282
rect 1470 -6316 1638 -6282
rect 1728 -6316 1896 -6282
rect 1986 -6316 2154 -6282
rect 2244 -6316 2412 -6282
rect 1212 -6826 1380 -6792
rect 1470 -6826 1638 -6792
rect 1728 -6826 1896 -6792
rect 1986 -6826 2154 -6792
rect 2244 -6826 2412 -6792
rect 1212 -6934 1380 -6900
rect 1470 -6934 1638 -6900
rect 1728 -6934 1896 -6900
rect 1986 -6934 2154 -6900
rect 2244 -6934 2412 -6900
rect 1212 -7444 1380 -7410
rect 1470 -7444 1638 -7410
rect 1728 -7444 1896 -7410
rect 1986 -7444 2154 -7410
rect 2244 -7444 2412 -7410
rect 1212 -7552 1380 -7518
rect 1470 -7552 1638 -7518
rect 1728 -7552 1896 -7518
rect 1986 -7552 2154 -7518
rect 2244 -7552 2412 -7518
rect 1212 -8062 1380 -8028
rect 1470 -8062 1638 -8028
rect 1728 -8062 1896 -8028
rect 1986 -8062 2154 -8028
rect 2244 -8062 2412 -8028
rect 3012 -4462 3180 -4428
rect 3270 -4462 3438 -4428
rect 3528 -4462 3696 -4428
rect 3786 -4462 3954 -4428
rect 4044 -4462 4212 -4428
rect 3012 -4972 3180 -4938
rect 3270 -4972 3438 -4938
rect 3528 -4972 3696 -4938
rect 3786 -4972 3954 -4938
rect 4044 -4972 4212 -4938
rect 3012 -5080 3180 -5046
rect 3270 -5080 3438 -5046
rect 3528 -5080 3696 -5046
rect 3786 -5080 3954 -5046
rect 4044 -5080 4212 -5046
rect 3012 -5590 3180 -5556
rect 3270 -5590 3438 -5556
rect 3528 -5590 3696 -5556
rect 3786 -5590 3954 -5556
rect 4044 -5590 4212 -5556
rect 3012 -5698 3180 -5664
rect 3270 -5698 3438 -5664
rect 3528 -5698 3696 -5664
rect 3786 -5698 3954 -5664
rect 4044 -5698 4212 -5664
rect 3012 -6208 3180 -6174
rect 3270 -6208 3438 -6174
rect 3528 -6208 3696 -6174
rect 3786 -6208 3954 -6174
rect 4044 -6208 4212 -6174
rect 3012 -6316 3180 -6282
rect 3270 -6316 3438 -6282
rect 3528 -6316 3696 -6282
rect 3786 -6316 3954 -6282
rect 4044 -6316 4212 -6282
rect 3012 -6826 3180 -6792
rect 3270 -6826 3438 -6792
rect 3528 -6826 3696 -6792
rect 3786 -6826 3954 -6792
rect 4044 -6826 4212 -6792
rect 3012 -6934 3180 -6900
rect 3270 -6934 3438 -6900
rect 3528 -6934 3696 -6900
rect 3786 -6934 3954 -6900
rect 4044 -6934 4212 -6900
rect 3012 -7444 3180 -7410
rect 3270 -7444 3438 -7410
rect 3528 -7444 3696 -7410
rect 3786 -7444 3954 -7410
rect 4044 -7444 4212 -7410
rect 3012 -7552 3180 -7518
rect 3270 -7552 3438 -7518
rect 3528 -7552 3696 -7518
rect 3786 -7552 3954 -7518
rect 4044 -7552 4212 -7518
rect 3012 -8062 3180 -8028
rect 3270 -8062 3438 -8028
rect 3528 -8062 3696 -8028
rect 3786 -8062 3954 -8028
rect 4044 -8062 4212 -8028
<< xpolycontact >>
rect -74 1678 208 2110
rect -74 446 208 878
rect 304 1678 586 2110
rect 304 446 586 878
rect 682 1678 964 2110
rect 682 446 964 878
rect 1060 1678 1342 2110
rect 1060 446 1342 878
rect 1438 1678 1720 2110
rect 1438 446 1720 878
rect 1816 1678 2098 2110
rect 1816 446 2098 878
<< xpolyres >>
rect -74 878 208 1678
rect 304 878 586 1678
rect 682 878 964 1678
rect 1060 878 1342 1678
rect 1438 878 1720 1678
rect 1816 878 2098 1678
<< locali >>
rect -204 2206 -108 2240
rect 2132 2206 2228 2240
rect 3420 2238 3600 2380
rect -204 2144 -170 2206
rect 2194 2144 2228 2206
rect -204 350 -170 412
rect 2336 2204 2432 2238
rect 4422 2204 4518 2238
rect 2336 2142 2370 2204
rect 4484 2142 4518 2204
rect 2482 2102 2498 2136
rect 2532 2102 2548 2136
rect 2674 2102 2690 2136
rect 2724 2102 2740 2136
rect 2866 2102 2882 2136
rect 2916 2102 2932 2136
rect 3058 2102 3074 2136
rect 3108 2102 3124 2136
rect 3250 2102 3266 2136
rect 3300 2102 3316 2136
rect 3442 2102 3458 2136
rect 3492 2102 3508 2136
rect 3634 2102 3650 2136
rect 3684 2102 3700 2136
rect 3826 2102 3842 2136
rect 3876 2102 3892 2136
rect 4018 2102 4034 2136
rect 4068 2102 4084 2136
rect 4210 2102 4226 2136
rect 4260 2102 4276 2136
rect 2450 2043 2484 2059
rect 2450 1651 2484 1667
rect 2546 2043 2580 2059
rect 2546 1651 2580 1667
rect 2642 2043 2676 2059
rect 2642 1651 2676 1667
rect 2738 2043 2772 2059
rect 2738 1651 2772 1667
rect 2834 2043 2868 2059
rect 2834 1651 2868 1667
rect 2930 2043 2964 2059
rect 2930 1651 2964 1667
rect 3026 2043 3060 2059
rect 3026 1651 3060 1667
rect 3122 2043 3156 2059
rect 3122 1651 3156 1667
rect 3218 2043 3252 2059
rect 3218 1651 3252 1667
rect 3314 2043 3348 2059
rect 3314 1651 3348 1667
rect 3410 2043 3444 2059
rect 3410 1651 3444 1667
rect 3506 2043 3540 2059
rect 3506 1651 3540 1667
rect 3602 2043 3636 2059
rect 3602 1651 3636 1667
rect 3698 2043 3732 2059
rect 3698 1651 3732 1667
rect 3794 2043 3828 2059
rect 3794 1651 3828 1667
rect 3890 2043 3924 2059
rect 3890 1651 3924 1667
rect 3986 2043 4020 2059
rect 3986 1651 4020 1667
rect 4082 2043 4116 2059
rect 4082 1651 4116 1667
rect 4178 2043 4212 2059
rect 4178 1651 4212 1667
rect 4274 2043 4308 2059
rect 4274 1651 4308 1667
rect 4370 2043 4404 2059
rect 4370 1651 4404 1667
rect 2578 1574 2594 1608
rect 2628 1574 2644 1608
rect 2770 1574 2786 1608
rect 2820 1574 2836 1608
rect 2962 1574 2978 1608
rect 3012 1574 3028 1608
rect 3154 1574 3170 1608
rect 3204 1574 3220 1608
rect 3346 1574 3362 1608
rect 3396 1574 3412 1608
rect 3538 1574 3554 1608
rect 3588 1574 3604 1608
rect 3730 1574 3746 1608
rect 3780 1574 3796 1608
rect 3922 1574 3938 1608
rect 3972 1574 3988 1608
rect 4114 1574 4130 1608
rect 4164 1574 4180 1608
rect 4306 1574 4322 1608
rect 4356 1574 4372 1608
rect 2578 1466 2594 1500
rect 2628 1466 2644 1500
rect 2770 1466 2786 1500
rect 2820 1466 2836 1500
rect 2962 1466 2978 1500
rect 3012 1466 3028 1500
rect 3154 1466 3170 1500
rect 3204 1466 3220 1500
rect 3346 1466 3362 1500
rect 3396 1466 3412 1500
rect 3538 1466 3554 1500
rect 3588 1466 3604 1500
rect 3730 1466 3746 1500
rect 3780 1466 3796 1500
rect 3922 1466 3938 1500
rect 3972 1466 3988 1500
rect 4114 1466 4130 1500
rect 4164 1466 4180 1500
rect 4306 1466 4322 1500
rect 4356 1466 4372 1500
rect 2450 1407 2484 1423
rect 2450 1015 2484 1031
rect 2546 1407 2580 1423
rect 2546 1015 2580 1031
rect 2642 1407 2676 1423
rect 2642 1015 2676 1031
rect 2738 1407 2772 1423
rect 2738 1015 2772 1031
rect 2834 1407 2868 1423
rect 2834 1015 2868 1031
rect 2930 1407 2964 1423
rect 2930 1015 2964 1031
rect 3026 1407 3060 1423
rect 3026 1015 3060 1031
rect 3122 1407 3156 1423
rect 3122 1015 3156 1031
rect 3218 1407 3252 1423
rect 3218 1015 3252 1031
rect 3314 1407 3348 1423
rect 3314 1015 3348 1031
rect 3410 1407 3444 1423
rect 3410 1015 3444 1031
rect 3506 1407 3540 1423
rect 3506 1015 3540 1031
rect 3602 1407 3636 1423
rect 3602 1015 3636 1031
rect 3698 1407 3732 1423
rect 3698 1015 3732 1031
rect 3794 1407 3828 1423
rect 3794 1015 3828 1031
rect 3890 1407 3924 1423
rect 3890 1015 3924 1031
rect 3986 1407 4020 1423
rect 3986 1015 4020 1031
rect 4082 1407 4116 1423
rect 4082 1015 4116 1031
rect 4178 1407 4212 1423
rect 4178 1015 4212 1031
rect 4274 1407 4308 1423
rect 4274 1015 4308 1031
rect 4370 1407 4404 1423
rect 4370 1015 4404 1031
rect 2482 938 2498 972
rect 2532 938 2548 972
rect 2674 938 2690 972
rect 2724 938 2740 972
rect 2866 938 2882 972
rect 2916 938 2932 972
rect 3058 938 3074 972
rect 3108 938 3124 972
rect 3250 938 3266 972
rect 3300 938 3316 972
rect 3442 938 3458 972
rect 3492 938 3508 972
rect 3634 938 3650 972
rect 3684 938 3700 972
rect 3826 938 3842 972
rect 3876 938 3892 972
rect 4018 938 4034 972
rect 4068 938 4084 972
rect 4210 938 4226 972
rect 4260 938 4276 972
rect 2336 870 2370 932
rect 4484 870 4518 932
rect 2336 836 2432 870
rect 4422 836 4518 870
rect 4836 2174 4932 2208
rect 6922 2174 7018 2208
rect 4836 2112 4870 2174
rect 2194 350 2228 412
rect -204 316 -108 350
rect 2132 316 2228 350
rect 2336 608 2432 642
rect 4422 608 4518 642
rect 2336 546 2370 608
rect 1400 200 1540 316
rect 16 166 112 200
rect 2102 166 2198 200
rect 16 104 50 166
rect 2164 104 2198 166
rect 258 64 274 98
rect 308 64 324 98
rect 450 64 466 98
rect 500 64 516 98
rect 642 64 658 98
rect 692 64 708 98
rect 834 64 850 98
rect 884 64 900 98
rect 1026 64 1042 98
rect 1076 64 1092 98
rect 1218 64 1234 98
rect 1268 64 1284 98
rect 1410 64 1426 98
rect 1460 64 1476 98
rect 1602 64 1618 98
rect 1652 64 1668 98
rect 1794 64 1810 98
rect 1844 64 1860 98
rect 1986 64 2002 98
rect 2036 64 2052 98
rect 130 14 164 30
rect 130 -378 164 -362
rect 226 14 260 30
rect 226 -378 260 -362
rect 322 14 356 30
rect 322 -378 356 -362
rect 418 14 452 30
rect 418 -378 452 -362
rect 514 14 548 30
rect 514 -378 548 -362
rect 610 14 644 30
rect 610 -378 644 -362
rect 706 14 740 30
rect 706 -378 740 -362
rect 802 14 836 30
rect 802 -378 836 -362
rect 898 14 932 30
rect 898 -378 932 -362
rect 994 14 1028 30
rect 994 -378 1028 -362
rect 1090 14 1124 30
rect 1090 -378 1124 -362
rect 1186 14 1220 30
rect 1186 -378 1220 -362
rect 1282 14 1316 30
rect 1282 -378 1316 -362
rect 1378 14 1412 30
rect 1378 -378 1412 -362
rect 1474 14 1508 30
rect 1474 -378 1508 -362
rect 1570 14 1604 30
rect 1570 -378 1604 -362
rect 1666 14 1700 30
rect 1666 -378 1700 -362
rect 1762 14 1796 30
rect 1762 -378 1796 -362
rect 1858 14 1892 30
rect 1858 -378 1892 -362
rect 1954 14 1988 30
rect 1954 -378 1988 -362
rect 2050 14 2084 30
rect 2050 -378 2084 -362
rect 162 -446 178 -412
rect 212 -446 228 -412
rect 354 -446 370 -412
rect 404 -446 420 -412
rect 546 -446 562 -412
rect 596 -446 612 -412
rect 738 -446 754 -412
rect 788 -446 804 -412
rect 930 -446 946 -412
rect 980 -446 996 -412
rect 1122 -446 1138 -412
rect 1172 -446 1188 -412
rect 1314 -446 1330 -412
rect 1364 -446 1380 -412
rect 1506 -446 1522 -412
rect 1556 -446 1572 -412
rect 1698 -446 1714 -412
rect 1748 -446 1764 -412
rect 1890 -446 1906 -412
rect 1940 -446 1956 -412
rect 162 -554 178 -520
rect 212 -554 228 -520
rect 354 -554 370 -520
rect 404 -554 420 -520
rect 546 -554 562 -520
rect 596 -554 612 -520
rect 738 -554 754 -520
rect 788 -554 804 -520
rect 930 -554 946 -520
rect 980 -554 996 -520
rect 1122 -554 1138 -520
rect 1172 -554 1188 -520
rect 1314 -554 1330 -520
rect 1364 -554 1380 -520
rect 1506 -554 1522 -520
rect 1556 -554 1572 -520
rect 1698 -554 1714 -520
rect 1748 -554 1764 -520
rect 1890 -554 1906 -520
rect 1940 -554 1956 -520
rect 130 -604 164 -588
rect 130 -996 164 -980
rect 226 -604 260 -588
rect 226 -996 260 -980
rect 322 -604 356 -588
rect 322 -996 356 -980
rect 418 -604 452 -588
rect 418 -996 452 -980
rect 514 -604 548 -588
rect 514 -996 548 -980
rect 610 -604 644 -588
rect 610 -996 644 -980
rect 706 -604 740 -588
rect 706 -996 740 -980
rect 802 -604 836 -588
rect 802 -996 836 -980
rect 898 -604 932 -588
rect 898 -996 932 -980
rect 994 -604 1028 -588
rect 994 -996 1028 -980
rect 1090 -604 1124 -588
rect 1090 -996 1124 -980
rect 1186 -604 1220 -588
rect 1186 -996 1220 -980
rect 1282 -604 1316 -588
rect 1282 -996 1316 -980
rect 1378 -604 1412 -588
rect 1378 -996 1412 -980
rect 1474 -604 1508 -588
rect 1474 -996 1508 -980
rect 1570 -604 1604 -588
rect 1570 -996 1604 -980
rect 1666 -604 1700 -588
rect 1666 -996 1700 -980
rect 1762 -604 1796 -588
rect 1762 -996 1796 -980
rect 1858 -604 1892 -588
rect 1858 -996 1892 -980
rect 1954 -604 1988 -588
rect 1954 -996 1988 -980
rect 2050 -604 2084 -588
rect 2050 -996 2084 -980
rect 258 -1064 274 -1030
rect 308 -1064 324 -1030
rect 450 -1064 466 -1030
rect 500 -1064 516 -1030
rect 642 -1064 658 -1030
rect 692 -1064 708 -1030
rect 834 -1064 850 -1030
rect 884 -1064 900 -1030
rect 1026 -1064 1042 -1030
rect 1076 -1064 1092 -1030
rect 1218 -1064 1234 -1030
rect 1268 -1064 1284 -1030
rect 1410 -1064 1426 -1030
rect 1460 -1064 1476 -1030
rect 1602 -1064 1618 -1030
rect 1652 -1064 1668 -1030
rect 1794 -1064 1810 -1030
rect 1844 -1064 1860 -1030
rect 1986 -1064 2002 -1030
rect 2036 -1064 2052 -1030
rect 258 -1172 274 -1138
rect 308 -1172 324 -1138
rect 450 -1172 466 -1138
rect 500 -1172 516 -1138
rect 642 -1172 658 -1138
rect 692 -1172 708 -1138
rect 834 -1172 850 -1138
rect 884 -1172 900 -1138
rect 1026 -1172 1042 -1138
rect 1076 -1172 1092 -1138
rect 1218 -1172 1234 -1138
rect 1268 -1172 1284 -1138
rect 1410 -1172 1426 -1138
rect 1460 -1172 1476 -1138
rect 1602 -1172 1618 -1138
rect 1652 -1172 1668 -1138
rect 1794 -1172 1810 -1138
rect 1844 -1172 1860 -1138
rect 1986 -1172 2002 -1138
rect 2036 -1172 2052 -1138
rect 130 -1222 164 -1206
rect 130 -1614 164 -1598
rect 226 -1222 260 -1206
rect 226 -1614 260 -1598
rect 322 -1222 356 -1206
rect 322 -1614 356 -1598
rect 418 -1222 452 -1206
rect 418 -1614 452 -1598
rect 514 -1222 548 -1206
rect 514 -1614 548 -1598
rect 610 -1222 644 -1206
rect 610 -1614 644 -1598
rect 706 -1222 740 -1206
rect 706 -1614 740 -1598
rect 802 -1222 836 -1206
rect 802 -1614 836 -1598
rect 898 -1222 932 -1206
rect 898 -1614 932 -1598
rect 994 -1222 1028 -1206
rect 994 -1614 1028 -1598
rect 1090 -1222 1124 -1206
rect 1090 -1614 1124 -1598
rect 1186 -1222 1220 -1206
rect 1186 -1614 1220 -1598
rect 1282 -1222 1316 -1206
rect 1282 -1614 1316 -1598
rect 1378 -1222 1412 -1206
rect 1378 -1614 1412 -1598
rect 1474 -1222 1508 -1206
rect 1474 -1614 1508 -1598
rect 1570 -1222 1604 -1206
rect 1570 -1614 1604 -1598
rect 1666 -1222 1700 -1206
rect 1666 -1614 1700 -1598
rect 1762 -1222 1796 -1206
rect 1762 -1614 1796 -1598
rect 1858 -1222 1892 -1206
rect 1858 -1614 1892 -1598
rect 1954 -1222 1988 -1206
rect 1954 -1614 1988 -1598
rect 2050 -1222 2084 -1206
rect 2050 -1614 2084 -1598
rect 162 -1682 178 -1648
rect 212 -1682 228 -1648
rect 354 -1682 370 -1648
rect 404 -1682 420 -1648
rect 546 -1682 562 -1648
rect 596 -1682 612 -1648
rect 738 -1682 754 -1648
rect 788 -1682 804 -1648
rect 930 -1682 946 -1648
rect 980 -1682 996 -1648
rect 1122 -1682 1138 -1648
rect 1172 -1682 1188 -1648
rect 1314 -1682 1330 -1648
rect 1364 -1682 1380 -1648
rect 1506 -1682 1522 -1648
rect 1556 -1682 1572 -1648
rect 1698 -1682 1714 -1648
rect 1748 -1682 1764 -1648
rect 1890 -1682 1906 -1648
rect 1940 -1682 1956 -1648
rect 16 -1750 50 -1688
rect 2198 -360 2336 -200
rect 4484 546 4518 608
rect 2482 506 2498 540
rect 2532 506 2548 540
rect 2674 506 2690 540
rect 2724 506 2740 540
rect 2866 506 2882 540
rect 2916 506 2932 540
rect 3058 506 3074 540
rect 3108 506 3124 540
rect 3250 506 3266 540
rect 3300 506 3316 540
rect 3442 506 3458 540
rect 3492 506 3508 540
rect 3634 506 3650 540
rect 3684 506 3700 540
rect 3826 506 3842 540
rect 3876 506 3892 540
rect 4018 506 4034 540
rect 4068 506 4084 540
rect 4210 506 4226 540
rect 4260 506 4276 540
rect 2450 456 2484 472
rect 2450 64 2484 80
rect 2546 456 2580 472
rect 2546 64 2580 80
rect 2642 456 2676 472
rect 2642 64 2676 80
rect 2738 456 2772 472
rect 2738 64 2772 80
rect 2834 456 2868 472
rect 2834 64 2868 80
rect 2930 456 2964 472
rect 2930 64 2964 80
rect 3026 456 3060 472
rect 3026 64 3060 80
rect 3122 456 3156 472
rect 3122 64 3156 80
rect 3218 456 3252 472
rect 3218 64 3252 80
rect 3314 456 3348 472
rect 3314 64 3348 80
rect 3410 456 3444 472
rect 3410 64 3444 80
rect 3506 456 3540 472
rect 3506 64 3540 80
rect 3602 456 3636 472
rect 3602 64 3636 80
rect 3698 456 3732 472
rect 3698 64 3732 80
rect 3794 456 3828 472
rect 3794 64 3828 80
rect 3890 456 3924 472
rect 3890 64 3924 80
rect 3986 456 4020 472
rect 3986 64 4020 80
rect 4082 456 4116 472
rect 4082 64 4116 80
rect 4178 456 4212 472
rect 4178 64 4212 80
rect 4274 456 4308 472
rect 4274 64 4308 80
rect 4370 456 4404 472
rect 4370 64 4404 80
rect 2578 -4 2594 30
rect 2628 -4 2644 30
rect 2770 -4 2786 30
rect 2820 -4 2836 30
rect 2962 -4 2978 30
rect 3012 -4 3028 30
rect 3154 -4 3170 30
rect 3204 -4 3220 30
rect 3346 -4 3362 30
rect 3396 -4 3412 30
rect 3538 -4 3554 30
rect 3588 -4 3604 30
rect 3730 -4 3746 30
rect 3780 -4 3796 30
rect 3922 -4 3938 30
rect 3972 -4 3988 30
rect 4114 -4 4130 30
rect 4164 -4 4180 30
rect 4306 -4 4322 30
rect 4356 -4 4372 30
rect 2578 -112 2594 -78
rect 2628 -112 2644 -78
rect 2770 -112 2786 -78
rect 2820 -112 2836 -78
rect 2962 -112 2978 -78
rect 3012 -112 3028 -78
rect 3154 -112 3170 -78
rect 3204 -112 3220 -78
rect 3346 -112 3362 -78
rect 3396 -112 3412 -78
rect 3538 -112 3554 -78
rect 3588 -112 3604 -78
rect 3730 -112 3746 -78
rect 3780 -112 3796 -78
rect 3922 -112 3938 -78
rect 3972 -112 3988 -78
rect 4114 -112 4130 -78
rect 4164 -112 4180 -78
rect 4306 -112 4322 -78
rect 4356 -112 4372 -78
rect 2450 -162 2484 -146
rect 2450 -554 2484 -538
rect 2546 -162 2580 -146
rect 2546 -554 2580 -538
rect 2642 -162 2676 -146
rect 2642 -554 2676 -538
rect 2738 -162 2772 -146
rect 2738 -554 2772 -538
rect 2834 -162 2868 -146
rect 2834 -554 2868 -538
rect 2930 -162 2964 -146
rect 2930 -554 2964 -538
rect 3026 -162 3060 -146
rect 3026 -554 3060 -538
rect 3122 -162 3156 -146
rect 3122 -554 3156 -538
rect 3218 -162 3252 -146
rect 3218 -554 3252 -538
rect 3314 -162 3348 -146
rect 3314 -554 3348 -538
rect 3410 -162 3444 -146
rect 3410 -554 3444 -538
rect 3506 -162 3540 -146
rect 3506 -554 3540 -538
rect 3602 -162 3636 -146
rect 3602 -554 3636 -538
rect 3698 -162 3732 -146
rect 3698 -554 3732 -538
rect 3794 -162 3828 -146
rect 3794 -554 3828 -538
rect 3890 -162 3924 -146
rect 3890 -554 3924 -538
rect 3986 -162 4020 -146
rect 3986 -554 4020 -538
rect 4082 -162 4116 -146
rect 4082 -554 4116 -538
rect 4178 -162 4212 -146
rect 4178 -554 4212 -538
rect 4274 -162 4308 -146
rect 4274 -554 4308 -538
rect 4370 -162 4404 -146
rect 4370 -554 4404 -538
rect 2482 -622 2498 -588
rect 2532 -622 2548 -588
rect 2674 -622 2690 -588
rect 2724 -622 2740 -588
rect 2866 -622 2882 -588
rect 2916 -622 2932 -588
rect 3058 -622 3074 -588
rect 3108 -622 3124 -588
rect 3250 -622 3266 -588
rect 3300 -622 3316 -588
rect 3442 -622 3458 -588
rect 3492 -622 3508 -588
rect 3634 -622 3650 -588
rect 3684 -622 3700 -588
rect 3826 -622 3842 -588
rect 3876 -622 3892 -588
rect 4018 -622 4034 -588
rect 4068 -622 4084 -588
rect 4210 -622 4226 -588
rect 4260 -622 4276 -588
rect 2336 -690 2370 -628
rect 4484 -690 4518 -628
rect 2336 -724 2432 -690
rect 4422 -724 4518 -690
rect 2164 -1750 2198 -1688
rect 16 -1784 112 -1750
rect 2102 -1784 2198 -1750
rect 1260 -2180 1460 -1784
rect -2564 -2214 -2468 -2180
rect -1438 -2214 -1342 -2180
rect -2564 -2276 -2530 -2214
rect -1376 -2276 -1342 -2214
rect -2322 -2316 -2306 -2282
rect -2272 -2316 -2256 -2282
rect -2130 -2316 -2114 -2282
rect -2080 -2316 -2064 -2282
rect -1938 -2316 -1922 -2282
rect -1888 -2316 -1872 -2282
rect -1746 -2316 -1730 -2282
rect -1696 -2316 -1680 -2282
rect -1554 -2316 -1538 -2282
rect -1504 -2316 -1488 -2282
rect -2450 -2366 -2416 -2350
rect -2450 -2758 -2416 -2742
rect -2354 -2366 -2320 -2350
rect -2354 -2758 -2320 -2742
rect -2258 -2366 -2224 -2350
rect -2258 -2758 -2224 -2742
rect -2162 -2366 -2128 -2350
rect -2162 -2758 -2128 -2742
rect -2066 -2366 -2032 -2350
rect -2066 -2758 -2032 -2742
rect -1970 -2366 -1936 -2350
rect -1970 -2758 -1936 -2742
rect -1874 -2366 -1840 -2350
rect -1874 -2758 -1840 -2742
rect -1778 -2366 -1744 -2350
rect -1778 -2758 -1744 -2742
rect -1682 -2366 -1648 -2350
rect -1682 -2758 -1648 -2742
rect -1586 -2366 -1552 -2350
rect -1586 -2758 -1552 -2742
rect -1490 -2366 -1456 -2350
rect -1490 -2758 -1456 -2742
rect -2418 -2826 -2402 -2792
rect -2368 -2826 -2352 -2792
rect -2226 -2826 -2210 -2792
rect -2176 -2826 -2160 -2792
rect -2034 -2826 -2018 -2792
rect -1984 -2826 -1968 -2792
rect -1842 -2826 -1826 -2792
rect -1792 -2826 -1776 -2792
rect -1650 -2826 -1634 -2792
rect -1600 -2826 -1584 -2792
rect -2418 -2934 -2402 -2900
rect -2368 -2934 -2352 -2900
rect -2226 -2934 -2210 -2900
rect -2176 -2934 -2160 -2900
rect -2034 -2934 -2018 -2900
rect -1984 -2934 -1968 -2900
rect -1842 -2934 -1826 -2900
rect -1792 -2934 -1776 -2900
rect -1650 -2934 -1634 -2900
rect -1600 -2934 -1584 -2900
rect -2450 -2984 -2416 -2968
rect -2450 -3376 -2416 -3360
rect -2354 -2984 -2320 -2968
rect -2354 -3376 -2320 -3360
rect -2258 -2984 -2224 -2968
rect -2258 -3376 -2224 -3360
rect -2162 -2984 -2128 -2968
rect -2162 -3376 -2128 -3360
rect -2066 -2984 -2032 -2968
rect -2066 -3376 -2032 -3360
rect -1970 -2984 -1936 -2968
rect -1970 -3376 -1936 -3360
rect -1874 -2984 -1840 -2968
rect -1874 -3376 -1840 -3360
rect -1778 -2984 -1744 -2968
rect -1778 -3376 -1744 -3360
rect -1682 -2984 -1648 -2968
rect -1682 -3376 -1648 -3360
rect -1586 -2984 -1552 -2968
rect -1586 -3376 -1552 -3360
rect -1490 -2984 -1456 -2968
rect -1490 -3376 -1456 -3360
rect -2322 -3444 -2306 -3410
rect -2272 -3444 -2256 -3410
rect -2130 -3444 -2114 -3410
rect -2080 -3444 -2064 -3410
rect -1938 -3444 -1922 -3410
rect -1888 -3444 -1872 -3410
rect -1746 -3444 -1730 -3410
rect -1696 -3444 -1680 -3410
rect -1554 -3444 -1538 -3410
rect -1504 -3444 -1488 -3410
rect -2322 -3552 -2306 -3518
rect -2272 -3552 -2256 -3518
rect -2130 -3552 -2114 -3518
rect -2080 -3552 -2064 -3518
rect -1938 -3552 -1922 -3518
rect -1888 -3552 -1872 -3518
rect -1746 -3552 -1730 -3518
rect -1696 -3552 -1680 -3518
rect -1554 -3552 -1538 -3518
rect -1504 -3552 -1488 -3518
rect -2450 -3602 -2416 -3586
rect -2450 -3994 -2416 -3978
rect -2354 -3602 -2320 -3586
rect -2354 -3994 -2320 -3978
rect -2258 -3602 -2224 -3586
rect -2258 -3994 -2224 -3978
rect -2162 -3602 -2128 -3586
rect -2162 -3994 -2128 -3978
rect -2066 -3602 -2032 -3586
rect -2066 -3994 -2032 -3978
rect -1970 -3602 -1936 -3586
rect -1970 -3994 -1936 -3978
rect -1874 -3602 -1840 -3586
rect -1874 -3994 -1840 -3978
rect -1778 -3602 -1744 -3586
rect -1778 -3994 -1744 -3978
rect -1682 -3602 -1648 -3586
rect -1682 -3994 -1648 -3978
rect -1586 -3602 -1552 -3586
rect -1586 -3994 -1552 -3978
rect -1490 -3602 -1456 -3586
rect -1490 -3994 -1456 -3978
rect -2418 -4062 -2402 -4028
rect -2368 -4062 -2352 -4028
rect -2226 -4062 -2210 -4028
rect -2176 -4062 -2160 -4028
rect -2034 -4062 -2018 -4028
rect -1984 -4062 -1968 -4028
rect -1842 -4062 -1826 -4028
rect -1792 -4062 -1776 -4028
rect -1650 -4062 -1634 -4028
rect -1600 -4062 -1584 -4028
rect -2564 -4130 -2530 -4068
rect -1376 -4130 -1342 -4068
rect -2564 -4164 -2468 -4130
rect -1438 -4164 -1342 -4130
rect -764 -2214 -668 -2180
rect 362 -2214 458 -2180
rect -764 -2276 -730 -2214
rect 424 -2276 458 -2214
rect -522 -2316 -506 -2282
rect -472 -2316 -456 -2282
rect -330 -2316 -314 -2282
rect -280 -2316 -264 -2282
rect -138 -2316 -122 -2282
rect -88 -2316 -72 -2282
rect 54 -2316 70 -2282
rect 104 -2316 120 -2282
rect 246 -2316 262 -2282
rect 296 -2316 312 -2282
rect -650 -2366 -616 -2350
rect -650 -2758 -616 -2742
rect -554 -2366 -520 -2350
rect -554 -2758 -520 -2742
rect -458 -2366 -424 -2350
rect -458 -2758 -424 -2742
rect -362 -2366 -328 -2350
rect -362 -2758 -328 -2742
rect -266 -2366 -232 -2350
rect -266 -2758 -232 -2742
rect -170 -2366 -136 -2350
rect -170 -2758 -136 -2742
rect -74 -2366 -40 -2350
rect -74 -2758 -40 -2742
rect 22 -2366 56 -2350
rect 22 -2758 56 -2742
rect 118 -2366 152 -2350
rect 118 -2758 152 -2742
rect 214 -2366 248 -2350
rect 214 -2758 248 -2742
rect 310 -2366 344 -2350
rect 310 -2758 344 -2742
rect -618 -2826 -602 -2792
rect -568 -2826 -552 -2792
rect -426 -2826 -410 -2792
rect -376 -2826 -360 -2792
rect -234 -2826 -218 -2792
rect -184 -2826 -168 -2792
rect -42 -2826 -26 -2792
rect 8 -2826 24 -2792
rect 150 -2826 166 -2792
rect 200 -2826 216 -2792
rect -618 -2934 -602 -2900
rect -568 -2934 -552 -2900
rect -426 -2934 -410 -2900
rect -376 -2934 -360 -2900
rect -234 -2934 -218 -2900
rect -184 -2934 -168 -2900
rect -42 -2934 -26 -2900
rect 8 -2934 24 -2900
rect 150 -2934 166 -2900
rect 200 -2934 216 -2900
rect -650 -2984 -616 -2968
rect -650 -3376 -616 -3360
rect -554 -2984 -520 -2968
rect -554 -3376 -520 -3360
rect -458 -2984 -424 -2968
rect -458 -3376 -424 -3360
rect -362 -2984 -328 -2968
rect -362 -3376 -328 -3360
rect -266 -2984 -232 -2968
rect -266 -3376 -232 -3360
rect -170 -2984 -136 -2968
rect -170 -3376 -136 -3360
rect -74 -2984 -40 -2968
rect -74 -3376 -40 -3360
rect 22 -2984 56 -2968
rect 22 -3376 56 -3360
rect 118 -2984 152 -2968
rect 118 -3376 152 -3360
rect 214 -2984 248 -2968
rect 214 -3376 248 -3360
rect 310 -2984 344 -2968
rect 310 -3376 344 -3360
rect -522 -3444 -506 -3410
rect -472 -3444 -456 -3410
rect -330 -3444 -314 -3410
rect -280 -3444 -264 -3410
rect -138 -3444 -122 -3410
rect -88 -3444 -72 -3410
rect 54 -3444 70 -3410
rect 104 -3444 120 -3410
rect 246 -3444 262 -3410
rect 296 -3444 312 -3410
rect -522 -3552 -506 -3518
rect -472 -3552 -456 -3518
rect -330 -3552 -314 -3518
rect -280 -3552 -264 -3518
rect -138 -3552 -122 -3518
rect -88 -3552 -72 -3518
rect 54 -3552 70 -3518
rect 104 -3552 120 -3518
rect 246 -3552 262 -3518
rect 296 -3552 312 -3518
rect -650 -3602 -616 -3586
rect -650 -3994 -616 -3978
rect -554 -3602 -520 -3586
rect -554 -3994 -520 -3978
rect -458 -3602 -424 -3586
rect -458 -3994 -424 -3978
rect -362 -3602 -328 -3586
rect -362 -3994 -328 -3978
rect -266 -3602 -232 -3586
rect -266 -3994 -232 -3978
rect -170 -3602 -136 -3586
rect -170 -3994 -136 -3978
rect -74 -3602 -40 -3586
rect -74 -3994 -40 -3978
rect 22 -3602 56 -3586
rect 22 -3994 56 -3978
rect 118 -3602 152 -3586
rect 118 -3994 152 -3978
rect 214 -3602 248 -3586
rect 214 -3994 248 -3978
rect 310 -3602 344 -3586
rect 310 -3994 344 -3978
rect -618 -4062 -602 -4028
rect -568 -4062 -552 -4028
rect -426 -4062 -410 -4028
rect -376 -4062 -360 -4028
rect -234 -4062 -218 -4028
rect -184 -4062 -168 -4028
rect -42 -4062 -26 -4028
rect 8 -4062 24 -4028
rect 150 -4062 166 -4028
rect 200 -4062 216 -4028
rect -764 -4130 -730 -4068
rect 424 -4130 458 -4068
rect -764 -4164 -668 -4130
rect 362 -4164 458 -4130
rect 1036 -2214 1132 -2180
rect 2162 -2214 2258 -2180
rect 1036 -2276 1070 -2214
rect 2224 -2276 2258 -2214
rect 1278 -2316 1294 -2282
rect 1328 -2316 1344 -2282
rect 1470 -2316 1486 -2282
rect 1520 -2316 1536 -2282
rect 1662 -2316 1678 -2282
rect 1712 -2316 1728 -2282
rect 1854 -2316 1870 -2282
rect 1904 -2316 1920 -2282
rect 2046 -2316 2062 -2282
rect 2096 -2316 2112 -2282
rect 1150 -2366 1184 -2350
rect 1150 -2758 1184 -2742
rect 1246 -2366 1280 -2350
rect 1246 -2758 1280 -2742
rect 1342 -2366 1376 -2350
rect 1342 -2758 1376 -2742
rect 1438 -2366 1472 -2350
rect 1438 -2758 1472 -2742
rect 1534 -2366 1568 -2350
rect 1534 -2758 1568 -2742
rect 1630 -2366 1664 -2350
rect 1630 -2758 1664 -2742
rect 1726 -2366 1760 -2350
rect 1726 -2758 1760 -2742
rect 1822 -2366 1856 -2350
rect 1822 -2758 1856 -2742
rect 1918 -2366 1952 -2350
rect 1918 -2758 1952 -2742
rect 2014 -2366 2048 -2350
rect 2014 -2758 2048 -2742
rect 2110 -2366 2144 -2350
rect 2110 -2758 2144 -2742
rect 1182 -2826 1198 -2792
rect 1232 -2826 1248 -2792
rect 1374 -2826 1390 -2792
rect 1424 -2826 1440 -2792
rect 1566 -2826 1582 -2792
rect 1616 -2826 1632 -2792
rect 1758 -2826 1774 -2792
rect 1808 -2826 1824 -2792
rect 1950 -2826 1966 -2792
rect 2000 -2826 2016 -2792
rect 1182 -2934 1198 -2900
rect 1232 -2934 1248 -2900
rect 1374 -2934 1390 -2900
rect 1424 -2934 1440 -2900
rect 1566 -2934 1582 -2900
rect 1616 -2934 1632 -2900
rect 1758 -2934 1774 -2900
rect 1808 -2934 1824 -2900
rect 1950 -2934 1966 -2900
rect 2000 -2934 2016 -2900
rect 1150 -2984 1184 -2968
rect 1150 -3376 1184 -3360
rect 1246 -2984 1280 -2968
rect 1246 -3376 1280 -3360
rect 1342 -2984 1376 -2968
rect 1342 -3376 1376 -3360
rect 1438 -2984 1472 -2968
rect 1438 -3376 1472 -3360
rect 1534 -2984 1568 -2968
rect 1534 -3376 1568 -3360
rect 1630 -2984 1664 -2968
rect 1630 -3376 1664 -3360
rect 1726 -2984 1760 -2968
rect 1726 -3376 1760 -3360
rect 1822 -2984 1856 -2968
rect 1822 -3376 1856 -3360
rect 1918 -2984 1952 -2968
rect 1918 -3376 1952 -3360
rect 2014 -2984 2048 -2968
rect 2014 -3376 2048 -3360
rect 2110 -2984 2144 -2968
rect 2110 -3376 2144 -3360
rect 1278 -3444 1294 -3410
rect 1328 -3444 1344 -3410
rect 1470 -3444 1486 -3410
rect 1520 -3444 1536 -3410
rect 1662 -3444 1678 -3410
rect 1712 -3444 1728 -3410
rect 1854 -3444 1870 -3410
rect 1904 -3444 1920 -3410
rect 2046 -3444 2062 -3410
rect 2096 -3444 2112 -3410
rect 1278 -3552 1294 -3518
rect 1328 -3552 1344 -3518
rect 1470 -3552 1486 -3518
rect 1520 -3552 1536 -3518
rect 1662 -3552 1678 -3518
rect 1712 -3552 1728 -3518
rect 1854 -3552 1870 -3518
rect 1904 -3552 1920 -3518
rect 2046 -3552 2062 -3518
rect 2096 -3552 2112 -3518
rect 1150 -3602 1184 -3586
rect 1150 -3994 1184 -3978
rect 1246 -3602 1280 -3586
rect 1246 -3994 1280 -3978
rect 1342 -3602 1376 -3586
rect 1342 -3994 1376 -3978
rect 1438 -3602 1472 -3586
rect 1438 -3994 1472 -3978
rect 1534 -3602 1568 -3586
rect 1534 -3994 1568 -3978
rect 1630 -3602 1664 -3586
rect 1630 -3994 1664 -3978
rect 1726 -3602 1760 -3586
rect 1726 -3994 1760 -3978
rect 1822 -3602 1856 -3586
rect 1822 -3994 1856 -3978
rect 1918 -3602 1952 -3586
rect 1918 -3994 1952 -3978
rect 2014 -3602 2048 -3586
rect 2014 -3994 2048 -3978
rect 2110 -3602 2144 -3586
rect 2110 -3994 2144 -3978
rect 1182 -4062 1198 -4028
rect 1232 -4062 1248 -4028
rect 1374 -4062 1390 -4028
rect 1424 -4062 1440 -4028
rect 1566 -4062 1582 -4028
rect 1616 -4062 1632 -4028
rect 1758 -4062 1774 -4028
rect 1808 -4062 1824 -4028
rect 1950 -4062 1966 -4028
rect 2000 -4062 2016 -4028
rect 1036 -4130 1070 -4068
rect 2224 -4130 2258 -4068
rect 1036 -4164 1132 -4130
rect 2162 -4164 2258 -4130
rect 2836 -2214 2932 -2180
rect 3962 -2214 4058 -2180
rect 2836 -2276 2870 -2214
rect 4024 -2276 4058 -2214
rect 3078 -2316 3094 -2282
rect 3128 -2316 3144 -2282
rect 3270 -2316 3286 -2282
rect 3320 -2316 3336 -2282
rect 3462 -2316 3478 -2282
rect 3512 -2316 3528 -2282
rect 3654 -2316 3670 -2282
rect 3704 -2316 3720 -2282
rect 3846 -2316 3862 -2282
rect 3896 -2316 3912 -2282
rect 2950 -2366 2984 -2350
rect 2950 -2758 2984 -2742
rect 3046 -2366 3080 -2350
rect 3046 -2758 3080 -2742
rect 3142 -2366 3176 -2350
rect 3142 -2758 3176 -2742
rect 3238 -2366 3272 -2350
rect 3238 -2758 3272 -2742
rect 3334 -2366 3368 -2350
rect 3334 -2758 3368 -2742
rect 3430 -2366 3464 -2350
rect 3430 -2758 3464 -2742
rect 3526 -2366 3560 -2350
rect 3526 -2758 3560 -2742
rect 3622 -2366 3656 -2350
rect 3622 -2758 3656 -2742
rect 3718 -2366 3752 -2350
rect 3718 -2758 3752 -2742
rect 3814 -2366 3848 -2350
rect 3814 -2758 3848 -2742
rect 3910 -2366 3944 -2350
rect 3910 -2758 3944 -2742
rect 2982 -2826 2998 -2792
rect 3032 -2826 3048 -2792
rect 3174 -2826 3190 -2792
rect 3224 -2826 3240 -2792
rect 3366 -2826 3382 -2792
rect 3416 -2826 3432 -2792
rect 3558 -2826 3574 -2792
rect 3608 -2826 3624 -2792
rect 3750 -2826 3766 -2792
rect 3800 -2826 3816 -2792
rect 2982 -2934 2998 -2900
rect 3032 -2934 3048 -2900
rect 3174 -2934 3190 -2900
rect 3224 -2934 3240 -2900
rect 3366 -2934 3382 -2900
rect 3416 -2934 3432 -2900
rect 3558 -2934 3574 -2900
rect 3608 -2934 3624 -2900
rect 3750 -2934 3766 -2900
rect 3800 -2934 3816 -2900
rect 2950 -2984 2984 -2968
rect 2950 -3376 2984 -3360
rect 3046 -2984 3080 -2968
rect 3046 -3376 3080 -3360
rect 3142 -2984 3176 -2968
rect 3142 -3376 3176 -3360
rect 3238 -2984 3272 -2968
rect 3238 -3376 3272 -3360
rect 3334 -2984 3368 -2968
rect 3334 -3376 3368 -3360
rect 3430 -2984 3464 -2968
rect 3430 -3376 3464 -3360
rect 3526 -2984 3560 -2968
rect 3526 -3376 3560 -3360
rect 3622 -2984 3656 -2968
rect 3622 -3376 3656 -3360
rect 3718 -2984 3752 -2968
rect 3718 -3376 3752 -3360
rect 3814 -2984 3848 -2968
rect 3814 -3376 3848 -3360
rect 3910 -2984 3944 -2968
rect 3910 -3376 3944 -3360
rect 3078 -3444 3094 -3410
rect 3128 -3444 3144 -3410
rect 3270 -3444 3286 -3410
rect 3320 -3444 3336 -3410
rect 3462 -3444 3478 -3410
rect 3512 -3444 3528 -3410
rect 3654 -3444 3670 -3410
rect 3704 -3444 3720 -3410
rect 3846 -3444 3862 -3410
rect 3896 -3444 3912 -3410
rect 3078 -3552 3094 -3518
rect 3128 -3552 3144 -3518
rect 3270 -3552 3286 -3518
rect 3320 -3552 3336 -3518
rect 3462 -3552 3478 -3518
rect 3512 -3552 3528 -3518
rect 3654 -3552 3670 -3518
rect 3704 -3552 3720 -3518
rect 3846 -3552 3862 -3518
rect 3896 -3552 3912 -3518
rect 2950 -3602 2984 -3586
rect 2950 -3994 2984 -3978
rect 3046 -3602 3080 -3586
rect 3046 -3994 3080 -3978
rect 3142 -3602 3176 -3586
rect 3142 -3994 3176 -3978
rect 3238 -3602 3272 -3586
rect 3238 -3994 3272 -3978
rect 3334 -3602 3368 -3586
rect 3334 -3994 3368 -3978
rect 3430 -3602 3464 -3586
rect 3430 -3994 3464 -3978
rect 3526 -3602 3560 -3586
rect 3526 -3994 3560 -3978
rect 3622 -3602 3656 -3586
rect 3622 -3994 3656 -3978
rect 3718 -3602 3752 -3586
rect 3718 -3994 3752 -3978
rect 3814 -3602 3848 -3586
rect 3814 -3994 3848 -3978
rect 3910 -3602 3944 -3586
rect 3910 -3994 3944 -3978
rect 2982 -4062 2998 -4028
rect 3032 -4062 3048 -4028
rect 3174 -4062 3190 -4028
rect 3224 -4062 3240 -4028
rect 3366 -4062 3382 -4028
rect 3416 -4062 3432 -4028
rect 3558 -4062 3574 -4028
rect 3608 -4062 3624 -4028
rect 3750 -4062 3766 -4028
rect 3800 -4062 3816 -4028
rect 2836 -4130 2870 -4068
rect 4058 -3240 4836 -3040
rect 6984 2112 7018 2174
rect 5078 2072 5094 2106
rect 5128 2072 5144 2106
rect 5270 2072 5286 2106
rect 5320 2072 5336 2106
rect 5462 2072 5478 2106
rect 5512 2072 5528 2106
rect 5654 2072 5670 2106
rect 5704 2072 5720 2106
rect 5846 2072 5862 2106
rect 5896 2072 5912 2106
rect 6038 2072 6054 2106
rect 6088 2072 6104 2106
rect 6230 2072 6246 2106
rect 6280 2072 6296 2106
rect 6422 2072 6438 2106
rect 6472 2072 6488 2106
rect 6614 2072 6630 2106
rect 6664 2072 6680 2106
rect 6806 2072 6822 2106
rect 6856 2072 6872 2106
rect 4950 2022 4984 2038
rect 4950 1630 4984 1646
rect 5046 2022 5080 2038
rect 5046 1630 5080 1646
rect 5142 2022 5176 2038
rect 5142 1630 5176 1646
rect 5238 2022 5272 2038
rect 5238 1630 5272 1646
rect 5334 2022 5368 2038
rect 5334 1630 5368 1646
rect 5430 2022 5464 2038
rect 5430 1630 5464 1646
rect 5526 2022 5560 2038
rect 5526 1630 5560 1646
rect 5622 2022 5656 2038
rect 5622 1630 5656 1646
rect 5718 2022 5752 2038
rect 5718 1630 5752 1646
rect 5814 2022 5848 2038
rect 5814 1630 5848 1646
rect 5910 2022 5944 2038
rect 5910 1630 5944 1646
rect 6006 2022 6040 2038
rect 6006 1630 6040 1646
rect 6102 2022 6136 2038
rect 6102 1630 6136 1646
rect 6198 2022 6232 2038
rect 6198 1630 6232 1646
rect 6294 2022 6328 2038
rect 6294 1630 6328 1646
rect 6390 2022 6424 2038
rect 6390 1630 6424 1646
rect 6486 2022 6520 2038
rect 6486 1630 6520 1646
rect 6582 2022 6616 2038
rect 6582 1630 6616 1646
rect 6678 2022 6712 2038
rect 6678 1630 6712 1646
rect 6774 2022 6808 2038
rect 6774 1630 6808 1646
rect 6870 2022 6904 2038
rect 6870 1630 6904 1646
rect 4982 1562 4998 1596
rect 5032 1562 5048 1596
rect 5174 1562 5190 1596
rect 5224 1562 5240 1596
rect 5366 1562 5382 1596
rect 5416 1562 5432 1596
rect 5558 1562 5574 1596
rect 5608 1562 5624 1596
rect 5750 1562 5766 1596
rect 5800 1562 5816 1596
rect 5942 1562 5958 1596
rect 5992 1562 6008 1596
rect 6134 1562 6150 1596
rect 6184 1562 6200 1596
rect 6326 1562 6342 1596
rect 6376 1562 6392 1596
rect 6518 1562 6534 1596
rect 6568 1562 6584 1596
rect 6710 1562 6726 1596
rect 6760 1562 6776 1596
rect 4982 1454 4998 1488
rect 5032 1454 5048 1488
rect 5174 1454 5190 1488
rect 5224 1454 5240 1488
rect 5366 1454 5382 1488
rect 5416 1454 5432 1488
rect 5558 1454 5574 1488
rect 5608 1454 5624 1488
rect 5750 1454 5766 1488
rect 5800 1454 5816 1488
rect 5942 1454 5958 1488
rect 5992 1454 6008 1488
rect 6134 1454 6150 1488
rect 6184 1454 6200 1488
rect 6326 1454 6342 1488
rect 6376 1454 6392 1488
rect 6518 1454 6534 1488
rect 6568 1454 6584 1488
rect 6710 1454 6726 1488
rect 6760 1454 6776 1488
rect 4950 1404 4984 1420
rect 4950 1012 4984 1028
rect 5046 1404 5080 1420
rect 5046 1012 5080 1028
rect 5142 1404 5176 1420
rect 5142 1012 5176 1028
rect 5238 1404 5272 1420
rect 5238 1012 5272 1028
rect 5334 1404 5368 1420
rect 5334 1012 5368 1028
rect 5430 1404 5464 1420
rect 5430 1012 5464 1028
rect 5526 1404 5560 1420
rect 5526 1012 5560 1028
rect 5622 1404 5656 1420
rect 5622 1012 5656 1028
rect 5718 1404 5752 1420
rect 5718 1012 5752 1028
rect 5814 1404 5848 1420
rect 5814 1012 5848 1028
rect 5910 1404 5944 1420
rect 5910 1012 5944 1028
rect 6006 1404 6040 1420
rect 6006 1012 6040 1028
rect 6102 1404 6136 1420
rect 6102 1012 6136 1028
rect 6198 1404 6232 1420
rect 6198 1012 6232 1028
rect 6294 1404 6328 1420
rect 6294 1012 6328 1028
rect 6390 1404 6424 1420
rect 6390 1012 6424 1028
rect 6486 1404 6520 1420
rect 6486 1012 6520 1028
rect 6582 1404 6616 1420
rect 6582 1012 6616 1028
rect 6678 1404 6712 1420
rect 6678 1012 6712 1028
rect 6774 1404 6808 1420
rect 6774 1012 6808 1028
rect 6870 1404 6904 1420
rect 6870 1012 6904 1028
rect 5078 944 5094 978
rect 5128 944 5144 978
rect 5270 944 5286 978
rect 5320 944 5336 978
rect 5462 944 5478 978
rect 5512 944 5528 978
rect 5654 944 5670 978
rect 5704 944 5720 978
rect 5846 944 5862 978
rect 5896 944 5912 978
rect 6038 944 6054 978
rect 6088 944 6104 978
rect 6230 944 6246 978
rect 6280 944 6296 978
rect 6422 944 6438 978
rect 6472 944 6488 978
rect 6614 944 6630 978
rect 6664 944 6680 978
rect 6806 944 6822 978
rect 6856 944 6872 978
rect 5078 836 5094 870
rect 5128 836 5144 870
rect 5270 836 5286 870
rect 5320 836 5336 870
rect 5462 836 5478 870
rect 5512 836 5528 870
rect 5654 836 5670 870
rect 5704 836 5720 870
rect 5846 836 5862 870
rect 5896 836 5912 870
rect 6038 836 6054 870
rect 6088 836 6104 870
rect 6230 836 6246 870
rect 6280 836 6296 870
rect 6422 836 6438 870
rect 6472 836 6488 870
rect 6614 836 6630 870
rect 6664 836 6680 870
rect 6806 836 6822 870
rect 6856 836 6872 870
rect 4950 786 4984 802
rect 4950 394 4984 410
rect 5046 786 5080 802
rect 5046 394 5080 410
rect 5142 786 5176 802
rect 5142 394 5176 410
rect 5238 786 5272 802
rect 5238 394 5272 410
rect 5334 786 5368 802
rect 5334 394 5368 410
rect 5430 786 5464 802
rect 5430 394 5464 410
rect 5526 786 5560 802
rect 5526 394 5560 410
rect 5622 786 5656 802
rect 5622 394 5656 410
rect 5718 786 5752 802
rect 5718 394 5752 410
rect 5814 786 5848 802
rect 5814 394 5848 410
rect 5910 786 5944 802
rect 5910 394 5944 410
rect 6006 786 6040 802
rect 6006 394 6040 410
rect 6102 786 6136 802
rect 6102 394 6136 410
rect 6198 786 6232 802
rect 6198 394 6232 410
rect 6294 786 6328 802
rect 6294 394 6328 410
rect 6390 786 6424 802
rect 6390 394 6424 410
rect 6486 786 6520 802
rect 6486 394 6520 410
rect 6582 786 6616 802
rect 6582 394 6616 410
rect 6678 786 6712 802
rect 6678 394 6712 410
rect 6774 786 6808 802
rect 6774 394 6808 410
rect 6870 786 6904 802
rect 6870 394 6904 410
rect 4982 326 4998 360
rect 5032 326 5048 360
rect 5174 326 5190 360
rect 5224 326 5240 360
rect 5366 326 5382 360
rect 5416 326 5432 360
rect 5558 326 5574 360
rect 5608 326 5624 360
rect 5750 326 5766 360
rect 5800 326 5816 360
rect 5942 326 5958 360
rect 5992 326 6008 360
rect 6134 326 6150 360
rect 6184 326 6200 360
rect 6326 326 6342 360
rect 6376 326 6392 360
rect 6518 326 6534 360
rect 6568 326 6584 360
rect 6710 326 6726 360
rect 6760 326 6776 360
rect 4982 218 4998 252
rect 5032 218 5048 252
rect 5174 218 5190 252
rect 5224 218 5240 252
rect 5366 218 5382 252
rect 5416 218 5432 252
rect 5558 218 5574 252
rect 5608 218 5624 252
rect 5750 218 5766 252
rect 5800 218 5816 252
rect 5942 218 5958 252
rect 5992 218 6008 252
rect 6134 218 6150 252
rect 6184 218 6200 252
rect 6326 218 6342 252
rect 6376 218 6392 252
rect 6518 218 6534 252
rect 6568 218 6584 252
rect 6710 218 6726 252
rect 6760 218 6776 252
rect 4950 168 4984 184
rect 4950 -224 4984 -208
rect 5046 168 5080 184
rect 5046 -224 5080 -208
rect 5142 168 5176 184
rect 5142 -224 5176 -208
rect 5238 168 5272 184
rect 5238 -224 5272 -208
rect 5334 168 5368 184
rect 5334 -224 5368 -208
rect 5430 168 5464 184
rect 5430 -224 5464 -208
rect 5526 168 5560 184
rect 5526 -224 5560 -208
rect 5622 168 5656 184
rect 5622 -224 5656 -208
rect 5718 168 5752 184
rect 5718 -224 5752 -208
rect 5814 168 5848 184
rect 5814 -224 5848 -208
rect 5910 168 5944 184
rect 5910 -224 5944 -208
rect 6006 168 6040 184
rect 6006 -224 6040 -208
rect 6102 168 6136 184
rect 6102 -224 6136 -208
rect 6198 168 6232 184
rect 6198 -224 6232 -208
rect 6294 168 6328 184
rect 6294 -224 6328 -208
rect 6390 168 6424 184
rect 6390 -224 6424 -208
rect 6486 168 6520 184
rect 6486 -224 6520 -208
rect 6582 168 6616 184
rect 6582 -224 6616 -208
rect 6678 168 6712 184
rect 6678 -224 6712 -208
rect 6774 168 6808 184
rect 6774 -224 6808 -208
rect 6870 168 6904 184
rect 6870 -224 6904 -208
rect 5078 -292 5094 -258
rect 5128 -292 5144 -258
rect 5270 -292 5286 -258
rect 5320 -292 5336 -258
rect 5462 -292 5478 -258
rect 5512 -292 5528 -258
rect 5654 -292 5670 -258
rect 5704 -292 5720 -258
rect 5846 -292 5862 -258
rect 5896 -292 5912 -258
rect 6038 -292 6054 -258
rect 6088 -292 6104 -258
rect 6230 -292 6246 -258
rect 6280 -292 6296 -258
rect 6422 -292 6438 -258
rect 6472 -292 6488 -258
rect 6614 -292 6630 -258
rect 6664 -292 6680 -258
rect 6806 -292 6822 -258
rect 6856 -292 6872 -258
rect 5078 -400 5094 -366
rect 5128 -400 5144 -366
rect 5270 -400 5286 -366
rect 5320 -400 5336 -366
rect 5462 -400 5478 -366
rect 5512 -400 5528 -366
rect 5654 -400 5670 -366
rect 5704 -400 5720 -366
rect 5846 -400 5862 -366
rect 5896 -400 5912 -366
rect 6038 -400 6054 -366
rect 6088 -400 6104 -366
rect 6230 -400 6246 -366
rect 6280 -400 6296 -366
rect 6422 -400 6438 -366
rect 6472 -400 6488 -366
rect 6614 -400 6630 -366
rect 6664 -400 6680 -366
rect 6806 -400 6822 -366
rect 6856 -400 6872 -366
rect 4950 -450 4984 -434
rect 4950 -842 4984 -826
rect 5046 -450 5080 -434
rect 5046 -842 5080 -826
rect 5142 -450 5176 -434
rect 5142 -842 5176 -826
rect 5238 -450 5272 -434
rect 5238 -842 5272 -826
rect 5334 -450 5368 -434
rect 5334 -842 5368 -826
rect 5430 -450 5464 -434
rect 5430 -842 5464 -826
rect 5526 -450 5560 -434
rect 5526 -842 5560 -826
rect 5622 -450 5656 -434
rect 5622 -842 5656 -826
rect 5718 -450 5752 -434
rect 5718 -842 5752 -826
rect 5814 -450 5848 -434
rect 5814 -842 5848 -826
rect 5910 -450 5944 -434
rect 5910 -842 5944 -826
rect 6006 -450 6040 -434
rect 6006 -842 6040 -826
rect 6102 -450 6136 -434
rect 6102 -842 6136 -826
rect 6198 -450 6232 -434
rect 6198 -842 6232 -826
rect 6294 -450 6328 -434
rect 6294 -842 6328 -826
rect 6390 -450 6424 -434
rect 6390 -842 6424 -826
rect 6486 -450 6520 -434
rect 6486 -842 6520 -826
rect 6582 -450 6616 -434
rect 6582 -842 6616 -826
rect 6678 -450 6712 -434
rect 6678 -842 6712 -826
rect 6774 -450 6808 -434
rect 6774 -842 6808 -826
rect 6870 -450 6904 -434
rect 6870 -842 6904 -826
rect 4982 -910 4998 -876
rect 5032 -910 5048 -876
rect 5174 -910 5190 -876
rect 5224 -910 5240 -876
rect 5366 -910 5382 -876
rect 5416 -910 5432 -876
rect 5558 -910 5574 -876
rect 5608 -910 5624 -876
rect 5750 -910 5766 -876
rect 5800 -910 5816 -876
rect 5942 -910 5958 -876
rect 5992 -910 6008 -876
rect 6134 -910 6150 -876
rect 6184 -910 6200 -876
rect 6326 -910 6342 -876
rect 6376 -910 6392 -876
rect 6518 -910 6534 -876
rect 6568 -910 6584 -876
rect 6710 -910 6726 -876
rect 6760 -910 6776 -876
rect 4982 -1018 4998 -984
rect 5032 -1018 5048 -984
rect 5174 -1018 5190 -984
rect 5224 -1018 5240 -984
rect 5366 -1018 5382 -984
rect 5416 -1018 5432 -984
rect 5558 -1018 5574 -984
rect 5608 -1018 5624 -984
rect 5750 -1018 5766 -984
rect 5800 -1018 5816 -984
rect 5942 -1018 5958 -984
rect 5992 -1018 6008 -984
rect 6134 -1018 6150 -984
rect 6184 -1018 6200 -984
rect 6326 -1018 6342 -984
rect 6376 -1018 6392 -984
rect 6518 -1018 6534 -984
rect 6568 -1018 6584 -984
rect 6710 -1018 6726 -984
rect 6760 -1018 6776 -984
rect 4950 -1068 4984 -1052
rect 4950 -1460 4984 -1444
rect 5046 -1068 5080 -1052
rect 5046 -1460 5080 -1444
rect 5142 -1068 5176 -1052
rect 5142 -1460 5176 -1444
rect 5238 -1068 5272 -1052
rect 5238 -1460 5272 -1444
rect 5334 -1068 5368 -1052
rect 5334 -1460 5368 -1444
rect 5430 -1068 5464 -1052
rect 5430 -1460 5464 -1444
rect 5526 -1068 5560 -1052
rect 5526 -1460 5560 -1444
rect 5622 -1068 5656 -1052
rect 5622 -1460 5656 -1444
rect 5718 -1068 5752 -1052
rect 5718 -1460 5752 -1444
rect 5814 -1068 5848 -1052
rect 5814 -1460 5848 -1444
rect 5910 -1068 5944 -1052
rect 5910 -1460 5944 -1444
rect 6006 -1068 6040 -1052
rect 6006 -1460 6040 -1444
rect 6102 -1068 6136 -1052
rect 6102 -1460 6136 -1444
rect 6198 -1068 6232 -1052
rect 6198 -1460 6232 -1444
rect 6294 -1068 6328 -1052
rect 6294 -1460 6328 -1444
rect 6390 -1068 6424 -1052
rect 6390 -1460 6424 -1444
rect 6486 -1068 6520 -1052
rect 6486 -1460 6520 -1444
rect 6582 -1068 6616 -1052
rect 6582 -1460 6616 -1444
rect 6678 -1068 6712 -1052
rect 6678 -1460 6712 -1444
rect 6774 -1068 6808 -1052
rect 6774 -1460 6808 -1444
rect 6870 -1068 6904 -1052
rect 6870 -1460 6904 -1444
rect 5078 -1528 5094 -1494
rect 5128 -1528 5144 -1494
rect 5270 -1528 5286 -1494
rect 5320 -1528 5336 -1494
rect 5462 -1528 5478 -1494
rect 5512 -1528 5528 -1494
rect 5654 -1528 5670 -1494
rect 5704 -1528 5720 -1494
rect 5846 -1528 5862 -1494
rect 5896 -1528 5912 -1494
rect 6038 -1528 6054 -1494
rect 6088 -1528 6104 -1494
rect 6230 -1528 6246 -1494
rect 6280 -1528 6296 -1494
rect 6422 -1528 6438 -1494
rect 6472 -1528 6488 -1494
rect 6614 -1528 6630 -1494
rect 6664 -1528 6680 -1494
rect 6806 -1528 6822 -1494
rect 6856 -1528 6872 -1494
rect 5078 -1636 5094 -1602
rect 5128 -1636 5144 -1602
rect 5270 -1636 5286 -1602
rect 5320 -1636 5336 -1602
rect 5462 -1636 5478 -1602
rect 5512 -1636 5528 -1602
rect 5654 -1636 5670 -1602
rect 5704 -1636 5720 -1602
rect 5846 -1636 5862 -1602
rect 5896 -1636 5912 -1602
rect 6038 -1636 6054 -1602
rect 6088 -1636 6104 -1602
rect 6230 -1636 6246 -1602
rect 6280 -1636 6296 -1602
rect 6422 -1636 6438 -1602
rect 6472 -1636 6488 -1602
rect 6614 -1636 6630 -1602
rect 6664 -1636 6680 -1602
rect 6806 -1636 6822 -1602
rect 6856 -1636 6872 -1602
rect 4950 -1686 4984 -1670
rect 4950 -2078 4984 -2062
rect 5046 -1686 5080 -1670
rect 5046 -2078 5080 -2062
rect 5142 -1686 5176 -1670
rect 5142 -2078 5176 -2062
rect 5238 -1686 5272 -1670
rect 5238 -2078 5272 -2062
rect 5334 -1686 5368 -1670
rect 5334 -2078 5368 -2062
rect 5430 -1686 5464 -1670
rect 5430 -2078 5464 -2062
rect 5526 -1686 5560 -1670
rect 5526 -2078 5560 -2062
rect 5622 -1686 5656 -1670
rect 5622 -2078 5656 -2062
rect 5718 -1686 5752 -1670
rect 5718 -2078 5752 -2062
rect 5814 -1686 5848 -1670
rect 5814 -2078 5848 -2062
rect 5910 -1686 5944 -1670
rect 5910 -2078 5944 -2062
rect 6006 -1686 6040 -1670
rect 6006 -2078 6040 -2062
rect 6102 -1686 6136 -1670
rect 6102 -2078 6136 -2062
rect 6198 -1686 6232 -1670
rect 6198 -2078 6232 -2062
rect 6294 -1686 6328 -1670
rect 6294 -2078 6328 -2062
rect 6390 -1686 6424 -1670
rect 6390 -2078 6424 -2062
rect 6486 -1686 6520 -1670
rect 6486 -2078 6520 -2062
rect 6582 -1686 6616 -1670
rect 6582 -2078 6616 -2062
rect 6678 -1686 6712 -1670
rect 6678 -2078 6712 -2062
rect 6774 -1686 6808 -1670
rect 6774 -2078 6808 -2062
rect 6870 -1686 6904 -1670
rect 6870 -2078 6904 -2062
rect 4982 -2146 4998 -2112
rect 5032 -2146 5048 -2112
rect 5174 -2146 5190 -2112
rect 5224 -2146 5240 -2112
rect 5366 -2146 5382 -2112
rect 5416 -2146 5432 -2112
rect 5558 -2146 5574 -2112
rect 5608 -2146 5624 -2112
rect 5750 -2146 5766 -2112
rect 5800 -2146 5816 -2112
rect 5942 -2146 5958 -2112
rect 5992 -2146 6008 -2112
rect 6134 -2146 6150 -2112
rect 6184 -2146 6200 -2112
rect 6326 -2146 6342 -2112
rect 6376 -2146 6392 -2112
rect 6518 -2146 6534 -2112
rect 6568 -2146 6584 -2112
rect 6710 -2146 6726 -2112
rect 6760 -2146 6776 -2112
rect 4982 -2254 4998 -2220
rect 5032 -2254 5048 -2220
rect 5174 -2254 5190 -2220
rect 5224 -2254 5240 -2220
rect 5366 -2254 5382 -2220
rect 5416 -2254 5432 -2220
rect 5558 -2254 5574 -2220
rect 5608 -2254 5624 -2220
rect 5750 -2254 5766 -2220
rect 5800 -2254 5816 -2220
rect 5942 -2254 5958 -2220
rect 5992 -2254 6008 -2220
rect 6134 -2254 6150 -2220
rect 6184 -2254 6200 -2220
rect 6326 -2254 6342 -2220
rect 6376 -2254 6392 -2220
rect 6518 -2254 6534 -2220
rect 6568 -2254 6584 -2220
rect 6710 -2254 6726 -2220
rect 6760 -2254 6776 -2220
rect 4950 -2304 4984 -2288
rect 4950 -2696 4984 -2680
rect 5046 -2304 5080 -2288
rect 5046 -2696 5080 -2680
rect 5142 -2304 5176 -2288
rect 5142 -2696 5176 -2680
rect 5238 -2304 5272 -2288
rect 5238 -2696 5272 -2680
rect 5334 -2304 5368 -2288
rect 5334 -2696 5368 -2680
rect 5430 -2304 5464 -2288
rect 5430 -2696 5464 -2680
rect 5526 -2304 5560 -2288
rect 5526 -2696 5560 -2680
rect 5622 -2304 5656 -2288
rect 5622 -2696 5656 -2680
rect 5718 -2304 5752 -2288
rect 5718 -2696 5752 -2680
rect 5814 -2304 5848 -2288
rect 5814 -2696 5848 -2680
rect 5910 -2304 5944 -2288
rect 5910 -2696 5944 -2680
rect 6006 -2304 6040 -2288
rect 6006 -2696 6040 -2680
rect 6102 -2304 6136 -2288
rect 6102 -2696 6136 -2680
rect 6198 -2304 6232 -2288
rect 6198 -2696 6232 -2680
rect 6294 -2304 6328 -2288
rect 6294 -2696 6328 -2680
rect 6390 -2304 6424 -2288
rect 6390 -2696 6424 -2680
rect 6486 -2304 6520 -2288
rect 6486 -2696 6520 -2680
rect 6582 -2304 6616 -2288
rect 6582 -2696 6616 -2680
rect 6678 -2304 6712 -2288
rect 6678 -2696 6712 -2680
rect 6774 -2304 6808 -2288
rect 6774 -2696 6808 -2680
rect 6870 -2304 6904 -2288
rect 6870 -2696 6904 -2680
rect 5078 -2764 5094 -2730
rect 5128 -2764 5144 -2730
rect 5270 -2764 5286 -2730
rect 5320 -2764 5336 -2730
rect 5462 -2764 5478 -2730
rect 5512 -2764 5528 -2730
rect 5654 -2764 5670 -2730
rect 5704 -2764 5720 -2730
rect 5846 -2764 5862 -2730
rect 5896 -2764 5912 -2730
rect 6038 -2764 6054 -2730
rect 6088 -2764 6104 -2730
rect 6230 -2764 6246 -2730
rect 6280 -2764 6296 -2730
rect 6422 -2764 6438 -2730
rect 6472 -2764 6488 -2730
rect 6614 -2764 6630 -2730
rect 6664 -2764 6680 -2730
rect 6806 -2764 6822 -2730
rect 6856 -2764 6872 -2730
rect 5078 -2872 5094 -2838
rect 5128 -2872 5144 -2838
rect 5270 -2872 5286 -2838
rect 5320 -2872 5336 -2838
rect 5462 -2872 5478 -2838
rect 5512 -2872 5528 -2838
rect 5654 -2872 5670 -2838
rect 5704 -2872 5720 -2838
rect 5846 -2872 5862 -2838
rect 5896 -2872 5912 -2838
rect 6038 -2872 6054 -2838
rect 6088 -2872 6104 -2838
rect 6230 -2872 6246 -2838
rect 6280 -2872 6296 -2838
rect 6422 -2872 6438 -2838
rect 6472 -2872 6488 -2838
rect 6614 -2872 6630 -2838
rect 6664 -2872 6680 -2838
rect 6806 -2872 6822 -2838
rect 6856 -2872 6872 -2838
rect 4950 -2922 4984 -2906
rect 4950 -3314 4984 -3298
rect 5046 -2922 5080 -2906
rect 5046 -3314 5080 -3298
rect 5142 -2922 5176 -2906
rect 5142 -3314 5176 -3298
rect 5238 -2922 5272 -2906
rect 5238 -3314 5272 -3298
rect 5334 -2922 5368 -2906
rect 5334 -3314 5368 -3298
rect 5430 -2922 5464 -2906
rect 5430 -3314 5464 -3298
rect 5526 -2922 5560 -2906
rect 5526 -3314 5560 -3298
rect 5622 -2922 5656 -2906
rect 5622 -3314 5656 -3298
rect 5718 -2922 5752 -2906
rect 5718 -3314 5752 -3298
rect 5814 -2922 5848 -2906
rect 5814 -3314 5848 -3298
rect 5910 -2922 5944 -2906
rect 5910 -3314 5944 -3298
rect 6006 -2922 6040 -2906
rect 6006 -3314 6040 -3298
rect 6102 -2922 6136 -2906
rect 6102 -3314 6136 -3298
rect 6198 -2922 6232 -2906
rect 6198 -3314 6232 -3298
rect 6294 -2922 6328 -2906
rect 6294 -3314 6328 -3298
rect 6390 -2922 6424 -2906
rect 6390 -3314 6424 -3298
rect 6486 -2922 6520 -2906
rect 6486 -3314 6520 -3298
rect 6582 -2922 6616 -2906
rect 6582 -3314 6616 -3298
rect 6678 -2922 6712 -2906
rect 6678 -3314 6712 -3298
rect 6774 -2922 6808 -2906
rect 6774 -3314 6808 -3298
rect 6870 -2922 6904 -2906
rect 6870 -3314 6904 -3298
rect 4982 -3382 4998 -3348
rect 5032 -3382 5048 -3348
rect 5174 -3382 5190 -3348
rect 5224 -3382 5240 -3348
rect 5366 -3382 5382 -3348
rect 5416 -3382 5432 -3348
rect 5558 -3382 5574 -3348
rect 5608 -3382 5624 -3348
rect 5750 -3382 5766 -3348
rect 5800 -3382 5816 -3348
rect 5942 -3382 5958 -3348
rect 5992 -3382 6008 -3348
rect 6134 -3382 6150 -3348
rect 6184 -3382 6200 -3348
rect 6326 -3382 6342 -3348
rect 6376 -3382 6392 -3348
rect 6518 -3382 6534 -3348
rect 6568 -3382 6584 -3348
rect 6710 -3382 6726 -3348
rect 6760 -3382 6776 -3348
rect 4836 -3450 4870 -3388
rect 6984 -3450 7018 -3388
rect 4836 -3484 4932 -3450
rect 6922 -3484 7018 -3450
rect 4024 -4130 4058 -4068
rect 2836 -4164 2932 -4130
rect 3962 -4164 4058 -4130
rect -2560 -4326 -2260 -4164
rect -760 -4326 -460 -4164
rect 1040 -4326 1340 -4164
rect 2840 -4326 3140 -4164
rect -2564 -4360 -2468 -4326
rect -1108 -4360 -1012 -4326
rect -2564 -4422 -2530 -4360
rect -1046 -4422 -1012 -4360
rect -2404 -4462 -2388 -4428
rect -2220 -4462 -2204 -4428
rect -2146 -4462 -2130 -4428
rect -1962 -4462 -1946 -4428
rect -1888 -4462 -1872 -4428
rect -1704 -4462 -1688 -4428
rect -1630 -4462 -1614 -4428
rect -1446 -4462 -1430 -4428
rect -1372 -4462 -1356 -4428
rect -1188 -4462 -1172 -4428
rect -2450 -4512 -2416 -4496
rect -2450 -4904 -2416 -4888
rect -2192 -4512 -2158 -4496
rect -2192 -4904 -2158 -4888
rect -1934 -4512 -1900 -4496
rect -1934 -4904 -1900 -4888
rect -1676 -4512 -1642 -4496
rect -1676 -4904 -1642 -4888
rect -1418 -4512 -1384 -4496
rect -1418 -4904 -1384 -4888
rect -1160 -4512 -1126 -4496
rect -1160 -4904 -1126 -4888
rect -2404 -4972 -2388 -4938
rect -2220 -4972 -2204 -4938
rect -2146 -4972 -2130 -4938
rect -1962 -4972 -1946 -4938
rect -1888 -4972 -1872 -4938
rect -1704 -4972 -1688 -4938
rect -1630 -4972 -1614 -4938
rect -1446 -4972 -1430 -4938
rect -1372 -4972 -1356 -4938
rect -1188 -4972 -1172 -4938
rect -2404 -5080 -2388 -5046
rect -2220 -5080 -2204 -5046
rect -2146 -5080 -2130 -5046
rect -1962 -5080 -1946 -5046
rect -1888 -5080 -1872 -5046
rect -1704 -5080 -1688 -5046
rect -1630 -5080 -1614 -5046
rect -1446 -5080 -1430 -5046
rect -1372 -5080 -1356 -5046
rect -1188 -5080 -1172 -5046
rect -2450 -5130 -2416 -5114
rect -2450 -5522 -2416 -5506
rect -2192 -5130 -2158 -5114
rect -2192 -5522 -2158 -5506
rect -1934 -5130 -1900 -5114
rect -1934 -5522 -1900 -5506
rect -1676 -5130 -1642 -5114
rect -1676 -5522 -1642 -5506
rect -1418 -5130 -1384 -5114
rect -1418 -5522 -1384 -5506
rect -1160 -5130 -1126 -5114
rect -1160 -5522 -1126 -5506
rect -2404 -5590 -2388 -5556
rect -2220 -5590 -2204 -5556
rect -2146 -5590 -2130 -5556
rect -1962 -5590 -1946 -5556
rect -1888 -5590 -1872 -5556
rect -1704 -5590 -1688 -5556
rect -1630 -5590 -1614 -5556
rect -1446 -5590 -1430 -5556
rect -1372 -5590 -1356 -5556
rect -1188 -5590 -1172 -5556
rect -2404 -5698 -2388 -5664
rect -2220 -5698 -2204 -5664
rect -2146 -5698 -2130 -5664
rect -1962 -5698 -1946 -5664
rect -1888 -5698 -1872 -5664
rect -1704 -5698 -1688 -5664
rect -1630 -5698 -1614 -5664
rect -1446 -5698 -1430 -5664
rect -1372 -5698 -1356 -5664
rect -1188 -5698 -1172 -5664
rect -2450 -5748 -2416 -5732
rect -2450 -6140 -2416 -6124
rect -2192 -5748 -2158 -5732
rect -2192 -6140 -2158 -6124
rect -1934 -5748 -1900 -5732
rect -1934 -6140 -1900 -6124
rect -1676 -5748 -1642 -5732
rect -1676 -6140 -1642 -6124
rect -1418 -5748 -1384 -5732
rect -1418 -6140 -1384 -6124
rect -1160 -5748 -1126 -5732
rect -1160 -6140 -1126 -6124
rect -2404 -6208 -2388 -6174
rect -2220 -6208 -2204 -6174
rect -2146 -6208 -2130 -6174
rect -1962 -6208 -1946 -6174
rect -1888 -6208 -1872 -6174
rect -1704 -6208 -1688 -6174
rect -1630 -6208 -1614 -6174
rect -1446 -6208 -1430 -6174
rect -1372 -6208 -1356 -6174
rect -1188 -6208 -1172 -6174
rect -2404 -6316 -2388 -6282
rect -2220 -6316 -2204 -6282
rect -2146 -6316 -2130 -6282
rect -1962 -6316 -1946 -6282
rect -1888 -6316 -1872 -6282
rect -1704 -6316 -1688 -6282
rect -1630 -6316 -1614 -6282
rect -1446 -6316 -1430 -6282
rect -1372 -6316 -1356 -6282
rect -1188 -6316 -1172 -6282
rect -2450 -6366 -2416 -6350
rect -2450 -6758 -2416 -6742
rect -2192 -6366 -2158 -6350
rect -2192 -6758 -2158 -6742
rect -1934 -6366 -1900 -6350
rect -1934 -6758 -1900 -6742
rect -1676 -6366 -1642 -6350
rect -1676 -6758 -1642 -6742
rect -1418 -6366 -1384 -6350
rect -1418 -6758 -1384 -6742
rect -1160 -6366 -1126 -6350
rect -1160 -6758 -1126 -6742
rect -2404 -6826 -2388 -6792
rect -2220 -6826 -2204 -6792
rect -2146 -6826 -2130 -6792
rect -1962 -6826 -1946 -6792
rect -1888 -6826 -1872 -6792
rect -1704 -6826 -1688 -6792
rect -1630 -6826 -1614 -6792
rect -1446 -6826 -1430 -6792
rect -1372 -6826 -1356 -6792
rect -1188 -6826 -1172 -6792
rect -2404 -6934 -2388 -6900
rect -2220 -6934 -2204 -6900
rect -2146 -6934 -2130 -6900
rect -1962 -6934 -1946 -6900
rect -1888 -6934 -1872 -6900
rect -1704 -6934 -1688 -6900
rect -1630 -6934 -1614 -6900
rect -1446 -6934 -1430 -6900
rect -1372 -6934 -1356 -6900
rect -1188 -6934 -1172 -6900
rect -2450 -6984 -2416 -6968
rect -2450 -7376 -2416 -7360
rect -2192 -6984 -2158 -6968
rect -2192 -7376 -2158 -7360
rect -1934 -6984 -1900 -6968
rect -1934 -7376 -1900 -7360
rect -1676 -6984 -1642 -6968
rect -1676 -7376 -1642 -7360
rect -1418 -6984 -1384 -6968
rect -1418 -7376 -1384 -7360
rect -1160 -6984 -1126 -6968
rect -1160 -7376 -1126 -7360
rect -2404 -7444 -2388 -7410
rect -2220 -7444 -2204 -7410
rect -2146 -7444 -2130 -7410
rect -1962 -7444 -1946 -7410
rect -1888 -7444 -1872 -7410
rect -1704 -7444 -1688 -7410
rect -1630 -7444 -1614 -7410
rect -1446 -7444 -1430 -7410
rect -1372 -7444 -1356 -7410
rect -1188 -7444 -1172 -7410
rect -2404 -7552 -2388 -7518
rect -2220 -7552 -2204 -7518
rect -2146 -7552 -2130 -7518
rect -1962 -7552 -1946 -7518
rect -1888 -7552 -1872 -7518
rect -1704 -7552 -1688 -7518
rect -1630 -7552 -1614 -7518
rect -1446 -7552 -1430 -7518
rect -1372 -7552 -1356 -7518
rect -1188 -7552 -1172 -7518
rect -2450 -7602 -2416 -7586
rect -2450 -7994 -2416 -7978
rect -2192 -7602 -2158 -7586
rect -2192 -7994 -2158 -7978
rect -1934 -7602 -1900 -7586
rect -1934 -7994 -1900 -7978
rect -1676 -7602 -1642 -7586
rect -1676 -7994 -1642 -7978
rect -1418 -7602 -1384 -7586
rect -1418 -7994 -1384 -7978
rect -1160 -7602 -1126 -7586
rect -1160 -7994 -1126 -7978
rect -2404 -8062 -2388 -8028
rect -2220 -8062 -2204 -8028
rect -2146 -8062 -2130 -8028
rect -1962 -8062 -1946 -8028
rect -1888 -8062 -1872 -8028
rect -1704 -8062 -1688 -8028
rect -1630 -8062 -1614 -8028
rect -1446 -8062 -1430 -8028
rect -1372 -8062 -1356 -8028
rect -1188 -8062 -1172 -8028
rect -2564 -8130 -2530 -8068
rect -764 -4360 -668 -4326
rect 692 -4360 788 -4326
rect -764 -4422 -730 -4360
rect -1012 -8068 -980 -7960
rect -1046 -8130 -980 -8068
rect -2564 -8164 -2468 -8130
rect -1108 -8160 -980 -8130
rect -800 -8068 -764 -7960
rect 754 -4422 788 -4360
rect -604 -4462 -588 -4428
rect -420 -4462 -404 -4428
rect -346 -4462 -330 -4428
rect -162 -4462 -146 -4428
rect -88 -4462 -72 -4428
rect 96 -4462 112 -4428
rect 170 -4462 186 -4428
rect 354 -4462 370 -4428
rect 428 -4462 444 -4428
rect 612 -4462 628 -4428
rect -650 -4512 -616 -4496
rect -650 -4904 -616 -4888
rect -392 -4512 -358 -4496
rect -392 -4904 -358 -4888
rect -134 -4512 -100 -4496
rect -134 -4904 -100 -4888
rect 124 -4512 158 -4496
rect 124 -4904 158 -4888
rect 382 -4512 416 -4496
rect 382 -4904 416 -4888
rect 640 -4512 674 -4496
rect 640 -4904 674 -4888
rect -604 -4972 -588 -4938
rect -420 -4972 -404 -4938
rect -346 -4972 -330 -4938
rect -162 -4972 -146 -4938
rect -88 -4972 -72 -4938
rect 96 -4972 112 -4938
rect 170 -4972 186 -4938
rect 354 -4972 370 -4938
rect 428 -4972 444 -4938
rect 612 -4972 628 -4938
rect -604 -5080 -588 -5046
rect -420 -5080 -404 -5046
rect -346 -5080 -330 -5046
rect -162 -5080 -146 -5046
rect -88 -5080 -72 -5046
rect 96 -5080 112 -5046
rect 170 -5080 186 -5046
rect 354 -5080 370 -5046
rect 428 -5080 444 -5046
rect 612 -5080 628 -5046
rect -650 -5130 -616 -5114
rect -650 -5522 -616 -5506
rect -392 -5130 -358 -5114
rect -392 -5522 -358 -5506
rect -134 -5130 -100 -5114
rect -134 -5522 -100 -5506
rect 124 -5130 158 -5114
rect 124 -5522 158 -5506
rect 382 -5130 416 -5114
rect 382 -5522 416 -5506
rect 640 -5130 674 -5114
rect 640 -5522 674 -5506
rect -604 -5590 -588 -5556
rect -420 -5590 -404 -5556
rect -346 -5590 -330 -5556
rect -162 -5590 -146 -5556
rect -88 -5590 -72 -5556
rect 96 -5590 112 -5556
rect 170 -5590 186 -5556
rect 354 -5590 370 -5556
rect 428 -5590 444 -5556
rect 612 -5590 628 -5556
rect -604 -5698 -588 -5664
rect -420 -5698 -404 -5664
rect -346 -5698 -330 -5664
rect -162 -5698 -146 -5664
rect -88 -5698 -72 -5664
rect 96 -5698 112 -5664
rect 170 -5698 186 -5664
rect 354 -5698 370 -5664
rect 428 -5698 444 -5664
rect 612 -5698 628 -5664
rect -650 -5748 -616 -5732
rect -650 -6140 -616 -6124
rect -392 -5748 -358 -5732
rect -392 -6140 -358 -6124
rect -134 -5748 -100 -5732
rect -134 -6140 -100 -6124
rect 124 -5748 158 -5732
rect 124 -6140 158 -6124
rect 382 -5748 416 -5732
rect 382 -6140 416 -6124
rect 640 -5748 674 -5732
rect 640 -6140 674 -6124
rect -604 -6208 -588 -6174
rect -420 -6208 -404 -6174
rect -346 -6208 -330 -6174
rect -162 -6208 -146 -6174
rect -88 -6208 -72 -6174
rect 96 -6208 112 -6174
rect 170 -6208 186 -6174
rect 354 -6208 370 -6174
rect 428 -6208 444 -6174
rect 612 -6208 628 -6174
rect -604 -6316 -588 -6282
rect -420 -6316 -404 -6282
rect -346 -6316 -330 -6282
rect -162 -6316 -146 -6282
rect -88 -6316 -72 -6282
rect 96 -6316 112 -6282
rect 170 -6316 186 -6282
rect 354 -6316 370 -6282
rect 428 -6316 444 -6282
rect 612 -6316 628 -6282
rect -650 -6366 -616 -6350
rect -650 -6758 -616 -6742
rect -392 -6366 -358 -6350
rect -392 -6758 -358 -6742
rect -134 -6366 -100 -6350
rect -134 -6758 -100 -6742
rect 124 -6366 158 -6350
rect 124 -6758 158 -6742
rect 382 -6366 416 -6350
rect 382 -6758 416 -6742
rect 640 -6366 674 -6350
rect 640 -6758 674 -6742
rect -604 -6826 -588 -6792
rect -420 -6826 -404 -6792
rect -346 -6826 -330 -6792
rect -162 -6826 -146 -6792
rect -88 -6826 -72 -6792
rect 96 -6826 112 -6792
rect 170 -6826 186 -6792
rect 354 -6826 370 -6792
rect 428 -6826 444 -6792
rect 612 -6826 628 -6792
rect -604 -6934 -588 -6900
rect -420 -6934 -404 -6900
rect -346 -6934 -330 -6900
rect -162 -6934 -146 -6900
rect -88 -6934 -72 -6900
rect 96 -6934 112 -6900
rect 170 -6934 186 -6900
rect 354 -6934 370 -6900
rect 428 -6934 444 -6900
rect 612 -6934 628 -6900
rect -650 -6984 -616 -6968
rect -650 -7376 -616 -7360
rect -392 -6984 -358 -6968
rect -392 -7376 -358 -7360
rect -134 -6984 -100 -6968
rect -134 -7376 -100 -7360
rect 124 -6984 158 -6968
rect 124 -7376 158 -7360
rect 382 -6984 416 -6968
rect 382 -7376 416 -7360
rect 640 -6984 674 -6968
rect 640 -7376 674 -7360
rect -604 -7444 -588 -7410
rect -420 -7444 -404 -7410
rect -346 -7444 -330 -7410
rect -162 -7444 -146 -7410
rect -88 -7444 -72 -7410
rect 96 -7444 112 -7410
rect 170 -7444 186 -7410
rect 354 -7444 370 -7410
rect 428 -7444 444 -7410
rect 612 -7444 628 -7410
rect -604 -7552 -588 -7518
rect -420 -7552 -404 -7518
rect -346 -7552 -330 -7518
rect -162 -7552 -146 -7518
rect -88 -7552 -72 -7518
rect 96 -7552 112 -7518
rect 170 -7552 186 -7518
rect 354 -7552 370 -7518
rect 428 -7552 444 -7518
rect 612 -7552 628 -7518
rect -650 -7602 -616 -7586
rect -650 -7994 -616 -7978
rect -392 -7602 -358 -7586
rect -392 -7994 -358 -7978
rect -134 -7602 -100 -7586
rect -134 -7994 -100 -7978
rect 124 -7602 158 -7586
rect 124 -7994 158 -7978
rect 382 -7602 416 -7586
rect 382 -7994 416 -7978
rect 640 -7602 674 -7586
rect 640 -7994 674 -7978
rect -604 -8062 -588 -8028
rect -420 -8062 -404 -8028
rect -346 -8062 -330 -8028
rect -162 -8062 -146 -8028
rect -88 -8062 -72 -8028
rect 96 -8062 112 -8028
rect 170 -8062 186 -8028
rect 354 -8062 370 -8028
rect 428 -8062 444 -8028
rect 612 -8062 628 -8028
rect -800 -8130 -730 -8068
rect 1036 -4360 1132 -4326
rect 2492 -4360 2588 -4326
rect 1036 -4422 1070 -4360
rect 788 -8068 1036 -7960
rect 2554 -4422 2588 -4360
rect 1196 -4462 1212 -4428
rect 1380 -4462 1396 -4428
rect 1454 -4462 1470 -4428
rect 1638 -4462 1654 -4428
rect 1712 -4462 1728 -4428
rect 1896 -4462 1912 -4428
rect 1970 -4462 1986 -4428
rect 2154 -4462 2170 -4428
rect 2228 -4462 2244 -4428
rect 2412 -4462 2428 -4428
rect 1150 -4512 1184 -4496
rect 1150 -4904 1184 -4888
rect 1408 -4512 1442 -4496
rect 1408 -4904 1442 -4888
rect 1666 -4512 1700 -4496
rect 1666 -4904 1700 -4888
rect 1924 -4512 1958 -4496
rect 1924 -4904 1958 -4888
rect 2182 -4512 2216 -4496
rect 2182 -4904 2216 -4888
rect 2440 -4512 2474 -4496
rect 2440 -4904 2474 -4888
rect 1196 -4972 1212 -4938
rect 1380 -4972 1396 -4938
rect 1454 -4972 1470 -4938
rect 1638 -4972 1654 -4938
rect 1712 -4972 1728 -4938
rect 1896 -4972 1912 -4938
rect 1970 -4972 1986 -4938
rect 2154 -4972 2170 -4938
rect 2228 -4972 2244 -4938
rect 2412 -4972 2428 -4938
rect 1196 -5080 1212 -5046
rect 1380 -5080 1396 -5046
rect 1454 -5080 1470 -5046
rect 1638 -5080 1654 -5046
rect 1712 -5080 1728 -5046
rect 1896 -5080 1912 -5046
rect 1970 -5080 1986 -5046
rect 2154 -5080 2170 -5046
rect 2228 -5080 2244 -5046
rect 2412 -5080 2428 -5046
rect 1150 -5130 1184 -5114
rect 1150 -5522 1184 -5506
rect 1408 -5130 1442 -5114
rect 1408 -5522 1442 -5506
rect 1666 -5130 1700 -5114
rect 1666 -5522 1700 -5506
rect 1924 -5130 1958 -5114
rect 1924 -5522 1958 -5506
rect 2182 -5130 2216 -5114
rect 2182 -5522 2216 -5506
rect 2440 -5130 2474 -5114
rect 2440 -5522 2474 -5506
rect 1196 -5590 1212 -5556
rect 1380 -5590 1396 -5556
rect 1454 -5590 1470 -5556
rect 1638 -5590 1654 -5556
rect 1712 -5590 1728 -5556
rect 1896 -5590 1912 -5556
rect 1970 -5590 1986 -5556
rect 2154 -5590 2170 -5556
rect 2228 -5590 2244 -5556
rect 2412 -5590 2428 -5556
rect 1196 -5698 1212 -5664
rect 1380 -5698 1396 -5664
rect 1454 -5698 1470 -5664
rect 1638 -5698 1654 -5664
rect 1712 -5698 1728 -5664
rect 1896 -5698 1912 -5664
rect 1970 -5698 1986 -5664
rect 2154 -5698 2170 -5664
rect 2228 -5698 2244 -5664
rect 2412 -5698 2428 -5664
rect 1150 -5748 1184 -5732
rect 1150 -6140 1184 -6124
rect 1408 -5748 1442 -5732
rect 1408 -6140 1442 -6124
rect 1666 -5748 1700 -5732
rect 1666 -6140 1700 -6124
rect 1924 -5748 1958 -5732
rect 1924 -6140 1958 -6124
rect 2182 -5748 2216 -5732
rect 2182 -6140 2216 -6124
rect 2440 -5748 2474 -5732
rect 2440 -6140 2474 -6124
rect 1196 -6208 1212 -6174
rect 1380 -6208 1396 -6174
rect 1454 -6208 1470 -6174
rect 1638 -6208 1654 -6174
rect 1712 -6208 1728 -6174
rect 1896 -6208 1912 -6174
rect 1970 -6208 1986 -6174
rect 2154 -6208 2170 -6174
rect 2228 -6208 2244 -6174
rect 2412 -6208 2428 -6174
rect 1196 -6316 1212 -6282
rect 1380 -6316 1396 -6282
rect 1454 -6316 1470 -6282
rect 1638 -6316 1654 -6282
rect 1712 -6316 1728 -6282
rect 1896 -6316 1912 -6282
rect 1970 -6316 1986 -6282
rect 2154 -6316 2170 -6282
rect 2228 -6316 2244 -6282
rect 2412 -6316 2428 -6282
rect 1150 -6366 1184 -6350
rect 1150 -6758 1184 -6742
rect 1408 -6366 1442 -6350
rect 1408 -6758 1442 -6742
rect 1666 -6366 1700 -6350
rect 1666 -6758 1700 -6742
rect 1924 -6366 1958 -6350
rect 1924 -6758 1958 -6742
rect 2182 -6366 2216 -6350
rect 2182 -6758 2216 -6742
rect 2440 -6366 2474 -6350
rect 2440 -6758 2474 -6742
rect 1196 -6826 1212 -6792
rect 1380 -6826 1396 -6792
rect 1454 -6826 1470 -6792
rect 1638 -6826 1654 -6792
rect 1712 -6826 1728 -6792
rect 1896 -6826 1912 -6792
rect 1970 -6826 1986 -6792
rect 2154 -6826 2170 -6792
rect 2228 -6826 2244 -6792
rect 2412 -6826 2428 -6792
rect 1196 -6934 1212 -6900
rect 1380 -6934 1396 -6900
rect 1454 -6934 1470 -6900
rect 1638 -6934 1654 -6900
rect 1712 -6934 1728 -6900
rect 1896 -6934 1912 -6900
rect 1970 -6934 1986 -6900
rect 2154 -6934 2170 -6900
rect 2228 -6934 2244 -6900
rect 2412 -6934 2428 -6900
rect 1150 -6984 1184 -6968
rect 1150 -7376 1184 -7360
rect 1408 -6984 1442 -6968
rect 1408 -7376 1442 -7360
rect 1666 -6984 1700 -6968
rect 1666 -7376 1700 -7360
rect 1924 -6984 1958 -6968
rect 1924 -7376 1958 -7360
rect 2182 -6984 2216 -6968
rect 2182 -7376 2216 -7360
rect 2440 -6984 2474 -6968
rect 2440 -7376 2474 -7360
rect 1196 -7444 1212 -7410
rect 1380 -7444 1396 -7410
rect 1454 -7444 1470 -7410
rect 1638 -7444 1654 -7410
rect 1712 -7444 1728 -7410
rect 1896 -7444 1912 -7410
rect 1970 -7444 1986 -7410
rect 2154 -7444 2170 -7410
rect 2228 -7444 2244 -7410
rect 2412 -7444 2428 -7410
rect 1196 -7552 1212 -7518
rect 1380 -7552 1396 -7518
rect 1454 -7552 1470 -7518
rect 1638 -7552 1654 -7518
rect 1712 -7552 1728 -7518
rect 1896 -7552 1912 -7518
rect 1970 -7552 1986 -7518
rect 2154 -7552 2170 -7518
rect 2228 -7552 2244 -7518
rect 2412 -7552 2428 -7518
rect 1150 -7602 1184 -7586
rect 1150 -7994 1184 -7978
rect 1408 -7602 1442 -7586
rect 1408 -7994 1442 -7978
rect 1666 -7602 1700 -7586
rect 1666 -7994 1700 -7978
rect 1924 -7602 1958 -7586
rect 1924 -7994 1958 -7978
rect 2182 -7602 2216 -7586
rect 2182 -7994 2216 -7978
rect 2440 -7602 2474 -7586
rect 2440 -7994 2474 -7978
rect 1196 -8062 1212 -8028
rect 1380 -8062 1396 -8028
rect 1454 -8062 1470 -8028
rect 1638 -8062 1654 -8028
rect 1712 -8062 1728 -8028
rect 1896 -8062 1912 -8028
rect 1970 -8062 1986 -8028
rect 2154 -8062 2170 -8028
rect 2228 -8062 2244 -8028
rect 2412 -8062 2428 -8028
rect 754 -8130 1070 -8068
rect 2836 -4360 2932 -4326
rect 4292 -4360 4388 -4326
rect 2836 -4422 2870 -4360
rect 2588 -8068 2836 -7960
rect 4354 -4422 4388 -4360
rect 2996 -4462 3012 -4428
rect 3180 -4462 3196 -4428
rect 3254 -4462 3270 -4428
rect 3438 -4462 3454 -4428
rect 3512 -4462 3528 -4428
rect 3696 -4462 3712 -4428
rect 3770 -4462 3786 -4428
rect 3954 -4462 3970 -4428
rect 4028 -4462 4044 -4428
rect 4212 -4462 4228 -4428
rect 2950 -4512 2984 -4496
rect 2950 -4904 2984 -4888
rect 3208 -4512 3242 -4496
rect 3208 -4904 3242 -4888
rect 3466 -4512 3500 -4496
rect 3466 -4904 3500 -4888
rect 3724 -4512 3758 -4496
rect 3724 -4904 3758 -4888
rect 3982 -4512 4016 -4496
rect 3982 -4904 4016 -4888
rect 4240 -4512 4274 -4496
rect 4240 -4904 4274 -4888
rect 2996 -4972 3012 -4938
rect 3180 -4972 3196 -4938
rect 3254 -4972 3270 -4938
rect 3438 -4972 3454 -4938
rect 3512 -4972 3528 -4938
rect 3696 -4972 3712 -4938
rect 3770 -4972 3786 -4938
rect 3954 -4972 3970 -4938
rect 4028 -4972 4044 -4938
rect 4212 -4972 4228 -4938
rect 2996 -5080 3012 -5046
rect 3180 -5080 3196 -5046
rect 3254 -5080 3270 -5046
rect 3438 -5080 3454 -5046
rect 3512 -5080 3528 -5046
rect 3696 -5080 3712 -5046
rect 3770 -5080 3786 -5046
rect 3954 -5080 3970 -5046
rect 4028 -5080 4044 -5046
rect 4212 -5080 4228 -5046
rect 2950 -5130 2984 -5114
rect 2950 -5522 2984 -5506
rect 3208 -5130 3242 -5114
rect 3208 -5522 3242 -5506
rect 3466 -5130 3500 -5114
rect 3466 -5522 3500 -5506
rect 3724 -5130 3758 -5114
rect 3724 -5522 3758 -5506
rect 3982 -5130 4016 -5114
rect 3982 -5522 4016 -5506
rect 4240 -5130 4274 -5114
rect 4240 -5522 4274 -5506
rect 2996 -5590 3012 -5556
rect 3180 -5590 3196 -5556
rect 3254 -5590 3270 -5556
rect 3438 -5590 3454 -5556
rect 3512 -5590 3528 -5556
rect 3696 -5590 3712 -5556
rect 3770 -5590 3786 -5556
rect 3954 -5590 3970 -5556
rect 4028 -5590 4044 -5556
rect 4212 -5590 4228 -5556
rect 2996 -5698 3012 -5664
rect 3180 -5698 3196 -5664
rect 3254 -5698 3270 -5664
rect 3438 -5698 3454 -5664
rect 3512 -5698 3528 -5664
rect 3696 -5698 3712 -5664
rect 3770 -5698 3786 -5664
rect 3954 -5698 3970 -5664
rect 4028 -5698 4044 -5664
rect 4212 -5698 4228 -5664
rect 2950 -5748 2984 -5732
rect 2950 -6140 2984 -6124
rect 3208 -5748 3242 -5732
rect 3208 -6140 3242 -6124
rect 3466 -5748 3500 -5732
rect 3466 -6140 3500 -6124
rect 3724 -5748 3758 -5732
rect 3724 -6140 3758 -6124
rect 3982 -5748 4016 -5732
rect 3982 -6140 4016 -6124
rect 4240 -5748 4274 -5732
rect 4240 -6140 4274 -6124
rect 2996 -6208 3012 -6174
rect 3180 -6208 3196 -6174
rect 3254 -6208 3270 -6174
rect 3438 -6208 3454 -6174
rect 3512 -6208 3528 -6174
rect 3696 -6208 3712 -6174
rect 3770 -6208 3786 -6174
rect 3954 -6208 3970 -6174
rect 4028 -6208 4044 -6174
rect 4212 -6208 4228 -6174
rect 2996 -6316 3012 -6282
rect 3180 -6316 3196 -6282
rect 3254 -6316 3270 -6282
rect 3438 -6316 3454 -6282
rect 3512 -6316 3528 -6282
rect 3696 -6316 3712 -6282
rect 3770 -6316 3786 -6282
rect 3954 -6316 3970 -6282
rect 4028 -6316 4044 -6282
rect 4212 -6316 4228 -6282
rect 2950 -6366 2984 -6350
rect 2950 -6758 2984 -6742
rect 3208 -6366 3242 -6350
rect 3208 -6758 3242 -6742
rect 3466 -6366 3500 -6350
rect 3466 -6758 3500 -6742
rect 3724 -6366 3758 -6350
rect 3724 -6758 3758 -6742
rect 3982 -6366 4016 -6350
rect 3982 -6758 4016 -6742
rect 4240 -6366 4274 -6350
rect 4240 -6758 4274 -6742
rect 2996 -6826 3012 -6792
rect 3180 -6826 3196 -6792
rect 3254 -6826 3270 -6792
rect 3438 -6826 3454 -6792
rect 3512 -6826 3528 -6792
rect 3696 -6826 3712 -6792
rect 3770 -6826 3786 -6792
rect 3954 -6826 3970 -6792
rect 4028 -6826 4044 -6792
rect 4212 -6826 4228 -6792
rect 2996 -6934 3012 -6900
rect 3180 -6934 3196 -6900
rect 3254 -6934 3270 -6900
rect 3438 -6934 3454 -6900
rect 3512 -6934 3528 -6900
rect 3696 -6934 3712 -6900
rect 3770 -6934 3786 -6900
rect 3954 -6934 3970 -6900
rect 4028 -6934 4044 -6900
rect 4212 -6934 4228 -6900
rect 2950 -6984 2984 -6968
rect 2950 -7376 2984 -7360
rect 3208 -6984 3242 -6968
rect 3208 -7376 3242 -7360
rect 3466 -6984 3500 -6968
rect 3466 -7376 3500 -7360
rect 3724 -6984 3758 -6968
rect 3724 -7376 3758 -7360
rect 3982 -6984 4016 -6968
rect 3982 -7376 4016 -7360
rect 4240 -6984 4274 -6968
rect 4240 -7376 4274 -7360
rect 2996 -7444 3012 -7410
rect 3180 -7444 3196 -7410
rect 3254 -7444 3270 -7410
rect 3438 -7444 3454 -7410
rect 3512 -7444 3528 -7410
rect 3696 -7444 3712 -7410
rect 3770 -7444 3786 -7410
rect 3954 -7444 3970 -7410
rect 4028 -7444 4044 -7410
rect 4212 -7444 4228 -7410
rect 2996 -7552 3012 -7518
rect 3180 -7552 3196 -7518
rect 3254 -7552 3270 -7518
rect 3438 -7552 3454 -7518
rect 3512 -7552 3528 -7518
rect 3696 -7552 3712 -7518
rect 3770 -7552 3786 -7518
rect 3954 -7552 3970 -7518
rect 4028 -7552 4044 -7518
rect 4212 -7552 4228 -7518
rect 2950 -7602 2984 -7586
rect 2950 -7994 2984 -7978
rect 3208 -7602 3242 -7586
rect 3208 -7994 3242 -7978
rect 3466 -7602 3500 -7586
rect 3466 -7994 3500 -7978
rect 3724 -7602 3758 -7586
rect 3724 -7994 3758 -7978
rect 3982 -7602 4016 -7586
rect 3982 -7994 4016 -7978
rect 4240 -7602 4274 -7586
rect 4240 -7994 4274 -7978
rect 2996 -8062 3012 -8028
rect 3180 -8062 3196 -8028
rect 3254 -8062 3270 -8028
rect 3438 -8062 3454 -8028
rect 3512 -8062 3528 -8028
rect 3696 -8062 3712 -8028
rect 3770 -8062 3786 -8028
rect 3954 -8062 3970 -8028
rect 4028 -8062 4044 -8028
rect 4212 -8062 4228 -8028
rect 2554 -8130 2870 -8068
rect 4354 -8130 4388 -8068
rect -800 -8160 -668 -8130
rect -1108 -8164 -1012 -8160
rect -764 -8164 -668 -8160
rect 692 -8160 1132 -8130
rect 692 -8164 788 -8160
rect 1036 -8164 1132 -8160
rect 2492 -8160 2932 -8130
rect 2492 -8164 2588 -8160
rect 2836 -8164 2932 -8160
rect 4292 -8164 4388 -8130
rect -5460 -9416 -5444 -8610
rect -4636 -9416 -4620 -8610
<< viali >>
rect 3420 2380 3600 2580
rect -58 1695 192 2092
rect 320 1695 570 2092
rect 698 1695 948 2092
rect 1076 1695 1326 2092
rect 1454 1695 1704 2092
rect 1832 1695 2082 2092
rect -58 464 192 861
rect 320 464 570 861
rect 698 464 948 861
rect 1076 464 1326 861
rect 1454 464 1704 861
rect 1832 464 2082 861
rect 2498 2102 2532 2136
rect 2690 2102 2724 2136
rect 2882 2102 2916 2136
rect 3074 2102 3108 2136
rect 3266 2102 3300 2136
rect 3458 2102 3492 2136
rect 3650 2102 3684 2136
rect 3842 2102 3876 2136
rect 4034 2102 4068 2136
rect 4226 2102 4260 2136
rect 2450 1667 2484 2043
rect 2546 1667 2580 2043
rect 2642 1667 2676 2043
rect 2738 1667 2772 2043
rect 2834 1667 2868 2043
rect 2930 1667 2964 2043
rect 3026 1667 3060 2043
rect 3122 1667 3156 2043
rect 3218 1667 3252 2043
rect 3314 1667 3348 2043
rect 3410 1667 3444 2043
rect 3506 1667 3540 2043
rect 3602 1667 3636 2043
rect 3698 1667 3732 2043
rect 3794 1667 3828 2043
rect 3890 1667 3924 2043
rect 3986 1667 4020 2043
rect 4082 1667 4116 2043
rect 4178 1667 4212 2043
rect 4274 1667 4308 2043
rect 4370 1667 4404 2043
rect 2594 1574 2628 1608
rect 2786 1574 2820 1608
rect 2978 1574 3012 1608
rect 3170 1574 3204 1608
rect 3362 1574 3396 1608
rect 3554 1574 3588 1608
rect 3746 1574 3780 1608
rect 3938 1574 3972 1608
rect 4130 1574 4164 1608
rect 4322 1574 4356 1608
rect 2594 1466 2628 1500
rect 2786 1466 2820 1500
rect 2978 1466 3012 1500
rect 3170 1466 3204 1500
rect 3362 1466 3396 1500
rect 3554 1466 3588 1500
rect 3746 1466 3780 1500
rect 3938 1466 3972 1500
rect 4130 1466 4164 1500
rect 4322 1466 4356 1500
rect 2450 1031 2484 1407
rect 2546 1031 2580 1407
rect 2642 1031 2676 1407
rect 2738 1031 2772 1407
rect 2834 1031 2868 1407
rect 2930 1031 2964 1407
rect 3026 1031 3060 1407
rect 3122 1031 3156 1407
rect 3218 1031 3252 1407
rect 3314 1031 3348 1407
rect 3410 1031 3444 1407
rect 3506 1031 3540 1407
rect 3602 1031 3636 1407
rect 3698 1031 3732 1407
rect 3794 1031 3828 1407
rect 3890 1031 3924 1407
rect 3986 1031 4020 1407
rect 4082 1031 4116 1407
rect 4178 1031 4212 1407
rect 4274 1031 4308 1407
rect 4370 1031 4404 1407
rect 2498 938 2532 972
rect 2690 938 2724 972
rect 2882 938 2916 972
rect 3074 938 3108 972
rect 3266 938 3300 972
rect 3458 938 3492 972
rect 3650 938 3684 972
rect 3842 938 3876 972
rect 4034 938 4068 972
rect 4226 938 4260 972
rect 274 64 308 98
rect 466 64 500 98
rect 658 64 692 98
rect 850 64 884 98
rect 1042 64 1076 98
rect 1234 64 1268 98
rect 1426 64 1460 98
rect 1618 64 1652 98
rect 1810 64 1844 98
rect 2002 64 2036 98
rect 130 -362 164 14
rect 226 -362 260 14
rect 322 -362 356 14
rect 418 -362 452 14
rect 514 -362 548 14
rect 610 -362 644 14
rect 706 -362 740 14
rect 802 -362 836 14
rect 898 -362 932 14
rect 994 -362 1028 14
rect 1090 -362 1124 14
rect 1186 -362 1220 14
rect 1282 -362 1316 14
rect 1378 -362 1412 14
rect 1474 -362 1508 14
rect 1570 -362 1604 14
rect 1666 -362 1700 14
rect 1762 -362 1796 14
rect 1858 -362 1892 14
rect 1954 -362 1988 14
rect 2050 -362 2084 14
rect 178 -446 212 -412
rect 370 -446 404 -412
rect 562 -446 596 -412
rect 754 -446 788 -412
rect 946 -446 980 -412
rect 1138 -446 1172 -412
rect 1330 -446 1364 -412
rect 1522 -446 1556 -412
rect 1714 -446 1748 -412
rect 1906 -446 1940 -412
rect 178 -554 212 -520
rect 370 -554 404 -520
rect 562 -554 596 -520
rect 754 -554 788 -520
rect 946 -554 980 -520
rect 1138 -554 1172 -520
rect 1330 -554 1364 -520
rect 1522 -554 1556 -520
rect 1714 -554 1748 -520
rect 1906 -554 1940 -520
rect 130 -980 164 -604
rect 226 -980 260 -604
rect 322 -980 356 -604
rect 418 -980 452 -604
rect 514 -980 548 -604
rect 610 -980 644 -604
rect 706 -980 740 -604
rect 802 -980 836 -604
rect 898 -980 932 -604
rect 994 -980 1028 -604
rect 1090 -980 1124 -604
rect 1186 -980 1220 -604
rect 1282 -980 1316 -604
rect 1378 -980 1412 -604
rect 1474 -980 1508 -604
rect 1570 -980 1604 -604
rect 1666 -980 1700 -604
rect 1762 -980 1796 -604
rect 1858 -980 1892 -604
rect 1954 -980 1988 -604
rect 2050 -980 2084 -604
rect 274 -1064 308 -1030
rect 466 -1064 500 -1030
rect 658 -1064 692 -1030
rect 850 -1064 884 -1030
rect 1042 -1064 1076 -1030
rect 1234 -1064 1268 -1030
rect 1426 -1064 1460 -1030
rect 1618 -1064 1652 -1030
rect 1810 -1064 1844 -1030
rect 2002 -1064 2036 -1030
rect 274 -1172 308 -1138
rect 466 -1172 500 -1138
rect 658 -1172 692 -1138
rect 850 -1172 884 -1138
rect 1042 -1172 1076 -1138
rect 1234 -1172 1268 -1138
rect 1426 -1172 1460 -1138
rect 1618 -1172 1652 -1138
rect 1810 -1172 1844 -1138
rect 2002 -1172 2036 -1138
rect 130 -1598 164 -1222
rect 226 -1598 260 -1222
rect 322 -1598 356 -1222
rect 418 -1598 452 -1222
rect 514 -1598 548 -1222
rect 610 -1598 644 -1222
rect 706 -1598 740 -1222
rect 802 -1598 836 -1222
rect 898 -1598 932 -1222
rect 994 -1598 1028 -1222
rect 1090 -1598 1124 -1222
rect 1186 -1598 1220 -1222
rect 1282 -1598 1316 -1222
rect 1378 -1598 1412 -1222
rect 1474 -1598 1508 -1222
rect 1570 -1598 1604 -1222
rect 1666 -1598 1700 -1222
rect 1762 -1598 1796 -1222
rect 1858 -1598 1892 -1222
rect 1954 -1598 1988 -1222
rect 2050 -1598 2084 -1222
rect 178 -1682 212 -1648
rect 370 -1682 404 -1648
rect 562 -1682 596 -1648
rect 754 -1682 788 -1648
rect 946 -1682 980 -1648
rect 1138 -1682 1172 -1648
rect 1330 -1682 1364 -1648
rect 1522 -1682 1556 -1648
rect 1714 -1682 1748 -1648
rect 1906 -1682 1940 -1648
rect 2498 506 2532 540
rect 2690 506 2724 540
rect 2882 506 2916 540
rect 3074 506 3108 540
rect 3266 506 3300 540
rect 3458 506 3492 540
rect 3650 506 3684 540
rect 3842 506 3876 540
rect 4034 506 4068 540
rect 4226 506 4260 540
rect 2450 80 2484 456
rect 2546 80 2580 456
rect 2642 80 2676 456
rect 2738 80 2772 456
rect 2834 80 2868 456
rect 2930 80 2964 456
rect 3026 80 3060 456
rect 3122 80 3156 456
rect 3218 80 3252 456
rect 3314 80 3348 456
rect 3410 80 3444 456
rect 3506 80 3540 456
rect 3602 80 3636 456
rect 3698 80 3732 456
rect 3794 80 3828 456
rect 3890 80 3924 456
rect 3986 80 4020 456
rect 4082 80 4116 456
rect 4178 80 4212 456
rect 4274 80 4308 456
rect 4370 80 4404 456
rect 2594 -4 2628 30
rect 2786 -4 2820 30
rect 2978 -4 3012 30
rect 3170 -4 3204 30
rect 3362 -4 3396 30
rect 3554 -4 3588 30
rect 3746 -4 3780 30
rect 3938 -4 3972 30
rect 4130 -4 4164 30
rect 4322 -4 4356 30
rect 2594 -112 2628 -78
rect 2786 -112 2820 -78
rect 2978 -112 3012 -78
rect 3170 -112 3204 -78
rect 3362 -112 3396 -78
rect 3554 -112 3588 -78
rect 3746 -112 3780 -78
rect 3938 -112 3972 -78
rect 4130 -112 4164 -78
rect 4322 -112 4356 -78
rect 2450 -538 2484 -162
rect 2546 -538 2580 -162
rect 2642 -538 2676 -162
rect 2738 -538 2772 -162
rect 2834 -538 2868 -162
rect 2930 -538 2964 -162
rect 3026 -538 3060 -162
rect 3122 -538 3156 -162
rect 3218 -538 3252 -162
rect 3314 -538 3348 -162
rect 3410 -538 3444 -162
rect 3506 -538 3540 -162
rect 3602 -538 3636 -162
rect 3698 -538 3732 -162
rect 3794 -538 3828 -162
rect 3890 -538 3924 -162
rect 3986 -538 4020 -162
rect 4082 -538 4116 -162
rect 4178 -538 4212 -162
rect 4274 -538 4308 -162
rect 4370 -538 4404 -162
rect 2498 -622 2532 -588
rect 2690 -622 2724 -588
rect 2882 -622 2916 -588
rect 3074 -622 3108 -588
rect 3266 -622 3300 -588
rect 3458 -622 3492 -588
rect 3650 -622 3684 -588
rect 3842 -622 3876 -588
rect 4034 -622 4068 -588
rect 4226 -622 4260 -588
rect -2306 -2316 -2272 -2282
rect -2114 -2316 -2080 -2282
rect -1922 -2316 -1888 -2282
rect -1730 -2316 -1696 -2282
rect -1538 -2316 -1504 -2282
rect -2450 -2742 -2416 -2366
rect -2354 -2742 -2320 -2366
rect -2258 -2742 -2224 -2366
rect -2162 -2742 -2128 -2366
rect -2066 -2742 -2032 -2366
rect -1970 -2742 -1936 -2366
rect -1874 -2742 -1840 -2366
rect -1778 -2742 -1744 -2366
rect -1682 -2742 -1648 -2366
rect -1586 -2742 -1552 -2366
rect -1490 -2742 -1456 -2366
rect -2402 -2826 -2368 -2792
rect -2210 -2826 -2176 -2792
rect -2018 -2826 -1984 -2792
rect -1826 -2826 -1792 -2792
rect -1634 -2826 -1600 -2792
rect -2402 -2934 -2368 -2900
rect -2210 -2934 -2176 -2900
rect -2018 -2934 -1984 -2900
rect -1826 -2934 -1792 -2900
rect -1634 -2934 -1600 -2900
rect -2450 -3360 -2416 -2984
rect -2354 -3360 -2320 -2984
rect -2258 -3360 -2224 -2984
rect -2162 -3360 -2128 -2984
rect -2066 -3360 -2032 -2984
rect -1970 -3360 -1936 -2984
rect -1874 -3360 -1840 -2984
rect -1778 -3360 -1744 -2984
rect -1682 -3360 -1648 -2984
rect -1586 -3360 -1552 -2984
rect -1490 -3360 -1456 -2984
rect -2306 -3444 -2272 -3410
rect -2114 -3444 -2080 -3410
rect -1922 -3444 -1888 -3410
rect -1730 -3444 -1696 -3410
rect -1538 -3444 -1504 -3410
rect -2306 -3552 -2272 -3518
rect -2114 -3552 -2080 -3518
rect -1922 -3552 -1888 -3518
rect -1730 -3552 -1696 -3518
rect -1538 -3552 -1504 -3518
rect -2450 -3978 -2416 -3602
rect -2354 -3978 -2320 -3602
rect -2258 -3978 -2224 -3602
rect -2162 -3978 -2128 -3602
rect -2066 -3978 -2032 -3602
rect -1970 -3978 -1936 -3602
rect -1874 -3978 -1840 -3602
rect -1778 -3978 -1744 -3602
rect -1682 -3978 -1648 -3602
rect -1586 -3978 -1552 -3602
rect -1490 -3978 -1456 -3602
rect -2402 -4062 -2368 -4028
rect -2210 -4062 -2176 -4028
rect -2018 -4062 -1984 -4028
rect -1826 -4062 -1792 -4028
rect -1634 -4062 -1600 -4028
rect -506 -2316 -472 -2282
rect -314 -2316 -280 -2282
rect -122 -2316 -88 -2282
rect 70 -2316 104 -2282
rect 262 -2316 296 -2282
rect -650 -2742 -616 -2366
rect -554 -2742 -520 -2366
rect -458 -2742 -424 -2366
rect -362 -2742 -328 -2366
rect -266 -2742 -232 -2366
rect -170 -2742 -136 -2366
rect -74 -2742 -40 -2366
rect 22 -2742 56 -2366
rect 118 -2742 152 -2366
rect 214 -2742 248 -2366
rect 310 -2742 344 -2366
rect -602 -2826 -568 -2792
rect -410 -2826 -376 -2792
rect -218 -2826 -184 -2792
rect -26 -2826 8 -2792
rect 166 -2826 200 -2792
rect -602 -2934 -568 -2900
rect -410 -2934 -376 -2900
rect -218 -2934 -184 -2900
rect -26 -2934 8 -2900
rect 166 -2934 200 -2900
rect -650 -3360 -616 -2984
rect -554 -3360 -520 -2984
rect -458 -3360 -424 -2984
rect -362 -3360 -328 -2984
rect -266 -3360 -232 -2984
rect -170 -3360 -136 -2984
rect -74 -3360 -40 -2984
rect 22 -3360 56 -2984
rect 118 -3360 152 -2984
rect 214 -3360 248 -2984
rect 310 -3360 344 -2984
rect -506 -3444 -472 -3410
rect -314 -3444 -280 -3410
rect -122 -3444 -88 -3410
rect 70 -3444 104 -3410
rect 262 -3444 296 -3410
rect -506 -3552 -472 -3518
rect -314 -3552 -280 -3518
rect -122 -3552 -88 -3518
rect 70 -3552 104 -3518
rect 262 -3552 296 -3518
rect -650 -3978 -616 -3602
rect -554 -3978 -520 -3602
rect -458 -3978 -424 -3602
rect -362 -3978 -328 -3602
rect -266 -3978 -232 -3602
rect -170 -3978 -136 -3602
rect -74 -3978 -40 -3602
rect 22 -3978 56 -3602
rect 118 -3978 152 -3602
rect 214 -3978 248 -3602
rect 310 -3978 344 -3602
rect -602 -4062 -568 -4028
rect -410 -4062 -376 -4028
rect -218 -4062 -184 -4028
rect -26 -4062 8 -4028
rect 166 -4062 200 -4028
rect 1294 -2316 1328 -2282
rect 1486 -2316 1520 -2282
rect 1678 -2316 1712 -2282
rect 1870 -2316 1904 -2282
rect 2062 -2316 2096 -2282
rect 1150 -2742 1184 -2366
rect 1246 -2742 1280 -2366
rect 1342 -2742 1376 -2366
rect 1438 -2742 1472 -2366
rect 1534 -2742 1568 -2366
rect 1630 -2742 1664 -2366
rect 1726 -2742 1760 -2366
rect 1822 -2742 1856 -2366
rect 1918 -2742 1952 -2366
rect 2014 -2742 2048 -2366
rect 2110 -2742 2144 -2366
rect 1198 -2826 1232 -2792
rect 1390 -2826 1424 -2792
rect 1582 -2826 1616 -2792
rect 1774 -2826 1808 -2792
rect 1966 -2826 2000 -2792
rect 1198 -2934 1232 -2900
rect 1390 -2934 1424 -2900
rect 1582 -2934 1616 -2900
rect 1774 -2934 1808 -2900
rect 1966 -2934 2000 -2900
rect 1150 -3360 1184 -2984
rect 1246 -3360 1280 -2984
rect 1342 -3360 1376 -2984
rect 1438 -3360 1472 -2984
rect 1534 -3360 1568 -2984
rect 1630 -3360 1664 -2984
rect 1726 -3360 1760 -2984
rect 1822 -3360 1856 -2984
rect 1918 -3360 1952 -2984
rect 2014 -3360 2048 -2984
rect 2110 -3360 2144 -2984
rect 1294 -3444 1328 -3410
rect 1486 -3444 1520 -3410
rect 1678 -3444 1712 -3410
rect 1870 -3444 1904 -3410
rect 2062 -3444 2096 -3410
rect 1294 -3552 1328 -3518
rect 1486 -3552 1520 -3518
rect 1678 -3552 1712 -3518
rect 1870 -3552 1904 -3518
rect 2062 -3552 2096 -3518
rect 1150 -3978 1184 -3602
rect 1246 -3978 1280 -3602
rect 1342 -3978 1376 -3602
rect 1438 -3978 1472 -3602
rect 1534 -3978 1568 -3602
rect 1630 -3978 1664 -3602
rect 1726 -3978 1760 -3602
rect 1822 -3978 1856 -3602
rect 1918 -3978 1952 -3602
rect 2014 -3978 2048 -3602
rect 2110 -3978 2144 -3602
rect 1198 -4062 1232 -4028
rect 1390 -4062 1424 -4028
rect 1582 -4062 1616 -4028
rect 1774 -4062 1808 -4028
rect 1966 -4062 2000 -4028
rect 3094 -2316 3128 -2282
rect 3286 -2316 3320 -2282
rect 3478 -2316 3512 -2282
rect 3670 -2316 3704 -2282
rect 3862 -2316 3896 -2282
rect 2950 -2742 2984 -2366
rect 3046 -2742 3080 -2366
rect 3142 -2742 3176 -2366
rect 3238 -2742 3272 -2366
rect 3334 -2742 3368 -2366
rect 3430 -2742 3464 -2366
rect 3526 -2742 3560 -2366
rect 3622 -2742 3656 -2366
rect 3718 -2742 3752 -2366
rect 3814 -2742 3848 -2366
rect 3910 -2742 3944 -2366
rect 2998 -2826 3032 -2792
rect 3190 -2826 3224 -2792
rect 3382 -2826 3416 -2792
rect 3574 -2826 3608 -2792
rect 3766 -2826 3800 -2792
rect 2998 -2934 3032 -2900
rect 3190 -2934 3224 -2900
rect 3382 -2934 3416 -2900
rect 3574 -2934 3608 -2900
rect 3766 -2934 3800 -2900
rect 2950 -3360 2984 -2984
rect 3046 -3360 3080 -2984
rect 3142 -3360 3176 -2984
rect 3238 -3360 3272 -2984
rect 3334 -3360 3368 -2984
rect 3430 -3360 3464 -2984
rect 3526 -3360 3560 -2984
rect 3622 -3360 3656 -2984
rect 3718 -3360 3752 -2984
rect 3814 -3360 3848 -2984
rect 3910 -3360 3944 -2984
rect 3094 -3444 3128 -3410
rect 3286 -3444 3320 -3410
rect 3478 -3444 3512 -3410
rect 3670 -3444 3704 -3410
rect 3862 -3444 3896 -3410
rect 3094 -3552 3128 -3518
rect 3286 -3552 3320 -3518
rect 3478 -3552 3512 -3518
rect 3670 -3552 3704 -3518
rect 3862 -3552 3896 -3518
rect 2950 -3978 2984 -3602
rect 3046 -3978 3080 -3602
rect 3142 -3978 3176 -3602
rect 3238 -3978 3272 -3602
rect 3334 -3978 3368 -3602
rect 3430 -3978 3464 -3602
rect 3526 -3978 3560 -3602
rect 3622 -3978 3656 -3602
rect 3718 -3978 3752 -3602
rect 3814 -3978 3848 -3602
rect 3910 -3978 3944 -3602
rect 2998 -4062 3032 -4028
rect 3190 -4062 3224 -4028
rect 3382 -4062 3416 -4028
rect 3574 -4062 3608 -4028
rect 3766 -4062 3800 -4028
rect 5094 2072 5128 2106
rect 5286 2072 5320 2106
rect 5478 2072 5512 2106
rect 5670 2072 5704 2106
rect 5862 2072 5896 2106
rect 6054 2072 6088 2106
rect 6246 2072 6280 2106
rect 6438 2072 6472 2106
rect 6630 2072 6664 2106
rect 6822 2072 6856 2106
rect 4950 1646 4984 2022
rect 5046 1646 5080 2022
rect 5142 1646 5176 2022
rect 5238 1646 5272 2022
rect 5334 1646 5368 2022
rect 5430 1646 5464 2022
rect 5526 1646 5560 2022
rect 5622 1646 5656 2022
rect 5718 1646 5752 2022
rect 5814 1646 5848 2022
rect 5910 1646 5944 2022
rect 6006 1646 6040 2022
rect 6102 1646 6136 2022
rect 6198 1646 6232 2022
rect 6294 1646 6328 2022
rect 6390 1646 6424 2022
rect 6486 1646 6520 2022
rect 6582 1646 6616 2022
rect 6678 1646 6712 2022
rect 6774 1646 6808 2022
rect 6870 1646 6904 2022
rect 4998 1562 5032 1596
rect 5190 1562 5224 1596
rect 5382 1562 5416 1596
rect 5574 1562 5608 1596
rect 5766 1562 5800 1596
rect 5958 1562 5992 1596
rect 6150 1562 6184 1596
rect 6342 1562 6376 1596
rect 6534 1562 6568 1596
rect 6726 1562 6760 1596
rect 4998 1454 5032 1488
rect 5190 1454 5224 1488
rect 5382 1454 5416 1488
rect 5574 1454 5608 1488
rect 5766 1454 5800 1488
rect 5958 1454 5992 1488
rect 6150 1454 6184 1488
rect 6342 1454 6376 1488
rect 6534 1454 6568 1488
rect 6726 1454 6760 1488
rect 4950 1028 4984 1404
rect 5046 1028 5080 1404
rect 5142 1028 5176 1404
rect 5238 1028 5272 1404
rect 5334 1028 5368 1404
rect 5430 1028 5464 1404
rect 5526 1028 5560 1404
rect 5622 1028 5656 1404
rect 5718 1028 5752 1404
rect 5814 1028 5848 1404
rect 5910 1028 5944 1404
rect 6006 1028 6040 1404
rect 6102 1028 6136 1404
rect 6198 1028 6232 1404
rect 6294 1028 6328 1404
rect 6390 1028 6424 1404
rect 6486 1028 6520 1404
rect 6582 1028 6616 1404
rect 6678 1028 6712 1404
rect 6774 1028 6808 1404
rect 6870 1028 6904 1404
rect 5094 944 5128 978
rect 5286 944 5320 978
rect 5478 944 5512 978
rect 5670 944 5704 978
rect 5862 944 5896 978
rect 6054 944 6088 978
rect 6246 944 6280 978
rect 6438 944 6472 978
rect 6630 944 6664 978
rect 6822 944 6856 978
rect 5094 836 5128 870
rect 5286 836 5320 870
rect 5478 836 5512 870
rect 5670 836 5704 870
rect 5862 836 5896 870
rect 6054 836 6088 870
rect 6246 836 6280 870
rect 6438 836 6472 870
rect 6630 836 6664 870
rect 6822 836 6856 870
rect 4950 410 4984 786
rect 5046 410 5080 786
rect 5142 410 5176 786
rect 5238 410 5272 786
rect 5334 410 5368 786
rect 5430 410 5464 786
rect 5526 410 5560 786
rect 5622 410 5656 786
rect 5718 410 5752 786
rect 5814 410 5848 786
rect 5910 410 5944 786
rect 6006 410 6040 786
rect 6102 410 6136 786
rect 6198 410 6232 786
rect 6294 410 6328 786
rect 6390 410 6424 786
rect 6486 410 6520 786
rect 6582 410 6616 786
rect 6678 410 6712 786
rect 6774 410 6808 786
rect 6870 410 6904 786
rect 4998 326 5032 360
rect 5190 326 5224 360
rect 5382 326 5416 360
rect 5574 326 5608 360
rect 5766 326 5800 360
rect 5958 326 5992 360
rect 6150 326 6184 360
rect 6342 326 6376 360
rect 6534 326 6568 360
rect 6726 326 6760 360
rect 4998 218 5032 252
rect 5190 218 5224 252
rect 5382 218 5416 252
rect 5574 218 5608 252
rect 5766 218 5800 252
rect 5958 218 5992 252
rect 6150 218 6184 252
rect 6342 218 6376 252
rect 6534 218 6568 252
rect 6726 218 6760 252
rect 4950 -208 4984 168
rect 5046 -208 5080 168
rect 5142 -208 5176 168
rect 5238 -208 5272 168
rect 5334 -208 5368 168
rect 5430 -208 5464 168
rect 5526 -208 5560 168
rect 5622 -208 5656 168
rect 5718 -208 5752 168
rect 5814 -208 5848 168
rect 5910 -208 5944 168
rect 6006 -208 6040 168
rect 6102 -208 6136 168
rect 6198 -208 6232 168
rect 6294 -208 6328 168
rect 6390 -208 6424 168
rect 6486 -208 6520 168
rect 6582 -208 6616 168
rect 6678 -208 6712 168
rect 6774 -208 6808 168
rect 6870 -208 6904 168
rect 5094 -292 5128 -258
rect 5286 -292 5320 -258
rect 5478 -292 5512 -258
rect 5670 -292 5704 -258
rect 5862 -292 5896 -258
rect 6054 -292 6088 -258
rect 6246 -292 6280 -258
rect 6438 -292 6472 -258
rect 6630 -292 6664 -258
rect 6822 -292 6856 -258
rect 5094 -400 5128 -366
rect 5286 -400 5320 -366
rect 5478 -400 5512 -366
rect 5670 -400 5704 -366
rect 5862 -400 5896 -366
rect 6054 -400 6088 -366
rect 6246 -400 6280 -366
rect 6438 -400 6472 -366
rect 6630 -400 6664 -366
rect 6822 -400 6856 -366
rect 4950 -826 4984 -450
rect 5046 -826 5080 -450
rect 5142 -826 5176 -450
rect 5238 -826 5272 -450
rect 5334 -826 5368 -450
rect 5430 -826 5464 -450
rect 5526 -826 5560 -450
rect 5622 -826 5656 -450
rect 5718 -826 5752 -450
rect 5814 -826 5848 -450
rect 5910 -826 5944 -450
rect 6006 -826 6040 -450
rect 6102 -826 6136 -450
rect 6198 -826 6232 -450
rect 6294 -826 6328 -450
rect 6390 -826 6424 -450
rect 6486 -826 6520 -450
rect 6582 -826 6616 -450
rect 6678 -826 6712 -450
rect 6774 -826 6808 -450
rect 6870 -826 6904 -450
rect 4998 -910 5032 -876
rect 5190 -910 5224 -876
rect 5382 -910 5416 -876
rect 5574 -910 5608 -876
rect 5766 -910 5800 -876
rect 5958 -910 5992 -876
rect 6150 -910 6184 -876
rect 6342 -910 6376 -876
rect 6534 -910 6568 -876
rect 6726 -910 6760 -876
rect 4998 -1018 5032 -984
rect 5190 -1018 5224 -984
rect 5382 -1018 5416 -984
rect 5574 -1018 5608 -984
rect 5766 -1018 5800 -984
rect 5958 -1018 5992 -984
rect 6150 -1018 6184 -984
rect 6342 -1018 6376 -984
rect 6534 -1018 6568 -984
rect 6726 -1018 6760 -984
rect 4950 -1444 4984 -1068
rect 5046 -1444 5080 -1068
rect 5142 -1444 5176 -1068
rect 5238 -1444 5272 -1068
rect 5334 -1444 5368 -1068
rect 5430 -1444 5464 -1068
rect 5526 -1444 5560 -1068
rect 5622 -1444 5656 -1068
rect 5718 -1444 5752 -1068
rect 5814 -1444 5848 -1068
rect 5910 -1444 5944 -1068
rect 6006 -1444 6040 -1068
rect 6102 -1444 6136 -1068
rect 6198 -1444 6232 -1068
rect 6294 -1444 6328 -1068
rect 6390 -1444 6424 -1068
rect 6486 -1444 6520 -1068
rect 6582 -1444 6616 -1068
rect 6678 -1444 6712 -1068
rect 6774 -1444 6808 -1068
rect 6870 -1444 6904 -1068
rect 5094 -1528 5128 -1494
rect 5286 -1528 5320 -1494
rect 5478 -1528 5512 -1494
rect 5670 -1528 5704 -1494
rect 5862 -1528 5896 -1494
rect 6054 -1528 6088 -1494
rect 6246 -1528 6280 -1494
rect 6438 -1528 6472 -1494
rect 6630 -1528 6664 -1494
rect 6822 -1528 6856 -1494
rect 5094 -1636 5128 -1602
rect 5286 -1636 5320 -1602
rect 5478 -1636 5512 -1602
rect 5670 -1636 5704 -1602
rect 5862 -1636 5896 -1602
rect 6054 -1636 6088 -1602
rect 6246 -1636 6280 -1602
rect 6438 -1636 6472 -1602
rect 6630 -1636 6664 -1602
rect 6822 -1636 6856 -1602
rect 4950 -2062 4984 -1686
rect 5046 -2062 5080 -1686
rect 5142 -2062 5176 -1686
rect 5238 -2062 5272 -1686
rect 5334 -2062 5368 -1686
rect 5430 -2062 5464 -1686
rect 5526 -2062 5560 -1686
rect 5622 -2062 5656 -1686
rect 5718 -2062 5752 -1686
rect 5814 -2062 5848 -1686
rect 5910 -2062 5944 -1686
rect 6006 -2062 6040 -1686
rect 6102 -2062 6136 -1686
rect 6198 -2062 6232 -1686
rect 6294 -2062 6328 -1686
rect 6390 -2062 6424 -1686
rect 6486 -2062 6520 -1686
rect 6582 -2062 6616 -1686
rect 6678 -2062 6712 -1686
rect 6774 -2062 6808 -1686
rect 6870 -2062 6904 -1686
rect 4998 -2146 5032 -2112
rect 5190 -2146 5224 -2112
rect 5382 -2146 5416 -2112
rect 5574 -2146 5608 -2112
rect 5766 -2146 5800 -2112
rect 5958 -2146 5992 -2112
rect 6150 -2146 6184 -2112
rect 6342 -2146 6376 -2112
rect 6534 -2146 6568 -2112
rect 6726 -2146 6760 -2112
rect 4998 -2254 5032 -2220
rect 5190 -2254 5224 -2220
rect 5382 -2254 5416 -2220
rect 5574 -2254 5608 -2220
rect 5766 -2254 5800 -2220
rect 5958 -2254 5992 -2220
rect 6150 -2254 6184 -2220
rect 6342 -2254 6376 -2220
rect 6534 -2254 6568 -2220
rect 6726 -2254 6760 -2220
rect 4950 -2680 4984 -2304
rect 5046 -2680 5080 -2304
rect 5142 -2680 5176 -2304
rect 5238 -2680 5272 -2304
rect 5334 -2680 5368 -2304
rect 5430 -2680 5464 -2304
rect 5526 -2680 5560 -2304
rect 5622 -2680 5656 -2304
rect 5718 -2680 5752 -2304
rect 5814 -2680 5848 -2304
rect 5910 -2680 5944 -2304
rect 6006 -2680 6040 -2304
rect 6102 -2680 6136 -2304
rect 6198 -2680 6232 -2304
rect 6294 -2680 6328 -2304
rect 6390 -2680 6424 -2304
rect 6486 -2680 6520 -2304
rect 6582 -2680 6616 -2304
rect 6678 -2680 6712 -2304
rect 6774 -2680 6808 -2304
rect 6870 -2680 6904 -2304
rect 5094 -2764 5128 -2730
rect 5286 -2764 5320 -2730
rect 5478 -2764 5512 -2730
rect 5670 -2764 5704 -2730
rect 5862 -2764 5896 -2730
rect 6054 -2764 6088 -2730
rect 6246 -2764 6280 -2730
rect 6438 -2764 6472 -2730
rect 6630 -2764 6664 -2730
rect 6822 -2764 6856 -2730
rect 5094 -2872 5128 -2838
rect 5286 -2872 5320 -2838
rect 5478 -2872 5512 -2838
rect 5670 -2872 5704 -2838
rect 5862 -2872 5896 -2838
rect 6054 -2872 6088 -2838
rect 6246 -2872 6280 -2838
rect 6438 -2872 6472 -2838
rect 6630 -2872 6664 -2838
rect 6822 -2872 6856 -2838
rect 4950 -3298 4984 -2922
rect 5046 -3298 5080 -2922
rect 5142 -3298 5176 -2922
rect 5238 -3298 5272 -2922
rect 5334 -3298 5368 -2922
rect 5430 -3298 5464 -2922
rect 5526 -3298 5560 -2922
rect 5622 -3298 5656 -2922
rect 5718 -3298 5752 -2922
rect 5814 -3298 5848 -2922
rect 5910 -3298 5944 -2922
rect 6006 -3298 6040 -2922
rect 6102 -3298 6136 -2922
rect 6198 -3298 6232 -2922
rect 6294 -3298 6328 -2922
rect 6390 -3298 6424 -2922
rect 6486 -3298 6520 -2922
rect 6582 -3298 6616 -2922
rect 6678 -3298 6712 -2922
rect 6774 -3298 6808 -2922
rect 6870 -3298 6904 -2922
rect 4998 -3382 5032 -3348
rect 5190 -3382 5224 -3348
rect 5382 -3382 5416 -3348
rect 5574 -3382 5608 -3348
rect 5766 -3382 5800 -3348
rect 5958 -3382 5992 -3348
rect 6150 -3382 6184 -3348
rect 6342 -3382 6376 -3348
rect 6534 -3382 6568 -3348
rect 6726 -3382 6760 -3348
rect -2388 -4462 -2220 -4428
rect -2130 -4462 -1962 -4428
rect -1872 -4462 -1704 -4428
rect -1614 -4462 -1446 -4428
rect -1356 -4462 -1188 -4428
rect -2450 -4888 -2416 -4512
rect -2192 -4888 -2158 -4512
rect -1934 -4888 -1900 -4512
rect -1676 -4888 -1642 -4512
rect -1418 -4888 -1384 -4512
rect -1160 -4888 -1126 -4512
rect -2388 -4972 -2220 -4938
rect -2130 -4972 -1962 -4938
rect -1872 -4972 -1704 -4938
rect -1614 -4972 -1446 -4938
rect -1356 -4972 -1188 -4938
rect -2388 -5080 -2220 -5046
rect -2130 -5080 -1962 -5046
rect -1872 -5080 -1704 -5046
rect -1614 -5080 -1446 -5046
rect -1356 -5080 -1188 -5046
rect -2450 -5506 -2416 -5130
rect -2192 -5506 -2158 -5130
rect -1934 -5506 -1900 -5130
rect -1676 -5506 -1642 -5130
rect -1418 -5506 -1384 -5130
rect -1160 -5506 -1126 -5130
rect -2388 -5590 -2220 -5556
rect -2130 -5590 -1962 -5556
rect -1872 -5590 -1704 -5556
rect -1614 -5590 -1446 -5556
rect -1356 -5590 -1188 -5556
rect -2388 -5698 -2220 -5664
rect -2130 -5698 -1962 -5664
rect -1872 -5698 -1704 -5664
rect -1614 -5698 -1446 -5664
rect -1356 -5698 -1188 -5664
rect -2450 -6124 -2416 -5748
rect -2192 -6124 -2158 -5748
rect -1934 -6124 -1900 -5748
rect -1676 -6124 -1642 -5748
rect -1418 -6124 -1384 -5748
rect -1160 -6124 -1126 -5748
rect -2388 -6208 -2220 -6174
rect -2130 -6208 -1962 -6174
rect -1872 -6208 -1704 -6174
rect -1614 -6208 -1446 -6174
rect -1356 -6208 -1188 -6174
rect -2388 -6316 -2220 -6282
rect -2130 -6316 -1962 -6282
rect -1872 -6316 -1704 -6282
rect -1614 -6316 -1446 -6282
rect -1356 -6316 -1188 -6282
rect -2450 -6742 -2416 -6366
rect -2192 -6742 -2158 -6366
rect -1934 -6742 -1900 -6366
rect -1676 -6742 -1642 -6366
rect -1418 -6742 -1384 -6366
rect -1160 -6742 -1126 -6366
rect -2388 -6826 -2220 -6792
rect -2130 -6826 -1962 -6792
rect -1872 -6826 -1704 -6792
rect -1614 -6826 -1446 -6792
rect -1356 -6826 -1188 -6792
rect -2388 -6934 -2220 -6900
rect -2130 -6934 -1962 -6900
rect -1872 -6934 -1704 -6900
rect -1614 -6934 -1446 -6900
rect -1356 -6934 -1188 -6900
rect -2450 -7360 -2416 -6984
rect -2192 -7360 -2158 -6984
rect -1934 -7360 -1900 -6984
rect -1676 -7360 -1642 -6984
rect -1418 -7360 -1384 -6984
rect -1160 -7360 -1126 -6984
rect -2388 -7444 -2220 -7410
rect -2130 -7444 -1962 -7410
rect -1872 -7444 -1704 -7410
rect -1614 -7444 -1446 -7410
rect -1356 -7444 -1188 -7410
rect -2388 -7552 -2220 -7518
rect -2130 -7552 -1962 -7518
rect -1872 -7552 -1704 -7518
rect -1614 -7552 -1446 -7518
rect -1356 -7552 -1188 -7518
rect -2450 -7978 -2416 -7602
rect -2192 -7978 -2158 -7602
rect -1934 -7978 -1900 -7602
rect -1676 -7978 -1642 -7602
rect -1418 -7978 -1384 -7602
rect -1160 -7978 -1126 -7602
rect -2388 -8062 -2220 -8028
rect -2130 -8062 -1962 -8028
rect -1872 -8062 -1704 -8028
rect -1614 -8062 -1446 -8028
rect -1356 -8062 -1188 -8028
rect -980 -8160 -800 -7960
rect -588 -4462 -420 -4428
rect -330 -4462 -162 -4428
rect -72 -4462 96 -4428
rect 186 -4462 354 -4428
rect 444 -4462 612 -4428
rect -650 -4888 -616 -4512
rect -392 -4888 -358 -4512
rect -134 -4888 -100 -4512
rect 124 -4888 158 -4512
rect 382 -4888 416 -4512
rect 640 -4888 674 -4512
rect -588 -4972 -420 -4938
rect -330 -4972 -162 -4938
rect -72 -4972 96 -4938
rect 186 -4972 354 -4938
rect 444 -4972 612 -4938
rect -588 -5080 -420 -5046
rect -330 -5080 -162 -5046
rect -72 -5080 96 -5046
rect 186 -5080 354 -5046
rect 444 -5080 612 -5046
rect -650 -5506 -616 -5130
rect -392 -5506 -358 -5130
rect -134 -5506 -100 -5130
rect 124 -5506 158 -5130
rect 382 -5506 416 -5130
rect 640 -5506 674 -5130
rect -588 -5590 -420 -5556
rect -330 -5590 -162 -5556
rect -72 -5590 96 -5556
rect 186 -5590 354 -5556
rect 444 -5590 612 -5556
rect -588 -5698 -420 -5664
rect -330 -5698 -162 -5664
rect -72 -5698 96 -5664
rect 186 -5698 354 -5664
rect 444 -5698 612 -5664
rect -650 -6124 -616 -5748
rect -392 -6124 -358 -5748
rect -134 -6124 -100 -5748
rect 124 -6124 158 -5748
rect 382 -6124 416 -5748
rect 640 -6124 674 -5748
rect -588 -6208 -420 -6174
rect -330 -6208 -162 -6174
rect -72 -6208 96 -6174
rect 186 -6208 354 -6174
rect 444 -6208 612 -6174
rect -588 -6316 -420 -6282
rect -330 -6316 -162 -6282
rect -72 -6316 96 -6282
rect 186 -6316 354 -6282
rect 444 -6316 612 -6282
rect -650 -6742 -616 -6366
rect -392 -6742 -358 -6366
rect -134 -6742 -100 -6366
rect 124 -6742 158 -6366
rect 382 -6742 416 -6366
rect 640 -6742 674 -6366
rect -588 -6826 -420 -6792
rect -330 -6826 -162 -6792
rect -72 -6826 96 -6792
rect 186 -6826 354 -6792
rect 444 -6826 612 -6792
rect -588 -6934 -420 -6900
rect -330 -6934 -162 -6900
rect -72 -6934 96 -6900
rect 186 -6934 354 -6900
rect 444 -6934 612 -6900
rect -650 -7360 -616 -6984
rect -392 -7360 -358 -6984
rect -134 -7360 -100 -6984
rect 124 -7360 158 -6984
rect 382 -7360 416 -6984
rect 640 -7360 674 -6984
rect -588 -7444 -420 -7410
rect -330 -7444 -162 -7410
rect -72 -7444 96 -7410
rect 186 -7444 354 -7410
rect 444 -7444 612 -7410
rect -588 -7552 -420 -7518
rect -330 -7552 -162 -7518
rect -72 -7552 96 -7518
rect 186 -7552 354 -7518
rect 444 -7552 612 -7518
rect -650 -7978 -616 -7602
rect -392 -7978 -358 -7602
rect -134 -7978 -100 -7602
rect 124 -7978 158 -7602
rect 382 -7978 416 -7602
rect 640 -7978 674 -7602
rect -588 -8062 -420 -8028
rect -330 -8062 -162 -8028
rect -72 -8062 96 -8028
rect 186 -8062 354 -8028
rect 444 -8062 612 -8028
rect 1212 -4462 1380 -4428
rect 1470 -4462 1638 -4428
rect 1728 -4462 1896 -4428
rect 1986 -4462 2154 -4428
rect 2244 -4462 2412 -4428
rect 1150 -4888 1184 -4512
rect 1408 -4888 1442 -4512
rect 1666 -4888 1700 -4512
rect 1924 -4888 1958 -4512
rect 2182 -4888 2216 -4512
rect 2440 -4888 2474 -4512
rect 1212 -4972 1380 -4938
rect 1470 -4972 1638 -4938
rect 1728 -4972 1896 -4938
rect 1986 -4972 2154 -4938
rect 2244 -4972 2412 -4938
rect 1212 -5080 1380 -5046
rect 1470 -5080 1638 -5046
rect 1728 -5080 1896 -5046
rect 1986 -5080 2154 -5046
rect 2244 -5080 2412 -5046
rect 1150 -5506 1184 -5130
rect 1408 -5506 1442 -5130
rect 1666 -5506 1700 -5130
rect 1924 -5506 1958 -5130
rect 2182 -5506 2216 -5130
rect 2440 -5506 2474 -5130
rect 1212 -5590 1380 -5556
rect 1470 -5590 1638 -5556
rect 1728 -5590 1896 -5556
rect 1986 -5590 2154 -5556
rect 2244 -5590 2412 -5556
rect 1212 -5698 1380 -5664
rect 1470 -5698 1638 -5664
rect 1728 -5698 1896 -5664
rect 1986 -5698 2154 -5664
rect 2244 -5698 2412 -5664
rect 1150 -6124 1184 -5748
rect 1408 -6124 1442 -5748
rect 1666 -6124 1700 -5748
rect 1924 -6124 1958 -5748
rect 2182 -6124 2216 -5748
rect 2440 -6124 2474 -5748
rect 1212 -6208 1380 -6174
rect 1470 -6208 1638 -6174
rect 1728 -6208 1896 -6174
rect 1986 -6208 2154 -6174
rect 2244 -6208 2412 -6174
rect 1212 -6316 1380 -6282
rect 1470 -6316 1638 -6282
rect 1728 -6316 1896 -6282
rect 1986 -6316 2154 -6282
rect 2244 -6316 2412 -6282
rect 1150 -6742 1184 -6366
rect 1408 -6742 1442 -6366
rect 1666 -6742 1700 -6366
rect 1924 -6742 1958 -6366
rect 2182 -6742 2216 -6366
rect 2440 -6742 2474 -6366
rect 1212 -6826 1380 -6792
rect 1470 -6826 1638 -6792
rect 1728 -6826 1896 -6792
rect 1986 -6826 2154 -6792
rect 2244 -6826 2412 -6792
rect 1212 -6934 1380 -6900
rect 1470 -6934 1638 -6900
rect 1728 -6934 1896 -6900
rect 1986 -6934 2154 -6900
rect 2244 -6934 2412 -6900
rect 1150 -7360 1184 -6984
rect 1408 -7360 1442 -6984
rect 1666 -7360 1700 -6984
rect 1924 -7360 1958 -6984
rect 2182 -7360 2216 -6984
rect 2440 -7360 2474 -6984
rect 1212 -7444 1380 -7410
rect 1470 -7444 1638 -7410
rect 1728 -7444 1896 -7410
rect 1986 -7444 2154 -7410
rect 2244 -7444 2412 -7410
rect 1212 -7552 1380 -7518
rect 1470 -7552 1638 -7518
rect 1728 -7552 1896 -7518
rect 1986 -7552 2154 -7518
rect 2244 -7552 2412 -7518
rect 1150 -7978 1184 -7602
rect 1408 -7978 1442 -7602
rect 1666 -7978 1700 -7602
rect 1924 -7978 1958 -7602
rect 2182 -7978 2216 -7602
rect 2440 -7978 2474 -7602
rect 1212 -8062 1380 -8028
rect 1470 -8062 1638 -8028
rect 1728 -8062 1896 -8028
rect 1986 -8062 2154 -8028
rect 2244 -8062 2412 -8028
rect 3012 -4462 3180 -4428
rect 3270 -4462 3438 -4428
rect 3528 -4462 3696 -4428
rect 3786 -4462 3954 -4428
rect 4044 -4462 4212 -4428
rect 2950 -4888 2984 -4512
rect 3208 -4888 3242 -4512
rect 3466 -4888 3500 -4512
rect 3724 -4888 3758 -4512
rect 3982 -4888 4016 -4512
rect 4240 -4888 4274 -4512
rect 3012 -4972 3180 -4938
rect 3270 -4972 3438 -4938
rect 3528 -4972 3696 -4938
rect 3786 -4972 3954 -4938
rect 4044 -4972 4212 -4938
rect 3012 -5080 3180 -5046
rect 3270 -5080 3438 -5046
rect 3528 -5080 3696 -5046
rect 3786 -5080 3954 -5046
rect 4044 -5080 4212 -5046
rect 2950 -5506 2984 -5130
rect 3208 -5506 3242 -5130
rect 3466 -5506 3500 -5130
rect 3724 -5506 3758 -5130
rect 3982 -5506 4016 -5130
rect 4240 -5506 4274 -5130
rect 3012 -5590 3180 -5556
rect 3270 -5590 3438 -5556
rect 3528 -5590 3696 -5556
rect 3786 -5590 3954 -5556
rect 4044 -5590 4212 -5556
rect 3012 -5698 3180 -5664
rect 3270 -5698 3438 -5664
rect 3528 -5698 3696 -5664
rect 3786 -5698 3954 -5664
rect 4044 -5698 4212 -5664
rect 2950 -6124 2984 -5748
rect 3208 -6124 3242 -5748
rect 3466 -6124 3500 -5748
rect 3724 -6124 3758 -5748
rect 3982 -6124 4016 -5748
rect 4240 -6124 4274 -5748
rect 3012 -6208 3180 -6174
rect 3270 -6208 3438 -6174
rect 3528 -6208 3696 -6174
rect 3786 -6208 3954 -6174
rect 4044 -6208 4212 -6174
rect 3012 -6316 3180 -6282
rect 3270 -6316 3438 -6282
rect 3528 -6316 3696 -6282
rect 3786 -6316 3954 -6282
rect 4044 -6316 4212 -6282
rect 2950 -6742 2984 -6366
rect 3208 -6742 3242 -6366
rect 3466 -6742 3500 -6366
rect 3724 -6742 3758 -6366
rect 3982 -6742 4016 -6366
rect 4240 -6742 4274 -6366
rect 3012 -6826 3180 -6792
rect 3270 -6826 3438 -6792
rect 3528 -6826 3696 -6792
rect 3786 -6826 3954 -6792
rect 4044 -6826 4212 -6792
rect 3012 -6934 3180 -6900
rect 3270 -6934 3438 -6900
rect 3528 -6934 3696 -6900
rect 3786 -6934 3954 -6900
rect 4044 -6934 4212 -6900
rect 2950 -7360 2984 -6984
rect 3208 -7360 3242 -6984
rect 3466 -7360 3500 -6984
rect 3724 -7360 3758 -6984
rect 3982 -7360 4016 -6984
rect 4240 -7360 4274 -6984
rect 3012 -7444 3180 -7410
rect 3270 -7444 3438 -7410
rect 3528 -7444 3696 -7410
rect 3786 -7444 3954 -7410
rect 4044 -7444 4212 -7410
rect 3012 -7552 3180 -7518
rect 3270 -7552 3438 -7518
rect 3528 -7552 3696 -7518
rect 3786 -7552 3954 -7518
rect 4044 -7552 4212 -7518
rect 2950 -7978 2984 -7602
rect 3208 -7978 3242 -7602
rect 3466 -7978 3500 -7602
rect 3724 -7978 3758 -7602
rect 3982 -7978 4016 -7602
rect 4240 -7978 4274 -7602
rect 3012 -8062 3180 -8028
rect 3270 -8062 3438 -8028
rect 3528 -8062 3696 -8028
rect 3786 -8062 3954 -8028
rect 4044 -8062 4212 -8028
<< metal1 >>
rect 3414 2580 3606 2592
rect 3410 2380 3420 2580
rect 3600 2380 3610 2580
rect 3414 2368 3606 2380
rect 4048 2200 4900 2208
rect 2480 2160 4900 2200
rect 2480 2136 6872 2160
rect -90 1676 -80 2112
rect 2096 1676 2106 2112
rect 2480 2102 2498 2136
rect 2532 2102 2690 2136
rect 2724 2102 2882 2136
rect 2916 2102 3074 2136
rect 3108 2102 3266 2136
rect 3300 2102 3458 2136
rect 3492 2102 3650 2136
rect 3684 2102 3842 2136
rect 3876 2102 4034 2136
rect 4068 2102 4226 2136
rect 4260 2106 6872 2136
rect 4260 2102 5094 2106
rect 2480 2096 5094 2102
rect 4480 2072 5094 2096
rect 5128 2072 5286 2106
rect 5320 2072 5478 2106
rect 5512 2072 5670 2106
rect 5704 2072 5862 2106
rect 5896 2072 6054 2106
rect 6088 2072 6246 2106
rect 6280 2072 6438 2106
rect 6472 2072 6630 2106
rect 6664 2072 6822 2106
rect 6856 2072 6872 2106
rect 4480 2064 6872 2072
rect 2444 2043 2490 2055
rect 2444 1832 2450 2043
rect 2484 1832 2490 2043
rect 2526 1876 2536 2056
rect 2592 1876 2602 2056
rect 2636 2043 2682 2055
rect 2430 1652 2440 1832
rect 2496 1652 2506 1832
rect 2540 1667 2546 1876
rect 2580 1667 2586 1876
rect 2636 1832 2642 2043
rect 2676 1832 2682 2043
rect 2718 1876 2728 2056
rect 2784 1876 2794 2056
rect 2828 2043 2874 2055
rect 2540 1655 2586 1667
rect 2622 1652 2632 1832
rect 2688 1652 2698 1832
rect 2732 1667 2738 1876
rect 2772 1667 2778 1876
rect 2828 1832 2834 2043
rect 2868 1832 2874 2043
rect 2910 1876 2920 2056
rect 2976 1876 2986 2056
rect 3020 2043 3066 2055
rect 2732 1655 2778 1667
rect 2814 1652 2824 1832
rect 2880 1652 2890 1832
rect 2924 1667 2930 1876
rect 2964 1667 2970 1876
rect 3020 1832 3026 2043
rect 3060 1832 3066 2043
rect 3102 1876 3112 2056
rect 3168 1876 3178 2056
rect 3212 2043 3258 2055
rect 2924 1655 2970 1667
rect 3006 1652 3016 1832
rect 3072 1652 3082 1832
rect 3116 1667 3122 1876
rect 3156 1667 3162 1876
rect 3212 1832 3218 2043
rect 3252 1832 3258 2043
rect 3294 1876 3304 2056
rect 3360 1876 3370 2056
rect 3404 2043 3450 2055
rect 3116 1655 3162 1667
rect 3198 1652 3208 1832
rect 3264 1652 3274 1832
rect 3308 1667 3314 1876
rect 3348 1667 3354 1876
rect 3404 1832 3410 2043
rect 3444 1832 3450 2043
rect 3486 1876 3496 2056
rect 3552 1876 3562 2056
rect 3596 2043 3642 2055
rect 3308 1655 3354 1667
rect 3390 1652 3400 1832
rect 3456 1652 3466 1832
rect 3500 1667 3506 1876
rect 3540 1667 3546 1876
rect 3596 1832 3602 2043
rect 3636 1832 3642 2043
rect 3678 1876 3688 2056
rect 3744 1876 3754 2056
rect 3788 2043 3834 2055
rect 3500 1655 3546 1667
rect 3582 1652 3592 1832
rect 3648 1652 3658 1832
rect 3692 1667 3698 1876
rect 3732 1667 3738 1876
rect 3788 1832 3794 2043
rect 3828 1832 3834 2043
rect 3870 1876 3880 2056
rect 3936 1876 3946 2056
rect 3980 2043 4026 2055
rect 3692 1655 3738 1667
rect 3774 1652 3784 1832
rect 3840 1652 3850 1832
rect 3884 1667 3890 1876
rect 3924 1667 3930 1876
rect 3980 1832 3986 2043
rect 4020 1832 4026 2043
rect 4062 1876 4072 2056
rect 4128 1876 4138 2056
rect 4172 2043 4218 2055
rect 3884 1655 3930 1667
rect 3966 1652 3976 1832
rect 4032 1652 4042 1832
rect 4076 1667 4082 1876
rect 4116 1667 4122 1876
rect 4172 1832 4178 2043
rect 4212 1832 4218 2043
rect 4254 1876 4264 2056
rect 4320 1876 4330 2056
rect 4364 2043 4410 2055
rect 4076 1655 4122 1667
rect 4158 1652 4168 1832
rect 4224 1652 4234 1832
rect 4268 1667 4274 1876
rect 4308 1667 4314 1876
rect 4364 1832 4370 2043
rect 4404 1832 4410 2043
rect 4268 1655 4314 1667
rect 4350 1652 4360 1832
rect 4416 1652 4426 1832
rect 4480 1616 4900 2064
rect 4944 2022 4990 2034
rect 4944 1816 4950 2022
rect 4984 1816 4990 2022
rect 5026 1852 5036 2036
rect 5092 1852 5102 2036
rect 5136 2022 5182 2034
rect 4930 1632 4940 1816
rect 4996 1632 5006 1816
rect 5040 1646 5046 1852
rect 5080 1646 5086 1852
rect 5136 1816 5142 2022
rect 5176 1816 5182 2022
rect 5218 1852 5228 2036
rect 5284 1852 5294 2036
rect 5328 2022 5374 2034
rect 5040 1634 5086 1646
rect 5122 1632 5132 1816
rect 5188 1632 5198 1816
rect 5232 1646 5238 1852
rect 5272 1646 5278 1852
rect 5328 1816 5334 2022
rect 5368 1816 5374 2022
rect 5410 1852 5420 2036
rect 5476 1852 5486 2036
rect 5520 2022 5566 2034
rect 5232 1634 5278 1646
rect 5314 1632 5324 1816
rect 5380 1632 5390 1816
rect 5424 1646 5430 1852
rect 5464 1646 5470 1852
rect 5520 1816 5526 2022
rect 5560 1816 5566 2022
rect 5602 1852 5612 2036
rect 5668 1852 5678 2036
rect 5712 2022 5758 2034
rect 5424 1634 5470 1646
rect 5506 1632 5516 1816
rect 5572 1632 5582 1816
rect 5616 1646 5622 1852
rect 5656 1646 5662 1852
rect 5712 1816 5718 2022
rect 5752 1816 5758 2022
rect 5794 1852 5804 2036
rect 5860 1852 5870 2036
rect 5904 2022 5950 2034
rect 5616 1634 5662 1646
rect 5698 1632 5708 1816
rect 5764 1632 5774 1816
rect 5808 1646 5814 1852
rect 5848 1646 5854 1852
rect 5904 1816 5910 2022
rect 5944 1816 5950 2022
rect 5986 1852 5996 2036
rect 6052 1852 6062 2036
rect 6096 2022 6142 2034
rect 5808 1634 5854 1646
rect 5890 1632 5900 1816
rect 5956 1632 5966 1816
rect 6000 1646 6006 1852
rect 6040 1646 6046 1852
rect 6096 1816 6102 2022
rect 6136 1816 6142 2022
rect 6178 1852 6188 2036
rect 6244 1852 6254 2036
rect 6288 2022 6334 2034
rect 6000 1634 6046 1646
rect 6082 1632 6092 1816
rect 6148 1632 6158 1816
rect 6192 1646 6198 1852
rect 6232 1646 6238 1852
rect 6288 1816 6294 2022
rect 6328 1816 6334 2022
rect 6370 1852 6380 2036
rect 6436 1852 6446 2036
rect 6480 2022 6526 2034
rect 6192 1634 6238 1646
rect 6274 1632 6284 1816
rect 6340 1632 6350 1816
rect 6384 1646 6390 1852
rect 6424 1646 6430 1852
rect 6480 1816 6486 2022
rect 6520 1816 6526 2022
rect 6562 1852 6572 2036
rect 6628 1852 6638 2036
rect 6672 2022 6718 2034
rect 6384 1634 6430 1646
rect 6466 1632 6476 1816
rect 6532 1632 6542 1816
rect 6576 1646 6582 1852
rect 6616 1646 6622 1852
rect 6672 1816 6678 2022
rect 6712 1816 6718 2022
rect 6754 1852 6764 2036
rect 6820 1852 6830 2036
rect 6864 2022 6910 2034
rect 6576 1634 6622 1646
rect 6658 1632 6668 1816
rect 6724 1632 6734 1816
rect 6768 1646 6774 1852
rect 6808 1646 6814 1852
rect 6864 1816 6870 2022
rect 6904 1816 6910 2022
rect 6768 1634 6814 1646
rect 6850 1632 6860 1816
rect 6916 1632 6926 1816
rect 2576 1608 4900 1616
rect 2576 1574 2594 1608
rect 2628 1574 2786 1608
rect 2820 1574 2978 1608
rect 3012 1574 3170 1608
rect 3204 1574 3362 1608
rect 3396 1574 3554 1608
rect 3588 1574 3746 1608
rect 3780 1574 3938 1608
rect 3972 1574 4130 1608
rect 4164 1574 4322 1608
rect 4356 1604 4900 1608
rect 4356 1596 6776 1604
rect 4356 1574 4998 1596
rect 2576 1562 4998 1574
rect 5032 1562 5190 1596
rect 5224 1562 5382 1596
rect 5416 1562 5574 1596
rect 5608 1562 5766 1596
rect 5800 1562 5958 1596
rect 5992 1562 6150 1596
rect 6184 1562 6342 1596
rect 6376 1562 6534 1596
rect 6568 1562 6726 1596
rect 6760 1562 6776 1596
rect 2576 1500 6776 1562
rect 2576 1466 2594 1500
rect 2628 1466 2786 1500
rect 2820 1466 2978 1500
rect 3012 1466 3170 1500
rect 3204 1466 3362 1500
rect 3396 1466 3554 1500
rect 3588 1466 3746 1500
rect 3780 1466 3938 1500
rect 3972 1466 4130 1500
rect 4164 1466 4322 1500
rect 4356 1488 6776 1500
rect 4356 1466 4998 1488
rect 2576 1460 4998 1466
rect 4480 1454 4998 1460
rect 5032 1454 5190 1488
rect 5224 1454 5382 1488
rect 5416 1454 5574 1488
rect 5608 1454 5766 1488
rect 5800 1454 5958 1488
rect 5992 1454 6150 1488
rect 6184 1454 6342 1488
rect 6376 1454 6534 1488
rect 6568 1454 6726 1488
rect 6760 1454 6776 1488
rect 4480 1448 6776 1454
rect 2444 1407 2490 1419
rect 2444 1200 2450 1407
rect 2484 1200 2490 1407
rect 2526 1244 2536 1424
rect 2592 1244 2602 1424
rect 2636 1407 2682 1419
rect 2430 1020 2440 1200
rect 2496 1020 2506 1200
rect 2540 1031 2546 1244
rect 2580 1031 2586 1244
rect 2636 1200 2642 1407
rect 2676 1200 2682 1407
rect 2718 1244 2728 1424
rect 2784 1244 2794 1424
rect 2828 1407 2874 1419
rect 2444 1019 2490 1020
rect 2540 1019 2586 1031
rect 2622 1020 2632 1200
rect 2688 1020 2698 1200
rect 2732 1031 2738 1244
rect 2772 1031 2778 1244
rect 2828 1200 2834 1407
rect 2868 1200 2874 1407
rect 2910 1244 2920 1424
rect 2976 1244 2986 1424
rect 3020 1407 3066 1419
rect 2636 1019 2682 1020
rect 2732 1019 2778 1031
rect 2814 1020 2824 1200
rect 2880 1020 2890 1200
rect 2924 1031 2930 1244
rect 2964 1031 2970 1244
rect 3020 1200 3026 1407
rect 3060 1200 3066 1407
rect 3102 1244 3112 1424
rect 3168 1244 3178 1424
rect 3212 1407 3258 1419
rect 2828 1019 2874 1020
rect 2924 1019 2970 1031
rect 3006 1020 3016 1200
rect 3072 1020 3082 1200
rect 3116 1031 3122 1244
rect 3156 1031 3162 1244
rect 3212 1200 3218 1407
rect 3252 1200 3258 1407
rect 3294 1244 3304 1424
rect 3360 1244 3370 1424
rect 3404 1407 3450 1419
rect 3020 1019 3066 1020
rect 3116 1019 3162 1031
rect 3198 1020 3208 1200
rect 3264 1020 3274 1200
rect 3308 1031 3314 1244
rect 3348 1031 3354 1244
rect 3404 1200 3410 1407
rect 3444 1200 3450 1407
rect 3486 1244 3496 1424
rect 3552 1244 3562 1424
rect 3596 1407 3642 1419
rect 3212 1019 3258 1020
rect 3308 1019 3354 1031
rect 3390 1020 3400 1200
rect 3456 1020 3466 1200
rect 3500 1031 3506 1244
rect 3540 1031 3546 1244
rect 3596 1200 3602 1407
rect 3636 1200 3642 1407
rect 3678 1244 3688 1424
rect 3744 1244 3754 1424
rect 3788 1407 3834 1419
rect 3404 1019 3450 1020
rect 3500 1019 3546 1031
rect 3582 1020 3592 1200
rect 3648 1020 3658 1200
rect 3692 1031 3698 1244
rect 3732 1031 3738 1244
rect 3788 1200 3794 1407
rect 3828 1200 3834 1407
rect 3870 1244 3880 1424
rect 3936 1244 3946 1424
rect 3980 1407 4026 1419
rect 3596 1019 3642 1020
rect 3692 1019 3738 1031
rect 3774 1020 3784 1200
rect 3840 1020 3850 1200
rect 3884 1031 3890 1244
rect 3924 1031 3930 1244
rect 3980 1200 3986 1407
rect 4020 1200 4026 1407
rect 4062 1244 4072 1424
rect 4128 1244 4138 1424
rect 4172 1407 4218 1419
rect 3788 1019 3834 1020
rect 3884 1019 3930 1031
rect 3966 1020 3976 1200
rect 4032 1020 4042 1200
rect 4076 1031 4082 1244
rect 4116 1031 4122 1244
rect 4172 1200 4178 1407
rect 4212 1200 4218 1407
rect 4254 1244 4264 1424
rect 4320 1244 4330 1424
rect 4364 1407 4410 1419
rect 3980 1019 4026 1020
rect 4076 1019 4122 1031
rect 4158 1020 4168 1200
rect 4224 1020 4234 1200
rect 4268 1031 4274 1244
rect 4308 1031 4314 1244
rect 4364 1200 4370 1407
rect 4404 1200 4410 1407
rect 4172 1019 4218 1020
rect 4268 1019 4314 1031
rect 4350 1020 4360 1200
rect 4416 1020 4426 1200
rect 4364 1019 4410 1020
rect 4480 984 4900 1448
rect 4944 1404 4990 1416
rect 4944 1200 4950 1404
rect 4984 1200 4990 1404
rect 5026 1236 5036 1420
rect 5092 1236 5102 1420
rect 5136 1404 5182 1416
rect 4930 1016 4940 1200
rect 4996 1016 5006 1200
rect 5040 1028 5046 1236
rect 5080 1028 5086 1236
rect 5136 1200 5142 1404
rect 5176 1200 5182 1404
rect 5218 1236 5228 1420
rect 5284 1236 5294 1420
rect 5328 1404 5374 1416
rect 5040 1016 5086 1028
rect 5122 1016 5132 1200
rect 5188 1016 5198 1200
rect 5232 1028 5238 1236
rect 5272 1028 5278 1236
rect 5328 1200 5334 1404
rect 5368 1200 5374 1404
rect 5410 1236 5420 1420
rect 5476 1236 5486 1420
rect 5520 1404 5566 1416
rect 5232 1016 5278 1028
rect 5314 1016 5324 1200
rect 5380 1016 5390 1200
rect 5424 1028 5430 1236
rect 5464 1028 5470 1236
rect 5520 1200 5526 1404
rect 5560 1200 5566 1404
rect 5602 1236 5612 1420
rect 5668 1236 5678 1420
rect 5712 1404 5758 1416
rect 5424 1016 5470 1028
rect 5506 1016 5516 1200
rect 5572 1016 5582 1200
rect 5616 1028 5622 1236
rect 5656 1028 5662 1236
rect 5712 1200 5718 1404
rect 5752 1200 5758 1404
rect 5794 1236 5804 1420
rect 5860 1236 5870 1420
rect 5904 1404 5950 1416
rect 5616 1016 5662 1028
rect 5698 1016 5708 1200
rect 5764 1016 5774 1200
rect 5808 1028 5814 1236
rect 5848 1028 5854 1236
rect 5904 1200 5910 1404
rect 5944 1200 5950 1404
rect 5986 1236 5996 1420
rect 6052 1236 6062 1420
rect 6096 1404 6142 1416
rect 5808 1016 5854 1028
rect 5890 1016 5900 1200
rect 5956 1016 5966 1200
rect 6000 1028 6006 1236
rect 6040 1028 6046 1236
rect 6096 1200 6102 1404
rect 6136 1200 6142 1404
rect 6178 1236 6188 1420
rect 6244 1236 6254 1420
rect 6288 1404 6334 1416
rect 6000 1016 6046 1028
rect 6082 1016 6092 1200
rect 6148 1016 6158 1200
rect 6192 1028 6198 1236
rect 6232 1028 6238 1236
rect 6288 1200 6294 1404
rect 6328 1200 6334 1404
rect 6370 1236 6380 1420
rect 6436 1236 6446 1420
rect 6480 1404 6526 1416
rect 6192 1016 6238 1028
rect 6274 1016 6284 1200
rect 6340 1016 6350 1200
rect 6384 1028 6390 1236
rect 6424 1028 6430 1236
rect 6480 1200 6486 1404
rect 6520 1200 6526 1404
rect 6562 1236 6572 1420
rect 6628 1236 6638 1420
rect 6672 1404 6718 1416
rect 6384 1016 6430 1028
rect 6466 1016 6476 1200
rect 6532 1016 6542 1200
rect 6576 1028 6582 1236
rect 6616 1028 6622 1236
rect 6672 1200 6678 1404
rect 6712 1200 6718 1404
rect 6754 1236 6764 1420
rect 6820 1236 6830 1420
rect 6864 1404 6910 1416
rect 6576 1016 6622 1028
rect 6658 1016 6668 1200
rect 6724 1016 6734 1200
rect 6768 1028 6774 1236
rect 6808 1028 6814 1236
rect 6864 1200 6870 1404
rect 6904 1200 6910 1404
rect 6768 1016 6814 1028
rect 6850 1016 6860 1200
rect 6916 1016 6926 1200
rect 4480 980 6872 984
rect 2480 978 6872 980
rect 2480 972 5094 978
rect 2480 938 2498 972
rect 2532 938 2690 972
rect 2724 938 2882 972
rect 2916 938 3074 972
rect 3108 938 3266 972
rect 3300 938 3458 972
rect 3492 938 3650 972
rect 3684 938 3842 972
rect 3876 938 4034 972
rect 4068 938 4226 972
rect 4260 944 5094 972
rect 5128 944 5286 978
rect 5320 944 5478 978
rect 5512 944 5670 978
rect 5704 944 5862 978
rect 5896 944 6054 978
rect 6088 944 6246 978
rect 6280 944 6438 978
rect 6472 944 6630 978
rect 6664 944 6822 978
rect 6856 944 6872 978
rect 4260 938 6872 944
rect -92 864 2100 888
rect 2480 876 6872 938
rect -92 861 300 864
rect 1760 861 2100 864
rect -92 464 -58 861
rect 192 464 300 861
rect 1760 464 1832 861
rect 2082 464 2100 861
rect 4480 870 6872 876
rect 4480 836 5094 870
rect 5128 836 5286 870
rect 5320 836 5478 870
rect 5512 836 5670 870
rect 5704 836 5862 870
rect 5896 836 6054 870
rect 6088 836 6246 870
rect 6280 836 6438 870
rect 6472 836 6630 870
rect 6664 836 6822 870
rect 6856 836 6872 870
rect 4480 828 6872 836
rect 4480 752 4900 828
rect 2476 540 4620 588
rect 2476 506 2498 540
rect 2532 506 2690 540
rect 2724 506 2882 540
rect 2916 506 3074 540
rect 3108 506 3266 540
rect 3300 506 3458 540
rect 3492 506 3650 540
rect 3684 506 3842 540
rect 3876 506 4034 540
rect 4068 506 4226 540
rect 4260 506 4620 540
rect 2476 500 4620 506
rect -92 448 300 464
rect 1760 448 2100 464
rect -92 436 2100 448
rect 2444 456 2490 468
rect 2144 420 2388 440
rect 2134 152 2144 420
rect 256 98 2140 152
rect 256 64 274 98
rect 308 64 466 98
rect 500 64 658 98
rect 692 64 850 98
rect 884 64 1042 98
rect 1076 64 1234 98
rect 1268 64 1426 98
rect 1460 64 1618 98
rect 1652 64 1810 98
rect 1844 64 2002 98
rect 2036 64 2140 98
rect 256 56 2140 64
rect 124 14 170 26
rect 124 -196 130 14
rect 164 -196 170 14
rect 206 -152 216 28
rect 272 -152 282 28
rect 316 14 362 26
rect 110 -376 120 -196
rect 176 -376 186 -196
rect 220 -362 226 -152
rect 260 -362 266 -152
rect 316 -196 322 14
rect 356 -196 362 14
rect 398 -152 408 28
rect 464 -152 474 28
rect 508 14 554 26
rect 220 -374 266 -362
rect 302 -376 312 -196
rect 368 -376 378 -196
rect 412 -362 418 -152
rect 452 -362 458 -152
rect 508 -196 514 14
rect 548 -196 554 14
rect 590 -152 600 28
rect 656 -152 666 28
rect 700 14 746 26
rect 412 -374 458 -362
rect 494 -376 504 -196
rect 560 -376 570 -196
rect 604 -362 610 -152
rect 644 -362 650 -152
rect 700 -196 706 14
rect 740 -196 746 14
rect 782 -152 792 28
rect 848 -152 858 28
rect 892 14 938 26
rect 604 -374 650 -362
rect 686 -376 696 -196
rect 752 -376 762 -196
rect 796 -362 802 -152
rect 836 -362 842 -152
rect 892 -196 898 14
rect 932 -196 938 14
rect 974 -152 984 28
rect 1040 -152 1050 28
rect 1084 14 1130 26
rect 796 -374 842 -362
rect 878 -376 888 -196
rect 944 -376 954 -196
rect 988 -362 994 -152
rect 1028 -362 1034 -152
rect 1084 -196 1090 14
rect 1124 -196 1130 14
rect 1166 -152 1176 28
rect 1232 -152 1242 28
rect 1276 14 1322 26
rect 988 -374 1034 -362
rect 1070 -376 1080 -196
rect 1136 -376 1146 -196
rect 1180 -362 1186 -152
rect 1220 -362 1226 -152
rect 1276 -196 1282 14
rect 1316 -196 1322 14
rect 1358 -152 1368 28
rect 1424 -152 1434 28
rect 1468 14 1514 26
rect 1180 -374 1226 -362
rect 1262 -376 1272 -196
rect 1328 -376 1338 -196
rect 1372 -362 1378 -152
rect 1412 -362 1418 -152
rect 1468 -196 1474 14
rect 1508 -196 1514 14
rect 1550 -152 1560 28
rect 1616 -152 1626 28
rect 1660 14 1706 26
rect 1372 -374 1418 -362
rect 1454 -376 1464 -196
rect 1520 -376 1530 -196
rect 1564 -362 1570 -152
rect 1604 -362 1610 -152
rect 1660 -196 1666 14
rect 1700 -196 1706 14
rect 1742 -152 1752 28
rect 1808 -152 1818 28
rect 1852 14 1898 26
rect 1564 -374 1610 -362
rect 1646 -376 1656 -196
rect 1712 -376 1722 -196
rect 1756 -362 1762 -152
rect 1796 -362 1802 -152
rect 1852 -196 1858 14
rect 1892 -196 1898 14
rect 1934 -152 1944 28
rect 2000 -152 2010 28
rect 2044 14 2090 26
rect 1756 -374 1802 -362
rect 1838 -376 1848 -196
rect 1904 -376 1914 -196
rect 1948 -362 1954 -152
rect 1988 -362 1994 -152
rect 2044 -196 2050 14
rect 2084 -196 2090 14
rect 2130 -120 2140 56
rect 2380 -120 2390 420
rect 2444 248 2450 456
rect 2484 248 2490 456
rect 2526 292 2536 472
rect 2592 292 2602 472
rect 2636 456 2682 468
rect 2430 68 2440 248
rect 2496 68 2506 248
rect 2540 80 2546 292
rect 2580 80 2586 292
rect 2636 248 2642 456
rect 2676 248 2682 456
rect 2718 292 2728 472
rect 2784 292 2794 472
rect 2828 456 2874 468
rect 2540 68 2586 80
rect 2622 68 2632 248
rect 2688 68 2698 248
rect 2732 80 2738 292
rect 2772 80 2778 292
rect 2828 248 2834 456
rect 2868 248 2874 456
rect 2910 292 2920 472
rect 2976 292 2986 472
rect 3020 456 3066 468
rect 2732 68 2778 80
rect 2814 68 2824 248
rect 2880 68 2890 248
rect 2924 80 2930 292
rect 2964 80 2970 292
rect 3020 248 3026 456
rect 3060 248 3066 456
rect 3102 292 3112 472
rect 3168 292 3178 472
rect 3212 456 3258 468
rect 2924 68 2970 80
rect 3006 68 3016 248
rect 3072 68 3082 248
rect 3116 80 3122 292
rect 3156 80 3162 292
rect 3212 248 3218 456
rect 3252 248 3258 456
rect 3294 292 3304 472
rect 3360 292 3370 472
rect 3404 456 3450 468
rect 3116 68 3162 80
rect 3198 68 3208 248
rect 3264 68 3274 248
rect 3308 80 3314 292
rect 3348 80 3354 292
rect 3404 248 3410 456
rect 3444 248 3450 456
rect 3486 292 3496 472
rect 3552 292 3562 472
rect 3596 456 3642 468
rect 3308 68 3354 80
rect 3390 68 3400 248
rect 3456 68 3466 248
rect 3500 80 3506 292
rect 3540 80 3546 292
rect 3596 248 3602 456
rect 3636 248 3642 456
rect 3678 292 3688 472
rect 3744 292 3754 472
rect 3788 456 3834 468
rect 3500 68 3546 80
rect 3582 68 3592 248
rect 3648 68 3658 248
rect 3692 80 3698 292
rect 3732 80 3738 292
rect 3788 248 3794 456
rect 3828 248 3834 456
rect 3870 292 3880 472
rect 3936 292 3946 472
rect 3980 456 4026 468
rect 3692 68 3738 80
rect 3774 68 3784 248
rect 3840 68 3850 248
rect 3884 80 3890 292
rect 3924 80 3930 292
rect 3980 248 3986 456
rect 4020 248 4026 456
rect 4062 292 4072 472
rect 4128 292 4138 472
rect 4172 456 4218 468
rect 3884 68 3930 80
rect 3966 68 3976 248
rect 4032 68 4042 248
rect 4076 80 4082 292
rect 4116 80 4122 292
rect 4172 248 4178 456
rect 4212 248 4218 456
rect 4254 292 4264 472
rect 4320 292 4330 472
rect 4364 456 4410 468
rect 4076 68 4122 80
rect 4158 68 4168 248
rect 4224 68 4234 248
rect 4268 80 4274 292
rect 4308 80 4314 292
rect 4364 248 4370 456
rect 4404 248 4410 456
rect 4268 68 4314 80
rect 4350 68 4360 248
rect 4416 68 4424 248
rect 4452 36 4620 500
rect 2576 30 4620 36
rect 2576 -4 2594 30
rect 2628 -4 2786 30
rect 2820 -4 2978 30
rect 3012 -4 3170 30
rect 3204 -4 3362 30
rect 3396 -4 3554 30
rect 3588 -4 3746 30
rect 3780 -4 3938 30
rect 3972 -4 4130 30
rect 4164 -4 4322 30
rect 4356 -4 4620 30
rect 2576 -78 4620 -4
rect 2576 -112 2594 -78
rect 2628 -112 2786 -78
rect 2820 -112 2978 -78
rect 3012 -112 3170 -78
rect 3204 -112 3362 -78
rect 3396 -112 3554 -78
rect 3588 -112 3746 -78
rect 3780 -112 3938 -78
rect 3972 -112 4130 -78
rect 4164 -112 4322 -78
rect 4356 -112 4620 -78
rect 2576 -120 4620 -112
rect 1948 -374 1994 -362
rect 2030 -376 2040 -196
rect 2096 -376 2106 -196
rect 166 -408 224 -406
rect 358 -408 416 -406
rect 550 -408 608 -406
rect 742 -408 800 -406
rect 934 -408 992 -406
rect 1126 -408 1184 -406
rect 1318 -408 1376 -406
rect 1510 -408 1568 -406
rect 1702 -408 1760 -406
rect 1894 -408 1952 -406
rect 2140 -408 2388 -120
rect 2444 -162 2490 -150
rect 2444 -372 2450 -162
rect 2484 -372 2490 -162
rect 2526 -328 2536 -148
rect 2592 -328 2602 -148
rect 2636 -162 2682 -150
rect 160 -412 2388 -408
rect 160 -446 178 -412
rect 212 -446 370 -412
rect 404 -446 562 -412
rect 596 -446 754 -412
rect 788 -446 946 -412
rect 980 -446 1138 -412
rect 1172 -446 1330 -412
rect 1364 -446 1522 -412
rect 1556 -446 1714 -412
rect 1748 -446 1906 -412
rect 1940 -446 2388 -412
rect 160 -520 2388 -446
rect 160 -554 178 -520
rect 212 -554 370 -520
rect 404 -554 562 -520
rect 596 -554 754 -520
rect 788 -554 946 -520
rect 980 -554 1138 -520
rect 1172 -554 1330 -520
rect 1364 -554 1522 -520
rect 1556 -554 1714 -520
rect 1748 -554 1906 -520
rect 1940 -554 2388 -520
rect 2430 -552 2440 -372
rect 2496 -552 2506 -372
rect 2540 -538 2546 -328
rect 2580 -538 2586 -328
rect 2636 -372 2642 -162
rect 2676 -372 2682 -162
rect 2718 -328 2728 -148
rect 2784 -328 2794 -148
rect 2828 -162 2874 -150
rect 2540 -550 2586 -538
rect 2622 -552 2632 -372
rect 2688 -552 2698 -372
rect 2732 -538 2738 -328
rect 2772 -538 2778 -328
rect 2828 -372 2834 -162
rect 2868 -372 2874 -162
rect 2910 -328 2920 -148
rect 2976 -328 2986 -148
rect 3020 -162 3066 -150
rect 2732 -550 2778 -538
rect 2814 -552 2824 -372
rect 2880 -552 2890 -372
rect 2924 -538 2930 -328
rect 2964 -538 2970 -328
rect 3020 -372 3026 -162
rect 3060 -372 3066 -162
rect 3102 -328 3112 -148
rect 3168 -328 3178 -148
rect 3212 -162 3258 -150
rect 2924 -550 2970 -538
rect 3006 -552 3016 -372
rect 3072 -552 3082 -372
rect 3116 -538 3122 -328
rect 3156 -538 3162 -328
rect 3212 -372 3218 -162
rect 3252 -372 3258 -162
rect 3294 -328 3304 -148
rect 3360 -328 3370 -148
rect 3404 -162 3450 -150
rect 3116 -550 3162 -538
rect 3198 -552 3208 -372
rect 3264 -552 3274 -372
rect 3308 -538 3314 -328
rect 3348 -538 3354 -328
rect 3404 -372 3410 -162
rect 3444 -372 3450 -162
rect 3486 -328 3496 -148
rect 3552 -328 3562 -148
rect 3596 -162 3642 -150
rect 3308 -550 3354 -538
rect 3390 -552 3400 -372
rect 3456 -552 3466 -372
rect 3500 -538 3506 -328
rect 3540 -538 3546 -328
rect 3596 -372 3602 -162
rect 3636 -372 3642 -162
rect 3678 -328 3688 -148
rect 3744 -328 3754 -148
rect 3788 -162 3834 -150
rect 3500 -550 3546 -538
rect 3582 -552 3592 -372
rect 3648 -552 3658 -372
rect 3692 -538 3698 -328
rect 3732 -538 3738 -328
rect 3788 -372 3794 -162
rect 3828 -372 3834 -162
rect 3870 -328 3880 -148
rect 3936 -328 3946 -148
rect 3980 -162 4026 -150
rect 3692 -550 3738 -538
rect 3774 -552 3784 -372
rect 3840 -552 3850 -372
rect 3884 -538 3890 -328
rect 3924 -538 3930 -328
rect 3980 -372 3986 -162
rect 4020 -372 4026 -162
rect 4062 -328 4072 -148
rect 4128 -328 4138 -148
rect 4172 -162 4218 -150
rect 3884 -550 3930 -538
rect 3966 -552 3976 -372
rect 4032 -552 4042 -372
rect 4076 -538 4082 -328
rect 4116 -538 4122 -328
rect 4172 -372 4178 -162
rect 4212 -372 4218 -162
rect 4254 -328 4264 -148
rect 4320 -328 4330 -148
rect 4364 -162 4410 -150
rect 4076 -550 4122 -538
rect 4158 -552 4168 -372
rect 4224 -552 4234 -372
rect 4268 -538 4274 -328
rect 4308 -538 4314 -328
rect 4364 -372 4370 -162
rect 4404 -372 4410 -162
rect 4268 -550 4314 -538
rect 4350 -552 4360 -372
rect 4416 -552 4424 -372
rect 160 -560 2388 -554
rect 124 -604 170 -592
rect 124 -812 130 -604
rect 164 -812 170 -604
rect 206 -768 216 -588
rect 272 -768 282 -588
rect 316 -604 362 -592
rect 110 -992 120 -812
rect 176 -992 186 -812
rect 220 -980 226 -768
rect 260 -980 266 -768
rect 316 -812 322 -604
rect 356 -812 362 -604
rect 398 -768 408 -588
rect 464 -768 474 -588
rect 508 -604 554 -592
rect 220 -992 266 -980
rect 302 -992 312 -812
rect 368 -992 378 -812
rect 412 -980 418 -768
rect 452 -980 458 -768
rect 508 -812 514 -604
rect 548 -812 554 -604
rect 590 -768 600 -588
rect 656 -768 666 -588
rect 700 -604 746 -592
rect 412 -992 458 -980
rect 494 -992 504 -812
rect 560 -992 570 -812
rect 604 -980 610 -768
rect 644 -980 650 -768
rect 700 -812 706 -604
rect 740 -812 746 -604
rect 782 -768 792 -588
rect 848 -768 858 -588
rect 892 -604 938 -592
rect 604 -992 650 -980
rect 686 -992 696 -812
rect 752 -992 762 -812
rect 796 -980 802 -768
rect 836 -980 842 -768
rect 892 -812 898 -604
rect 932 -812 938 -604
rect 974 -768 984 -588
rect 1040 -768 1050 -588
rect 1084 -604 1130 -592
rect 796 -992 842 -980
rect 878 -992 888 -812
rect 944 -992 954 -812
rect 988 -980 994 -768
rect 1028 -980 1034 -768
rect 1084 -812 1090 -604
rect 1124 -812 1130 -604
rect 1166 -768 1176 -588
rect 1232 -768 1242 -588
rect 1276 -604 1322 -592
rect 988 -992 1034 -980
rect 1070 -992 1080 -812
rect 1136 -992 1146 -812
rect 1180 -980 1186 -768
rect 1220 -980 1226 -768
rect 1276 -812 1282 -604
rect 1316 -812 1322 -604
rect 1358 -768 1368 -588
rect 1424 -768 1434 -588
rect 1468 -604 1514 -592
rect 1180 -992 1226 -980
rect 1262 -992 1272 -812
rect 1328 -992 1338 -812
rect 1372 -980 1378 -768
rect 1412 -980 1418 -768
rect 1468 -812 1474 -604
rect 1508 -812 1514 -604
rect 1550 -768 1560 -588
rect 1616 -768 1626 -588
rect 1660 -604 1706 -592
rect 1372 -992 1418 -980
rect 1454 -992 1464 -812
rect 1520 -992 1530 -812
rect 1564 -980 1570 -768
rect 1604 -980 1610 -768
rect 1660 -812 1666 -604
rect 1700 -812 1706 -604
rect 1742 -768 1752 -588
rect 1808 -768 1818 -588
rect 1852 -604 1898 -592
rect 1564 -992 1610 -980
rect 1646 -992 1656 -812
rect 1712 -992 1722 -812
rect 1756 -980 1762 -768
rect 1796 -980 1802 -768
rect 1852 -812 1858 -604
rect 1892 -812 1898 -604
rect 1934 -768 1944 -588
rect 2000 -768 2010 -588
rect 2044 -604 2090 -592
rect 1756 -992 1802 -980
rect 1838 -992 1848 -812
rect 1904 -992 1914 -812
rect 1948 -980 1954 -768
rect 1988 -980 1994 -768
rect 2044 -812 2050 -604
rect 2084 -812 2090 -604
rect 2140 -756 2388 -560
rect 4452 -580 4620 -120
rect 2480 -588 4620 -580
rect 2480 -622 2498 -588
rect 2532 -622 2690 -588
rect 2724 -622 2882 -588
rect 2916 -622 3074 -588
rect 3108 -622 3266 -588
rect 3300 -622 3458 -588
rect 3492 -622 3650 -588
rect 3684 -622 3842 -588
rect 3876 -622 4034 -588
rect 4068 -622 4226 -588
rect 4260 -622 4620 -588
rect 2480 -676 4620 -622
rect 3696 -716 3892 -676
rect 4244 -716 4620 -676
rect 1948 -992 1994 -980
rect 2030 -992 2040 -812
rect 2096 -992 2106 -812
rect 2140 -1024 2460 -756
rect 256 -1028 2460 -1024
rect 2688 -1028 2698 -756
rect 3696 -844 3708 -716
rect 256 -1030 2588 -1028
rect 256 -1064 274 -1030
rect 308 -1064 466 -1030
rect 500 -1064 658 -1030
rect 692 -1064 850 -1030
rect 884 -1064 1042 -1030
rect 1076 -1064 1234 -1030
rect 1268 -1064 1426 -1030
rect 1460 -1064 1618 -1030
rect 1652 -1064 1810 -1030
rect 1844 -1064 2002 -1030
rect 2036 -1064 2588 -1030
rect 256 -1138 2588 -1064
rect 256 -1172 274 -1138
rect 308 -1172 466 -1138
rect 500 -1172 658 -1138
rect 692 -1172 850 -1138
rect 884 -1172 1042 -1138
rect 1076 -1172 1234 -1138
rect 1268 -1172 1426 -1138
rect 1460 -1172 1618 -1138
rect 1652 -1172 1810 -1138
rect 1844 -1172 2002 -1138
rect 2036 -1172 2588 -1138
rect 256 -1176 2588 -1172
rect 262 -1178 320 -1176
rect 454 -1178 512 -1176
rect 646 -1178 704 -1176
rect 838 -1178 896 -1176
rect 1030 -1178 1088 -1176
rect 1222 -1178 1280 -1176
rect 1414 -1178 1472 -1176
rect 1606 -1178 1664 -1176
rect 1798 -1178 1856 -1176
rect 1990 -1178 2048 -1176
rect 124 -1222 170 -1210
rect 124 -1432 130 -1222
rect 164 -1432 170 -1222
rect 206 -1388 216 -1208
rect 272 -1388 282 -1208
rect 316 -1222 362 -1210
rect 110 -1612 120 -1432
rect 176 -1612 186 -1432
rect 220 -1598 226 -1388
rect 260 -1598 266 -1388
rect 316 -1432 322 -1222
rect 356 -1432 362 -1222
rect 398 -1388 408 -1208
rect 464 -1388 474 -1208
rect 508 -1222 554 -1210
rect 220 -1610 266 -1598
rect 302 -1612 312 -1432
rect 368 -1612 378 -1432
rect 412 -1598 418 -1388
rect 452 -1598 458 -1388
rect 508 -1432 514 -1222
rect 548 -1432 554 -1222
rect 590 -1388 600 -1208
rect 656 -1388 666 -1208
rect 700 -1222 746 -1210
rect 412 -1610 458 -1598
rect 494 -1612 504 -1432
rect 560 -1612 570 -1432
rect 604 -1598 610 -1388
rect 644 -1598 650 -1388
rect 700 -1432 706 -1222
rect 740 -1432 746 -1222
rect 782 -1388 792 -1208
rect 848 -1388 858 -1208
rect 892 -1222 938 -1210
rect 604 -1610 650 -1598
rect 686 -1612 696 -1432
rect 752 -1612 762 -1432
rect 796 -1598 802 -1388
rect 836 -1598 842 -1388
rect 892 -1432 898 -1222
rect 932 -1432 938 -1222
rect 974 -1388 984 -1208
rect 1040 -1388 1050 -1208
rect 1084 -1222 1130 -1210
rect 796 -1610 842 -1598
rect 878 -1612 888 -1432
rect 944 -1612 954 -1432
rect 988 -1598 994 -1388
rect 1028 -1598 1034 -1388
rect 1084 -1432 1090 -1222
rect 1124 -1432 1130 -1222
rect 1166 -1388 1176 -1208
rect 1232 -1388 1242 -1208
rect 1276 -1222 1322 -1210
rect 988 -1610 1034 -1598
rect 1070 -1612 1080 -1432
rect 1136 -1612 1146 -1432
rect 1180 -1598 1186 -1388
rect 1220 -1598 1226 -1388
rect 1276 -1432 1282 -1222
rect 1316 -1432 1322 -1222
rect 1358 -1388 1368 -1208
rect 1424 -1388 1434 -1208
rect 1468 -1222 1514 -1210
rect 1180 -1610 1226 -1598
rect 1262 -1612 1272 -1432
rect 1328 -1612 1338 -1432
rect 1372 -1598 1378 -1388
rect 1412 -1598 1418 -1388
rect 1468 -1432 1474 -1222
rect 1508 -1432 1514 -1222
rect 1550 -1388 1560 -1208
rect 1616 -1388 1626 -1208
rect 1660 -1222 1706 -1210
rect 1372 -1610 1418 -1598
rect 1454 -1612 1464 -1432
rect 1520 -1612 1530 -1432
rect 1564 -1598 1570 -1388
rect 1604 -1598 1610 -1388
rect 1660 -1432 1666 -1222
rect 1700 -1432 1706 -1222
rect 1742 -1388 1752 -1208
rect 1808 -1388 1818 -1208
rect 1852 -1222 1898 -1210
rect 1564 -1610 1610 -1598
rect 1646 -1612 1656 -1432
rect 1712 -1612 1722 -1432
rect 1756 -1598 1762 -1388
rect 1796 -1598 1802 -1388
rect 1852 -1432 1858 -1222
rect 1892 -1432 1898 -1222
rect 1934 -1388 1944 -1208
rect 2000 -1388 2010 -1208
rect 2044 -1222 2090 -1210
rect 1756 -1610 1802 -1598
rect 1838 -1612 1848 -1432
rect 1904 -1612 1914 -1432
rect 1948 -1598 1954 -1388
rect 1988 -1598 1994 -1388
rect 2044 -1432 2050 -1222
rect 2084 -1432 2090 -1222
rect 1948 -1610 1994 -1598
rect 2030 -1612 2040 -1432
rect 2096 -1612 2106 -1432
rect 2140 -1640 2588 -1176
rect 3698 -1228 3708 -844
rect 4400 -836 4620 -716
rect 4648 368 4900 752
rect 4944 786 4990 798
rect 4944 580 4950 786
rect 4984 580 4990 786
rect 5026 616 5036 800
rect 5092 616 5102 800
rect 5136 786 5182 798
rect 4930 396 4940 580
rect 4996 396 5006 580
rect 5040 410 5046 616
rect 5080 410 5086 616
rect 5136 580 5142 786
rect 5176 580 5182 786
rect 5218 616 5228 800
rect 5284 616 5294 800
rect 5328 786 5374 798
rect 5040 398 5086 410
rect 5122 396 5132 580
rect 5188 396 5198 580
rect 5232 410 5238 616
rect 5272 410 5278 616
rect 5328 580 5334 786
rect 5368 580 5374 786
rect 5410 616 5420 800
rect 5476 616 5486 800
rect 5520 786 5566 798
rect 5232 398 5278 410
rect 5314 396 5324 580
rect 5380 396 5390 580
rect 5424 410 5430 616
rect 5464 410 5470 616
rect 5520 580 5526 786
rect 5560 580 5566 786
rect 5602 616 5612 800
rect 5668 616 5678 800
rect 5712 786 5758 798
rect 5424 398 5470 410
rect 5506 396 5516 580
rect 5572 396 5582 580
rect 5616 410 5622 616
rect 5656 410 5662 616
rect 5712 580 5718 786
rect 5752 580 5758 786
rect 5794 616 5804 800
rect 5860 616 5870 800
rect 5904 786 5950 798
rect 5616 398 5662 410
rect 5698 396 5708 580
rect 5764 396 5774 580
rect 5808 410 5814 616
rect 5848 410 5854 616
rect 5904 580 5910 786
rect 5944 580 5950 786
rect 5986 616 5996 800
rect 6052 616 6062 800
rect 6096 786 6142 798
rect 5808 398 5854 410
rect 5890 396 5900 580
rect 5956 396 5966 580
rect 6000 410 6006 616
rect 6040 410 6046 616
rect 6096 580 6102 786
rect 6136 580 6142 786
rect 6178 616 6188 800
rect 6244 616 6254 800
rect 6288 786 6334 798
rect 6000 398 6046 410
rect 6082 396 6092 580
rect 6148 396 6158 580
rect 6192 410 6198 616
rect 6232 410 6238 616
rect 6288 580 6294 786
rect 6328 580 6334 786
rect 6370 616 6380 800
rect 6436 616 6446 800
rect 6480 786 6526 798
rect 6192 398 6238 410
rect 6274 396 6284 580
rect 6340 396 6350 580
rect 6384 410 6390 616
rect 6424 410 6430 616
rect 6480 580 6486 786
rect 6520 580 6526 786
rect 6562 616 6572 800
rect 6628 616 6638 800
rect 6672 786 6718 798
rect 6384 398 6430 410
rect 6466 396 6476 580
rect 6532 396 6542 580
rect 6576 410 6582 616
rect 6616 410 6622 616
rect 6672 580 6678 786
rect 6712 580 6718 786
rect 6754 616 6764 800
rect 6820 616 6830 800
rect 6864 786 6910 798
rect 6576 398 6622 410
rect 6658 396 6668 580
rect 6724 396 6734 580
rect 6768 410 6774 616
rect 6808 410 6814 616
rect 6864 580 6870 786
rect 6904 580 6910 786
rect 6768 398 6814 410
rect 6850 396 6860 580
rect 6916 396 6926 580
rect 4648 360 6776 368
rect 4648 326 4998 360
rect 5032 326 5190 360
rect 5224 326 5382 360
rect 5416 326 5574 360
rect 5608 326 5766 360
rect 5800 326 5958 360
rect 5992 326 6150 360
rect 6184 326 6342 360
rect 6376 326 6534 360
rect 6568 326 6726 360
rect 6760 326 6776 360
rect 4648 252 6776 326
rect 4648 218 4998 252
rect 5032 218 5190 252
rect 5224 218 5382 252
rect 5416 218 5574 252
rect 5608 218 5766 252
rect 5800 218 5958 252
rect 5992 218 6150 252
rect 6184 218 6342 252
rect 6376 218 6534 252
rect 6568 218 6726 252
rect 6760 218 6776 252
rect 4648 212 6776 218
rect 4648 -252 4900 212
rect 4944 168 4990 180
rect 4944 -36 4950 168
rect 4984 -36 4990 168
rect 5026 0 5036 184
rect 5092 0 5102 184
rect 5136 168 5182 180
rect 4930 -220 4940 -36
rect 4996 -220 5006 -36
rect 5040 -208 5046 0
rect 5080 -208 5086 0
rect 5136 -36 5142 168
rect 5176 -36 5182 168
rect 5218 0 5228 184
rect 5284 0 5294 184
rect 5328 168 5374 180
rect 5040 -220 5086 -208
rect 5122 -220 5132 -36
rect 5188 -220 5198 -36
rect 5232 -208 5238 0
rect 5272 -208 5278 0
rect 5328 -36 5334 168
rect 5368 -36 5374 168
rect 5410 0 5420 184
rect 5476 0 5486 184
rect 5520 168 5566 180
rect 5232 -220 5278 -208
rect 5314 -220 5324 -36
rect 5380 -220 5390 -36
rect 5424 -208 5430 0
rect 5464 -208 5470 0
rect 5520 -36 5526 168
rect 5560 -36 5566 168
rect 5602 0 5612 184
rect 5668 0 5678 184
rect 5712 168 5758 180
rect 5424 -220 5470 -208
rect 5506 -220 5516 -36
rect 5572 -220 5582 -36
rect 5616 -208 5622 0
rect 5656 -208 5662 0
rect 5712 -36 5718 168
rect 5752 -36 5758 168
rect 5794 0 5804 184
rect 5860 0 5870 184
rect 5904 168 5950 180
rect 5616 -220 5662 -208
rect 5698 -220 5708 -36
rect 5764 -220 5774 -36
rect 5808 -208 5814 0
rect 5848 -208 5854 0
rect 5904 -36 5910 168
rect 5944 -36 5950 168
rect 5986 0 5996 184
rect 6052 0 6062 184
rect 6096 168 6142 180
rect 5808 -220 5854 -208
rect 5890 -220 5900 -36
rect 5956 -220 5966 -36
rect 6000 -208 6006 0
rect 6040 -208 6046 0
rect 6096 -36 6102 168
rect 6136 -36 6142 168
rect 6178 0 6188 184
rect 6244 0 6254 184
rect 6288 168 6334 180
rect 6000 -220 6046 -208
rect 6082 -220 6092 -36
rect 6148 -220 6158 -36
rect 6192 -208 6198 0
rect 6232 -208 6238 0
rect 6288 -36 6294 168
rect 6328 -36 6334 168
rect 6370 0 6380 184
rect 6436 0 6446 184
rect 6480 168 6526 180
rect 6192 -220 6238 -208
rect 6274 -220 6284 -36
rect 6340 -220 6350 -36
rect 6384 -208 6390 0
rect 6424 -208 6430 0
rect 6480 -36 6486 168
rect 6520 -36 6526 168
rect 6562 0 6572 184
rect 6628 0 6638 184
rect 6672 168 6718 180
rect 6384 -220 6430 -208
rect 6466 -220 6476 -36
rect 6532 -220 6542 -36
rect 6576 -208 6582 0
rect 6616 -208 6622 0
rect 6672 -36 6678 168
rect 6712 -36 6718 168
rect 6754 0 6764 184
rect 6820 0 6830 184
rect 6864 168 6910 180
rect 6576 -220 6622 -208
rect 6658 -220 6668 -36
rect 6724 -220 6734 -36
rect 6768 -208 6774 0
rect 6808 -208 6814 0
rect 6864 -36 6870 168
rect 6904 -36 6910 168
rect 6768 -220 6814 -208
rect 6850 -220 6860 -36
rect 6916 -220 6926 -36
rect 4648 -258 6872 -252
rect 4648 -292 5094 -258
rect 5128 -292 5286 -258
rect 5320 -292 5478 -258
rect 5512 -292 5670 -258
rect 5704 -292 5862 -258
rect 5896 -292 6054 -258
rect 6088 -292 6246 -258
rect 6280 -292 6438 -258
rect 6472 -292 6630 -258
rect 6664 -292 6822 -258
rect 6856 -292 6872 -258
rect 4648 -366 6872 -292
rect 4648 -400 5094 -366
rect 5128 -400 5286 -366
rect 5320 -400 5478 -366
rect 5512 -400 5670 -366
rect 5704 -400 5862 -366
rect 5896 -400 6054 -366
rect 6088 -400 6246 -366
rect 6280 -400 6438 -366
rect 6472 -400 6630 -366
rect 6664 -400 6822 -366
rect 6856 -400 6872 -366
rect 4648 -408 6872 -400
rect 4400 -1228 4410 -836
rect 4648 -868 4900 -408
rect 4944 -450 4990 -438
rect 4944 -656 4950 -450
rect 4984 -656 4990 -450
rect 5026 -620 5036 -436
rect 5092 -620 5102 -436
rect 5136 -450 5182 -438
rect 4930 -840 4940 -656
rect 4996 -840 5006 -656
rect 5040 -826 5046 -620
rect 5080 -826 5086 -620
rect 5136 -656 5142 -450
rect 5176 -656 5182 -450
rect 5218 -620 5228 -436
rect 5284 -620 5294 -436
rect 5328 -450 5374 -438
rect 5040 -838 5086 -826
rect 5122 -840 5132 -656
rect 5188 -840 5198 -656
rect 5232 -826 5238 -620
rect 5272 -826 5278 -620
rect 5328 -656 5334 -450
rect 5368 -656 5374 -450
rect 5410 -620 5420 -436
rect 5476 -620 5486 -436
rect 5520 -450 5566 -438
rect 5232 -838 5278 -826
rect 5314 -840 5324 -656
rect 5380 -840 5390 -656
rect 5424 -826 5430 -620
rect 5464 -826 5470 -620
rect 5520 -656 5526 -450
rect 5560 -656 5566 -450
rect 5602 -620 5612 -436
rect 5668 -620 5678 -436
rect 5712 -450 5758 -438
rect 5424 -838 5470 -826
rect 5506 -840 5516 -656
rect 5572 -840 5582 -656
rect 5616 -826 5622 -620
rect 5656 -826 5662 -620
rect 5712 -656 5718 -450
rect 5752 -656 5758 -450
rect 5794 -620 5804 -436
rect 5860 -620 5870 -436
rect 5904 -450 5950 -438
rect 5616 -838 5662 -826
rect 5698 -840 5708 -656
rect 5764 -840 5774 -656
rect 5808 -826 5814 -620
rect 5848 -826 5854 -620
rect 5904 -656 5910 -450
rect 5944 -656 5950 -450
rect 5986 -620 5996 -436
rect 6052 -620 6062 -436
rect 6096 -450 6142 -438
rect 5808 -838 5854 -826
rect 5890 -840 5900 -656
rect 5956 -840 5966 -656
rect 6000 -826 6006 -620
rect 6040 -826 6046 -620
rect 6096 -656 6102 -450
rect 6136 -656 6142 -450
rect 6178 -620 6188 -436
rect 6244 -620 6254 -436
rect 6288 -450 6334 -438
rect 6000 -838 6046 -826
rect 6082 -840 6092 -656
rect 6148 -840 6158 -656
rect 6192 -826 6198 -620
rect 6232 -826 6238 -620
rect 6288 -656 6294 -450
rect 6328 -656 6334 -450
rect 6370 -620 6380 -436
rect 6436 -620 6446 -436
rect 6480 -450 6526 -438
rect 6192 -838 6238 -826
rect 6274 -840 6284 -656
rect 6340 -840 6350 -656
rect 6384 -826 6390 -620
rect 6424 -826 6430 -620
rect 6480 -656 6486 -450
rect 6520 -656 6526 -450
rect 6562 -620 6572 -436
rect 6628 -620 6638 -436
rect 6672 -450 6718 -438
rect 6384 -838 6430 -826
rect 6466 -840 6476 -656
rect 6532 -840 6542 -656
rect 6576 -826 6582 -620
rect 6616 -826 6622 -620
rect 6672 -656 6678 -450
rect 6712 -656 6718 -450
rect 6754 -620 6764 -436
rect 6820 -620 6830 -436
rect 6864 -450 6910 -438
rect 6576 -838 6622 -826
rect 6658 -840 6668 -656
rect 6724 -840 6734 -656
rect 6768 -826 6774 -620
rect 6808 -826 6814 -620
rect 6864 -656 6870 -450
rect 6904 -656 6910 -450
rect 6768 -838 6814 -826
rect 6850 -840 6860 -656
rect 6916 -840 6926 -656
rect 4480 -876 6776 -868
rect 4480 -910 4998 -876
rect 5032 -910 5190 -876
rect 5224 -910 5382 -876
rect 5416 -910 5574 -876
rect 5608 -910 5766 -876
rect 5800 -910 5958 -876
rect 5992 -910 6150 -876
rect 6184 -910 6342 -876
rect 6376 -910 6534 -876
rect 6568 -910 6726 -876
rect 6760 -910 6776 -876
rect 4480 -984 6776 -910
rect 4480 -1018 4998 -984
rect 5032 -1018 5190 -984
rect 5224 -1018 5382 -984
rect 5416 -1018 5574 -984
rect 5608 -1018 5766 -984
rect 5800 -1018 5958 -984
rect 5992 -1018 6150 -984
rect 6184 -1018 6342 -984
rect 6376 -1018 6534 -984
rect 6568 -1018 6726 -984
rect 6760 -1018 6776 -984
rect 4480 -1024 6776 -1018
rect 4480 -1300 4900 -1024
rect 4944 -1068 4990 -1056
rect 4944 -1272 4950 -1068
rect 4984 -1272 4990 -1068
rect 5026 -1236 5036 -1052
rect 5092 -1236 5102 -1052
rect 5136 -1068 5182 -1056
rect 4314 -1628 4324 -1300
rect 4852 -1488 4900 -1300
rect 4930 -1456 4940 -1272
rect 4996 -1456 5006 -1272
rect 5040 -1444 5046 -1236
rect 5080 -1444 5086 -1236
rect 5136 -1272 5142 -1068
rect 5176 -1272 5182 -1068
rect 5218 -1236 5228 -1052
rect 5284 -1236 5294 -1052
rect 5328 -1068 5374 -1056
rect 5040 -1456 5086 -1444
rect 5122 -1456 5132 -1272
rect 5188 -1456 5198 -1272
rect 5232 -1444 5238 -1236
rect 5272 -1444 5278 -1236
rect 5328 -1272 5334 -1068
rect 5368 -1272 5374 -1068
rect 5410 -1236 5420 -1052
rect 5476 -1236 5486 -1052
rect 5520 -1068 5566 -1056
rect 5232 -1456 5278 -1444
rect 5314 -1456 5324 -1272
rect 5380 -1456 5390 -1272
rect 5424 -1444 5430 -1236
rect 5464 -1444 5470 -1236
rect 5520 -1272 5526 -1068
rect 5560 -1272 5566 -1068
rect 5602 -1236 5612 -1052
rect 5668 -1236 5678 -1052
rect 5712 -1068 5758 -1056
rect 5424 -1456 5470 -1444
rect 5506 -1456 5516 -1272
rect 5572 -1456 5582 -1272
rect 5616 -1444 5622 -1236
rect 5656 -1444 5662 -1236
rect 5712 -1272 5718 -1068
rect 5752 -1272 5758 -1068
rect 5794 -1236 5804 -1052
rect 5860 -1236 5870 -1052
rect 5904 -1068 5950 -1056
rect 5616 -1456 5662 -1444
rect 5698 -1456 5708 -1272
rect 5764 -1456 5774 -1272
rect 5808 -1444 5814 -1236
rect 5848 -1444 5854 -1236
rect 5904 -1272 5910 -1068
rect 5944 -1272 5950 -1068
rect 5986 -1236 5996 -1052
rect 6052 -1236 6062 -1052
rect 6096 -1068 6142 -1056
rect 5808 -1456 5854 -1444
rect 5890 -1456 5900 -1272
rect 5956 -1456 5966 -1272
rect 6000 -1444 6006 -1236
rect 6040 -1444 6046 -1236
rect 6096 -1272 6102 -1068
rect 6136 -1272 6142 -1068
rect 6178 -1236 6188 -1052
rect 6244 -1236 6254 -1052
rect 6288 -1068 6334 -1056
rect 6000 -1456 6046 -1444
rect 6082 -1456 6092 -1272
rect 6148 -1456 6158 -1272
rect 6192 -1444 6198 -1236
rect 6232 -1444 6238 -1236
rect 6288 -1272 6294 -1068
rect 6328 -1272 6334 -1068
rect 6370 -1236 6380 -1052
rect 6436 -1236 6446 -1052
rect 6480 -1068 6526 -1056
rect 6192 -1456 6238 -1444
rect 6274 -1456 6284 -1272
rect 6340 -1456 6350 -1272
rect 6384 -1444 6390 -1236
rect 6424 -1444 6430 -1236
rect 6480 -1272 6486 -1068
rect 6520 -1272 6526 -1068
rect 6562 -1236 6572 -1052
rect 6628 -1236 6638 -1052
rect 6672 -1068 6718 -1056
rect 6384 -1456 6430 -1444
rect 6466 -1456 6476 -1272
rect 6532 -1456 6542 -1272
rect 6576 -1444 6582 -1236
rect 6616 -1444 6622 -1236
rect 6672 -1272 6678 -1068
rect 6712 -1272 6718 -1068
rect 6754 -1236 6764 -1052
rect 6820 -1236 6830 -1052
rect 6864 -1068 6910 -1056
rect 6576 -1456 6622 -1444
rect 6658 -1456 6668 -1272
rect 6724 -1456 6734 -1272
rect 6768 -1444 6774 -1236
rect 6808 -1444 6814 -1236
rect 6864 -1272 6870 -1068
rect 6904 -1272 6910 -1068
rect 6768 -1456 6814 -1444
rect 6850 -1456 6860 -1272
rect 6916 -1456 6926 -1272
rect 4852 -1494 6872 -1488
rect 4852 -1528 5094 -1494
rect 5128 -1528 5286 -1494
rect 5320 -1528 5478 -1494
rect 5512 -1528 5670 -1494
rect 5704 -1528 5862 -1494
rect 5896 -1528 6054 -1494
rect 6088 -1528 6246 -1494
rect 6280 -1528 6438 -1494
rect 6472 -1528 6630 -1494
rect 6664 -1528 6822 -1494
rect 6856 -1528 6872 -1494
rect 4852 -1602 6872 -1528
rect 4852 -1628 5094 -1602
rect 144 -1648 2588 -1640
rect 144 -1682 178 -1648
rect 212 -1682 370 -1648
rect 404 -1682 562 -1648
rect 596 -1682 754 -1648
rect 788 -1682 946 -1648
rect 980 -1682 1138 -1648
rect 1172 -1682 1330 -1648
rect 1364 -1682 1522 -1648
rect 1556 -1682 1714 -1648
rect 1748 -1682 1906 -1648
rect 1940 -1682 2588 -1648
rect 144 -1736 2588 -1682
rect 4480 -1636 5094 -1628
rect 5128 -1636 5286 -1602
rect 5320 -1636 5478 -1602
rect 5512 -1636 5670 -1602
rect 5704 -1636 5862 -1602
rect 5896 -1636 6054 -1602
rect 6088 -1636 6246 -1602
rect 6280 -1636 6438 -1602
rect 6472 -1636 6630 -1602
rect 6664 -1636 6822 -1602
rect 6856 -1636 6872 -1602
rect 4480 -1644 6872 -1636
rect 4480 -1756 4900 -1644
rect 4274 -2072 4284 -1756
rect 4780 -2072 4900 -1756
rect 4944 -1686 4990 -1674
rect 4944 -1892 4950 -1686
rect 4984 -1892 4990 -1686
rect 5026 -1856 5036 -1672
rect 5092 -1856 5102 -1672
rect 5136 -1686 5182 -1674
rect 4480 -2104 4900 -2072
rect 4930 -2076 4940 -1892
rect 4996 -2076 5006 -1892
rect 5040 -2062 5046 -1856
rect 5080 -2062 5086 -1856
rect 5136 -1892 5142 -1686
rect 5176 -1892 5182 -1686
rect 5218 -1856 5228 -1672
rect 5284 -1856 5294 -1672
rect 5328 -1686 5374 -1674
rect 5040 -2074 5086 -2062
rect 5122 -2076 5132 -1892
rect 5188 -2076 5198 -1892
rect 5232 -2062 5238 -1856
rect 5272 -2062 5278 -1856
rect 5328 -1892 5334 -1686
rect 5368 -1892 5374 -1686
rect 5410 -1856 5420 -1672
rect 5476 -1856 5486 -1672
rect 5520 -1686 5566 -1674
rect 5232 -2074 5278 -2062
rect 5314 -2076 5324 -1892
rect 5380 -2076 5390 -1892
rect 5424 -2062 5430 -1856
rect 5464 -2062 5470 -1856
rect 5520 -1892 5526 -1686
rect 5560 -1892 5566 -1686
rect 5602 -1856 5612 -1672
rect 5668 -1856 5678 -1672
rect 5712 -1686 5758 -1674
rect 5424 -2074 5470 -2062
rect 5506 -2076 5516 -1892
rect 5572 -2076 5582 -1892
rect 5616 -2062 5622 -1856
rect 5656 -2062 5662 -1856
rect 5712 -1892 5718 -1686
rect 5752 -1892 5758 -1686
rect 5794 -1856 5804 -1672
rect 5860 -1856 5870 -1672
rect 5904 -1686 5950 -1674
rect 5616 -2074 5662 -2062
rect 5698 -2076 5708 -1892
rect 5764 -2076 5774 -1892
rect 5808 -2062 5814 -1856
rect 5848 -2062 5854 -1856
rect 5904 -1892 5910 -1686
rect 5944 -1892 5950 -1686
rect 5986 -1856 5996 -1672
rect 6052 -1856 6062 -1672
rect 6096 -1686 6142 -1674
rect 5808 -2074 5854 -2062
rect 5890 -2076 5900 -1892
rect 5956 -2076 5966 -1892
rect 6000 -2062 6006 -1856
rect 6040 -2062 6046 -1856
rect 6096 -1892 6102 -1686
rect 6136 -1892 6142 -1686
rect 6178 -1856 6188 -1672
rect 6244 -1856 6254 -1672
rect 6288 -1686 6334 -1674
rect 6000 -2074 6046 -2062
rect 6082 -2076 6092 -1892
rect 6148 -2076 6158 -1892
rect 6192 -2062 6198 -1856
rect 6232 -2062 6238 -1856
rect 6288 -1892 6294 -1686
rect 6328 -1892 6334 -1686
rect 6370 -1856 6380 -1672
rect 6436 -1856 6446 -1672
rect 6480 -1686 6526 -1674
rect 6192 -2074 6238 -2062
rect 6274 -2076 6284 -1892
rect 6340 -2076 6350 -1892
rect 6384 -2062 6390 -1856
rect 6424 -2062 6430 -1856
rect 6480 -1892 6486 -1686
rect 6520 -1892 6526 -1686
rect 6562 -1856 6572 -1672
rect 6628 -1856 6638 -1672
rect 6672 -1686 6718 -1674
rect 6384 -2074 6430 -2062
rect 6466 -2076 6476 -1892
rect 6532 -2076 6542 -1892
rect 6576 -2062 6582 -1856
rect 6616 -2062 6622 -1856
rect 6672 -1892 6678 -1686
rect 6712 -1892 6718 -1686
rect 6754 -1856 6764 -1672
rect 6820 -1856 6830 -1672
rect 6864 -1686 6910 -1674
rect 6576 -2074 6622 -2062
rect 6658 -2076 6668 -1892
rect 6724 -2076 6734 -1892
rect 6768 -2062 6774 -1856
rect 6808 -2062 6814 -1856
rect 6864 -1892 6870 -1686
rect 6904 -1892 6910 -1686
rect 6768 -2074 6814 -2062
rect 6850 -2076 6860 -1892
rect 6916 -2076 6926 -1892
rect 4480 -2112 6776 -2104
rect 4480 -2146 4998 -2112
rect 5032 -2146 5190 -2112
rect 5224 -2146 5382 -2112
rect 5416 -2146 5574 -2112
rect 5608 -2146 5766 -2112
rect 5800 -2146 5958 -2112
rect 5992 -2146 6150 -2112
rect 6184 -2146 6342 -2112
rect 6376 -2146 6534 -2112
rect 6568 -2146 6726 -2112
rect 6760 -2146 6776 -2112
rect 4480 -2148 6776 -2146
rect -3072 -2240 3988 -2176
rect -3072 -2244 4092 -2240
rect -3072 -2282 4228 -2244
rect -3072 -2316 -2306 -2282
rect -2272 -2316 -2114 -2282
rect -2080 -2316 -1922 -2282
rect -1888 -2316 -1730 -2282
rect -1696 -2316 -1538 -2282
rect -1504 -2316 -506 -2282
rect -472 -2316 -314 -2282
rect -280 -2316 -122 -2282
rect -88 -2316 70 -2282
rect 104 -2316 262 -2282
rect 296 -2316 1294 -2282
rect 1328 -2316 1486 -2282
rect 1520 -2316 1678 -2282
rect 1712 -2316 1870 -2282
rect 1904 -2316 2062 -2282
rect 2096 -2316 3094 -2282
rect 3128 -2316 3286 -2282
rect 3320 -2316 3478 -2282
rect 3512 -2316 3670 -2282
rect 3704 -2316 3862 -2282
rect 3896 -2316 4228 -2282
rect -3072 -2320 4228 -2316
rect -3072 -2792 -2592 -2320
rect -2318 -2322 -2260 -2320
rect -2126 -2322 -2068 -2320
rect -1934 -2322 -1876 -2320
rect -1742 -2322 -1684 -2320
rect -1550 -2322 -1492 -2320
rect -2456 -2366 -2410 -2354
rect -2456 -2576 -2450 -2366
rect -2416 -2576 -2410 -2366
rect -2374 -2532 -2364 -2352
rect -2312 -2532 -2302 -2352
rect -2264 -2366 -2218 -2354
rect -2470 -2756 -2460 -2576
rect -2408 -2756 -2398 -2576
rect -2360 -2742 -2354 -2532
rect -2320 -2742 -2314 -2532
rect -2264 -2576 -2258 -2366
rect -2224 -2576 -2218 -2366
rect -2182 -2532 -2172 -2352
rect -2120 -2532 -2110 -2352
rect -2072 -2366 -2026 -2354
rect -2360 -2754 -2314 -2742
rect -2278 -2756 -2268 -2576
rect -2216 -2756 -2206 -2576
rect -2168 -2742 -2162 -2532
rect -2128 -2742 -2122 -2532
rect -2072 -2576 -2066 -2366
rect -2032 -2576 -2026 -2366
rect -1990 -2532 -1980 -2352
rect -1928 -2532 -1918 -2352
rect -1880 -2366 -1834 -2354
rect -2168 -2754 -2122 -2742
rect -2086 -2756 -2076 -2576
rect -2024 -2756 -2014 -2576
rect -1976 -2742 -1970 -2532
rect -1936 -2742 -1930 -2532
rect -1880 -2576 -1874 -2366
rect -1840 -2576 -1834 -2366
rect -1798 -2532 -1788 -2352
rect -1736 -2532 -1726 -2352
rect -1688 -2366 -1642 -2354
rect -1976 -2754 -1930 -2742
rect -1894 -2756 -1884 -2576
rect -1832 -2756 -1822 -2576
rect -1784 -2742 -1778 -2532
rect -1744 -2742 -1738 -2532
rect -1688 -2576 -1682 -2366
rect -1648 -2576 -1642 -2366
rect -1606 -2532 -1596 -2352
rect -1544 -2532 -1534 -2352
rect -1496 -2366 -1450 -2354
rect -1784 -2754 -1738 -2742
rect -1702 -2756 -1692 -2576
rect -1640 -2756 -1630 -2576
rect -1592 -2742 -1586 -2532
rect -1552 -2742 -1546 -2532
rect -1496 -2576 -1490 -2366
rect -1456 -2576 -1450 -2366
rect -1592 -2754 -1546 -2742
rect -1510 -2756 -1500 -2576
rect -1448 -2756 -1438 -2576
rect -2414 -2792 -2356 -2786
rect -2222 -2792 -2164 -2786
rect -2030 -2792 -1972 -2786
rect -1838 -2792 -1780 -2786
rect -1646 -2792 -1588 -2786
rect -1408 -2792 -1176 -2320
rect -518 -2322 -460 -2320
rect -326 -2322 -268 -2320
rect -134 -2322 -76 -2320
rect 58 -2322 116 -2320
rect 250 -2322 308 -2320
rect -656 -2366 -610 -2354
rect -656 -2576 -650 -2366
rect -616 -2576 -610 -2366
rect -574 -2532 -564 -2352
rect -512 -2532 -502 -2352
rect -464 -2366 -418 -2354
rect -670 -2756 -660 -2576
rect -608 -2756 -598 -2576
rect -560 -2742 -554 -2532
rect -520 -2742 -514 -2532
rect -464 -2576 -458 -2366
rect -424 -2576 -418 -2366
rect -382 -2532 -372 -2352
rect -320 -2532 -310 -2352
rect -272 -2366 -226 -2354
rect -560 -2754 -514 -2742
rect -478 -2756 -468 -2576
rect -416 -2756 -406 -2576
rect -368 -2742 -362 -2532
rect -328 -2742 -322 -2532
rect -272 -2576 -266 -2366
rect -232 -2576 -226 -2366
rect -190 -2532 -180 -2352
rect -128 -2532 -118 -2352
rect -80 -2366 -34 -2354
rect -368 -2754 -322 -2742
rect -286 -2756 -276 -2576
rect -224 -2756 -214 -2576
rect -176 -2742 -170 -2532
rect -136 -2742 -130 -2532
rect -80 -2576 -74 -2366
rect -40 -2576 -34 -2366
rect 2 -2532 12 -2352
rect 64 -2532 74 -2352
rect 112 -2366 158 -2354
rect -176 -2754 -130 -2742
rect -94 -2756 -84 -2576
rect -32 -2756 -22 -2576
rect 16 -2742 22 -2532
rect 56 -2742 62 -2532
rect 112 -2576 118 -2366
rect 152 -2576 158 -2366
rect 194 -2532 204 -2352
rect 256 -2532 266 -2352
rect 304 -2366 350 -2354
rect 16 -2754 62 -2742
rect 98 -2756 108 -2576
rect 160 -2756 170 -2576
rect 208 -2742 214 -2532
rect 248 -2742 254 -2532
rect 304 -2576 310 -2366
rect 344 -2576 350 -2366
rect 208 -2754 254 -2742
rect 290 -2756 300 -2576
rect 352 -2756 362 -2576
rect -614 -2792 -556 -2786
rect -422 -2792 -364 -2786
rect -230 -2792 -172 -2786
rect -38 -2792 20 -2786
rect 154 -2792 212 -2786
rect 392 -2792 628 -2320
rect 1282 -2322 1340 -2320
rect 1474 -2322 1532 -2320
rect 1666 -2322 1724 -2320
rect 1858 -2322 1916 -2320
rect 2050 -2322 2108 -2320
rect 1144 -2366 1190 -2354
rect 1144 -2576 1150 -2366
rect 1184 -2576 1190 -2366
rect 1226 -2532 1236 -2352
rect 1288 -2532 1298 -2352
rect 1336 -2366 1382 -2354
rect 1130 -2756 1140 -2576
rect 1192 -2756 1202 -2576
rect 1240 -2742 1246 -2532
rect 1280 -2742 1286 -2532
rect 1336 -2576 1342 -2366
rect 1376 -2576 1382 -2366
rect 1418 -2532 1428 -2352
rect 1480 -2532 1490 -2352
rect 1528 -2366 1574 -2354
rect 1240 -2754 1286 -2742
rect 1322 -2756 1332 -2576
rect 1384 -2756 1394 -2576
rect 1432 -2742 1438 -2532
rect 1472 -2742 1478 -2532
rect 1528 -2576 1534 -2366
rect 1568 -2576 1574 -2366
rect 1610 -2532 1620 -2352
rect 1672 -2532 1682 -2352
rect 1720 -2366 1766 -2354
rect 1432 -2754 1478 -2742
rect 1514 -2756 1524 -2576
rect 1576 -2756 1586 -2576
rect 1624 -2742 1630 -2532
rect 1664 -2742 1670 -2532
rect 1720 -2576 1726 -2366
rect 1760 -2576 1766 -2366
rect 1802 -2532 1812 -2352
rect 1864 -2532 1874 -2352
rect 1912 -2366 1958 -2354
rect 1624 -2754 1670 -2742
rect 1706 -2756 1716 -2576
rect 1768 -2756 1778 -2576
rect 1816 -2742 1822 -2532
rect 1856 -2742 1862 -2532
rect 1912 -2576 1918 -2366
rect 1952 -2576 1958 -2366
rect 1994 -2532 2004 -2352
rect 2056 -2532 2066 -2352
rect 2104 -2366 2150 -2354
rect 1816 -2754 1862 -2742
rect 1898 -2756 1908 -2576
rect 1960 -2756 1970 -2576
rect 2008 -2742 2014 -2532
rect 2048 -2742 2054 -2532
rect 2104 -2576 2110 -2366
rect 2144 -2576 2150 -2366
rect 2008 -2754 2054 -2742
rect 2090 -2756 2100 -2576
rect 2152 -2756 2162 -2576
rect 1186 -2792 1244 -2786
rect 1378 -2792 1436 -2786
rect 1570 -2792 1628 -2786
rect 1762 -2792 1820 -2786
rect 1954 -2792 2012 -2786
rect 2192 -2792 2428 -2320
rect 3082 -2322 3140 -2320
rect 3274 -2322 3332 -2320
rect 3466 -2322 3524 -2320
rect 3658 -2322 3716 -2320
rect 3850 -2322 3908 -2320
rect 2944 -2366 2990 -2354
rect 2944 -2576 2950 -2366
rect 2984 -2576 2990 -2366
rect 3026 -2532 3036 -2352
rect 3088 -2532 3098 -2352
rect 3136 -2366 3182 -2354
rect 2930 -2756 2940 -2576
rect 2992 -2756 3002 -2576
rect 3040 -2742 3046 -2532
rect 3080 -2742 3086 -2532
rect 3136 -2576 3142 -2366
rect 3176 -2576 3182 -2366
rect 3218 -2532 3228 -2352
rect 3280 -2532 3290 -2352
rect 3328 -2366 3374 -2354
rect 3040 -2754 3086 -2742
rect 3122 -2756 3132 -2576
rect 3184 -2756 3194 -2576
rect 3232 -2742 3238 -2532
rect 3272 -2742 3278 -2532
rect 3328 -2576 3334 -2366
rect 3368 -2576 3374 -2366
rect 3410 -2532 3420 -2352
rect 3472 -2532 3482 -2352
rect 3520 -2366 3566 -2354
rect 3232 -2754 3278 -2742
rect 3314 -2756 3324 -2576
rect 3376 -2756 3386 -2576
rect 3424 -2742 3430 -2532
rect 3464 -2742 3470 -2532
rect 3520 -2576 3526 -2366
rect 3560 -2576 3566 -2366
rect 3602 -2532 3612 -2352
rect 3664 -2532 3674 -2352
rect 3712 -2366 3758 -2354
rect 3424 -2754 3470 -2742
rect 3506 -2756 3516 -2576
rect 3568 -2756 3578 -2576
rect 3616 -2742 3622 -2532
rect 3656 -2742 3662 -2532
rect 3712 -2576 3718 -2366
rect 3752 -2576 3758 -2366
rect 3794 -2532 3804 -2352
rect 3856 -2532 3866 -2352
rect 3904 -2366 3950 -2354
rect 3616 -2754 3662 -2742
rect 3698 -2756 3708 -2576
rect 3760 -2756 3770 -2576
rect 3808 -2742 3814 -2532
rect 3848 -2742 3854 -2532
rect 3904 -2576 3910 -2366
rect 3944 -2576 3950 -2366
rect 3808 -2754 3854 -2742
rect 3890 -2756 3900 -2576
rect 3952 -2756 3962 -2576
rect 2986 -2792 3044 -2786
rect 3178 -2792 3236 -2786
rect 3370 -2792 3428 -2786
rect 3562 -2792 3620 -2786
rect 3754 -2792 3812 -2786
rect 3992 -2792 4228 -2320
rect 4402 -2648 4412 -2148
rect 4696 -2220 6776 -2148
rect 4696 -2254 4998 -2220
rect 5032 -2254 5190 -2220
rect 5224 -2254 5382 -2220
rect 5416 -2254 5574 -2220
rect 5608 -2254 5766 -2220
rect 5800 -2254 5958 -2220
rect 5992 -2254 6150 -2220
rect 6184 -2254 6342 -2220
rect 6376 -2254 6534 -2220
rect 6568 -2254 6726 -2220
rect 6760 -2254 6776 -2220
rect 4696 -2260 6776 -2254
rect 4696 -2648 4900 -2260
rect 4944 -2304 4990 -2292
rect 4944 -2508 4950 -2304
rect 4984 -2508 4990 -2304
rect 5026 -2472 5036 -2288
rect 5092 -2472 5102 -2288
rect 5136 -2304 5182 -2292
rect -3072 -2826 -2402 -2792
rect -2368 -2826 -2210 -2792
rect -2176 -2826 -2018 -2792
rect -1984 -2826 -1826 -2792
rect -1792 -2826 -1634 -2792
rect -1600 -2826 -602 -2792
rect -568 -2826 -410 -2792
rect -376 -2826 -218 -2792
rect -184 -2826 -26 -2792
rect 8 -2826 166 -2792
rect 200 -2826 1198 -2792
rect 1232 -2826 1390 -2792
rect 1424 -2826 1582 -2792
rect 1616 -2826 1774 -2792
rect 1808 -2826 1966 -2792
rect 2000 -2826 2998 -2792
rect 3032 -2826 3190 -2792
rect 3224 -2826 3382 -2792
rect 3416 -2826 3574 -2792
rect 3608 -2826 3766 -2792
rect 3800 -2826 4228 -2792
rect -3072 -2900 4228 -2826
rect -3072 -2934 -2402 -2900
rect -2368 -2934 -2210 -2900
rect -2176 -2934 -2018 -2900
rect -1984 -2934 -1826 -2900
rect -1792 -2934 -1634 -2900
rect -1600 -2934 -602 -2900
rect -568 -2934 -410 -2900
rect -376 -2934 -218 -2900
rect -184 -2934 -26 -2900
rect 8 -2934 166 -2900
rect 200 -2934 1198 -2900
rect 1232 -2934 1390 -2900
rect 1424 -2934 1582 -2900
rect 1616 -2934 1774 -2900
rect 1808 -2934 1966 -2900
rect 2000 -2934 2998 -2900
rect 3032 -2934 3190 -2900
rect 3224 -2934 3382 -2900
rect 3416 -2934 3574 -2900
rect 3608 -2934 3766 -2900
rect 3800 -2934 4228 -2900
rect -3072 -2936 4228 -2934
rect -3072 -3136 -2592 -2936
rect -2414 -2940 -2356 -2936
rect -2222 -2940 -2164 -2936
rect -2030 -2940 -1972 -2936
rect -1838 -2940 -1780 -2936
rect -1646 -2940 -1588 -2936
rect -3090 -3828 -3080 -3136
rect -2648 -3408 -2592 -3136
rect -2456 -2984 -2410 -2972
rect -2456 -3192 -2450 -2984
rect -2416 -3192 -2410 -2984
rect -2374 -3148 -2364 -2968
rect -2312 -3148 -2302 -2968
rect -2264 -2984 -2218 -2972
rect -2470 -3372 -2460 -3192
rect -2408 -3372 -2398 -3192
rect -2360 -3360 -2354 -3148
rect -2320 -3360 -2314 -3148
rect -2264 -3192 -2258 -2984
rect -2224 -3192 -2218 -2984
rect -2182 -3148 -2172 -2968
rect -2120 -3148 -2110 -2968
rect -2072 -2984 -2026 -2972
rect -2360 -3372 -2314 -3360
rect -2278 -3372 -2268 -3192
rect -2216 -3372 -2206 -3192
rect -2168 -3360 -2162 -3148
rect -2128 -3360 -2122 -3148
rect -2072 -3192 -2066 -2984
rect -2032 -3192 -2026 -2984
rect -1990 -3148 -1980 -2968
rect -1928 -3148 -1918 -2968
rect -1880 -2984 -1834 -2972
rect -2168 -3372 -2122 -3360
rect -2086 -3372 -2076 -3192
rect -2024 -3372 -2014 -3192
rect -1976 -3360 -1970 -3148
rect -1936 -3360 -1930 -3148
rect -1880 -3192 -1874 -2984
rect -1840 -3192 -1834 -2984
rect -1798 -3148 -1788 -2968
rect -1736 -3148 -1726 -2968
rect -1688 -2984 -1642 -2972
rect -1976 -3372 -1930 -3360
rect -1894 -3372 -1884 -3192
rect -1832 -3372 -1822 -3192
rect -1784 -3360 -1778 -3148
rect -1744 -3360 -1738 -3148
rect -1688 -3192 -1682 -2984
rect -1648 -3192 -1642 -2984
rect -1606 -3148 -1596 -2968
rect -1544 -3148 -1534 -2968
rect -1496 -2984 -1450 -2972
rect -1784 -3372 -1738 -3360
rect -1702 -3372 -1692 -3192
rect -1640 -3372 -1630 -3192
rect -1592 -3360 -1586 -3148
rect -1552 -3360 -1546 -3148
rect -1496 -3192 -1490 -2984
rect -1456 -3192 -1450 -2984
rect -1592 -3372 -1546 -3360
rect -1510 -3372 -1500 -3192
rect -1448 -3372 -1438 -3192
rect -2318 -3408 -2260 -3404
rect -2126 -3408 -2068 -3404
rect -1934 -3408 -1876 -3404
rect -1742 -3408 -1684 -3404
rect -1550 -3408 -1492 -3404
rect -1408 -3408 -1176 -2936
rect -614 -2940 -556 -2936
rect -422 -2940 -364 -2936
rect -230 -2940 -172 -2936
rect -38 -2940 20 -2936
rect 154 -2940 212 -2936
rect -656 -2984 -610 -2972
rect -656 -3192 -650 -2984
rect -616 -3192 -610 -2984
rect -574 -3148 -564 -2968
rect -512 -3148 -502 -2968
rect -464 -2984 -418 -2972
rect -670 -3372 -660 -3192
rect -608 -3372 -598 -3192
rect -560 -3360 -554 -3148
rect -520 -3360 -514 -3148
rect -464 -3192 -458 -2984
rect -424 -3192 -418 -2984
rect -382 -3148 -372 -2968
rect -320 -3148 -310 -2968
rect -272 -2984 -226 -2972
rect -560 -3372 -514 -3360
rect -478 -3372 -468 -3192
rect -416 -3372 -406 -3192
rect -368 -3360 -362 -3148
rect -328 -3360 -322 -3148
rect -272 -3192 -266 -2984
rect -232 -3192 -226 -2984
rect -190 -3148 -180 -2968
rect -128 -3148 -118 -2968
rect -80 -2984 -34 -2972
rect -368 -3372 -322 -3360
rect -286 -3372 -276 -3192
rect -224 -3372 -214 -3192
rect -176 -3360 -170 -3148
rect -136 -3360 -130 -3148
rect -80 -3192 -74 -2984
rect -40 -3192 -34 -2984
rect 2 -3148 12 -2968
rect 64 -3148 74 -2968
rect 112 -2984 158 -2972
rect -176 -3372 -130 -3360
rect -94 -3372 -84 -3192
rect -32 -3372 -22 -3192
rect 16 -3360 22 -3148
rect 56 -3360 62 -3148
rect 112 -3192 118 -2984
rect 152 -3192 158 -2984
rect 194 -3148 204 -2968
rect 256 -3148 266 -2968
rect 304 -2984 350 -2972
rect 16 -3372 62 -3360
rect 98 -3372 108 -3192
rect 160 -3372 170 -3192
rect 208 -3360 214 -3148
rect 248 -3360 254 -3148
rect 304 -3192 310 -2984
rect 344 -3192 350 -2984
rect 208 -3372 254 -3360
rect 290 -3372 300 -3192
rect 352 -3372 362 -3192
rect -518 -3408 -460 -3404
rect -326 -3408 -268 -3404
rect -134 -3408 -76 -3404
rect 58 -3408 116 -3404
rect 250 -3408 308 -3404
rect 392 -3408 628 -2936
rect 1186 -2940 1244 -2936
rect 1378 -2940 1436 -2936
rect 1570 -2940 1628 -2936
rect 1762 -2940 1820 -2936
rect 1954 -2940 2012 -2936
rect 1144 -2984 1190 -2972
rect 1144 -3192 1150 -2984
rect 1184 -3192 1190 -2984
rect 1226 -3148 1236 -2968
rect 1288 -3148 1298 -2968
rect 1336 -2984 1382 -2972
rect 1130 -3372 1140 -3192
rect 1192 -3372 1202 -3192
rect 1240 -3360 1246 -3148
rect 1280 -3360 1286 -3148
rect 1336 -3192 1342 -2984
rect 1376 -3192 1382 -2984
rect 1418 -3148 1428 -2968
rect 1480 -3148 1490 -2968
rect 1528 -2984 1574 -2972
rect 1240 -3372 1286 -3360
rect 1322 -3372 1332 -3192
rect 1384 -3372 1394 -3192
rect 1432 -3360 1438 -3148
rect 1472 -3360 1478 -3148
rect 1528 -3192 1534 -2984
rect 1568 -3192 1574 -2984
rect 1610 -3148 1620 -2968
rect 1672 -3148 1682 -2968
rect 1720 -2984 1766 -2972
rect 1432 -3372 1478 -3360
rect 1514 -3372 1524 -3192
rect 1576 -3372 1586 -3192
rect 1624 -3360 1630 -3148
rect 1664 -3360 1670 -3148
rect 1720 -3192 1726 -2984
rect 1760 -3192 1766 -2984
rect 1802 -3148 1812 -2968
rect 1864 -3148 1874 -2968
rect 1912 -2984 1958 -2972
rect 1624 -3372 1670 -3360
rect 1706 -3372 1716 -3192
rect 1768 -3372 1778 -3192
rect 1816 -3360 1822 -3148
rect 1856 -3360 1862 -3148
rect 1912 -3192 1918 -2984
rect 1952 -3192 1958 -2984
rect 1994 -3148 2004 -2968
rect 2056 -3148 2066 -2968
rect 2104 -2984 2150 -2972
rect 1816 -3372 1862 -3360
rect 1898 -3372 1908 -3192
rect 1960 -3372 1970 -3192
rect 2008 -3360 2014 -3148
rect 2048 -3360 2054 -3148
rect 2104 -3192 2110 -2984
rect 2144 -3192 2150 -2984
rect 2008 -3372 2054 -3360
rect 2090 -3372 2100 -3192
rect 2152 -3372 2162 -3192
rect 1282 -3408 1340 -3404
rect 1474 -3408 1532 -3404
rect 1666 -3408 1724 -3404
rect 1858 -3408 1916 -3404
rect 2050 -3408 2108 -3404
rect 2192 -3408 2428 -2936
rect 2986 -2940 3044 -2936
rect 3178 -2940 3236 -2936
rect 3370 -2940 3428 -2936
rect 3562 -2940 3620 -2936
rect 3754 -2940 3812 -2936
rect 2944 -2984 2990 -2972
rect 2944 -3192 2950 -2984
rect 2984 -3192 2990 -2984
rect 3026 -3148 3036 -2968
rect 3088 -3148 3098 -2968
rect 3136 -2984 3182 -2972
rect 2930 -3372 2940 -3192
rect 2992 -3372 3002 -3192
rect 3040 -3360 3046 -3148
rect 3080 -3360 3086 -3148
rect 3136 -3192 3142 -2984
rect 3176 -3192 3182 -2984
rect 3218 -3148 3228 -2968
rect 3280 -3148 3290 -2968
rect 3328 -2984 3374 -2972
rect 3040 -3372 3086 -3360
rect 3122 -3372 3132 -3192
rect 3184 -3372 3194 -3192
rect 3232 -3360 3238 -3148
rect 3272 -3360 3278 -3148
rect 3328 -3192 3334 -2984
rect 3368 -3192 3374 -2984
rect 3410 -3148 3420 -2968
rect 3472 -3148 3482 -2968
rect 3520 -2984 3566 -2972
rect 3232 -3372 3278 -3360
rect 3314 -3372 3324 -3192
rect 3376 -3372 3386 -3192
rect 3424 -3360 3430 -3148
rect 3464 -3360 3470 -3148
rect 3520 -3192 3526 -2984
rect 3560 -3192 3566 -2984
rect 3602 -3148 3612 -2968
rect 3664 -3148 3674 -2968
rect 3712 -2984 3758 -2972
rect 3424 -3372 3470 -3360
rect 3506 -3372 3516 -3192
rect 3568 -3372 3578 -3192
rect 3616 -3360 3622 -3148
rect 3656 -3360 3662 -3148
rect 3712 -3192 3718 -2984
rect 3752 -3192 3758 -2984
rect 3794 -3148 3804 -2968
rect 3856 -3148 3866 -2968
rect 3904 -2984 3950 -2972
rect 3616 -3372 3662 -3360
rect 3698 -3372 3708 -3192
rect 3760 -3372 3770 -3192
rect 3808 -3360 3814 -3148
rect 3848 -3360 3854 -3148
rect 3904 -3192 3910 -2984
rect 3944 -3192 3950 -2984
rect 3808 -3372 3854 -3360
rect 3890 -3372 3900 -3192
rect 3952 -3372 3962 -3192
rect 3082 -3408 3140 -3404
rect 3274 -3408 3332 -3404
rect 3466 -3408 3524 -3404
rect 3658 -3408 3716 -3404
rect 3850 -3408 3908 -3404
rect 3992 -3408 4228 -2936
rect -2648 -3410 4228 -3408
rect -2648 -3444 -2306 -3410
rect -2272 -3444 -2114 -3410
rect -2080 -3444 -1922 -3410
rect -1888 -3444 -1730 -3410
rect -1696 -3444 -1538 -3410
rect -1504 -3444 -506 -3410
rect -472 -3444 -314 -3410
rect -280 -3444 -122 -3410
rect -88 -3444 70 -3410
rect 104 -3444 262 -3410
rect 296 -3444 1294 -3410
rect 1328 -3444 1486 -3410
rect 1520 -3444 1678 -3410
rect 1712 -3444 1870 -3410
rect 1904 -3444 2062 -3410
rect 2096 -3444 3094 -3410
rect 3128 -3444 3286 -3410
rect 3320 -3444 3478 -3410
rect 3512 -3444 3670 -3410
rect 3704 -3444 3862 -3410
rect 3896 -3444 4228 -3410
rect 4480 -2724 4900 -2648
rect 4930 -2692 4940 -2508
rect 4996 -2692 5006 -2508
rect 5040 -2680 5046 -2472
rect 5080 -2680 5086 -2472
rect 5136 -2508 5142 -2304
rect 5176 -2508 5182 -2304
rect 5218 -2472 5228 -2288
rect 5284 -2472 5294 -2288
rect 5328 -2304 5374 -2292
rect 5040 -2692 5086 -2680
rect 5122 -2692 5132 -2508
rect 5188 -2692 5198 -2508
rect 5232 -2680 5238 -2472
rect 5272 -2680 5278 -2472
rect 5328 -2508 5334 -2304
rect 5368 -2508 5374 -2304
rect 5410 -2472 5420 -2288
rect 5476 -2472 5486 -2288
rect 5520 -2304 5566 -2292
rect 5232 -2692 5278 -2680
rect 5314 -2692 5324 -2508
rect 5380 -2692 5390 -2508
rect 5424 -2680 5430 -2472
rect 5464 -2680 5470 -2472
rect 5520 -2508 5526 -2304
rect 5560 -2508 5566 -2304
rect 5602 -2472 5612 -2288
rect 5668 -2472 5678 -2288
rect 5712 -2304 5758 -2292
rect 5424 -2692 5470 -2680
rect 5506 -2692 5516 -2508
rect 5572 -2692 5582 -2508
rect 5616 -2680 5622 -2472
rect 5656 -2680 5662 -2472
rect 5712 -2508 5718 -2304
rect 5752 -2508 5758 -2304
rect 5794 -2472 5804 -2288
rect 5860 -2472 5870 -2288
rect 5904 -2304 5950 -2292
rect 5616 -2692 5662 -2680
rect 5698 -2692 5708 -2508
rect 5764 -2692 5774 -2508
rect 5808 -2680 5814 -2472
rect 5848 -2680 5854 -2472
rect 5904 -2508 5910 -2304
rect 5944 -2508 5950 -2304
rect 5986 -2472 5996 -2288
rect 6052 -2472 6062 -2288
rect 6096 -2304 6142 -2292
rect 5808 -2692 5854 -2680
rect 5890 -2692 5900 -2508
rect 5956 -2692 5966 -2508
rect 6000 -2680 6006 -2472
rect 6040 -2680 6046 -2472
rect 6096 -2508 6102 -2304
rect 6136 -2508 6142 -2304
rect 6178 -2472 6188 -2288
rect 6244 -2472 6254 -2288
rect 6288 -2304 6334 -2292
rect 6000 -2692 6046 -2680
rect 6082 -2692 6092 -2508
rect 6148 -2692 6158 -2508
rect 6192 -2680 6198 -2472
rect 6232 -2680 6238 -2472
rect 6288 -2508 6294 -2304
rect 6328 -2508 6334 -2304
rect 6370 -2472 6380 -2288
rect 6436 -2472 6446 -2288
rect 6480 -2304 6526 -2292
rect 6192 -2692 6238 -2680
rect 6274 -2692 6284 -2508
rect 6340 -2692 6350 -2508
rect 6384 -2680 6390 -2472
rect 6424 -2680 6430 -2472
rect 6480 -2508 6486 -2304
rect 6520 -2508 6526 -2304
rect 6562 -2472 6572 -2288
rect 6628 -2472 6638 -2288
rect 6672 -2304 6718 -2292
rect 6384 -2692 6430 -2680
rect 6466 -2692 6476 -2508
rect 6532 -2692 6542 -2508
rect 6576 -2680 6582 -2472
rect 6616 -2680 6622 -2472
rect 6672 -2508 6678 -2304
rect 6712 -2508 6718 -2304
rect 6754 -2472 6764 -2288
rect 6820 -2472 6830 -2288
rect 6864 -2304 6910 -2292
rect 6576 -2692 6622 -2680
rect 6658 -2692 6668 -2508
rect 6724 -2692 6734 -2508
rect 6768 -2680 6774 -2472
rect 6808 -2680 6814 -2472
rect 6864 -2508 6870 -2304
rect 6904 -2508 6910 -2304
rect 6768 -2692 6814 -2680
rect 6850 -2692 6860 -2508
rect 6916 -2692 6926 -2508
rect 4480 -2730 6872 -2724
rect 4480 -2764 5094 -2730
rect 5128 -2764 5286 -2730
rect 5320 -2764 5478 -2730
rect 5512 -2764 5670 -2730
rect 5704 -2764 5862 -2730
rect 5896 -2764 6054 -2730
rect 6088 -2764 6246 -2730
rect 6280 -2764 6438 -2730
rect 6472 -2764 6630 -2730
rect 6664 -2764 6822 -2730
rect 6856 -2764 6872 -2730
rect 4480 -2838 6872 -2764
rect 4480 -2872 5094 -2838
rect 5128 -2872 5286 -2838
rect 5320 -2872 5478 -2838
rect 5512 -2872 5670 -2838
rect 5704 -2872 5862 -2838
rect 5896 -2872 6054 -2838
rect 6088 -2872 6246 -2838
rect 6280 -2872 6438 -2838
rect 6472 -2872 6630 -2838
rect 6664 -2872 6822 -2838
rect 6856 -2872 6872 -2838
rect 4480 -2880 6872 -2872
rect 4480 -3340 4900 -2880
rect 4944 -2922 4990 -2910
rect 4944 -3128 4950 -2922
rect 4984 -3128 4990 -2922
rect 5026 -3092 5036 -2908
rect 5092 -3092 5102 -2908
rect 5136 -2922 5182 -2910
rect 4930 -3312 4940 -3128
rect 4996 -3312 5006 -3128
rect 5040 -3298 5046 -3092
rect 5080 -3298 5086 -3092
rect 5136 -3128 5142 -2922
rect 5176 -3128 5182 -2922
rect 5218 -3092 5228 -2908
rect 5284 -3092 5294 -2908
rect 5328 -2922 5374 -2910
rect 5040 -3310 5086 -3298
rect 5122 -3312 5132 -3128
rect 5188 -3312 5198 -3128
rect 5232 -3298 5238 -3092
rect 5272 -3298 5278 -3092
rect 5328 -3128 5334 -2922
rect 5368 -3128 5374 -2922
rect 5410 -3092 5420 -2908
rect 5476 -3092 5486 -2908
rect 5520 -2922 5566 -2910
rect 5232 -3310 5278 -3298
rect 5314 -3312 5324 -3128
rect 5380 -3312 5390 -3128
rect 5424 -3298 5430 -3092
rect 5464 -3298 5470 -3092
rect 5520 -3128 5526 -2922
rect 5560 -3128 5566 -2922
rect 5602 -3092 5612 -2908
rect 5668 -3092 5678 -2908
rect 5712 -2922 5758 -2910
rect 5424 -3310 5470 -3298
rect 5506 -3312 5516 -3128
rect 5572 -3312 5582 -3128
rect 5616 -3298 5622 -3092
rect 5656 -3298 5662 -3092
rect 5712 -3128 5718 -2922
rect 5752 -3128 5758 -2922
rect 5794 -3092 5804 -2908
rect 5860 -3092 5870 -2908
rect 5904 -2922 5950 -2910
rect 5616 -3310 5662 -3298
rect 5698 -3312 5708 -3128
rect 5764 -3312 5774 -3128
rect 5808 -3298 5814 -3092
rect 5848 -3298 5854 -3092
rect 5904 -3128 5910 -2922
rect 5944 -3128 5950 -2922
rect 5986 -3092 5996 -2908
rect 6052 -3092 6062 -2908
rect 6096 -2922 6142 -2910
rect 5808 -3310 5854 -3298
rect 5890 -3312 5900 -3128
rect 5956 -3312 5966 -3128
rect 6000 -3298 6006 -3092
rect 6040 -3298 6046 -3092
rect 6096 -3128 6102 -2922
rect 6136 -3128 6142 -2922
rect 6178 -3092 6188 -2908
rect 6244 -3092 6254 -2908
rect 6288 -2922 6334 -2910
rect 6000 -3310 6046 -3298
rect 6082 -3312 6092 -3128
rect 6148 -3312 6158 -3128
rect 6192 -3298 6198 -3092
rect 6232 -3298 6238 -3092
rect 6288 -3128 6294 -2922
rect 6328 -3128 6334 -2922
rect 6370 -3092 6380 -2908
rect 6436 -3092 6446 -2908
rect 6480 -2922 6526 -2910
rect 6192 -3310 6238 -3298
rect 6274 -3312 6284 -3128
rect 6340 -3312 6350 -3128
rect 6384 -3298 6390 -3092
rect 6424 -3298 6430 -3092
rect 6480 -3128 6486 -2922
rect 6520 -3128 6526 -2922
rect 6562 -3092 6572 -2908
rect 6628 -3092 6638 -2908
rect 6672 -2922 6718 -2910
rect 6384 -3310 6430 -3298
rect 6466 -3312 6476 -3128
rect 6532 -3312 6542 -3128
rect 6576 -3298 6582 -3092
rect 6616 -3298 6622 -3092
rect 6672 -3128 6678 -2922
rect 6712 -3128 6718 -2922
rect 6754 -3092 6764 -2908
rect 6820 -3092 6830 -2908
rect 6864 -2922 6910 -2910
rect 6576 -3310 6622 -3298
rect 6658 -3312 6668 -3128
rect 6724 -3312 6734 -3128
rect 6768 -3298 6774 -3092
rect 6808 -3298 6814 -3092
rect 6864 -3128 6870 -2922
rect 6904 -3128 6910 -2922
rect 6768 -3310 6814 -3298
rect 6850 -3312 6860 -3128
rect 6916 -3312 6926 -3128
rect 4480 -3348 6776 -3340
rect 4480 -3382 4998 -3348
rect 5032 -3382 5190 -3348
rect 5224 -3382 5382 -3348
rect 5416 -3382 5574 -3348
rect 5608 -3382 5766 -3348
rect 5800 -3382 5958 -3348
rect 5992 -3382 6150 -3348
rect 6184 -3382 6342 -3348
rect 6376 -3382 6534 -3348
rect 6568 -3382 6726 -3348
rect 6760 -3382 6776 -3348
rect 4480 -3436 6776 -3382
rect -2648 -3518 4228 -3444
rect -2648 -3552 -2306 -3518
rect -2272 -3552 -2114 -3518
rect -2080 -3552 -1922 -3518
rect -1888 -3552 -1730 -3518
rect -1696 -3552 -1538 -3518
rect -1504 -3552 -506 -3518
rect -472 -3552 -314 -3518
rect -280 -3552 -122 -3518
rect -88 -3552 70 -3518
rect 104 -3552 262 -3518
rect 296 -3552 1294 -3518
rect 1328 -3552 1486 -3518
rect 1520 -3552 1678 -3518
rect 1712 -3552 1870 -3518
rect 1904 -3552 2062 -3518
rect 2096 -3552 3094 -3518
rect 3128 -3552 3286 -3518
rect 3320 -3552 3478 -3518
rect 3512 -3552 3670 -3518
rect 3704 -3552 3862 -3518
rect 3896 -3552 4228 -3518
rect -2648 -3828 -2592 -3552
rect -2318 -3558 -2260 -3552
rect -2126 -3558 -2068 -3552
rect -1934 -3558 -1876 -3552
rect -1742 -3558 -1684 -3552
rect -1550 -3558 -1492 -3552
rect -2456 -3602 -2410 -3590
rect -2456 -3812 -2450 -3602
rect -2416 -3812 -2410 -3602
rect -2374 -3768 -2364 -3588
rect -2312 -3768 -2302 -3588
rect -2264 -3602 -2218 -3590
rect -3072 -4032 -2592 -3828
rect -2470 -3992 -2460 -3812
rect -2408 -3992 -2398 -3812
rect -2360 -3978 -2354 -3768
rect -2320 -3978 -2314 -3768
rect -2264 -3812 -2258 -3602
rect -2224 -3812 -2218 -3602
rect -2182 -3768 -2172 -3588
rect -2120 -3768 -2110 -3588
rect -2072 -3602 -2026 -3590
rect -2360 -3990 -2314 -3978
rect -2278 -3992 -2268 -3812
rect -2216 -3992 -2206 -3812
rect -2168 -3978 -2162 -3768
rect -2128 -3978 -2122 -3768
rect -2072 -3812 -2066 -3602
rect -2032 -3812 -2026 -3602
rect -1990 -3768 -1980 -3588
rect -1928 -3768 -1918 -3588
rect -1880 -3602 -1834 -3590
rect -2168 -3990 -2122 -3978
rect -2086 -3992 -2076 -3812
rect -2024 -3992 -2014 -3812
rect -1976 -3978 -1970 -3768
rect -1936 -3978 -1930 -3768
rect -1880 -3812 -1874 -3602
rect -1840 -3812 -1834 -3602
rect -1798 -3768 -1788 -3588
rect -1736 -3768 -1726 -3588
rect -1688 -3602 -1642 -3590
rect -1976 -3990 -1930 -3978
rect -1894 -3992 -1884 -3812
rect -1832 -3992 -1822 -3812
rect -1784 -3978 -1778 -3768
rect -1744 -3978 -1738 -3768
rect -1688 -3812 -1682 -3602
rect -1648 -3812 -1642 -3602
rect -1606 -3768 -1596 -3588
rect -1544 -3768 -1534 -3588
rect -1496 -3602 -1450 -3590
rect -1784 -3990 -1738 -3978
rect -1702 -3992 -1692 -3812
rect -1640 -3992 -1630 -3812
rect -1592 -3978 -1586 -3768
rect -1552 -3978 -1546 -3768
rect -1496 -3812 -1490 -3602
rect -1456 -3812 -1450 -3602
rect -1592 -3990 -1546 -3978
rect -1510 -3992 -1500 -3812
rect -1448 -3992 -1438 -3812
rect -2414 -4028 -2356 -4022
rect -2222 -4028 -2164 -4022
rect -2030 -4028 -1972 -4022
rect -1838 -4028 -1780 -4022
rect -1646 -4028 -1588 -4022
rect -1408 -4028 -1176 -3552
rect -518 -3558 -460 -3552
rect -326 -3558 -268 -3552
rect -134 -3558 -76 -3552
rect 58 -3558 116 -3552
rect 250 -3558 308 -3552
rect -656 -3602 -610 -3590
rect -656 -3812 -650 -3602
rect -616 -3812 -610 -3602
rect -574 -3768 -564 -3588
rect -512 -3768 -502 -3588
rect -464 -3602 -418 -3590
rect -670 -3992 -660 -3812
rect -608 -3992 -598 -3812
rect -560 -3978 -554 -3768
rect -520 -3978 -514 -3768
rect -464 -3812 -458 -3602
rect -424 -3812 -418 -3602
rect -382 -3768 -372 -3588
rect -320 -3768 -310 -3588
rect -272 -3602 -226 -3590
rect -560 -3990 -514 -3978
rect -478 -3992 -468 -3812
rect -416 -3992 -406 -3812
rect -368 -3978 -362 -3768
rect -328 -3978 -322 -3768
rect -272 -3812 -266 -3602
rect -232 -3812 -226 -3602
rect -190 -3768 -180 -3588
rect -128 -3768 -118 -3588
rect -80 -3602 -34 -3590
rect -368 -3990 -322 -3978
rect -286 -3992 -276 -3812
rect -224 -3992 -214 -3812
rect -176 -3978 -170 -3768
rect -136 -3978 -130 -3768
rect -80 -3812 -74 -3602
rect -40 -3812 -34 -3602
rect 2 -3768 12 -3588
rect 64 -3768 74 -3588
rect 112 -3602 158 -3590
rect -176 -3990 -130 -3978
rect -94 -3992 -84 -3812
rect -32 -3992 -22 -3812
rect 16 -3978 22 -3768
rect 56 -3978 62 -3768
rect 112 -3812 118 -3602
rect 152 -3812 158 -3602
rect 194 -3768 204 -3588
rect 256 -3768 266 -3588
rect 304 -3602 350 -3590
rect 16 -3990 62 -3978
rect 98 -3992 108 -3812
rect 160 -3992 170 -3812
rect 208 -3978 214 -3768
rect 248 -3978 254 -3768
rect 304 -3812 310 -3602
rect 344 -3812 350 -3602
rect 208 -3990 254 -3978
rect 290 -3992 300 -3812
rect 352 -3992 362 -3812
rect -614 -4028 -556 -4022
rect -422 -4028 -364 -4022
rect -230 -4028 -172 -4022
rect -38 -4028 20 -4022
rect 154 -4028 212 -4022
rect 392 -4028 628 -3552
rect 1282 -3558 1340 -3552
rect 1474 -3558 1532 -3552
rect 1666 -3558 1724 -3552
rect 1858 -3558 1916 -3552
rect 2050 -3558 2108 -3552
rect 1144 -3602 1190 -3590
rect 1144 -3812 1150 -3602
rect 1184 -3812 1190 -3602
rect 1226 -3768 1236 -3588
rect 1288 -3768 1298 -3588
rect 1336 -3602 1382 -3590
rect 1130 -3992 1140 -3812
rect 1192 -3992 1202 -3812
rect 1240 -3978 1246 -3768
rect 1280 -3978 1286 -3768
rect 1336 -3812 1342 -3602
rect 1376 -3812 1382 -3602
rect 1418 -3768 1428 -3588
rect 1480 -3768 1490 -3588
rect 1528 -3602 1574 -3590
rect 1240 -3990 1286 -3978
rect 1322 -3992 1332 -3812
rect 1384 -3992 1394 -3812
rect 1432 -3978 1438 -3768
rect 1472 -3978 1478 -3768
rect 1528 -3812 1534 -3602
rect 1568 -3812 1574 -3602
rect 1610 -3768 1620 -3588
rect 1672 -3768 1682 -3588
rect 1720 -3602 1766 -3590
rect 1432 -3990 1478 -3978
rect 1514 -3992 1524 -3812
rect 1576 -3992 1586 -3812
rect 1624 -3978 1630 -3768
rect 1664 -3978 1670 -3768
rect 1720 -3812 1726 -3602
rect 1760 -3812 1766 -3602
rect 1802 -3768 1812 -3588
rect 1864 -3768 1874 -3588
rect 1912 -3602 1958 -3590
rect 1624 -3990 1670 -3978
rect 1706 -3992 1716 -3812
rect 1768 -3992 1778 -3812
rect 1816 -3978 1822 -3768
rect 1856 -3978 1862 -3768
rect 1912 -3812 1918 -3602
rect 1952 -3812 1958 -3602
rect 1994 -3768 2004 -3588
rect 2056 -3768 2066 -3588
rect 2104 -3602 2150 -3590
rect 1816 -3990 1862 -3978
rect 1898 -3992 1908 -3812
rect 1960 -3992 1970 -3812
rect 2008 -3978 2014 -3768
rect 2048 -3978 2054 -3768
rect 2104 -3812 2110 -3602
rect 2144 -3812 2150 -3602
rect 2008 -3990 2054 -3978
rect 2090 -3992 2100 -3812
rect 2152 -3992 2162 -3812
rect 1186 -4028 1244 -4022
rect 1378 -4028 1436 -4022
rect 1570 -4028 1628 -4022
rect 1762 -4028 1820 -4022
rect 1954 -4028 2012 -4022
rect 2192 -4028 2428 -3552
rect 3082 -3558 3140 -3552
rect 3274 -3558 3332 -3552
rect 3466 -3558 3524 -3552
rect 3658 -3558 3716 -3552
rect 3850 -3558 3908 -3552
rect 2944 -3602 2990 -3590
rect 2944 -3812 2950 -3602
rect 2984 -3812 2990 -3602
rect 3026 -3768 3036 -3588
rect 3088 -3768 3098 -3588
rect 3136 -3602 3182 -3590
rect 2930 -3992 2940 -3812
rect 2992 -3992 3002 -3812
rect 3040 -3978 3046 -3768
rect 3080 -3978 3086 -3768
rect 3136 -3812 3142 -3602
rect 3176 -3812 3182 -3602
rect 3218 -3768 3228 -3588
rect 3280 -3768 3290 -3588
rect 3328 -3602 3374 -3590
rect 3040 -3990 3086 -3978
rect 3122 -3992 3132 -3812
rect 3184 -3992 3194 -3812
rect 3232 -3978 3238 -3768
rect 3272 -3978 3278 -3768
rect 3328 -3812 3334 -3602
rect 3368 -3812 3374 -3602
rect 3410 -3768 3420 -3588
rect 3472 -3768 3482 -3588
rect 3520 -3602 3566 -3590
rect 3232 -3990 3278 -3978
rect 3314 -3992 3324 -3812
rect 3376 -3992 3386 -3812
rect 3424 -3978 3430 -3768
rect 3464 -3978 3470 -3768
rect 3520 -3812 3526 -3602
rect 3560 -3812 3566 -3602
rect 3602 -3768 3612 -3588
rect 3664 -3768 3674 -3588
rect 3712 -3602 3758 -3590
rect 3424 -3990 3470 -3978
rect 3506 -3992 3516 -3812
rect 3568 -3992 3578 -3812
rect 3616 -3978 3622 -3768
rect 3656 -3978 3662 -3768
rect 3712 -3812 3718 -3602
rect 3752 -3812 3758 -3602
rect 3794 -3768 3804 -3588
rect 3856 -3768 3866 -3588
rect 3904 -3602 3950 -3590
rect 3616 -3990 3662 -3978
rect 3698 -3992 3708 -3812
rect 3760 -3992 3770 -3812
rect 3808 -3978 3814 -3768
rect 3848 -3978 3854 -3768
rect 3904 -3812 3910 -3602
rect 3944 -3812 3950 -3602
rect 3808 -3990 3854 -3978
rect 3890 -3992 3900 -3812
rect 3952 -3992 3962 -3812
rect 2986 -4028 3044 -4022
rect 3178 -4028 3236 -4022
rect 3370 -4028 3428 -4022
rect 3562 -4028 3620 -4022
rect 3754 -4028 3812 -4022
rect 3992 -4028 4228 -3552
rect -2420 -4032 -2402 -4028
rect -3072 -4062 -2402 -4032
rect -2368 -4062 -2210 -4028
rect -2176 -4062 -2018 -4028
rect -1984 -4062 -1826 -4028
rect -1792 -4062 -1634 -4028
rect -1600 -4032 -1176 -4028
rect -620 -4032 -602 -4028
rect -1600 -4062 -602 -4032
rect -568 -4062 -410 -4028
rect -376 -4062 -218 -4028
rect -184 -4062 -26 -4028
rect 8 -4062 166 -4028
rect 200 -4032 628 -4028
rect 1180 -4032 1198 -4028
rect 200 -4062 1198 -4032
rect 1232 -4062 1390 -4028
rect 1424 -4062 1582 -4028
rect 1616 -4062 1774 -4028
rect 1808 -4062 1966 -4028
rect 2000 -4032 2428 -4028
rect 2980 -4032 2998 -4028
rect 2000 -4062 2998 -4032
rect 3032 -4062 3190 -4028
rect 3224 -4062 3382 -4028
rect 3416 -4062 3574 -4028
rect 3608 -4062 3766 -4028
rect 3800 -4032 4228 -4028
rect 3800 -4062 4460 -4032
rect -3072 -4428 4460 -4062
rect -3072 -4440 -2388 -4428
rect -2412 -4462 -2388 -4440
rect -2220 -4462 -2130 -4428
rect -1962 -4462 -1872 -4428
rect -1704 -4462 -1614 -4428
rect -1446 -4462 -1356 -4428
rect -1188 -4440 -588 -4428
rect -1188 -4462 -1172 -4440
rect -2412 -4468 -1172 -4462
rect -612 -4462 -588 -4440
rect -420 -4462 -330 -4428
rect -162 -4462 -72 -4428
rect 96 -4462 186 -4428
rect 354 -4462 444 -4428
rect 612 -4440 1212 -4428
rect 612 -4462 628 -4440
rect -612 -4468 628 -4462
rect 1188 -4462 1212 -4440
rect 1380 -4462 1470 -4428
rect 1638 -4462 1728 -4428
rect 1896 -4462 1986 -4428
rect 2154 -4462 2244 -4428
rect 2412 -4440 3012 -4428
rect 2412 -4462 2428 -4440
rect 1188 -4468 2428 -4462
rect 2988 -4462 3012 -4440
rect 3180 -4462 3270 -4428
rect 3438 -4462 3528 -4428
rect 3696 -4462 3786 -4428
rect 3954 -4462 4044 -4428
rect 4212 -4440 4460 -4428
rect 4212 -4462 4228 -4440
rect 2988 -4468 4228 -4462
rect -2470 -4680 -2460 -4500
rect -2408 -4680 -2398 -4500
rect -2198 -4512 -2152 -4500
rect -2456 -4888 -2450 -4680
rect -2416 -4888 -2410 -4680
rect -2198 -4720 -2192 -4512
rect -2158 -4720 -2152 -4512
rect -2456 -4900 -2410 -4888
rect -2210 -4900 -2200 -4720
rect -2148 -4900 -2138 -4720
rect -2108 -4932 -1988 -4468
rect -1954 -4680 -1944 -4500
rect -1892 -4680 -1882 -4500
rect -1940 -4888 -1934 -4680
rect -1900 -4888 -1894 -4680
rect -1940 -4900 -1894 -4888
rect -1848 -4932 -1728 -4468
rect -1682 -4512 -1636 -4500
rect -1682 -4720 -1676 -4512
rect -1642 -4720 -1636 -4512
rect -1694 -4900 -1684 -4720
rect -1632 -4900 -1622 -4720
rect -1588 -4932 -1468 -4468
rect -1438 -4680 -1428 -4500
rect -1376 -4680 -1366 -4500
rect -1166 -4512 -1120 -4500
rect -1424 -4888 -1418 -4680
rect -1384 -4888 -1378 -4680
rect -1166 -4720 -1160 -4512
rect -1126 -4720 -1120 -4512
rect -670 -4680 -660 -4500
rect -608 -4680 -598 -4500
rect -398 -4512 -352 -4500
rect -1424 -4900 -1378 -4888
rect -1178 -4900 -1168 -4720
rect -1116 -4900 -1106 -4720
rect -656 -4888 -650 -4680
rect -616 -4888 -610 -4680
rect -398 -4720 -392 -4512
rect -358 -4720 -352 -4512
rect -656 -4900 -610 -4888
rect -410 -4900 -400 -4720
rect -348 -4900 -338 -4720
rect -308 -4932 -188 -4468
rect -154 -4680 -144 -4500
rect -92 -4680 -82 -4500
rect -140 -4888 -134 -4680
rect -100 -4888 -94 -4680
rect -140 -4900 -94 -4888
rect -48 -4932 72 -4468
rect 118 -4512 164 -4500
rect 118 -4720 124 -4512
rect 158 -4720 164 -4512
rect 106 -4900 116 -4720
rect 168 -4900 178 -4720
rect 212 -4932 332 -4468
rect 362 -4680 372 -4500
rect 424 -4680 434 -4500
rect 634 -4512 680 -4500
rect 376 -4888 382 -4680
rect 416 -4888 422 -4680
rect 634 -4720 640 -4512
rect 674 -4720 680 -4512
rect 1130 -4680 1140 -4500
rect 1192 -4680 1202 -4500
rect 1402 -4512 1448 -4500
rect 376 -4900 422 -4888
rect 622 -4900 632 -4720
rect 684 -4900 694 -4720
rect 1144 -4888 1150 -4680
rect 1184 -4888 1190 -4680
rect 1402 -4720 1408 -4512
rect 1442 -4720 1448 -4512
rect 1144 -4900 1190 -4888
rect 1390 -4900 1400 -4720
rect 1452 -4900 1462 -4720
rect 1492 -4932 1612 -4468
rect 1646 -4680 1656 -4500
rect 1708 -4680 1718 -4500
rect 1660 -4888 1666 -4680
rect 1700 -4888 1706 -4680
rect 1660 -4900 1706 -4888
rect 1752 -4932 1872 -4468
rect 1918 -4512 1964 -4500
rect 1918 -4720 1924 -4512
rect 1958 -4720 1964 -4512
rect 1906 -4900 1916 -4720
rect 1968 -4900 1978 -4720
rect 2012 -4932 2132 -4468
rect 2162 -4680 2172 -4500
rect 2224 -4680 2234 -4500
rect 2434 -4512 2480 -4500
rect 2176 -4888 2182 -4680
rect 2216 -4888 2222 -4680
rect 2434 -4720 2440 -4512
rect 2474 -4720 2480 -4512
rect 2930 -4680 2940 -4500
rect 2992 -4680 3002 -4500
rect 3202 -4512 3248 -4500
rect 2176 -4900 2222 -4888
rect 2422 -4900 2432 -4720
rect 2484 -4900 2494 -4720
rect 2944 -4888 2950 -4680
rect 2984 -4888 2990 -4680
rect 3202 -4720 3208 -4512
rect 3242 -4720 3248 -4512
rect 2944 -4900 2990 -4888
rect 3190 -4900 3200 -4720
rect 3252 -4900 3262 -4720
rect 3292 -4932 3412 -4468
rect 3446 -4680 3456 -4500
rect 3508 -4680 3518 -4500
rect 3460 -4888 3466 -4680
rect 3500 -4888 3506 -4680
rect 3460 -4900 3506 -4888
rect 3552 -4932 3672 -4468
rect 3718 -4512 3764 -4500
rect 3718 -4720 3724 -4512
rect 3758 -4720 3764 -4512
rect 3706 -4900 3716 -4720
rect 3768 -4900 3778 -4720
rect 3812 -4932 3932 -4468
rect 3962 -4680 3972 -4500
rect 4024 -4680 4034 -4500
rect 4234 -4512 4280 -4500
rect 3976 -4888 3982 -4680
rect 4016 -4888 4022 -4680
rect 4234 -4720 4240 -4512
rect 4274 -4720 4280 -4512
rect 3976 -4900 4022 -4888
rect 4222 -4900 4232 -4720
rect 4284 -4900 4294 -4720
rect -2412 -4936 -1172 -4932
rect -612 -4936 628 -4932
rect 1188 -4936 2428 -4932
rect 2988 -4936 4228 -4932
rect -2416 -4938 -1172 -4936
rect -2416 -4972 -2388 -4938
rect -2220 -4972 -2130 -4938
rect -1962 -4972 -1872 -4938
rect -1704 -4972 -1614 -4938
rect -1446 -4972 -1356 -4938
rect -1188 -4972 -1172 -4938
rect -2416 -5046 -1172 -4972
rect -2416 -5080 -2388 -5046
rect -2220 -5080 -2130 -5046
rect -1962 -5080 -1872 -5046
rect -1704 -5080 -1614 -5046
rect -1446 -5080 -1356 -5046
rect -1188 -5080 -1172 -5046
rect -2416 -5084 -1172 -5080
rect -616 -4938 628 -4936
rect -616 -4972 -588 -4938
rect -420 -4972 -330 -4938
rect -162 -4972 -72 -4938
rect 96 -4972 186 -4938
rect 354 -4972 444 -4938
rect 612 -4972 628 -4938
rect -616 -5046 628 -4972
rect -616 -5080 -588 -5046
rect -420 -5080 -330 -5046
rect -162 -5080 -72 -5046
rect 96 -5080 186 -5046
rect 354 -5080 444 -5046
rect 612 -5080 628 -5046
rect -616 -5084 628 -5080
rect 1184 -4938 2428 -4936
rect 1184 -4972 1212 -4938
rect 1380 -4972 1470 -4938
rect 1638 -4972 1728 -4938
rect 1896 -4972 1986 -4938
rect 2154 -4972 2244 -4938
rect 2412 -4972 2428 -4938
rect 1184 -5046 2428 -4972
rect 1184 -5080 1212 -5046
rect 1380 -5080 1470 -5046
rect 1638 -5080 1728 -5046
rect 1896 -5080 1986 -5046
rect 2154 -5080 2244 -5046
rect 2412 -5080 2428 -5046
rect 1184 -5084 2428 -5080
rect 2984 -4938 4228 -4936
rect 2984 -4972 3012 -4938
rect 3180 -4972 3270 -4938
rect 3438 -4972 3528 -4938
rect 3696 -4972 3786 -4938
rect 3954 -4972 4044 -4938
rect 4212 -4972 4228 -4938
rect 2984 -5046 4228 -4972
rect 2984 -5080 3012 -5046
rect 3180 -5080 3270 -5046
rect 3438 -5080 3528 -5046
rect 3696 -5080 3786 -5046
rect 3954 -5080 4044 -5046
rect 4212 -5080 4228 -5046
rect 2984 -5084 4228 -5080
rect -2400 -5086 -2208 -5084
rect -2142 -5086 -1950 -5084
rect -1884 -5086 -1692 -5084
rect -1626 -5086 -1434 -5084
rect -1368 -5086 -1176 -5084
rect -600 -5086 -408 -5084
rect -342 -5086 -150 -5084
rect -84 -5086 108 -5084
rect 174 -5086 366 -5084
rect 432 -5086 624 -5084
rect 1200 -5086 1392 -5084
rect 1458 -5086 1650 -5084
rect 1716 -5086 1908 -5084
rect 1974 -5086 2166 -5084
rect 2232 -5086 2424 -5084
rect 3000 -5086 3192 -5084
rect 3258 -5086 3450 -5084
rect 3516 -5086 3708 -5084
rect 3774 -5086 3966 -5084
rect 4032 -5086 4224 -5084
rect -2470 -5296 -2460 -5116
rect -2408 -5296 -2398 -5116
rect -2198 -5130 -2152 -5118
rect -2456 -5506 -2450 -5296
rect -2416 -5506 -2410 -5296
rect -2198 -5336 -2192 -5130
rect -2158 -5336 -2152 -5130
rect -2456 -5518 -2410 -5506
rect -2210 -5516 -2200 -5336
rect -2148 -5516 -2138 -5336
rect -2198 -5518 -2152 -5516
rect -2108 -5550 -1988 -5086
rect -1954 -5296 -1944 -5116
rect -1892 -5296 -1882 -5116
rect -1940 -5506 -1934 -5296
rect -1900 -5506 -1894 -5296
rect -1940 -5518 -1894 -5506
rect -1848 -5548 -1728 -5086
rect -1682 -5130 -1636 -5118
rect -1682 -5336 -1676 -5130
rect -1642 -5336 -1636 -5130
rect -1694 -5516 -1684 -5336
rect -1632 -5516 -1622 -5336
rect -1682 -5518 -1636 -5516
rect -1860 -5550 -1716 -5548
rect -1588 -5550 -1468 -5086
rect -1438 -5296 -1428 -5116
rect -1376 -5296 -1366 -5116
rect -1166 -5130 -1120 -5118
rect -1424 -5506 -1418 -5296
rect -1384 -5506 -1378 -5296
rect -1166 -5336 -1160 -5130
rect -1126 -5336 -1120 -5130
rect -670 -5296 -660 -5116
rect -608 -5296 -598 -5116
rect -398 -5130 -352 -5118
rect -1424 -5518 -1378 -5506
rect -1178 -5516 -1168 -5336
rect -1116 -5516 -1106 -5336
rect -656 -5506 -650 -5296
rect -616 -5506 -610 -5296
rect -398 -5336 -392 -5130
rect -358 -5336 -352 -5130
rect -1166 -5518 -1120 -5516
rect -656 -5518 -610 -5506
rect -410 -5516 -400 -5336
rect -348 -5516 -338 -5336
rect -398 -5518 -352 -5516
rect -308 -5550 -188 -5086
rect -154 -5296 -144 -5116
rect -92 -5296 -82 -5116
rect -140 -5506 -134 -5296
rect -100 -5506 -94 -5296
rect -140 -5518 -94 -5506
rect -48 -5548 72 -5086
rect 118 -5130 164 -5118
rect 118 -5336 124 -5130
rect 158 -5336 164 -5130
rect 106 -5516 116 -5336
rect 168 -5516 178 -5336
rect 118 -5518 164 -5516
rect -60 -5550 84 -5548
rect 212 -5550 332 -5086
rect 362 -5296 372 -5116
rect 424 -5296 434 -5116
rect 634 -5130 680 -5118
rect 376 -5506 382 -5296
rect 416 -5506 422 -5296
rect 634 -5336 640 -5130
rect 674 -5336 680 -5130
rect 1130 -5296 1140 -5116
rect 1192 -5296 1202 -5116
rect 1402 -5130 1448 -5118
rect 376 -5518 422 -5506
rect 622 -5516 632 -5336
rect 684 -5516 694 -5336
rect 1144 -5506 1150 -5296
rect 1184 -5506 1190 -5296
rect 1402 -5336 1408 -5130
rect 1442 -5336 1448 -5130
rect 634 -5518 680 -5516
rect 1144 -5518 1190 -5506
rect 1390 -5516 1400 -5336
rect 1452 -5516 1462 -5336
rect 1402 -5518 1448 -5516
rect 1492 -5550 1612 -5086
rect 1646 -5296 1656 -5116
rect 1708 -5296 1718 -5116
rect 1660 -5506 1666 -5296
rect 1700 -5506 1706 -5296
rect 1660 -5518 1706 -5506
rect 1752 -5548 1872 -5086
rect 1918 -5130 1964 -5118
rect 1918 -5336 1924 -5130
rect 1958 -5336 1964 -5130
rect 1906 -5516 1916 -5336
rect 1968 -5516 1978 -5336
rect 1918 -5518 1964 -5516
rect 1740 -5550 1884 -5548
rect 2012 -5550 2132 -5086
rect 2162 -5296 2172 -5116
rect 2224 -5296 2234 -5116
rect 2434 -5130 2480 -5118
rect 2176 -5506 2182 -5296
rect 2216 -5506 2222 -5296
rect 2434 -5336 2440 -5130
rect 2474 -5336 2480 -5130
rect 2930 -5296 2940 -5116
rect 2992 -5296 3002 -5116
rect 3202 -5130 3248 -5118
rect 2176 -5518 2222 -5506
rect 2422 -5516 2432 -5336
rect 2484 -5516 2494 -5336
rect 2944 -5506 2950 -5296
rect 2984 -5506 2990 -5296
rect 3202 -5336 3208 -5130
rect 3242 -5336 3248 -5130
rect 2434 -5518 2480 -5516
rect 2944 -5518 2990 -5506
rect 3190 -5516 3200 -5336
rect 3252 -5516 3262 -5336
rect 3202 -5518 3248 -5516
rect 3292 -5550 3412 -5086
rect 3446 -5296 3456 -5116
rect 3508 -5296 3518 -5116
rect 3460 -5506 3466 -5296
rect 3500 -5506 3506 -5296
rect 3460 -5518 3506 -5506
rect 3552 -5548 3672 -5086
rect 3718 -5130 3764 -5118
rect 3718 -5336 3724 -5130
rect 3758 -5336 3764 -5130
rect 3706 -5516 3716 -5336
rect 3768 -5516 3778 -5336
rect 3718 -5518 3764 -5516
rect 3540 -5550 3684 -5548
rect 3812 -5550 3932 -5086
rect 3962 -5296 3972 -5116
rect 4024 -5296 4034 -5116
rect 4234 -5130 4280 -5118
rect 3976 -5506 3982 -5296
rect 4016 -5506 4022 -5296
rect 4234 -5336 4240 -5130
rect 4274 -5336 4280 -5130
rect 3976 -5518 4022 -5506
rect 4222 -5516 4232 -5336
rect 4284 -5516 4294 -5336
rect 4234 -5518 4280 -5516
rect -2400 -5552 -2208 -5550
rect -2142 -5552 -1950 -5550
rect -1884 -5552 -1692 -5550
rect -1626 -5552 -1434 -5550
rect -1368 -5552 -1176 -5550
rect -600 -5552 -408 -5550
rect -342 -5552 -150 -5550
rect -84 -5552 108 -5550
rect 174 -5552 366 -5550
rect 432 -5552 624 -5550
rect 1200 -5552 1392 -5550
rect 1458 -5552 1650 -5550
rect 1716 -5552 1908 -5550
rect 1974 -5552 2166 -5550
rect 2232 -5552 2424 -5550
rect 3000 -5552 3192 -5550
rect 3258 -5552 3450 -5550
rect 3516 -5552 3708 -5550
rect 3774 -5552 3966 -5550
rect 4032 -5552 4224 -5550
rect -2412 -5556 -1172 -5552
rect -612 -5556 628 -5552
rect 1188 -5556 2428 -5552
rect 2988 -5556 4228 -5552
rect -2412 -5590 -2388 -5556
rect -2220 -5590 -2130 -5556
rect -1962 -5590 -1872 -5556
rect -1704 -5590 -1614 -5556
rect -1446 -5590 -1356 -5556
rect -1188 -5590 -1168 -5556
rect -2412 -5664 -1168 -5590
rect -2412 -5698 -2388 -5664
rect -2220 -5698 -2130 -5664
rect -1962 -5698 -1872 -5664
rect -1704 -5698 -1614 -5664
rect -1446 -5698 -1356 -5664
rect -1188 -5698 -1168 -5664
rect -2412 -5704 -1168 -5698
rect -612 -5590 -588 -5556
rect -420 -5590 -330 -5556
rect -162 -5590 -72 -5556
rect 96 -5590 186 -5556
rect 354 -5590 444 -5556
rect 612 -5590 632 -5556
rect -612 -5664 632 -5590
rect -612 -5698 -588 -5664
rect -420 -5698 -330 -5664
rect -162 -5698 -72 -5664
rect 96 -5698 186 -5664
rect 354 -5698 444 -5664
rect 612 -5698 632 -5664
rect -612 -5704 632 -5698
rect 1188 -5590 1212 -5556
rect 1380 -5590 1470 -5556
rect 1638 -5590 1728 -5556
rect 1896 -5590 1986 -5556
rect 2154 -5590 2244 -5556
rect 2412 -5590 2432 -5556
rect 1188 -5664 2432 -5590
rect 1188 -5698 1212 -5664
rect 1380 -5698 1470 -5664
rect 1638 -5698 1728 -5664
rect 1896 -5698 1986 -5664
rect 2154 -5698 2244 -5664
rect 2412 -5698 2432 -5664
rect 1188 -5704 2432 -5698
rect 2988 -5590 3012 -5556
rect 3180 -5590 3270 -5556
rect 3438 -5590 3528 -5556
rect 3696 -5590 3786 -5556
rect 3954 -5590 4044 -5556
rect 4212 -5590 4232 -5556
rect 2988 -5664 4232 -5590
rect 2988 -5698 3012 -5664
rect 3180 -5698 3270 -5664
rect 3438 -5698 3528 -5664
rect 3696 -5698 3786 -5664
rect 3954 -5698 4044 -5664
rect 4212 -5698 4232 -5664
rect 2988 -5704 4232 -5698
rect -2470 -5916 -2460 -5736
rect -2408 -5916 -2398 -5736
rect -2198 -5748 -2152 -5736
rect -2456 -6124 -2450 -5916
rect -2416 -6124 -2410 -5916
rect -2198 -5956 -2192 -5748
rect -2158 -5956 -2152 -5748
rect -2456 -6136 -2410 -6124
rect -2210 -6136 -2200 -5956
rect -2148 -6136 -2138 -5956
rect -2108 -6168 -1988 -5704
rect -1954 -5916 -1944 -5736
rect -1892 -5916 -1882 -5736
rect -1940 -6124 -1934 -5916
rect -1900 -6124 -1894 -5916
rect -1940 -6136 -1894 -6124
rect -1848 -6168 -1728 -5704
rect -1682 -5748 -1636 -5736
rect -1682 -5956 -1676 -5748
rect -1642 -5956 -1636 -5748
rect -1694 -6136 -1684 -5956
rect -1632 -6136 -1622 -5956
rect -1588 -6168 -1468 -5704
rect -1438 -5916 -1428 -5736
rect -1376 -5916 -1366 -5736
rect -1166 -5748 -1120 -5736
rect -1424 -6124 -1418 -5916
rect -1384 -6124 -1378 -5916
rect -1166 -5956 -1160 -5748
rect -1126 -5956 -1120 -5748
rect -670 -5916 -660 -5736
rect -608 -5916 -598 -5736
rect -398 -5748 -352 -5736
rect -1424 -6136 -1378 -6124
rect -1178 -6136 -1168 -5956
rect -1116 -6136 -1106 -5956
rect -656 -6124 -650 -5916
rect -616 -6124 -610 -5916
rect -398 -5956 -392 -5748
rect -358 -5956 -352 -5748
rect -656 -6136 -610 -6124
rect -410 -6136 -400 -5956
rect -348 -6136 -338 -5956
rect -308 -6168 -188 -5704
rect -154 -5916 -144 -5736
rect -92 -5916 -82 -5736
rect -140 -6124 -134 -5916
rect -100 -6124 -94 -5916
rect -140 -6136 -94 -6124
rect -48 -6168 72 -5704
rect 118 -5748 164 -5736
rect 118 -5956 124 -5748
rect 158 -5956 164 -5748
rect 106 -6136 116 -5956
rect 168 -6136 178 -5956
rect 212 -6168 332 -5704
rect 362 -5916 372 -5736
rect 424 -5916 434 -5736
rect 634 -5748 680 -5736
rect 376 -6124 382 -5916
rect 416 -6124 422 -5916
rect 634 -5956 640 -5748
rect 674 -5956 680 -5748
rect 1130 -5916 1140 -5736
rect 1192 -5916 1202 -5736
rect 1402 -5748 1448 -5736
rect 376 -6136 422 -6124
rect 622 -6136 632 -5956
rect 684 -6136 694 -5956
rect 1144 -6124 1150 -5916
rect 1184 -6124 1190 -5916
rect 1402 -5956 1408 -5748
rect 1442 -5956 1448 -5748
rect 1144 -6136 1190 -6124
rect 1390 -6136 1400 -5956
rect 1452 -6136 1462 -5956
rect 1492 -6168 1612 -5704
rect 1646 -5916 1656 -5736
rect 1708 -5916 1718 -5736
rect 1660 -6124 1666 -5916
rect 1700 -6124 1706 -5916
rect 1660 -6136 1706 -6124
rect 1752 -6168 1872 -5704
rect 1918 -5748 1964 -5736
rect 1918 -5956 1924 -5748
rect 1958 -5956 1964 -5748
rect 1906 -6136 1916 -5956
rect 1968 -6136 1978 -5956
rect 2012 -6168 2132 -5704
rect 2162 -5916 2172 -5736
rect 2224 -5916 2234 -5736
rect 2434 -5748 2480 -5736
rect 2176 -6124 2182 -5916
rect 2216 -6124 2222 -5916
rect 2434 -5956 2440 -5748
rect 2474 -5956 2480 -5748
rect 2930 -5916 2940 -5736
rect 2992 -5916 3002 -5736
rect 3202 -5748 3248 -5736
rect 2176 -6136 2222 -6124
rect 2422 -6136 2432 -5956
rect 2484 -6136 2494 -5956
rect 2944 -6124 2950 -5916
rect 2984 -6124 2990 -5916
rect 3202 -5956 3208 -5748
rect 3242 -5956 3248 -5748
rect 2944 -6136 2990 -6124
rect 3190 -6136 3200 -5956
rect 3252 -6136 3262 -5956
rect 3292 -6168 3412 -5704
rect 3446 -5916 3456 -5736
rect 3508 -5916 3518 -5736
rect 3460 -6124 3466 -5916
rect 3500 -6124 3506 -5916
rect 3460 -6136 3506 -6124
rect 3552 -6168 3672 -5704
rect 3718 -5748 3764 -5736
rect 3718 -5956 3724 -5748
rect 3758 -5956 3764 -5748
rect 3706 -6136 3716 -5956
rect 3768 -6136 3778 -5956
rect 3812 -6168 3932 -5704
rect 3962 -5916 3972 -5736
rect 4024 -5916 4034 -5736
rect 4234 -5748 4280 -5736
rect 3976 -6124 3982 -5916
rect 4016 -6124 4022 -5916
rect 4234 -5956 4240 -5748
rect 4274 -5956 4280 -5748
rect 3976 -6136 4022 -6124
rect 4222 -6136 4232 -5956
rect 4284 -6136 4294 -5956
rect -2412 -6172 -2208 -6168
rect -2416 -6174 -2208 -6172
rect -2416 -6208 -2388 -6174
rect -2220 -6204 -2208 -6174
rect -2142 -6174 -1692 -6168
rect -2142 -6204 -2130 -6174
rect -2220 -6208 -2130 -6204
rect -1962 -6208 -1872 -6174
rect -1704 -6204 -1692 -6174
rect -1626 -6174 -1176 -6168
rect -612 -6172 -408 -6168
rect -1626 -6204 -1614 -6174
rect -1704 -6208 -1614 -6204
rect -1446 -6208 -1356 -6174
rect -1188 -6204 -1176 -6174
rect -616 -6174 -408 -6172
rect -1188 -6208 -1172 -6204
rect -2416 -6282 -1172 -6208
rect -2416 -6316 -2388 -6282
rect -2220 -6316 -2130 -6282
rect -1962 -6316 -1872 -6282
rect -1704 -6316 -1614 -6282
rect -1446 -6316 -1356 -6282
rect -1188 -6316 -1172 -6282
rect -2416 -6320 -1172 -6316
rect -616 -6208 -588 -6174
rect -420 -6204 -408 -6174
rect -342 -6174 108 -6168
rect -342 -6204 -330 -6174
rect -420 -6208 -330 -6204
rect -162 -6208 -72 -6174
rect 96 -6204 108 -6174
rect 174 -6174 624 -6168
rect 1188 -6172 1392 -6168
rect 174 -6204 186 -6174
rect 96 -6208 186 -6204
rect 354 -6208 444 -6174
rect 612 -6204 624 -6174
rect 1184 -6174 1392 -6172
rect 612 -6208 628 -6204
rect -616 -6282 628 -6208
rect -616 -6316 -588 -6282
rect -420 -6316 -330 -6282
rect -162 -6316 -72 -6282
rect 96 -6316 186 -6282
rect 354 -6316 444 -6282
rect 612 -6316 628 -6282
rect -616 -6320 628 -6316
rect 1184 -6208 1212 -6174
rect 1380 -6204 1392 -6174
rect 1458 -6174 1908 -6168
rect 1458 -6204 1470 -6174
rect 1380 -6208 1470 -6204
rect 1638 -6208 1728 -6174
rect 1896 -6204 1908 -6174
rect 1974 -6174 2424 -6168
rect 2988 -6172 3192 -6168
rect 1974 -6204 1986 -6174
rect 1896 -6208 1986 -6204
rect 2154 -6208 2244 -6174
rect 2412 -6204 2424 -6174
rect 2984 -6174 3192 -6172
rect 2412 -6208 2428 -6204
rect 1184 -6282 2428 -6208
rect 1184 -6316 1212 -6282
rect 1380 -6316 1470 -6282
rect 1638 -6316 1728 -6282
rect 1896 -6316 1986 -6282
rect 2154 -6316 2244 -6282
rect 2412 -6316 2428 -6282
rect 1184 -6320 2428 -6316
rect 2984 -6208 3012 -6174
rect 3180 -6204 3192 -6174
rect 3258 -6174 3708 -6168
rect 3258 -6204 3270 -6174
rect 3180 -6208 3270 -6204
rect 3438 -6208 3528 -6174
rect 3696 -6204 3708 -6174
rect 3774 -6174 4224 -6168
rect 3774 -6204 3786 -6174
rect 3696 -6208 3786 -6204
rect 3954 -6208 4044 -6174
rect 4212 -6204 4224 -6174
rect 4212 -6208 4228 -6204
rect 2984 -6282 4228 -6208
rect 2984 -6316 3012 -6282
rect 3180 -6316 3270 -6282
rect 3438 -6316 3528 -6282
rect 3696 -6316 3786 -6282
rect 3954 -6316 4044 -6282
rect 4212 -6316 4228 -6282
rect 2984 -6320 4228 -6316
rect -2400 -6322 -2208 -6320
rect -2142 -6322 -1950 -6320
rect -1884 -6322 -1692 -6320
rect -1626 -6322 -1434 -6320
rect -1368 -6322 -1176 -6320
rect -600 -6322 -408 -6320
rect -342 -6322 -150 -6320
rect -84 -6322 108 -6320
rect 174 -6322 366 -6320
rect 432 -6322 624 -6320
rect 1200 -6322 1392 -6320
rect 1458 -6322 1650 -6320
rect 1716 -6322 1908 -6320
rect 1974 -6322 2166 -6320
rect 2232 -6322 2424 -6320
rect 3000 -6322 3192 -6320
rect 3258 -6322 3450 -6320
rect 3516 -6322 3708 -6320
rect 3774 -6322 3966 -6320
rect 4032 -6322 4224 -6320
rect -2470 -6532 -2460 -6352
rect -2408 -6532 -2398 -6352
rect -2198 -6366 -2152 -6354
rect -2456 -6742 -2450 -6532
rect -2416 -6742 -2410 -6532
rect -2198 -6572 -2192 -6366
rect -2158 -6572 -2152 -6366
rect -2456 -6754 -2410 -6742
rect -2210 -6752 -2200 -6572
rect -2148 -6752 -2138 -6572
rect -2198 -6754 -2152 -6752
rect -2108 -6786 -1988 -6322
rect -1860 -6324 -1716 -6322
rect -1954 -6532 -1944 -6352
rect -1892 -6532 -1882 -6352
rect -1940 -6742 -1934 -6532
rect -1900 -6742 -1894 -6532
rect -1940 -6754 -1894 -6742
rect -1848 -6786 -1728 -6324
rect -1682 -6366 -1636 -6354
rect -1682 -6572 -1676 -6366
rect -1642 -6572 -1636 -6366
rect -1694 -6752 -1684 -6572
rect -1632 -6752 -1622 -6572
rect -1682 -6754 -1636 -6752
rect -1588 -6786 -1468 -6322
rect -1438 -6532 -1428 -6352
rect -1376 -6532 -1366 -6352
rect -1166 -6366 -1120 -6354
rect -1424 -6742 -1418 -6532
rect -1384 -6742 -1378 -6532
rect -1166 -6572 -1160 -6366
rect -1126 -6572 -1120 -6366
rect -670 -6532 -660 -6352
rect -608 -6532 -598 -6352
rect -398 -6366 -352 -6354
rect -1424 -6754 -1378 -6742
rect -1178 -6752 -1168 -6572
rect -1116 -6752 -1106 -6572
rect -656 -6742 -650 -6532
rect -616 -6742 -610 -6532
rect -398 -6572 -392 -6366
rect -358 -6572 -352 -6366
rect -1166 -6754 -1120 -6752
rect -656 -6754 -610 -6742
rect -410 -6752 -400 -6572
rect -348 -6752 -338 -6572
rect -398 -6754 -352 -6752
rect -308 -6786 -188 -6322
rect -60 -6324 84 -6322
rect -154 -6532 -144 -6352
rect -92 -6532 -82 -6352
rect -140 -6742 -134 -6532
rect -100 -6742 -94 -6532
rect -140 -6754 -94 -6742
rect -48 -6786 72 -6324
rect 118 -6366 164 -6354
rect 118 -6572 124 -6366
rect 158 -6572 164 -6366
rect 106 -6752 116 -6572
rect 168 -6752 178 -6572
rect 118 -6754 164 -6752
rect 212 -6786 332 -6322
rect 362 -6532 372 -6352
rect 424 -6532 434 -6352
rect 634 -6366 680 -6354
rect 376 -6742 382 -6532
rect 416 -6742 422 -6532
rect 634 -6572 640 -6366
rect 674 -6572 680 -6366
rect 1130 -6532 1140 -6352
rect 1192 -6532 1202 -6352
rect 1402 -6366 1448 -6354
rect 376 -6754 422 -6742
rect 622 -6752 632 -6572
rect 684 -6752 694 -6572
rect 1144 -6742 1150 -6532
rect 1184 -6742 1190 -6532
rect 1402 -6572 1408 -6366
rect 1442 -6572 1448 -6366
rect 634 -6754 680 -6752
rect 1144 -6754 1190 -6742
rect 1390 -6752 1400 -6572
rect 1452 -6752 1462 -6572
rect 1402 -6754 1448 -6752
rect 1492 -6786 1612 -6322
rect 1740 -6324 1884 -6322
rect 1646 -6532 1656 -6352
rect 1708 -6532 1718 -6352
rect 1660 -6742 1666 -6532
rect 1700 -6742 1706 -6532
rect 1660 -6754 1706 -6742
rect 1752 -6786 1872 -6324
rect 1918 -6366 1964 -6354
rect 1918 -6572 1924 -6366
rect 1958 -6572 1964 -6366
rect 1906 -6752 1916 -6572
rect 1968 -6752 1978 -6572
rect 1918 -6754 1964 -6752
rect 2012 -6786 2132 -6322
rect 2162 -6532 2172 -6352
rect 2224 -6532 2234 -6352
rect 2434 -6366 2480 -6354
rect 2176 -6742 2182 -6532
rect 2216 -6742 2222 -6532
rect 2434 -6572 2440 -6366
rect 2474 -6572 2480 -6366
rect 2930 -6532 2940 -6352
rect 2992 -6532 3002 -6352
rect 3202 -6366 3248 -6354
rect 2176 -6754 2222 -6742
rect 2422 -6752 2432 -6572
rect 2484 -6752 2494 -6572
rect 2944 -6742 2950 -6532
rect 2984 -6742 2990 -6532
rect 3202 -6572 3208 -6366
rect 3242 -6572 3248 -6366
rect 2434 -6754 2480 -6752
rect 2944 -6754 2990 -6742
rect 3190 -6752 3200 -6572
rect 3252 -6752 3262 -6572
rect 3202 -6754 3248 -6752
rect 3292 -6786 3412 -6322
rect 3540 -6324 3684 -6322
rect 3446 -6532 3456 -6352
rect 3508 -6532 3518 -6352
rect 3460 -6742 3466 -6532
rect 3500 -6742 3506 -6532
rect 3460 -6754 3506 -6742
rect 3552 -6786 3672 -6324
rect 3718 -6366 3764 -6354
rect 3718 -6572 3724 -6366
rect 3758 -6572 3764 -6366
rect 3706 -6752 3716 -6572
rect 3768 -6752 3778 -6572
rect 3718 -6754 3764 -6752
rect 3812 -6786 3932 -6322
rect 3962 -6532 3972 -6352
rect 4024 -6532 4034 -6352
rect 4234 -6366 4280 -6354
rect 3976 -6742 3982 -6532
rect 4016 -6742 4022 -6532
rect 4234 -6572 4240 -6366
rect 4274 -6572 4280 -6366
rect 3976 -6754 4022 -6742
rect 4222 -6752 4232 -6572
rect 4284 -6752 4294 -6572
rect 4234 -6754 4280 -6752
rect -2400 -6788 -2208 -6786
rect -2142 -6788 -1950 -6786
rect -1884 -6788 -1692 -6786
rect -1626 -6788 -1434 -6786
rect -1368 -6788 -1176 -6786
rect -600 -6788 -408 -6786
rect -342 -6788 -150 -6786
rect -84 -6788 108 -6786
rect 174 -6788 366 -6786
rect 432 -6788 624 -6786
rect 1200 -6788 1392 -6786
rect 1458 -6788 1650 -6786
rect 1716 -6788 1908 -6786
rect 1974 -6788 2166 -6786
rect 2232 -6788 2424 -6786
rect 3000 -6788 3192 -6786
rect 3258 -6788 3450 -6786
rect 3516 -6788 3708 -6786
rect 3774 -6788 3966 -6786
rect 4032 -6788 4224 -6786
rect -2412 -6792 -1172 -6788
rect -612 -6792 628 -6788
rect 1188 -6792 2428 -6788
rect 2988 -6792 4228 -6788
rect -2412 -6826 -2388 -6792
rect -2220 -6826 -2130 -6792
rect -1962 -6826 -1872 -6792
rect -1704 -6826 -1614 -6792
rect -1446 -6826 -1356 -6792
rect -1188 -6826 -1168 -6792
rect -2412 -6900 -1168 -6826
rect -2412 -6934 -2388 -6900
rect -2220 -6934 -2130 -6900
rect -1962 -6934 -1872 -6900
rect -1704 -6934 -1614 -6900
rect -1446 -6934 -1356 -6900
rect -1188 -6934 -1168 -6900
rect -2412 -6940 -1168 -6934
rect -612 -6826 -588 -6792
rect -420 -6826 -330 -6792
rect -162 -6826 -72 -6792
rect 96 -6826 186 -6792
rect 354 -6826 444 -6792
rect 612 -6826 632 -6792
rect -612 -6900 632 -6826
rect -612 -6934 -588 -6900
rect -420 -6934 -330 -6900
rect -162 -6934 -72 -6900
rect 96 -6934 186 -6900
rect 354 -6934 444 -6900
rect 612 -6934 632 -6900
rect -612 -6940 632 -6934
rect 1188 -6826 1212 -6792
rect 1380 -6826 1470 -6792
rect 1638 -6826 1728 -6792
rect 1896 -6826 1986 -6792
rect 2154 -6826 2244 -6792
rect 2412 -6826 2432 -6792
rect 1188 -6900 2432 -6826
rect 1188 -6934 1212 -6900
rect 1380 -6934 1470 -6900
rect 1638 -6934 1728 -6900
rect 1896 -6934 1986 -6900
rect 2154 -6934 2244 -6900
rect 2412 -6934 2432 -6900
rect 1188 -6940 2432 -6934
rect 2988 -6826 3012 -6792
rect 3180 -6826 3270 -6792
rect 3438 -6826 3528 -6792
rect 3696 -6826 3786 -6792
rect 3954 -6826 4044 -6792
rect 4212 -6826 4232 -6792
rect 2988 -6900 4232 -6826
rect 2988 -6934 3012 -6900
rect 3180 -6934 3270 -6900
rect 3438 -6934 3528 -6900
rect 3696 -6934 3786 -6900
rect 3954 -6934 4044 -6900
rect 4212 -6934 4232 -6900
rect 2988 -6940 4232 -6934
rect -2470 -7152 -2460 -6972
rect -2408 -7152 -2398 -6972
rect -2198 -6984 -2152 -6972
rect -2456 -7360 -2450 -7152
rect -2416 -7360 -2410 -7152
rect -2198 -7192 -2192 -6984
rect -2158 -7192 -2152 -6984
rect -2456 -7372 -2410 -7360
rect -2210 -7372 -2200 -7192
rect -2148 -7372 -2138 -7192
rect -2108 -7404 -1988 -6940
rect -1954 -7152 -1944 -6972
rect -1892 -7152 -1882 -6972
rect -1940 -7360 -1934 -7152
rect -1900 -7360 -1894 -7152
rect -1940 -7372 -1894 -7360
rect -1848 -7404 -1728 -6940
rect -1682 -6984 -1636 -6972
rect -1682 -7192 -1676 -6984
rect -1642 -7192 -1636 -6984
rect -1694 -7372 -1684 -7192
rect -1632 -7372 -1622 -7192
rect -1588 -7404 -1468 -6940
rect -1438 -7152 -1428 -6972
rect -1376 -7152 -1366 -6972
rect -1166 -6984 -1120 -6972
rect -1424 -7360 -1418 -7152
rect -1384 -7360 -1378 -7152
rect -1166 -7192 -1160 -6984
rect -1126 -7192 -1120 -6984
rect -670 -7152 -660 -6972
rect -608 -7152 -598 -6972
rect -398 -6984 -352 -6972
rect -1424 -7372 -1378 -7360
rect -1178 -7372 -1168 -7192
rect -1116 -7372 -1106 -7192
rect -656 -7360 -650 -7152
rect -616 -7360 -610 -7152
rect -398 -7192 -392 -6984
rect -358 -7192 -352 -6984
rect -656 -7372 -610 -7360
rect -410 -7372 -400 -7192
rect -348 -7372 -338 -7192
rect -308 -7404 -188 -6940
rect -154 -7152 -144 -6972
rect -92 -7152 -82 -6972
rect -140 -7360 -134 -7152
rect -100 -7360 -94 -7152
rect -140 -7372 -94 -7360
rect -48 -7404 72 -6940
rect 118 -6984 164 -6972
rect 118 -7192 124 -6984
rect 158 -7192 164 -6984
rect 106 -7372 116 -7192
rect 168 -7372 178 -7192
rect 212 -7404 332 -6940
rect 362 -7152 372 -6972
rect 424 -7152 434 -6972
rect 634 -6984 680 -6972
rect 376 -7360 382 -7152
rect 416 -7360 422 -7152
rect 634 -7192 640 -6984
rect 674 -7192 680 -6984
rect 1130 -7152 1140 -6972
rect 1192 -7152 1202 -6972
rect 1402 -6984 1448 -6972
rect 376 -7372 422 -7360
rect 622 -7372 632 -7192
rect 684 -7372 694 -7192
rect 1144 -7360 1150 -7152
rect 1184 -7360 1190 -7152
rect 1402 -7192 1408 -6984
rect 1442 -7192 1448 -6984
rect 1144 -7372 1190 -7360
rect 1390 -7372 1400 -7192
rect 1452 -7372 1462 -7192
rect 1492 -7404 1612 -6940
rect 1646 -7152 1656 -6972
rect 1708 -7152 1718 -6972
rect 1660 -7360 1666 -7152
rect 1700 -7360 1706 -7152
rect 1660 -7372 1706 -7360
rect 1752 -7404 1872 -6940
rect 1918 -6984 1964 -6972
rect 1918 -7192 1924 -6984
rect 1958 -7192 1964 -6984
rect 1906 -7372 1916 -7192
rect 1968 -7372 1978 -7192
rect 2012 -7404 2132 -6940
rect 2162 -7152 2172 -6972
rect 2224 -7152 2234 -6972
rect 2434 -6984 2480 -6972
rect 2176 -7360 2182 -7152
rect 2216 -7360 2222 -7152
rect 2434 -7192 2440 -6984
rect 2474 -7192 2480 -6984
rect 2930 -7152 2940 -6972
rect 2992 -7152 3002 -6972
rect 3202 -6984 3248 -6972
rect 2176 -7372 2222 -7360
rect 2422 -7372 2432 -7192
rect 2484 -7372 2494 -7192
rect 2944 -7360 2950 -7152
rect 2984 -7360 2990 -7152
rect 3202 -7192 3208 -6984
rect 3242 -7192 3248 -6984
rect 2944 -7372 2990 -7360
rect 3190 -7372 3200 -7192
rect 3252 -7372 3262 -7192
rect 3292 -7404 3412 -6940
rect 3446 -7152 3456 -6972
rect 3508 -7152 3518 -6972
rect 3460 -7360 3466 -7152
rect 3500 -7360 3506 -7152
rect 3460 -7372 3506 -7360
rect 3552 -7404 3672 -6940
rect 3718 -6984 3764 -6972
rect 3718 -7192 3724 -6984
rect 3758 -7192 3764 -6984
rect 3706 -7372 3716 -7192
rect 3768 -7372 3778 -7192
rect 3812 -7404 3932 -6940
rect 3962 -7152 3972 -6972
rect 4024 -7152 4034 -6972
rect 4234 -6984 4280 -6972
rect 3976 -7360 3982 -7152
rect 4016 -7360 4022 -7152
rect 4234 -7192 4240 -6984
rect 4274 -7192 4280 -6984
rect 3976 -7372 4022 -7360
rect 4222 -7372 4232 -7192
rect 4284 -7372 4294 -7192
rect -2412 -7410 -2208 -7404
rect -2412 -7444 -2388 -7410
rect -2220 -7420 -2208 -7410
rect -2142 -7410 -1692 -7404
rect -2142 -7420 -2130 -7410
rect -2220 -7444 -2130 -7420
rect -1962 -7444 -1872 -7410
rect -1704 -7420 -1692 -7410
rect -1626 -7410 -1176 -7404
rect -1626 -7420 -1614 -7410
rect -1704 -7444 -1614 -7420
rect -1446 -7444 -1356 -7410
rect -1188 -7420 -1176 -7410
rect -612 -7410 -408 -7404
rect -1188 -7444 -1168 -7420
rect -2412 -7518 -1168 -7444
rect -2412 -7552 -2388 -7518
rect -2220 -7552 -2130 -7518
rect -1962 -7552 -1872 -7518
rect -1704 -7552 -1614 -7518
rect -1446 -7552 -1356 -7518
rect -1188 -7552 -1168 -7518
rect -2412 -7556 -1168 -7552
rect -612 -7444 -588 -7410
rect -420 -7420 -408 -7410
rect -342 -7410 108 -7404
rect -342 -7420 -330 -7410
rect -420 -7444 -330 -7420
rect -162 -7444 -72 -7410
rect 96 -7420 108 -7410
rect 174 -7410 624 -7404
rect 174 -7420 186 -7410
rect 96 -7444 186 -7420
rect 354 -7444 444 -7410
rect 612 -7420 624 -7410
rect 1188 -7410 1392 -7404
rect 612 -7444 632 -7420
rect -612 -7518 632 -7444
rect -612 -7552 -588 -7518
rect -420 -7552 -330 -7518
rect -162 -7552 -72 -7518
rect 96 -7552 186 -7518
rect 354 -7552 444 -7518
rect 612 -7552 632 -7518
rect -612 -7556 632 -7552
rect 1188 -7444 1212 -7410
rect 1380 -7420 1392 -7410
rect 1458 -7410 1908 -7404
rect 1458 -7420 1470 -7410
rect 1380 -7444 1470 -7420
rect 1638 -7444 1728 -7410
rect 1896 -7420 1908 -7410
rect 1974 -7410 2424 -7404
rect 1974 -7420 1986 -7410
rect 1896 -7444 1986 -7420
rect 2154 -7444 2244 -7410
rect 2412 -7420 2424 -7410
rect 2988 -7410 3192 -7404
rect 2412 -7444 2432 -7420
rect 1188 -7518 2432 -7444
rect 1188 -7552 1212 -7518
rect 1380 -7552 1470 -7518
rect 1638 -7552 1728 -7518
rect 1896 -7552 1986 -7518
rect 2154 -7552 2244 -7518
rect 2412 -7552 2432 -7518
rect 1188 -7556 2432 -7552
rect 2988 -7444 3012 -7410
rect 3180 -7420 3192 -7410
rect 3258 -7410 3708 -7404
rect 3258 -7420 3270 -7410
rect 3180 -7444 3270 -7420
rect 3438 -7444 3528 -7410
rect 3696 -7420 3708 -7410
rect 3774 -7410 4224 -7404
rect 3774 -7420 3786 -7410
rect 3696 -7444 3786 -7420
rect 3954 -7444 4044 -7410
rect 4212 -7420 4224 -7410
rect 4212 -7444 4232 -7420
rect 2988 -7518 4232 -7444
rect 2988 -7552 3012 -7518
rect 3180 -7552 3270 -7518
rect 3438 -7552 3528 -7518
rect 3696 -7552 3786 -7518
rect 3954 -7552 4044 -7518
rect 4212 -7552 4232 -7518
rect 2988 -7556 4232 -7552
rect -2400 -7558 -2208 -7556
rect -2142 -7558 -1950 -7556
rect -1884 -7558 -1692 -7556
rect -1626 -7558 -1434 -7556
rect -1368 -7558 -1176 -7556
rect -600 -7558 -408 -7556
rect -342 -7558 -150 -7556
rect -84 -7558 108 -7556
rect 174 -7558 366 -7556
rect 432 -7558 624 -7556
rect 1200 -7558 1392 -7556
rect 1458 -7558 1650 -7556
rect 1716 -7558 1908 -7556
rect 1974 -7558 2166 -7556
rect 2232 -7558 2424 -7556
rect 3000 -7558 3192 -7556
rect 3258 -7558 3450 -7556
rect 3516 -7558 3708 -7556
rect 3774 -7558 3966 -7556
rect 4032 -7558 4224 -7556
rect -2470 -7768 -2460 -7588
rect -2408 -7768 -2398 -7588
rect -2198 -7602 -2152 -7590
rect -2456 -7978 -2450 -7768
rect -2416 -7978 -2410 -7768
rect -2198 -7808 -2192 -7602
rect -2158 -7808 -2152 -7602
rect -2456 -7990 -2410 -7978
rect -2210 -7988 -2200 -7808
rect -2148 -7988 -2138 -7808
rect -2198 -7990 -2152 -7988
rect -2108 -8020 -1988 -7558
rect -1954 -7768 -1944 -7588
rect -1892 -7768 -1882 -7588
rect -1940 -7978 -1934 -7768
rect -1900 -7978 -1894 -7768
rect -1940 -7990 -1894 -7978
rect -1848 -8020 -1728 -7558
rect -1682 -7602 -1636 -7590
rect -1682 -7808 -1676 -7602
rect -1642 -7808 -1636 -7602
rect -1694 -7988 -1684 -7808
rect -1632 -7988 -1622 -7808
rect -1682 -7990 -1636 -7988
rect -1588 -8020 -1468 -7558
rect -1438 -7768 -1428 -7588
rect -1376 -7768 -1366 -7588
rect -1166 -7602 -1120 -7590
rect -1424 -7978 -1418 -7768
rect -1384 -7978 -1378 -7768
rect -1166 -7808 -1160 -7602
rect -1126 -7808 -1120 -7602
rect -670 -7768 -660 -7588
rect -608 -7768 -598 -7588
rect -398 -7602 -352 -7590
rect -1424 -7990 -1378 -7978
rect -1178 -7988 -1168 -7808
rect -1116 -7988 -1106 -7808
rect -986 -7960 -794 -7948
rect -1166 -7990 -1120 -7988
rect -2412 -8028 -1172 -8020
rect -2412 -8062 -2388 -8028
rect -2220 -8062 -2130 -8028
rect -1962 -8062 -1872 -8028
rect -1704 -8062 -1614 -8028
rect -1446 -8062 -1356 -8028
rect -1188 -8062 -1172 -8028
rect -2412 -8080 -1172 -8062
rect -990 -8160 -980 -7960
rect -800 -8160 -790 -7960
rect -656 -7978 -650 -7768
rect -616 -7978 -610 -7768
rect -398 -7808 -392 -7602
rect -358 -7808 -352 -7602
rect -656 -7990 -610 -7978
rect -410 -7988 -400 -7808
rect -348 -7988 -338 -7808
rect -398 -7990 -352 -7988
rect -308 -8020 -188 -7558
rect -154 -7768 -144 -7588
rect -92 -7768 -82 -7588
rect -140 -7978 -134 -7768
rect -100 -7978 -94 -7768
rect -140 -7990 -94 -7978
rect -48 -8020 72 -7558
rect 118 -7602 164 -7590
rect 118 -7808 124 -7602
rect 158 -7808 164 -7602
rect 106 -7988 116 -7808
rect 168 -7988 178 -7808
rect 118 -7990 164 -7988
rect 212 -8020 332 -7558
rect 362 -7768 372 -7588
rect 424 -7768 434 -7588
rect 634 -7602 680 -7590
rect 376 -7978 382 -7768
rect 416 -7978 422 -7768
rect 634 -7808 640 -7602
rect 674 -7808 680 -7602
rect 1130 -7768 1140 -7588
rect 1192 -7768 1202 -7588
rect 1402 -7602 1448 -7590
rect 376 -7990 422 -7978
rect 622 -7988 632 -7808
rect 684 -7988 694 -7808
rect 1144 -7978 1150 -7768
rect 1184 -7978 1190 -7768
rect 1402 -7808 1408 -7602
rect 1442 -7808 1448 -7602
rect 634 -7990 680 -7988
rect 1144 -7990 1190 -7978
rect 1390 -7988 1400 -7808
rect 1452 -7988 1462 -7808
rect 1402 -7990 1448 -7988
rect 1492 -8020 1612 -7558
rect 1646 -7768 1656 -7588
rect 1708 -7768 1718 -7588
rect 1660 -7978 1666 -7768
rect 1700 -7978 1706 -7768
rect 1660 -7990 1706 -7978
rect 1752 -8020 1872 -7558
rect 1918 -7602 1964 -7590
rect 1918 -7808 1924 -7602
rect 1958 -7808 1964 -7602
rect 1906 -7988 1916 -7808
rect 1968 -7988 1978 -7808
rect 1918 -7990 1964 -7988
rect 2012 -8020 2132 -7558
rect 2162 -7768 2172 -7588
rect 2224 -7768 2234 -7588
rect 2434 -7602 2480 -7590
rect 2176 -7978 2182 -7768
rect 2216 -7978 2222 -7768
rect 2434 -7808 2440 -7602
rect 2474 -7808 2480 -7602
rect 2930 -7768 2940 -7588
rect 2992 -7768 3002 -7588
rect 3202 -7602 3248 -7590
rect 2176 -7990 2222 -7978
rect 2422 -7988 2432 -7808
rect 2484 -7988 2494 -7808
rect 2944 -7978 2950 -7768
rect 2984 -7978 2990 -7768
rect 3202 -7808 3208 -7602
rect 3242 -7808 3248 -7602
rect 2434 -7990 2480 -7988
rect 2944 -7990 2990 -7978
rect 3190 -7988 3200 -7808
rect 3252 -7988 3262 -7808
rect 3202 -7990 3248 -7988
rect 3292 -8020 3412 -7558
rect 3446 -7768 3456 -7588
rect 3508 -7768 3518 -7588
rect 3460 -7978 3466 -7768
rect 3500 -7978 3506 -7768
rect 3460 -7990 3506 -7978
rect 3552 -8020 3672 -7558
rect 3718 -7602 3764 -7590
rect 3718 -7808 3724 -7602
rect 3758 -7808 3764 -7602
rect 3706 -7988 3716 -7808
rect 3768 -7988 3778 -7808
rect 3718 -7990 3764 -7988
rect 3812 -8020 3932 -7558
rect 3962 -7768 3972 -7588
rect 4024 -7768 4034 -7588
rect 4234 -7602 4280 -7590
rect 3976 -7978 3982 -7768
rect 4016 -7978 4022 -7768
rect 4234 -7808 4240 -7602
rect 4274 -7808 4280 -7602
rect 3976 -7990 4022 -7978
rect 4222 -7988 4232 -7808
rect 4284 -7988 4294 -7808
rect 4234 -7990 4280 -7988
rect -612 -8028 628 -8020
rect -612 -8062 -588 -8028
rect -420 -8062 -330 -8028
rect -162 -8062 -72 -8028
rect 96 -8062 186 -8028
rect 354 -8062 444 -8028
rect 612 -8062 628 -8028
rect -612 -8080 628 -8062
rect 1188 -8028 2428 -8020
rect 1188 -8062 1212 -8028
rect 1380 -8062 1470 -8028
rect 1638 -8062 1728 -8028
rect 1896 -8062 1986 -8028
rect 2154 -8062 2244 -8028
rect 2412 -8062 2428 -8028
rect 1188 -8080 2428 -8062
rect 2988 -8028 4228 -8020
rect 2988 -8062 3012 -8028
rect 3180 -8062 3270 -8028
rect 3438 -8062 3528 -8028
rect 3696 -8062 3786 -8028
rect 3954 -8062 4044 -8028
rect 4212 -8062 4228 -8028
rect 2988 -8080 4228 -8062
rect -986 -8172 -794 -8160
rect -5454 -9416 -5444 -8610
rect -4636 -9416 -4626 -8610
<< via1 >>
rect 3420 2380 3600 2580
rect -80 2092 2096 2112
rect -80 1695 -58 2092
rect -58 1695 192 2092
rect 192 1695 320 2092
rect 320 1695 570 2092
rect 570 1695 698 2092
rect 698 1695 948 2092
rect 948 1695 1076 2092
rect 1076 1695 1326 2092
rect 1326 1695 1454 2092
rect 1454 1695 1704 2092
rect 1704 1695 1832 2092
rect 1832 1695 2082 2092
rect 2082 1695 2096 2092
rect -80 1676 2096 1695
rect 2536 2043 2592 2056
rect 2536 1876 2546 2043
rect 2546 1876 2580 2043
rect 2580 1876 2592 2043
rect 2440 1667 2450 1832
rect 2450 1667 2484 1832
rect 2484 1667 2496 1832
rect 2440 1652 2496 1667
rect 2728 2043 2784 2056
rect 2728 1876 2738 2043
rect 2738 1876 2772 2043
rect 2772 1876 2784 2043
rect 2632 1667 2642 1832
rect 2642 1667 2676 1832
rect 2676 1667 2688 1832
rect 2632 1652 2688 1667
rect 2920 2043 2976 2056
rect 2920 1876 2930 2043
rect 2930 1876 2964 2043
rect 2964 1876 2976 2043
rect 2824 1667 2834 1832
rect 2834 1667 2868 1832
rect 2868 1667 2880 1832
rect 2824 1652 2880 1667
rect 3112 2043 3168 2056
rect 3112 1876 3122 2043
rect 3122 1876 3156 2043
rect 3156 1876 3168 2043
rect 3016 1667 3026 1832
rect 3026 1667 3060 1832
rect 3060 1667 3072 1832
rect 3016 1652 3072 1667
rect 3304 2043 3360 2056
rect 3304 1876 3314 2043
rect 3314 1876 3348 2043
rect 3348 1876 3360 2043
rect 3208 1667 3218 1832
rect 3218 1667 3252 1832
rect 3252 1667 3264 1832
rect 3208 1652 3264 1667
rect 3496 2043 3552 2056
rect 3496 1876 3506 2043
rect 3506 1876 3540 2043
rect 3540 1876 3552 2043
rect 3400 1667 3410 1832
rect 3410 1667 3444 1832
rect 3444 1667 3456 1832
rect 3400 1652 3456 1667
rect 3688 2043 3744 2056
rect 3688 1876 3698 2043
rect 3698 1876 3732 2043
rect 3732 1876 3744 2043
rect 3592 1667 3602 1832
rect 3602 1667 3636 1832
rect 3636 1667 3648 1832
rect 3592 1652 3648 1667
rect 3880 2043 3936 2056
rect 3880 1876 3890 2043
rect 3890 1876 3924 2043
rect 3924 1876 3936 2043
rect 3784 1667 3794 1832
rect 3794 1667 3828 1832
rect 3828 1667 3840 1832
rect 3784 1652 3840 1667
rect 4072 2043 4128 2056
rect 4072 1876 4082 2043
rect 4082 1876 4116 2043
rect 4116 1876 4128 2043
rect 3976 1667 3986 1832
rect 3986 1667 4020 1832
rect 4020 1667 4032 1832
rect 3976 1652 4032 1667
rect 4264 2043 4320 2056
rect 4264 1876 4274 2043
rect 4274 1876 4308 2043
rect 4308 1876 4320 2043
rect 4168 1667 4178 1832
rect 4178 1667 4212 1832
rect 4212 1667 4224 1832
rect 4168 1652 4224 1667
rect 4360 1667 4370 1832
rect 4370 1667 4404 1832
rect 4404 1667 4416 1832
rect 4360 1652 4416 1667
rect 5036 2022 5092 2036
rect 5036 1852 5046 2022
rect 5046 1852 5080 2022
rect 5080 1852 5092 2022
rect 4940 1646 4950 1816
rect 4950 1646 4984 1816
rect 4984 1646 4996 1816
rect 4940 1632 4996 1646
rect 5228 2022 5284 2036
rect 5228 1852 5238 2022
rect 5238 1852 5272 2022
rect 5272 1852 5284 2022
rect 5132 1646 5142 1816
rect 5142 1646 5176 1816
rect 5176 1646 5188 1816
rect 5132 1632 5188 1646
rect 5420 2022 5476 2036
rect 5420 1852 5430 2022
rect 5430 1852 5464 2022
rect 5464 1852 5476 2022
rect 5324 1646 5334 1816
rect 5334 1646 5368 1816
rect 5368 1646 5380 1816
rect 5324 1632 5380 1646
rect 5612 2022 5668 2036
rect 5612 1852 5622 2022
rect 5622 1852 5656 2022
rect 5656 1852 5668 2022
rect 5516 1646 5526 1816
rect 5526 1646 5560 1816
rect 5560 1646 5572 1816
rect 5516 1632 5572 1646
rect 5804 2022 5860 2036
rect 5804 1852 5814 2022
rect 5814 1852 5848 2022
rect 5848 1852 5860 2022
rect 5708 1646 5718 1816
rect 5718 1646 5752 1816
rect 5752 1646 5764 1816
rect 5708 1632 5764 1646
rect 5996 2022 6052 2036
rect 5996 1852 6006 2022
rect 6006 1852 6040 2022
rect 6040 1852 6052 2022
rect 5900 1646 5910 1816
rect 5910 1646 5944 1816
rect 5944 1646 5956 1816
rect 5900 1632 5956 1646
rect 6188 2022 6244 2036
rect 6188 1852 6198 2022
rect 6198 1852 6232 2022
rect 6232 1852 6244 2022
rect 6092 1646 6102 1816
rect 6102 1646 6136 1816
rect 6136 1646 6148 1816
rect 6092 1632 6148 1646
rect 6380 2022 6436 2036
rect 6380 1852 6390 2022
rect 6390 1852 6424 2022
rect 6424 1852 6436 2022
rect 6284 1646 6294 1816
rect 6294 1646 6328 1816
rect 6328 1646 6340 1816
rect 6284 1632 6340 1646
rect 6572 2022 6628 2036
rect 6572 1852 6582 2022
rect 6582 1852 6616 2022
rect 6616 1852 6628 2022
rect 6476 1646 6486 1816
rect 6486 1646 6520 1816
rect 6520 1646 6532 1816
rect 6476 1632 6532 1646
rect 6764 2022 6820 2036
rect 6764 1852 6774 2022
rect 6774 1852 6808 2022
rect 6808 1852 6820 2022
rect 6668 1646 6678 1816
rect 6678 1646 6712 1816
rect 6712 1646 6724 1816
rect 6668 1632 6724 1646
rect 6860 1646 6870 1816
rect 6870 1646 6904 1816
rect 6904 1646 6916 1816
rect 6860 1632 6916 1646
rect 2536 1407 2592 1424
rect 2536 1244 2546 1407
rect 2546 1244 2580 1407
rect 2580 1244 2592 1407
rect 2440 1031 2450 1200
rect 2450 1031 2484 1200
rect 2484 1031 2496 1200
rect 2440 1020 2496 1031
rect 2728 1407 2784 1424
rect 2728 1244 2738 1407
rect 2738 1244 2772 1407
rect 2772 1244 2784 1407
rect 2632 1031 2642 1200
rect 2642 1031 2676 1200
rect 2676 1031 2688 1200
rect 2632 1020 2688 1031
rect 2920 1407 2976 1424
rect 2920 1244 2930 1407
rect 2930 1244 2964 1407
rect 2964 1244 2976 1407
rect 2824 1031 2834 1200
rect 2834 1031 2868 1200
rect 2868 1031 2880 1200
rect 2824 1020 2880 1031
rect 3112 1407 3168 1424
rect 3112 1244 3122 1407
rect 3122 1244 3156 1407
rect 3156 1244 3168 1407
rect 3016 1031 3026 1200
rect 3026 1031 3060 1200
rect 3060 1031 3072 1200
rect 3016 1020 3072 1031
rect 3304 1407 3360 1424
rect 3304 1244 3314 1407
rect 3314 1244 3348 1407
rect 3348 1244 3360 1407
rect 3208 1031 3218 1200
rect 3218 1031 3252 1200
rect 3252 1031 3264 1200
rect 3208 1020 3264 1031
rect 3496 1407 3552 1424
rect 3496 1244 3506 1407
rect 3506 1244 3540 1407
rect 3540 1244 3552 1407
rect 3400 1031 3410 1200
rect 3410 1031 3444 1200
rect 3444 1031 3456 1200
rect 3400 1020 3456 1031
rect 3688 1407 3744 1424
rect 3688 1244 3698 1407
rect 3698 1244 3732 1407
rect 3732 1244 3744 1407
rect 3592 1031 3602 1200
rect 3602 1031 3636 1200
rect 3636 1031 3648 1200
rect 3592 1020 3648 1031
rect 3880 1407 3936 1424
rect 3880 1244 3890 1407
rect 3890 1244 3924 1407
rect 3924 1244 3936 1407
rect 3784 1031 3794 1200
rect 3794 1031 3828 1200
rect 3828 1031 3840 1200
rect 3784 1020 3840 1031
rect 4072 1407 4128 1424
rect 4072 1244 4082 1407
rect 4082 1244 4116 1407
rect 4116 1244 4128 1407
rect 3976 1031 3986 1200
rect 3986 1031 4020 1200
rect 4020 1031 4032 1200
rect 3976 1020 4032 1031
rect 4264 1407 4320 1424
rect 4264 1244 4274 1407
rect 4274 1244 4308 1407
rect 4308 1244 4320 1407
rect 4168 1031 4178 1200
rect 4178 1031 4212 1200
rect 4212 1031 4224 1200
rect 4168 1020 4224 1031
rect 4360 1031 4370 1200
rect 4370 1031 4404 1200
rect 4404 1031 4416 1200
rect 4360 1020 4416 1031
rect 5036 1404 5092 1420
rect 5036 1236 5046 1404
rect 5046 1236 5080 1404
rect 5080 1236 5092 1404
rect 4940 1028 4950 1200
rect 4950 1028 4984 1200
rect 4984 1028 4996 1200
rect 4940 1016 4996 1028
rect 5228 1404 5284 1420
rect 5228 1236 5238 1404
rect 5238 1236 5272 1404
rect 5272 1236 5284 1404
rect 5132 1028 5142 1200
rect 5142 1028 5176 1200
rect 5176 1028 5188 1200
rect 5132 1016 5188 1028
rect 5420 1404 5476 1420
rect 5420 1236 5430 1404
rect 5430 1236 5464 1404
rect 5464 1236 5476 1404
rect 5324 1028 5334 1200
rect 5334 1028 5368 1200
rect 5368 1028 5380 1200
rect 5324 1016 5380 1028
rect 5612 1404 5668 1420
rect 5612 1236 5622 1404
rect 5622 1236 5656 1404
rect 5656 1236 5668 1404
rect 5516 1028 5526 1200
rect 5526 1028 5560 1200
rect 5560 1028 5572 1200
rect 5516 1016 5572 1028
rect 5804 1404 5860 1420
rect 5804 1236 5814 1404
rect 5814 1236 5848 1404
rect 5848 1236 5860 1404
rect 5708 1028 5718 1200
rect 5718 1028 5752 1200
rect 5752 1028 5764 1200
rect 5708 1016 5764 1028
rect 5996 1404 6052 1420
rect 5996 1236 6006 1404
rect 6006 1236 6040 1404
rect 6040 1236 6052 1404
rect 5900 1028 5910 1200
rect 5910 1028 5944 1200
rect 5944 1028 5956 1200
rect 5900 1016 5956 1028
rect 6188 1404 6244 1420
rect 6188 1236 6198 1404
rect 6198 1236 6232 1404
rect 6232 1236 6244 1404
rect 6092 1028 6102 1200
rect 6102 1028 6136 1200
rect 6136 1028 6148 1200
rect 6092 1016 6148 1028
rect 6380 1404 6436 1420
rect 6380 1236 6390 1404
rect 6390 1236 6424 1404
rect 6424 1236 6436 1404
rect 6284 1028 6294 1200
rect 6294 1028 6328 1200
rect 6328 1028 6340 1200
rect 6284 1016 6340 1028
rect 6572 1404 6628 1420
rect 6572 1236 6582 1404
rect 6582 1236 6616 1404
rect 6616 1236 6628 1404
rect 6476 1028 6486 1200
rect 6486 1028 6520 1200
rect 6520 1028 6532 1200
rect 6476 1016 6532 1028
rect 6764 1404 6820 1420
rect 6764 1236 6774 1404
rect 6774 1236 6808 1404
rect 6808 1236 6820 1404
rect 6668 1028 6678 1200
rect 6678 1028 6712 1200
rect 6712 1028 6724 1200
rect 6668 1016 6724 1028
rect 6860 1028 6870 1200
rect 6870 1028 6904 1200
rect 6904 1028 6916 1200
rect 6860 1016 6916 1028
rect 300 861 1760 864
rect 300 464 320 861
rect 320 464 570 861
rect 570 464 698 861
rect 698 464 948 861
rect 948 464 1076 861
rect 1076 464 1326 861
rect 1326 464 1454 861
rect 1454 464 1704 861
rect 1704 464 1760 861
rect 300 448 1760 464
rect 2144 152 2380 420
rect 216 14 272 28
rect 216 -152 226 14
rect 226 -152 260 14
rect 260 -152 272 14
rect 120 -362 130 -196
rect 130 -362 164 -196
rect 164 -362 176 -196
rect 120 -376 176 -362
rect 408 14 464 28
rect 408 -152 418 14
rect 418 -152 452 14
rect 452 -152 464 14
rect 312 -362 322 -196
rect 322 -362 356 -196
rect 356 -362 368 -196
rect 312 -376 368 -362
rect 600 14 656 28
rect 600 -152 610 14
rect 610 -152 644 14
rect 644 -152 656 14
rect 504 -362 514 -196
rect 514 -362 548 -196
rect 548 -362 560 -196
rect 504 -376 560 -362
rect 792 14 848 28
rect 792 -152 802 14
rect 802 -152 836 14
rect 836 -152 848 14
rect 696 -362 706 -196
rect 706 -362 740 -196
rect 740 -362 752 -196
rect 696 -376 752 -362
rect 984 14 1040 28
rect 984 -152 994 14
rect 994 -152 1028 14
rect 1028 -152 1040 14
rect 888 -362 898 -196
rect 898 -362 932 -196
rect 932 -362 944 -196
rect 888 -376 944 -362
rect 1176 14 1232 28
rect 1176 -152 1186 14
rect 1186 -152 1220 14
rect 1220 -152 1232 14
rect 1080 -362 1090 -196
rect 1090 -362 1124 -196
rect 1124 -362 1136 -196
rect 1080 -376 1136 -362
rect 1368 14 1424 28
rect 1368 -152 1378 14
rect 1378 -152 1412 14
rect 1412 -152 1424 14
rect 1272 -362 1282 -196
rect 1282 -362 1316 -196
rect 1316 -362 1328 -196
rect 1272 -376 1328 -362
rect 1560 14 1616 28
rect 1560 -152 1570 14
rect 1570 -152 1604 14
rect 1604 -152 1616 14
rect 1464 -362 1474 -196
rect 1474 -362 1508 -196
rect 1508 -362 1520 -196
rect 1464 -376 1520 -362
rect 1752 14 1808 28
rect 1752 -152 1762 14
rect 1762 -152 1796 14
rect 1796 -152 1808 14
rect 1656 -362 1666 -196
rect 1666 -362 1700 -196
rect 1700 -362 1712 -196
rect 1656 -376 1712 -362
rect 1944 14 2000 28
rect 1944 -152 1954 14
rect 1954 -152 1988 14
rect 1988 -152 2000 14
rect 1848 -362 1858 -196
rect 1858 -362 1892 -196
rect 1892 -362 1904 -196
rect 1848 -376 1904 -362
rect 2140 -120 2380 152
rect 2536 456 2592 472
rect 2536 292 2546 456
rect 2546 292 2580 456
rect 2580 292 2592 456
rect 2440 80 2450 248
rect 2450 80 2484 248
rect 2484 80 2496 248
rect 2440 68 2496 80
rect 2728 456 2784 472
rect 2728 292 2738 456
rect 2738 292 2772 456
rect 2772 292 2784 456
rect 2632 80 2642 248
rect 2642 80 2676 248
rect 2676 80 2688 248
rect 2632 68 2688 80
rect 2920 456 2976 472
rect 2920 292 2930 456
rect 2930 292 2964 456
rect 2964 292 2976 456
rect 2824 80 2834 248
rect 2834 80 2868 248
rect 2868 80 2880 248
rect 2824 68 2880 80
rect 3112 456 3168 472
rect 3112 292 3122 456
rect 3122 292 3156 456
rect 3156 292 3168 456
rect 3016 80 3026 248
rect 3026 80 3060 248
rect 3060 80 3072 248
rect 3016 68 3072 80
rect 3304 456 3360 472
rect 3304 292 3314 456
rect 3314 292 3348 456
rect 3348 292 3360 456
rect 3208 80 3218 248
rect 3218 80 3252 248
rect 3252 80 3264 248
rect 3208 68 3264 80
rect 3496 456 3552 472
rect 3496 292 3506 456
rect 3506 292 3540 456
rect 3540 292 3552 456
rect 3400 80 3410 248
rect 3410 80 3444 248
rect 3444 80 3456 248
rect 3400 68 3456 80
rect 3688 456 3744 472
rect 3688 292 3698 456
rect 3698 292 3732 456
rect 3732 292 3744 456
rect 3592 80 3602 248
rect 3602 80 3636 248
rect 3636 80 3648 248
rect 3592 68 3648 80
rect 3880 456 3936 472
rect 3880 292 3890 456
rect 3890 292 3924 456
rect 3924 292 3936 456
rect 3784 80 3794 248
rect 3794 80 3828 248
rect 3828 80 3840 248
rect 3784 68 3840 80
rect 4072 456 4128 472
rect 4072 292 4082 456
rect 4082 292 4116 456
rect 4116 292 4128 456
rect 3976 80 3986 248
rect 3986 80 4020 248
rect 4020 80 4032 248
rect 3976 68 4032 80
rect 4264 456 4320 472
rect 4264 292 4274 456
rect 4274 292 4308 456
rect 4308 292 4320 456
rect 4168 80 4178 248
rect 4178 80 4212 248
rect 4212 80 4224 248
rect 4168 68 4224 80
rect 4360 80 4370 248
rect 4370 80 4404 248
rect 4404 80 4416 248
rect 4360 68 4416 80
rect 2040 -362 2050 -196
rect 2050 -362 2084 -196
rect 2084 -362 2096 -196
rect 2040 -376 2096 -362
rect 2536 -162 2592 -148
rect 2536 -328 2546 -162
rect 2546 -328 2580 -162
rect 2580 -328 2592 -162
rect 2440 -538 2450 -372
rect 2450 -538 2484 -372
rect 2484 -538 2496 -372
rect 2440 -552 2496 -538
rect 2728 -162 2784 -148
rect 2728 -328 2738 -162
rect 2738 -328 2772 -162
rect 2772 -328 2784 -162
rect 2632 -538 2642 -372
rect 2642 -538 2676 -372
rect 2676 -538 2688 -372
rect 2632 -552 2688 -538
rect 2920 -162 2976 -148
rect 2920 -328 2930 -162
rect 2930 -328 2964 -162
rect 2964 -328 2976 -162
rect 2824 -538 2834 -372
rect 2834 -538 2868 -372
rect 2868 -538 2880 -372
rect 2824 -552 2880 -538
rect 3112 -162 3168 -148
rect 3112 -328 3122 -162
rect 3122 -328 3156 -162
rect 3156 -328 3168 -162
rect 3016 -538 3026 -372
rect 3026 -538 3060 -372
rect 3060 -538 3072 -372
rect 3016 -552 3072 -538
rect 3304 -162 3360 -148
rect 3304 -328 3314 -162
rect 3314 -328 3348 -162
rect 3348 -328 3360 -162
rect 3208 -538 3218 -372
rect 3218 -538 3252 -372
rect 3252 -538 3264 -372
rect 3208 -552 3264 -538
rect 3496 -162 3552 -148
rect 3496 -328 3506 -162
rect 3506 -328 3540 -162
rect 3540 -328 3552 -162
rect 3400 -538 3410 -372
rect 3410 -538 3444 -372
rect 3444 -538 3456 -372
rect 3400 -552 3456 -538
rect 3688 -162 3744 -148
rect 3688 -328 3698 -162
rect 3698 -328 3732 -162
rect 3732 -328 3744 -162
rect 3592 -538 3602 -372
rect 3602 -538 3636 -372
rect 3636 -538 3648 -372
rect 3592 -552 3648 -538
rect 3880 -162 3936 -148
rect 3880 -328 3890 -162
rect 3890 -328 3924 -162
rect 3924 -328 3936 -162
rect 3784 -538 3794 -372
rect 3794 -538 3828 -372
rect 3828 -538 3840 -372
rect 3784 -552 3840 -538
rect 4072 -162 4128 -148
rect 4072 -328 4082 -162
rect 4082 -328 4116 -162
rect 4116 -328 4128 -162
rect 3976 -538 3986 -372
rect 3986 -538 4020 -372
rect 4020 -538 4032 -372
rect 3976 -552 4032 -538
rect 4264 -162 4320 -148
rect 4264 -328 4274 -162
rect 4274 -328 4308 -162
rect 4308 -328 4320 -162
rect 4168 -538 4178 -372
rect 4178 -538 4212 -372
rect 4212 -538 4224 -372
rect 4168 -552 4224 -538
rect 4360 -538 4370 -372
rect 4370 -538 4404 -372
rect 4404 -538 4416 -372
rect 4360 -552 4416 -538
rect 216 -604 272 -588
rect 216 -768 226 -604
rect 226 -768 260 -604
rect 260 -768 272 -604
rect 120 -980 130 -812
rect 130 -980 164 -812
rect 164 -980 176 -812
rect 120 -992 176 -980
rect 408 -604 464 -588
rect 408 -768 418 -604
rect 418 -768 452 -604
rect 452 -768 464 -604
rect 312 -980 322 -812
rect 322 -980 356 -812
rect 356 -980 368 -812
rect 312 -992 368 -980
rect 600 -604 656 -588
rect 600 -768 610 -604
rect 610 -768 644 -604
rect 644 -768 656 -604
rect 504 -980 514 -812
rect 514 -980 548 -812
rect 548 -980 560 -812
rect 504 -992 560 -980
rect 792 -604 848 -588
rect 792 -768 802 -604
rect 802 -768 836 -604
rect 836 -768 848 -604
rect 696 -980 706 -812
rect 706 -980 740 -812
rect 740 -980 752 -812
rect 696 -992 752 -980
rect 984 -604 1040 -588
rect 984 -768 994 -604
rect 994 -768 1028 -604
rect 1028 -768 1040 -604
rect 888 -980 898 -812
rect 898 -980 932 -812
rect 932 -980 944 -812
rect 888 -992 944 -980
rect 1176 -604 1232 -588
rect 1176 -768 1186 -604
rect 1186 -768 1220 -604
rect 1220 -768 1232 -604
rect 1080 -980 1090 -812
rect 1090 -980 1124 -812
rect 1124 -980 1136 -812
rect 1080 -992 1136 -980
rect 1368 -604 1424 -588
rect 1368 -768 1378 -604
rect 1378 -768 1412 -604
rect 1412 -768 1424 -604
rect 1272 -980 1282 -812
rect 1282 -980 1316 -812
rect 1316 -980 1328 -812
rect 1272 -992 1328 -980
rect 1560 -604 1616 -588
rect 1560 -768 1570 -604
rect 1570 -768 1604 -604
rect 1604 -768 1616 -604
rect 1464 -980 1474 -812
rect 1474 -980 1508 -812
rect 1508 -980 1520 -812
rect 1464 -992 1520 -980
rect 1752 -604 1808 -588
rect 1752 -768 1762 -604
rect 1762 -768 1796 -604
rect 1796 -768 1808 -604
rect 1656 -980 1666 -812
rect 1666 -980 1700 -812
rect 1700 -980 1712 -812
rect 1656 -992 1712 -980
rect 1944 -604 2000 -588
rect 1944 -768 1954 -604
rect 1954 -768 1988 -604
rect 1988 -768 2000 -604
rect 1848 -980 1858 -812
rect 1858 -980 1892 -812
rect 1892 -980 1904 -812
rect 1848 -992 1904 -980
rect 2040 -980 2050 -812
rect 2050 -980 2084 -812
rect 2084 -980 2096 -812
rect 2040 -992 2096 -980
rect 2460 -1028 2688 -756
rect 216 -1222 272 -1208
rect 216 -1388 226 -1222
rect 226 -1388 260 -1222
rect 260 -1388 272 -1222
rect 120 -1598 130 -1432
rect 130 -1598 164 -1432
rect 164 -1598 176 -1432
rect 120 -1612 176 -1598
rect 408 -1222 464 -1208
rect 408 -1388 418 -1222
rect 418 -1388 452 -1222
rect 452 -1388 464 -1222
rect 312 -1598 322 -1432
rect 322 -1598 356 -1432
rect 356 -1598 368 -1432
rect 312 -1612 368 -1598
rect 600 -1222 656 -1208
rect 600 -1388 610 -1222
rect 610 -1388 644 -1222
rect 644 -1388 656 -1222
rect 504 -1598 514 -1432
rect 514 -1598 548 -1432
rect 548 -1598 560 -1432
rect 504 -1612 560 -1598
rect 792 -1222 848 -1208
rect 792 -1388 802 -1222
rect 802 -1388 836 -1222
rect 836 -1388 848 -1222
rect 696 -1598 706 -1432
rect 706 -1598 740 -1432
rect 740 -1598 752 -1432
rect 696 -1612 752 -1598
rect 984 -1222 1040 -1208
rect 984 -1388 994 -1222
rect 994 -1388 1028 -1222
rect 1028 -1388 1040 -1222
rect 888 -1598 898 -1432
rect 898 -1598 932 -1432
rect 932 -1598 944 -1432
rect 888 -1612 944 -1598
rect 1176 -1222 1232 -1208
rect 1176 -1388 1186 -1222
rect 1186 -1388 1220 -1222
rect 1220 -1388 1232 -1222
rect 1080 -1598 1090 -1432
rect 1090 -1598 1124 -1432
rect 1124 -1598 1136 -1432
rect 1080 -1612 1136 -1598
rect 1368 -1222 1424 -1208
rect 1368 -1388 1378 -1222
rect 1378 -1388 1412 -1222
rect 1412 -1388 1424 -1222
rect 1272 -1598 1282 -1432
rect 1282 -1598 1316 -1432
rect 1316 -1598 1328 -1432
rect 1272 -1612 1328 -1598
rect 1560 -1222 1616 -1208
rect 1560 -1388 1570 -1222
rect 1570 -1388 1604 -1222
rect 1604 -1388 1616 -1222
rect 1464 -1598 1474 -1432
rect 1474 -1598 1508 -1432
rect 1508 -1598 1520 -1432
rect 1464 -1612 1520 -1598
rect 1752 -1222 1808 -1208
rect 1752 -1388 1762 -1222
rect 1762 -1388 1796 -1222
rect 1796 -1388 1808 -1222
rect 1656 -1598 1666 -1432
rect 1666 -1598 1700 -1432
rect 1700 -1598 1712 -1432
rect 1656 -1612 1712 -1598
rect 1944 -1222 2000 -1208
rect 1944 -1388 1954 -1222
rect 1954 -1388 1988 -1222
rect 1988 -1388 2000 -1222
rect 1848 -1598 1858 -1432
rect 1858 -1598 1892 -1432
rect 1892 -1598 1904 -1432
rect 1848 -1612 1904 -1598
rect 2040 -1598 2050 -1432
rect 2050 -1598 2084 -1432
rect 2084 -1598 2096 -1432
rect 2040 -1612 2096 -1598
rect 3708 -1228 4400 -716
rect 5036 786 5092 800
rect 5036 616 5046 786
rect 5046 616 5080 786
rect 5080 616 5092 786
rect 4940 410 4950 580
rect 4950 410 4984 580
rect 4984 410 4996 580
rect 4940 396 4996 410
rect 5228 786 5284 800
rect 5228 616 5238 786
rect 5238 616 5272 786
rect 5272 616 5284 786
rect 5132 410 5142 580
rect 5142 410 5176 580
rect 5176 410 5188 580
rect 5132 396 5188 410
rect 5420 786 5476 800
rect 5420 616 5430 786
rect 5430 616 5464 786
rect 5464 616 5476 786
rect 5324 410 5334 580
rect 5334 410 5368 580
rect 5368 410 5380 580
rect 5324 396 5380 410
rect 5612 786 5668 800
rect 5612 616 5622 786
rect 5622 616 5656 786
rect 5656 616 5668 786
rect 5516 410 5526 580
rect 5526 410 5560 580
rect 5560 410 5572 580
rect 5516 396 5572 410
rect 5804 786 5860 800
rect 5804 616 5814 786
rect 5814 616 5848 786
rect 5848 616 5860 786
rect 5708 410 5718 580
rect 5718 410 5752 580
rect 5752 410 5764 580
rect 5708 396 5764 410
rect 5996 786 6052 800
rect 5996 616 6006 786
rect 6006 616 6040 786
rect 6040 616 6052 786
rect 5900 410 5910 580
rect 5910 410 5944 580
rect 5944 410 5956 580
rect 5900 396 5956 410
rect 6188 786 6244 800
rect 6188 616 6198 786
rect 6198 616 6232 786
rect 6232 616 6244 786
rect 6092 410 6102 580
rect 6102 410 6136 580
rect 6136 410 6148 580
rect 6092 396 6148 410
rect 6380 786 6436 800
rect 6380 616 6390 786
rect 6390 616 6424 786
rect 6424 616 6436 786
rect 6284 410 6294 580
rect 6294 410 6328 580
rect 6328 410 6340 580
rect 6284 396 6340 410
rect 6572 786 6628 800
rect 6572 616 6582 786
rect 6582 616 6616 786
rect 6616 616 6628 786
rect 6476 410 6486 580
rect 6486 410 6520 580
rect 6520 410 6532 580
rect 6476 396 6532 410
rect 6764 786 6820 800
rect 6764 616 6774 786
rect 6774 616 6808 786
rect 6808 616 6820 786
rect 6668 410 6678 580
rect 6678 410 6712 580
rect 6712 410 6724 580
rect 6668 396 6724 410
rect 6860 410 6870 580
rect 6870 410 6904 580
rect 6904 410 6916 580
rect 6860 396 6916 410
rect 5036 168 5092 184
rect 5036 0 5046 168
rect 5046 0 5080 168
rect 5080 0 5092 168
rect 4940 -208 4950 -36
rect 4950 -208 4984 -36
rect 4984 -208 4996 -36
rect 4940 -220 4996 -208
rect 5228 168 5284 184
rect 5228 0 5238 168
rect 5238 0 5272 168
rect 5272 0 5284 168
rect 5132 -208 5142 -36
rect 5142 -208 5176 -36
rect 5176 -208 5188 -36
rect 5132 -220 5188 -208
rect 5420 168 5476 184
rect 5420 0 5430 168
rect 5430 0 5464 168
rect 5464 0 5476 168
rect 5324 -208 5334 -36
rect 5334 -208 5368 -36
rect 5368 -208 5380 -36
rect 5324 -220 5380 -208
rect 5612 168 5668 184
rect 5612 0 5622 168
rect 5622 0 5656 168
rect 5656 0 5668 168
rect 5516 -208 5526 -36
rect 5526 -208 5560 -36
rect 5560 -208 5572 -36
rect 5516 -220 5572 -208
rect 5804 168 5860 184
rect 5804 0 5814 168
rect 5814 0 5848 168
rect 5848 0 5860 168
rect 5708 -208 5718 -36
rect 5718 -208 5752 -36
rect 5752 -208 5764 -36
rect 5708 -220 5764 -208
rect 5996 168 6052 184
rect 5996 0 6006 168
rect 6006 0 6040 168
rect 6040 0 6052 168
rect 5900 -208 5910 -36
rect 5910 -208 5944 -36
rect 5944 -208 5956 -36
rect 5900 -220 5956 -208
rect 6188 168 6244 184
rect 6188 0 6198 168
rect 6198 0 6232 168
rect 6232 0 6244 168
rect 6092 -208 6102 -36
rect 6102 -208 6136 -36
rect 6136 -208 6148 -36
rect 6092 -220 6148 -208
rect 6380 168 6436 184
rect 6380 0 6390 168
rect 6390 0 6424 168
rect 6424 0 6436 168
rect 6284 -208 6294 -36
rect 6294 -208 6328 -36
rect 6328 -208 6340 -36
rect 6284 -220 6340 -208
rect 6572 168 6628 184
rect 6572 0 6582 168
rect 6582 0 6616 168
rect 6616 0 6628 168
rect 6476 -208 6486 -36
rect 6486 -208 6520 -36
rect 6520 -208 6532 -36
rect 6476 -220 6532 -208
rect 6764 168 6820 184
rect 6764 0 6774 168
rect 6774 0 6808 168
rect 6808 0 6820 168
rect 6668 -208 6678 -36
rect 6678 -208 6712 -36
rect 6712 -208 6724 -36
rect 6668 -220 6724 -208
rect 6860 -208 6870 -36
rect 6870 -208 6904 -36
rect 6904 -208 6916 -36
rect 6860 -220 6916 -208
rect 5036 -450 5092 -436
rect 5036 -620 5046 -450
rect 5046 -620 5080 -450
rect 5080 -620 5092 -450
rect 4940 -826 4950 -656
rect 4950 -826 4984 -656
rect 4984 -826 4996 -656
rect 4940 -840 4996 -826
rect 5228 -450 5284 -436
rect 5228 -620 5238 -450
rect 5238 -620 5272 -450
rect 5272 -620 5284 -450
rect 5132 -826 5142 -656
rect 5142 -826 5176 -656
rect 5176 -826 5188 -656
rect 5132 -840 5188 -826
rect 5420 -450 5476 -436
rect 5420 -620 5430 -450
rect 5430 -620 5464 -450
rect 5464 -620 5476 -450
rect 5324 -826 5334 -656
rect 5334 -826 5368 -656
rect 5368 -826 5380 -656
rect 5324 -840 5380 -826
rect 5612 -450 5668 -436
rect 5612 -620 5622 -450
rect 5622 -620 5656 -450
rect 5656 -620 5668 -450
rect 5516 -826 5526 -656
rect 5526 -826 5560 -656
rect 5560 -826 5572 -656
rect 5516 -840 5572 -826
rect 5804 -450 5860 -436
rect 5804 -620 5814 -450
rect 5814 -620 5848 -450
rect 5848 -620 5860 -450
rect 5708 -826 5718 -656
rect 5718 -826 5752 -656
rect 5752 -826 5764 -656
rect 5708 -840 5764 -826
rect 5996 -450 6052 -436
rect 5996 -620 6006 -450
rect 6006 -620 6040 -450
rect 6040 -620 6052 -450
rect 5900 -826 5910 -656
rect 5910 -826 5944 -656
rect 5944 -826 5956 -656
rect 5900 -840 5956 -826
rect 6188 -450 6244 -436
rect 6188 -620 6198 -450
rect 6198 -620 6232 -450
rect 6232 -620 6244 -450
rect 6092 -826 6102 -656
rect 6102 -826 6136 -656
rect 6136 -826 6148 -656
rect 6092 -840 6148 -826
rect 6380 -450 6436 -436
rect 6380 -620 6390 -450
rect 6390 -620 6424 -450
rect 6424 -620 6436 -450
rect 6284 -826 6294 -656
rect 6294 -826 6328 -656
rect 6328 -826 6340 -656
rect 6284 -840 6340 -826
rect 6572 -450 6628 -436
rect 6572 -620 6582 -450
rect 6582 -620 6616 -450
rect 6616 -620 6628 -450
rect 6476 -826 6486 -656
rect 6486 -826 6520 -656
rect 6520 -826 6532 -656
rect 6476 -840 6532 -826
rect 6764 -450 6820 -436
rect 6764 -620 6774 -450
rect 6774 -620 6808 -450
rect 6808 -620 6820 -450
rect 6668 -826 6678 -656
rect 6678 -826 6712 -656
rect 6712 -826 6724 -656
rect 6668 -840 6724 -826
rect 6860 -826 6870 -656
rect 6870 -826 6904 -656
rect 6904 -826 6916 -656
rect 6860 -840 6916 -826
rect 5036 -1068 5092 -1052
rect 5036 -1236 5046 -1068
rect 5046 -1236 5080 -1068
rect 5080 -1236 5092 -1068
rect 4324 -1628 4852 -1300
rect 4940 -1444 4950 -1272
rect 4950 -1444 4984 -1272
rect 4984 -1444 4996 -1272
rect 4940 -1456 4996 -1444
rect 5228 -1068 5284 -1052
rect 5228 -1236 5238 -1068
rect 5238 -1236 5272 -1068
rect 5272 -1236 5284 -1068
rect 5132 -1444 5142 -1272
rect 5142 -1444 5176 -1272
rect 5176 -1444 5188 -1272
rect 5132 -1456 5188 -1444
rect 5420 -1068 5476 -1052
rect 5420 -1236 5430 -1068
rect 5430 -1236 5464 -1068
rect 5464 -1236 5476 -1068
rect 5324 -1444 5334 -1272
rect 5334 -1444 5368 -1272
rect 5368 -1444 5380 -1272
rect 5324 -1456 5380 -1444
rect 5612 -1068 5668 -1052
rect 5612 -1236 5622 -1068
rect 5622 -1236 5656 -1068
rect 5656 -1236 5668 -1068
rect 5516 -1444 5526 -1272
rect 5526 -1444 5560 -1272
rect 5560 -1444 5572 -1272
rect 5516 -1456 5572 -1444
rect 5804 -1068 5860 -1052
rect 5804 -1236 5814 -1068
rect 5814 -1236 5848 -1068
rect 5848 -1236 5860 -1068
rect 5708 -1444 5718 -1272
rect 5718 -1444 5752 -1272
rect 5752 -1444 5764 -1272
rect 5708 -1456 5764 -1444
rect 5996 -1068 6052 -1052
rect 5996 -1236 6006 -1068
rect 6006 -1236 6040 -1068
rect 6040 -1236 6052 -1068
rect 5900 -1444 5910 -1272
rect 5910 -1444 5944 -1272
rect 5944 -1444 5956 -1272
rect 5900 -1456 5956 -1444
rect 6188 -1068 6244 -1052
rect 6188 -1236 6198 -1068
rect 6198 -1236 6232 -1068
rect 6232 -1236 6244 -1068
rect 6092 -1444 6102 -1272
rect 6102 -1444 6136 -1272
rect 6136 -1444 6148 -1272
rect 6092 -1456 6148 -1444
rect 6380 -1068 6436 -1052
rect 6380 -1236 6390 -1068
rect 6390 -1236 6424 -1068
rect 6424 -1236 6436 -1068
rect 6284 -1444 6294 -1272
rect 6294 -1444 6328 -1272
rect 6328 -1444 6340 -1272
rect 6284 -1456 6340 -1444
rect 6572 -1068 6628 -1052
rect 6572 -1236 6582 -1068
rect 6582 -1236 6616 -1068
rect 6616 -1236 6628 -1068
rect 6476 -1444 6486 -1272
rect 6486 -1444 6520 -1272
rect 6520 -1444 6532 -1272
rect 6476 -1456 6532 -1444
rect 6764 -1068 6820 -1052
rect 6764 -1236 6774 -1068
rect 6774 -1236 6808 -1068
rect 6808 -1236 6820 -1068
rect 6668 -1444 6678 -1272
rect 6678 -1444 6712 -1272
rect 6712 -1444 6724 -1272
rect 6668 -1456 6724 -1444
rect 6860 -1444 6870 -1272
rect 6870 -1444 6904 -1272
rect 6904 -1444 6916 -1272
rect 6860 -1456 6916 -1444
rect 4284 -2072 4780 -1756
rect 5036 -1686 5092 -1672
rect 5036 -1856 5046 -1686
rect 5046 -1856 5080 -1686
rect 5080 -1856 5092 -1686
rect 4940 -2062 4950 -1892
rect 4950 -2062 4984 -1892
rect 4984 -2062 4996 -1892
rect 4940 -2076 4996 -2062
rect 5228 -1686 5284 -1672
rect 5228 -1856 5238 -1686
rect 5238 -1856 5272 -1686
rect 5272 -1856 5284 -1686
rect 5132 -2062 5142 -1892
rect 5142 -2062 5176 -1892
rect 5176 -2062 5188 -1892
rect 5132 -2076 5188 -2062
rect 5420 -1686 5476 -1672
rect 5420 -1856 5430 -1686
rect 5430 -1856 5464 -1686
rect 5464 -1856 5476 -1686
rect 5324 -2062 5334 -1892
rect 5334 -2062 5368 -1892
rect 5368 -2062 5380 -1892
rect 5324 -2076 5380 -2062
rect 5612 -1686 5668 -1672
rect 5612 -1856 5622 -1686
rect 5622 -1856 5656 -1686
rect 5656 -1856 5668 -1686
rect 5516 -2062 5526 -1892
rect 5526 -2062 5560 -1892
rect 5560 -2062 5572 -1892
rect 5516 -2076 5572 -2062
rect 5804 -1686 5860 -1672
rect 5804 -1856 5814 -1686
rect 5814 -1856 5848 -1686
rect 5848 -1856 5860 -1686
rect 5708 -2062 5718 -1892
rect 5718 -2062 5752 -1892
rect 5752 -2062 5764 -1892
rect 5708 -2076 5764 -2062
rect 5996 -1686 6052 -1672
rect 5996 -1856 6006 -1686
rect 6006 -1856 6040 -1686
rect 6040 -1856 6052 -1686
rect 5900 -2062 5910 -1892
rect 5910 -2062 5944 -1892
rect 5944 -2062 5956 -1892
rect 5900 -2076 5956 -2062
rect 6188 -1686 6244 -1672
rect 6188 -1856 6198 -1686
rect 6198 -1856 6232 -1686
rect 6232 -1856 6244 -1686
rect 6092 -2062 6102 -1892
rect 6102 -2062 6136 -1892
rect 6136 -2062 6148 -1892
rect 6092 -2076 6148 -2062
rect 6380 -1686 6436 -1672
rect 6380 -1856 6390 -1686
rect 6390 -1856 6424 -1686
rect 6424 -1856 6436 -1686
rect 6284 -2062 6294 -1892
rect 6294 -2062 6328 -1892
rect 6328 -2062 6340 -1892
rect 6284 -2076 6340 -2062
rect 6572 -1686 6628 -1672
rect 6572 -1856 6582 -1686
rect 6582 -1856 6616 -1686
rect 6616 -1856 6628 -1686
rect 6476 -2062 6486 -1892
rect 6486 -2062 6520 -1892
rect 6520 -2062 6532 -1892
rect 6476 -2076 6532 -2062
rect 6764 -1686 6820 -1672
rect 6764 -1856 6774 -1686
rect 6774 -1856 6808 -1686
rect 6808 -1856 6820 -1686
rect 6668 -2062 6678 -1892
rect 6678 -2062 6712 -1892
rect 6712 -2062 6724 -1892
rect 6668 -2076 6724 -2062
rect 6860 -2062 6870 -1892
rect 6870 -2062 6904 -1892
rect 6904 -2062 6916 -1892
rect 6860 -2076 6916 -2062
rect -2364 -2366 -2312 -2352
rect -2364 -2532 -2354 -2366
rect -2354 -2532 -2320 -2366
rect -2320 -2532 -2312 -2366
rect -2460 -2742 -2450 -2576
rect -2450 -2742 -2416 -2576
rect -2416 -2742 -2408 -2576
rect -2460 -2756 -2408 -2742
rect -2172 -2366 -2120 -2352
rect -2172 -2532 -2162 -2366
rect -2162 -2532 -2128 -2366
rect -2128 -2532 -2120 -2366
rect -2268 -2742 -2258 -2576
rect -2258 -2742 -2224 -2576
rect -2224 -2742 -2216 -2576
rect -2268 -2756 -2216 -2742
rect -1980 -2366 -1928 -2352
rect -1980 -2532 -1970 -2366
rect -1970 -2532 -1936 -2366
rect -1936 -2532 -1928 -2366
rect -2076 -2742 -2066 -2576
rect -2066 -2742 -2032 -2576
rect -2032 -2742 -2024 -2576
rect -2076 -2756 -2024 -2742
rect -1788 -2366 -1736 -2352
rect -1788 -2532 -1778 -2366
rect -1778 -2532 -1744 -2366
rect -1744 -2532 -1736 -2366
rect -1884 -2742 -1874 -2576
rect -1874 -2742 -1840 -2576
rect -1840 -2742 -1832 -2576
rect -1884 -2756 -1832 -2742
rect -1596 -2366 -1544 -2352
rect -1596 -2532 -1586 -2366
rect -1586 -2532 -1552 -2366
rect -1552 -2532 -1544 -2366
rect -1692 -2742 -1682 -2576
rect -1682 -2742 -1648 -2576
rect -1648 -2742 -1640 -2576
rect -1692 -2756 -1640 -2742
rect -1500 -2742 -1490 -2576
rect -1490 -2742 -1456 -2576
rect -1456 -2742 -1448 -2576
rect -1500 -2756 -1448 -2742
rect -564 -2366 -512 -2352
rect -564 -2532 -554 -2366
rect -554 -2532 -520 -2366
rect -520 -2532 -512 -2366
rect -660 -2742 -650 -2576
rect -650 -2742 -616 -2576
rect -616 -2742 -608 -2576
rect -660 -2756 -608 -2742
rect -372 -2366 -320 -2352
rect -372 -2532 -362 -2366
rect -362 -2532 -328 -2366
rect -328 -2532 -320 -2366
rect -468 -2742 -458 -2576
rect -458 -2742 -424 -2576
rect -424 -2742 -416 -2576
rect -468 -2756 -416 -2742
rect -180 -2366 -128 -2352
rect -180 -2532 -170 -2366
rect -170 -2532 -136 -2366
rect -136 -2532 -128 -2366
rect -276 -2742 -266 -2576
rect -266 -2742 -232 -2576
rect -232 -2742 -224 -2576
rect -276 -2756 -224 -2742
rect 12 -2366 64 -2352
rect 12 -2532 22 -2366
rect 22 -2532 56 -2366
rect 56 -2532 64 -2366
rect -84 -2742 -74 -2576
rect -74 -2742 -40 -2576
rect -40 -2742 -32 -2576
rect -84 -2756 -32 -2742
rect 204 -2366 256 -2352
rect 204 -2532 214 -2366
rect 214 -2532 248 -2366
rect 248 -2532 256 -2366
rect 108 -2742 118 -2576
rect 118 -2742 152 -2576
rect 152 -2742 160 -2576
rect 108 -2756 160 -2742
rect 300 -2742 310 -2576
rect 310 -2742 344 -2576
rect 344 -2742 352 -2576
rect 300 -2756 352 -2742
rect 1236 -2366 1288 -2352
rect 1236 -2532 1246 -2366
rect 1246 -2532 1280 -2366
rect 1280 -2532 1288 -2366
rect 1140 -2742 1150 -2576
rect 1150 -2742 1184 -2576
rect 1184 -2742 1192 -2576
rect 1140 -2756 1192 -2742
rect 1428 -2366 1480 -2352
rect 1428 -2532 1438 -2366
rect 1438 -2532 1472 -2366
rect 1472 -2532 1480 -2366
rect 1332 -2742 1342 -2576
rect 1342 -2742 1376 -2576
rect 1376 -2742 1384 -2576
rect 1332 -2756 1384 -2742
rect 1620 -2366 1672 -2352
rect 1620 -2532 1630 -2366
rect 1630 -2532 1664 -2366
rect 1664 -2532 1672 -2366
rect 1524 -2742 1534 -2576
rect 1534 -2742 1568 -2576
rect 1568 -2742 1576 -2576
rect 1524 -2756 1576 -2742
rect 1812 -2366 1864 -2352
rect 1812 -2532 1822 -2366
rect 1822 -2532 1856 -2366
rect 1856 -2532 1864 -2366
rect 1716 -2742 1726 -2576
rect 1726 -2742 1760 -2576
rect 1760 -2742 1768 -2576
rect 1716 -2756 1768 -2742
rect 2004 -2366 2056 -2352
rect 2004 -2532 2014 -2366
rect 2014 -2532 2048 -2366
rect 2048 -2532 2056 -2366
rect 1908 -2742 1918 -2576
rect 1918 -2742 1952 -2576
rect 1952 -2742 1960 -2576
rect 1908 -2756 1960 -2742
rect 2100 -2742 2110 -2576
rect 2110 -2742 2144 -2576
rect 2144 -2742 2152 -2576
rect 2100 -2756 2152 -2742
rect 3036 -2366 3088 -2352
rect 3036 -2532 3046 -2366
rect 3046 -2532 3080 -2366
rect 3080 -2532 3088 -2366
rect 2940 -2742 2950 -2576
rect 2950 -2742 2984 -2576
rect 2984 -2742 2992 -2576
rect 2940 -2756 2992 -2742
rect 3228 -2366 3280 -2352
rect 3228 -2532 3238 -2366
rect 3238 -2532 3272 -2366
rect 3272 -2532 3280 -2366
rect 3132 -2742 3142 -2576
rect 3142 -2742 3176 -2576
rect 3176 -2742 3184 -2576
rect 3132 -2756 3184 -2742
rect 3420 -2366 3472 -2352
rect 3420 -2532 3430 -2366
rect 3430 -2532 3464 -2366
rect 3464 -2532 3472 -2366
rect 3324 -2742 3334 -2576
rect 3334 -2742 3368 -2576
rect 3368 -2742 3376 -2576
rect 3324 -2756 3376 -2742
rect 3612 -2366 3664 -2352
rect 3612 -2532 3622 -2366
rect 3622 -2532 3656 -2366
rect 3656 -2532 3664 -2366
rect 3516 -2742 3526 -2576
rect 3526 -2742 3560 -2576
rect 3560 -2742 3568 -2576
rect 3516 -2756 3568 -2742
rect 3804 -2366 3856 -2352
rect 3804 -2532 3814 -2366
rect 3814 -2532 3848 -2366
rect 3848 -2532 3856 -2366
rect 3708 -2742 3718 -2576
rect 3718 -2742 3752 -2576
rect 3752 -2742 3760 -2576
rect 3708 -2756 3760 -2742
rect 3900 -2742 3910 -2576
rect 3910 -2742 3944 -2576
rect 3944 -2742 3952 -2576
rect 3900 -2756 3952 -2742
rect 4412 -2648 4696 -2148
rect 5036 -2304 5092 -2288
rect 5036 -2472 5046 -2304
rect 5046 -2472 5080 -2304
rect 5080 -2472 5092 -2304
rect -3080 -3828 -2648 -3136
rect -2364 -2984 -2312 -2968
rect -2364 -3148 -2354 -2984
rect -2354 -3148 -2320 -2984
rect -2320 -3148 -2312 -2984
rect -2460 -3360 -2450 -3192
rect -2450 -3360 -2416 -3192
rect -2416 -3360 -2408 -3192
rect -2460 -3372 -2408 -3360
rect -2172 -2984 -2120 -2968
rect -2172 -3148 -2162 -2984
rect -2162 -3148 -2128 -2984
rect -2128 -3148 -2120 -2984
rect -2268 -3360 -2258 -3192
rect -2258 -3360 -2224 -3192
rect -2224 -3360 -2216 -3192
rect -2268 -3372 -2216 -3360
rect -1980 -2984 -1928 -2968
rect -1980 -3148 -1970 -2984
rect -1970 -3148 -1936 -2984
rect -1936 -3148 -1928 -2984
rect -2076 -3360 -2066 -3192
rect -2066 -3360 -2032 -3192
rect -2032 -3360 -2024 -3192
rect -2076 -3372 -2024 -3360
rect -1788 -2984 -1736 -2968
rect -1788 -3148 -1778 -2984
rect -1778 -3148 -1744 -2984
rect -1744 -3148 -1736 -2984
rect -1884 -3360 -1874 -3192
rect -1874 -3360 -1840 -3192
rect -1840 -3360 -1832 -3192
rect -1884 -3372 -1832 -3360
rect -1596 -2984 -1544 -2968
rect -1596 -3148 -1586 -2984
rect -1586 -3148 -1552 -2984
rect -1552 -3148 -1544 -2984
rect -1692 -3360 -1682 -3192
rect -1682 -3360 -1648 -3192
rect -1648 -3360 -1640 -3192
rect -1692 -3372 -1640 -3360
rect -1500 -3360 -1490 -3192
rect -1490 -3360 -1456 -3192
rect -1456 -3360 -1448 -3192
rect -1500 -3372 -1448 -3360
rect -564 -2984 -512 -2968
rect -564 -3148 -554 -2984
rect -554 -3148 -520 -2984
rect -520 -3148 -512 -2984
rect -660 -3360 -650 -3192
rect -650 -3360 -616 -3192
rect -616 -3360 -608 -3192
rect -660 -3372 -608 -3360
rect -372 -2984 -320 -2968
rect -372 -3148 -362 -2984
rect -362 -3148 -328 -2984
rect -328 -3148 -320 -2984
rect -468 -3360 -458 -3192
rect -458 -3360 -424 -3192
rect -424 -3360 -416 -3192
rect -468 -3372 -416 -3360
rect -180 -2984 -128 -2968
rect -180 -3148 -170 -2984
rect -170 -3148 -136 -2984
rect -136 -3148 -128 -2984
rect -276 -3360 -266 -3192
rect -266 -3360 -232 -3192
rect -232 -3360 -224 -3192
rect -276 -3372 -224 -3360
rect 12 -2984 64 -2968
rect 12 -3148 22 -2984
rect 22 -3148 56 -2984
rect 56 -3148 64 -2984
rect -84 -3360 -74 -3192
rect -74 -3360 -40 -3192
rect -40 -3360 -32 -3192
rect -84 -3372 -32 -3360
rect 204 -2984 256 -2968
rect 204 -3148 214 -2984
rect 214 -3148 248 -2984
rect 248 -3148 256 -2984
rect 108 -3360 118 -3192
rect 118 -3360 152 -3192
rect 152 -3360 160 -3192
rect 108 -3372 160 -3360
rect 300 -3360 310 -3192
rect 310 -3360 344 -3192
rect 344 -3360 352 -3192
rect 300 -3372 352 -3360
rect 1236 -2984 1288 -2968
rect 1236 -3148 1246 -2984
rect 1246 -3148 1280 -2984
rect 1280 -3148 1288 -2984
rect 1140 -3360 1150 -3192
rect 1150 -3360 1184 -3192
rect 1184 -3360 1192 -3192
rect 1140 -3372 1192 -3360
rect 1428 -2984 1480 -2968
rect 1428 -3148 1438 -2984
rect 1438 -3148 1472 -2984
rect 1472 -3148 1480 -2984
rect 1332 -3360 1342 -3192
rect 1342 -3360 1376 -3192
rect 1376 -3360 1384 -3192
rect 1332 -3372 1384 -3360
rect 1620 -2984 1672 -2968
rect 1620 -3148 1630 -2984
rect 1630 -3148 1664 -2984
rect 1664 -3148 1672 -2984
rect 1524 -3360 1534 -3192
rect 1534 -3360 1568 -3192
rect 1568 -3360 1576 -3192
rect 1524 -3372 1576 -3360
rect 1812 -2984 1864 -2968
rect 1812 -3148 1822 -2984
rect 1822 -3148 1856 -2984
rect 1856 -3148 1864 -2984
rect 1716 -3360 1726 -3192
rect 1726 -3360 1760 -3192
rect 1760 -3360 1768 -3192
rect 1716 -3372 1768 -3360
rect 2004 -2984 2056 -2968
rect 2004 -3148 2014 -2984
rect 2014 -3148 2048 -2984
rect 2048 -3148 2056 -2984
rect 1908 -3360 1918 -3192
rect 1918 -3360 1952 -3192
rect 1952 -3360 1960 -3192
rect 1908 -3372 1960 -3360
rect 2100 -3360 2110 -3192
rect 2110 -3360 2144 -3192
rect 2144 -3360 2152 -3192
rect 2100 -3372 2152 -3360
rect 3036 -2984 3088 -2968
rect 3036 -3148 3046 -2984
rect 3046 -3148 3080 -2984
rect 3080 -3148 3088 -2984
rect 2940 -3360 2950 -3192
rect 2950 -3360 2984 -3192
rect 2984 -3360 2992 -3192
rect 2940 -3372 2992 -3360
rect 3228 -2984 3280 -2968
rect 3228 -3148 3238 -2984
rect 3238 -3148 3272 -2984
rect 3272 -3148 3280 -2984
rect 3132 -3360 3142 -3192
rect 3142 -3360 3176 -3192
rect 3176 -3360 3184 -3192
rect 3132 -3372 3184 -3360
rect 3420 -2984 3472 -2968
rect 3420 -3148 3430 -2984
rect 3430 -3148 3464 -2984
rect 3464 -3148 3472 -2984
rect 3324 -3360 3334 -3192
rect 3334 -3360 3368 -3192
rect 3368 -3360 3376 -3192
rect 3324 -3372 3376 -3360
rect 3612 -2984 3664 -2968
rect 3612 -3148 3622 -2984
rect 3622 -3148 3656 -2984
rect 3656 -3148 3664 -2984
rect 3516 -3360 3526 -3192
rect 3526 -3360 3560 -3192
rect 3560 -3360 3568 -3192
rect 3516 -3372 3568 -3360
rect 3804 -2984 3856 -2968
rect 3804 -3148 3814 -2984
rect 3814 -3148 3848 -2984
rect 3848 -3148 3856 -2984
rect 3708 -3360 3718 -3192
rect 3718 -3360 3752 -3192
rect 3752 -3360 3760 -3192
rect 3708 -3372 3760 -3360
rect 3900 -3360 3910 -3192
rect 3910 -3360 3944 -3192
rect 3944 -3360 3952 -3192
rect 3900 -3372 3952 -3360
rect 4940 -2680 4950 -2508
rect 4950 -2680 4984 -2508
rect 4984 -2680 4996 -2508
rect 4940 -2692 4996 -2680
rect 5228 -2304 5284 -2288
rect 5228 -2472 5238 -2304
rect 5238 -2472 5272 -2304
rect 5272 -2472 5284 -2304
rect 5132 -2680 5142 -2508
rect 5142 -2680 5176 -2508
rect 5176 -2680 5188 -2508
rect 5132 -2692 5188 -2680
rect 5420 -2304 5476 -2288
rect 5420 -2472 5430 -2304
rect 5430 -2472 5464 -2304
rect 5464 -2472 5476 -2304
rect 5324 -2680 5334 -2508
rect 5334 -2680 5368 -2508
rect 5368 -2680 5380 -2508
rect 5324 -2692 5380 -2680
rect 5612 -2304 5668 -2288
rect 5612 -2472 5622 -2304
rect 5622 -2472 5656 -2304
rect 5656 -2472 5668 -2304
rect 5516 -2680 5526 -2508
rect 5526 -2680 5560 -2508
rect 5560 -2680 5572 -2508
rect 5516 -2692 5572 -2680
rect 5804 -2304 5860 -2288
rect 5804 -2472 5814 -2304
rect 5814 -2472 5848 -2304
rect 5848 -2472 5860 -2304
rect 5708 -2680 5718 -2508
rect 5718 -2680 5752 -2508
rect 5752 -2680 5764 -2508
rect 5708 -2692 5764 -2680
rect 5996 -2304 6052 -2288
rect 5996 -2472 6006 -2304
rect 6006 -2472 6040 -2304
rect 6040 -2472 6052 -2304
rect 5900 -2680 5910 -2508
rect 5910 -2680 5944 -2508
rect 5944 -2680 5956 -2508
rect 5900 -2692 5956 -2680
rect 6188 -2304 6244 -2288
rect 6188 -2472 6198 -2304
rect 6198 -2472 6232 -2304
rect 6232 -2472 6244 -2304
rect 6092 -2680 6102 -2508
rect 6102 -2680 6136 -2508
rect 6136 -2680 6148 -2508
rect 6092 -2692 6148 -2680
rect 6380 -2304 6436 -2288
rect 6380 -2472 6390 -2304
rect 6390 -2472 6424 -2304
rect 6424 -2472 6436 -2304
rect 6284 -2680 6294 -2508
rect 6294 -2680 6328 -2508
rect 6328 -2680 6340 -2508
rect 6284 -2692 6340 -2680
rect 6572 -2304 6628 -2288
rect 6572 -2472 6582 -2304
rect 6582 -2472 6616 -2304
rect 6616 -2472 6628 -2304
rect 6476 -2680 6486 -2508
rect 6486 -2680 6520 -2508
rect 6520 -2680 6532 -2508
rect 6476 -2692 6532 -2680
rect 6764 -2304 6820 -2288
rect 6764 -2472 6774 -2304
rect 6774 -2472 6808 -2304
rect 6808 -2472 6820 -2304
rect 6668 -2680 6678 -2508
rect 6678 -2680 6712 -2508
rect 6712 -2680 6724 -2508
rect 6668 -2692 6724 -2680
rect 6860 -2680 6870 -2508
rect 6870 -2680 6904 -2508
rect 6904 -2680 6916 -2508
rect 6860 -2692 6916 -2680
rect 5036 -2922 5092 -2908
rect 5036 -3092 5046 -2922
rect 5046 -3092 5080 -2922
rect 5080 -3092 5092 -2922
rect 4940 -3298 4950 -3128
rect 4950 -3298 4984 -3128
rect 4984 -3298 4996 -3128
rect 4940 -3312 4996 -3298
rect 5228 -2922 5284 -2908
rect 5228 -3092 5238 -2922
rect 5238 -3092 5272 -2922
rect 5272 -3092 5284 -2922
rect 5132 -3298 5142 -3128
rect 5142 -3298 5176 -3128
rect 5176 -3298 5188 -3128
rect 5132 -3312 5188 -3298
rect 5420 -2922 5476 -2908
rect 5420 -3092 5430 -2922
rect 5430 -3092 5464 -2922
rect 5464 -3092 5476 -2922
rect 5324 -3298 5334 -3128
rect 5334 -3298 5368 -3128
rect 5368 -3298 5380 -3128
rect 5324 -3312 5380 -3298
rect 5612 -2922 5668 -2908
rect 5612 -3092 5622 -2922
rect 5622 -3092 5656 -2922
rect 5656 -3092 5668 -2922
rect 5516 -3298 5526 -3128
rect 5526 -3298 5560 -3128
rect 5560 -3298 5572 -3128
rect 5516 -3312 5572 -3298
rect 5804 -2922 5860 -2908
rect 5804 -3092 5814 -2922
rect 5814 -3092 5848 -2922
rect 5848 -3092 5860 -2922
rect 5708 -3298 5718 -3128
rect 5718 -3298 5752 -3128
rect 5752 -3298 5764 -3128
rect 5708 -3312 5764 -3298
rect 5996 -2922 6052 -2908
rect 5996 -3092 6006 -2922
rect 6006 -3092 6040 -2922
rect 6040 -3092 6052 -2922
rect 5900 -3298 5910 -3128
rect 5910 -3298 5944 -3128
rect 5944 -3298 5956 -3128
rect 5900 -3312 5956 -3298
rect 6188 -2922 6244 -2908
rect 6188 -3092 6198 -2922
rect 6198 -3092 6232 -2922
rect 6232 -3092 6244 -2922
rect 6092 -3298 6102 -3128
rect 6102 -3298 6136 -3128
rect 6136 -3298 6148 -3128
rect 6092 -3312 6148 -3298
rect 6380 -2922 6436 -2908
rect 6380 -3092 6390 -2922
rect 6390 -3092 6424 -2922
rect 6424 -3092 6436 -2922
rect 6284 -3298 6294 -3128
rect 6294 -3298 6328 -3128
rect 6328 -3298 6340 -3128
rect 6284 -3312 6340 -3298
rect 6572 -2922 6628 -2908
rect 6572 -3092 6582 -2922
rect 6582 -3092 6616 -2922
rect 6616 -3092 6628 -2922
rect 6476 -3298 6486 -3128
rect 6486 -3298 6520 -3128
rect 6520 -3298 6532 -3128
rect 6476 -3312 6532 -3298
rect 6764 -2922 6820 -2908
rect 6764 -3092 6774 -2922
rect 6774 -3092 6808 -2922
rect 6808 -3092 6820 -2922
rect 6668 -3298 6678 -3128
rect 6678 -3298 6712 -3128
rect 6712 -3298 6724 -3128
rect 6668 -3312 6724 -3298
rect 6860 -3298 6870 -3128
rect 6870 -3298 6904 -3128
rect 6904 -3298 6916 -3128
rect 6860 -3312 6916 -3298
rect -2364 -3602 -2312 -3588
rect -2364 -3768 -2354 -3602
rect -2354 -3768 -2320 -3602
rect -2320 -3768 -2312 -3602
rect -2460 -3978 -2450 -3812
rect -2450 -3978 -2416 -3812
rect -2416 -3978 -2408 -3812
rect -2460 -3992 -2408 -3978
rect -2172 -3602 -2120 -3588
rect -2172 -3768 -2162 -3602
rect -2162 -3768 -2128 -3602
rect -2128 -3768 -2120 -3602
rect -2268 -3978 -2258 -3812
rect -2258 -3978 -2224 -3812
rect -2224 -3978 -2216 -3812
rect -2268 -3992 -2216 -3978
rect -1980 -3602 -1928 -3588
rect -1980 -3768 -1970 -3602
rect -1970 -3768 -1936 -3602
rect -1936 -3768 -1928 -3602
rect -2076 -3978 -2066 -3812
rect -2066 -3978 -2032 -3812
rect -2032 -3978 -2024 -3812
rect -2076 -3992 -2024 -3978
rect -1788 -3602 -1736 -3588
rect -1788 -3768 -1778 -3602
rect -1778 -3768 -1744 -3602
rect -1744 -3768 -1736 -3602
rect -1884 -3978 -1874 -3812
rect -1874 -3978 -1840 -3812
rect -1840 -3978 -1832 -3812
rect -1884 -3992 -1832 -3978
rect -1596 -3602 -1544 -3588
rect -1596 -3768 -1586 -3602
rect -1586 -3768 -1552 -3602
rect -1552 -3768 -1544 -3602
rect -1692 -3978 -1682 -3812
rect -1682 -3978 -1648 -3812
rect -1648 -3978 -1640 -3812
rect -1692 -3992 -1640 -3978
rect -1500 -3978 -1490 -3812
rect -1490 -3978 -1456 -3812
rect -1456 -3978 -1448 -3812
rect -1500 -3992 -1448 -3978
rect -564 -3602 -512 -3588
rect -564 -3768 -554 -3602
rect -554 -3768 -520 -3602
rect -520 -3768 -512 -3602
rect -660 -3978 -650 -3812
rect -650 -3978 -616 -3812
rect -616 -3978 -608 -3812
rect -660 -3992 -608 -3978
rect -372 -3602 -320 -3588
rect -372 -3768 -362 -3602
rect -362 -3768 -328 -3602
rect -328 -3768 -320 -3602
rect -468 -3978 -458 -3812
rect -458 -3978 -424 -3812
rect -424 -3978 -416 -3812
rect -468 -3992 -416 -3978
rect -180 -3602 -128 -3588
rect -180 -3768 -170 -3602
rect -170 -3768 -136 -3602
rect -136 -3768 -128 -3602
rect -276 -3978 -266 -3812
rect -266 -3978 -232 -3812
rect -232 -3978 -224 -3812
rect -276 -3992 -224 -3978
rect 12 -3602 64 -3588
rect 12 -3768 22 -3602
rect 22 -3768 56 -3602
rect 56 -3768 64 -3602
rect -84 -3978 -74 -3812
rect -74 -3978 -40 -3812
rect -40 -3978 -32 -3812
rect -84 -3992 -32 -3978
rect 204 -3602 256 -3588
rect 204 -3768 214 -3602
rect 214 -3768 248 -3602
rect 248 -3768 256 -3602
rect 108 -3978 118 -3812
rect 118 -3978 152 -3812
rect 152 -3978 160 -3812
rect 108 -3992 160 -3978
rect 300 -3978 310 -3812
rect 310 -3978 344 -3812
rect 344 -3978 352 -3812
rect 300 -3992 352 -3978
rect 1236 -3602 1288 -3588
rect 1236 -3768 1246 -3602
rect 1246 -3768 1280 -3602
rect 1280 -3768 1288 -3602
rect 1140 -3978 1150 -3812
rect 1150 -3978 1184 -3812
rect 1184 -3978 1192 -3812
rect 1140 -3992 1192 -3978
rect 1428 -3602 1480 -3588
rect 1428 -3768 1438 -3602
rect 1438 -3768 1472 -3602
rect 1472 -3768 1480 -3602
rect 1332 -3978 1342 -3812
rect 1342 -3978 1376 -3812
rect 1376 -3978 1384 -3812
rect 1332 -3992 1384 -3978
rect 1620 -3602 1672 -3588
rect 1620 -3768 1630 -3602
rect 1630 -3768 1664 -3602
rect 1664 -3768 1672 -3602
rect 1524 -3978 1534 -3812
rect 1534 -3978 1568 -3812
rect 1568 -3978 1576 -3812
rect 1524 -3992 1576 -3978
rect 1812 -3602 1864 -3588
rect 1812 -3768 1822 -3602
rect 1822 -3768 1856 -3602
rect 1856 -3768 1864 -3602
rect 1716 -3978 1726 -3812
rect 1726 -3978 1760 -3812
rect 1760 -3978 1768 -3812
rect 1716 -3992 1768 -3978
rect 2004 -3602 2056 -3588
rect 2004 -3768 2014 -3602
rect 2014 -3768 2048 -3602
rect 2048 -3768 2056 -3602
rect 1908 -3978 1918 -3812
rect 1918 -3978 1952 -3812
rect 1952 -3978 1960 -3812
rect 1908 -3992 1960 -3978
rect 2100 -3978 2110 -3812
rect 2110 -3978 2144 -3812
rect 2144 -3978 2152 -3812
rect 2100 -3992 2152 -3978
rect 3036 -3602 3088 -3588
rect 3036 -3768 3046 -3602
rect 3046 -3768 3080 -3602
rect 3080 -3768 3088 -3602
rect 2940 -3978 2950 -3812
rect 2950 -3978 2984 -3812
rect 2984 -3978 2992 -3812
rect 2940 -3992 2992 -3978
rect 3228 -3602 3280 -3588
rect 3228 -3768 3238 -3602
rect 3238 -3768 3272 -3602
rect 3272 -3768 3280 -3602
rect 3132 -3978 3142 -3812
rect 3142 -3978 3176 -3812
rect 3176 -3978 3184 -3812
rect 3132 -3992 3184 -3978
rect 3420 -3602 3472 -3588
rect 3420 -3768 3430 -3602
rect 3430 -3768 3464 -3602
rect 3464 -3768 3472 -3602
rect 3324 -3978 3334 -3812
rect 3334 -3978 3368 -3812
rect 3368 -3978 3376 -3812
rect 3324 -3992 3376 -3978
rect 3612 -3602 3664 -3588
rect 3612 -3768 3622 -3602
rect 3622 -3768 3656 -3602
rect 3656 -3768 3664 -3602
rect 3516 -3978 3526 -3812
rect 3526 -3978 3560 -3812
rect 3560 -3978 3568 -3812
rect 3516 -3992 3568 -3978
rect 3804 -3602 3856 -3588
rect 3804 -3768 3814 -3602
rect 3814 -3768 3848 -3602
rect 3848 -3768 3856 -3602
rect 3708 -3978 3718 -3812
rect 3718 -3978 3752 -3812
rect 3752 -3978 3760 -3812
rect 3708 -3992 3760 -3978
rect 3900 -3978 3910 -3812
rect 3910 -3978 3944 -3812
rect 3944 -3978 3952 -3812
rect 3900 -3992 3952 -3978
rect -2460 -4512 -2408 -4500
rect -2460 -4680 -2450 -4512
rect -2450 -4680 -2416 -4512
rect -2416 -4680 -2408 -4512
rect -2200 -4888 -2192 -4720
rect -2192 -4888 -2158 -4720
rect -2158 -4888 -2148 -4720
rect -2200 -4900 -2148 -4888
rect -1944 -4512 -1892 -4500
rect -1944 -4680 -1934 -4512
rect -1934 -4680 -1900 -4512
rect -1900 -4680 -1892 -4512
rect -1684 -4888 -1676 -4720
rect -1676 -4888 -1642 -4720
rect -1642 -4888 -1632 -4720
rect -1684 -4900 -1632 -4888
rect -1428 -4512 -1376 -4500
rect -1428 -4680 -1418 -4512
rect -1418 -4680 -1384 -4512
rect -1384 -4680 -1376 -4512
rect -660 -4512 -608 -4500
rect -660 -4680 -650 -4512
rect -650 -4680 -616 -4512
rect -616 -4680 -608 -4512
rect -1168 -4888 -1160 -4720
rect -1160 -4888 -1126 -4720
rect -1126 -4888 -1116 -4720
rect -1168 -4900 -1116 -4888
rect -400 -4888 -392 -4720
rect -392 -4888 -358 -4720
rect -358 -4888 -348 -4720
rect -400 -4900 -348 -4888
rect -144 -4512 -92 -4500
rect -144 -4680 -134 -4512
rect -134 -4680 -100 -4512
rect -100 -4680 -92 -4512
rect 116 -4888 124 -4720
rect 124 -4888 158 -4720
rect 158 -4888 168 -4720
rect 116 -4900 168 -4888
rect 372 -4512 424 -4500
rect 372 -4680 382 -4512
rect 382 -4680 416 -4512
rect 416 -4680 424 -4512
rect 1140 -4512 1192 -4500
rect 1140 -4680 1150 -4512
rect 1150 -4680 1184 -4512
rect 1184 -4680 1192 -4512
rect 632 -4888 640 -4720
rect 640 -4888 674 -4720
rect 674 -4888 684 -4720
rect 632 -4900 684 -4888
rect 1400 -4888 1408 -4720
rect 1408 -4888 1442 -4720
rect 1442 -4888 1452 -4720
rect 1400 -4900 1452 -4888
rect 1656 -4512 1708 -4500
rect 1656 -4680 1666 -4512
rect 1666 -4680 1700 -4512
rect 1700 -4680 1708 -4512
rect 1916 -4888 1924 -4720
rect 1924 -4888 1958 -4720
rect 1958 -4888 1968 -4720
rect 1916 -4900 1968 -4888
rect 2172 -4512 2224 -4500
rect 2172 -4680 2182 -4512
rect 2182 -4680 2216 -4512
rect 2216 -4680 2224 -4512
rect 2940 -4512 2992 -4500
rect 2940 -4680 2950 -4512
rect 2950 -4680 2984 -4512
rect 2984 -4680 2992 -4512
rect 2432 -4888 2440 -4720
rect 2440 -4888 2474 -4720
rect 2474 -4888 2484 -4720
rect 2432 -4900 2484 -4888
rect 3200 -4888 3208 -4720
rect 3208 -4888 3242 -4720
rect 3242 -4888 3252 -4720
rect 3200 -4900 3252 -4888
rect 3456 -4512 3508 -4500
rect 3456 -4680 3466 -4512
rect 3466 -4680 3500 -4512
rect 3500 -4680 3508 -4512
rect 3716 -4888 3724 -4720
rect 3724 -4888 3758 -4720
rect 3758 -4888 3768 -4720
rect 3716 -4900 3768 -4888
rect 3972 -4512 4024 -4500
rect 3972 -4680 3982 -4512
rect 3982 -4680 4016 -4512
rect 4016 -4680 4024 -4512
rect 4232 -4888 4240 -4720
rect 4240 -4888 4274 -4720
rect 4274 -4888 4284 -4720
rect 4232 -4900 4284 -4888
rect -2460 -5130 -2408 -5116
rect -2460 -5296 -2450 -5130
rect -2450 -5296 -2416 -5130
rect -2416 -5296 -2408 -5130
rect -2200 -5506 -2192 -5336
rect -2192 -5506 -2158 -5336
rect -2158 -5506 -2148 -5336
rect -2200 -5516 -2148 -5506
rect -1944 -5130 -1892 -5116
rect -1944 -5296 -1934 -5130
rect -1934 -5296 -1900 -5130
rect -1900 -5296 -1892 -5130
rect -1684 -5506 -1676 -5336
rect -1676 -5506 -1642 -5336
rect -1642 -5506 -1632 -5336
rect -1684 -5516 -1632 -5506
rect -1428 -5130 -1376 -5116
rect -1428 -5296 -1418 -5130
rect -1418 -5296 -1384 -5130
rect -1384 -5296 -1376 -5130
rect -660 -5130 -608 -5116
rect -660 -5296 -650 -5130
rect -650 -5296 -616 -5130
rect -616 -5296 -608 -5130
rect -1168 -5506 -1160 -5336
rect -1160 -5506 -1126 -5336
rect -1126 -5506 -1116 -5336
rect -1168 -5516 -1116 -5506
rect -400 -5506 -392 -5336
rect -392 -5506 -358 -5336
rect -358 -5506 -348 -5336
rect -400 -5516 -348 -5506
rect -144 -5130 -92 -5116
rect -144 -5296 -134 -5130
rect -134 -5296 -100 -5130
rect -100 -5296 -92 -5130
rect 116 -5506 124 -5336
rect 124 -5506 158 -5336
rect 158 -5506 168 -5336
rect 116 -5516 168 -5506
rect 372 -5130 424 -5116
rect 372 -5296 382 -5130
rect 382 -5296 416 -5130
rect 416 -5296 424 -5130
rect 1140 -5130 1192 -5116
rect 1140 -5296 1150 -5130
rect 1150 -5296 1184 -5130
rect 1184 -5296 1192 -5130
rect 632 -5506 640 -5336
rect 640 -5506 674 -5336
rect 674 -5506 684 -5336
rect 632 -5516 684 -5506
rect 1400 -5506 1408 -5336
rect 1408 -5506 1442 -5336
rect 1442 -5506 1452 -5336
rect 1400 -5516 1452 -5506
rect 1656 -5130 1708 -5116
rect 1656 -5296 1666 -5130
rect 1666 -5296 1700 -5130
rect 1700 -5296 1708 -5130
rect 1916 -5506 1924 -5336
rect 1924 -5506 1958 -5336
rect 1958 -5506 1968 -5336
rect 1916 -5516 1968 -5506
rect 2172 -5130 2224 -5116
rect 2172 -5296 2182 -5130
rect 2182 -5296 2216 -5130
rect 2216 -5296 2224 -5130
rect 2940 -5130 2992 -5116
rect 2940 -5296 2950 -5130
rect 2950 -5296 2984 -5130
rect 2984 -5296 2992 -5130
rect 2432 -5506 2440 -5336
rect 2440 -5506 2474 -5336
rect 2474 -5506 2484 -5336
rect 2432 -5516 2484 -5506
rect 3200 -5506 3208 -5336
rect 3208 -5506 3242 -5336
rect 3242 -5506 3252 -5336
rect 3200 -5516 3252 -5506
rect 3456 -5130 3508 -5116
rect 3456 -5296 3466 -5130
rect 3466 -5296 3500 -5130
rect 3500 -5296 3508 -5130
rect 3716 -5506 3724 -5336
rect 3724 -5506 3758 -5336
rect 3758 -5506 3768 -5336
rect 3716 -5516 3768 -5506
rect 3972 -5130 4024 -5116
rect 3972 -5296 3982 -5130
rect 3982 -5296 4016 -5130
rect 4016 -5296 4024 -5130
rect 4232 -5506 4240 -5336
rect 4240 -5506 4274 -5336
rect 4274 -5506 4284 -5336
rect 4232 -5516 4284 -5506
rect -2460 -5748 -2408 -5736
rect -2460 -5916 -2450 -5748
rect -2450 -5916 -2416 -5748
rect -2416 -5916 -2408 -5748
rect -2200 -6124 -2192 -5956
rect -2192 -6124 -2158 -5956
rect -2158 -6124 -2148 -5956
rect -2200 -6136 -2148 -6124
rect -1944 -5748 -1892 -5736
rect -1944 -5916 -1934 -5748
rect -1934 -5916 -1900 -5748
rect -1900 -5916 -1892 -5748
rect -1684 -6124 -1676 -5956
rect -1676 -6124 -1642 -5956
rect -1642 -6124 -1632 -5956
rect -1684 -6136 -1632 -6124
rect -1428 -5748 -1376 -5736
rect -1428 -5916 -1418 -5748
rect -1418 -5916 -1384 -5748
rect -1384 -5916 -1376 -5748
rect -660 -5748 -608 -5736
rect -660 -5916 -650 -5748
rect -650 -5916 -616 -5748
rect -616 -5916 -608 -5748
rect -1168 -6124 -1160 -5956
rect -1160 -6124 -1126 -5956
rect -1126 -6124 -1116 -5956
rect -1168 -6136 -1116 -6124
rect -400 -6124 -392 -5956
rect -392 -6124 -358 -5956
rect -358 -6124 -348 -5956
rect -400 -6136 -348 -6124
rect -144 -5748 -92 -5736
rect -144 -5916 -134 -5748
rect -134 -5916 -100 -5748
rect -100 -5916 -92 -5748
rect 116 -6124 124 -5956
rect 124 -6124 158 -5956
rect 158 -6124 168 -5956
rect 116 -6136 168 -6124
rect 372 -5748 424 -5736
rect 372 -5916 382 -5748
rect 382 -5916 416 -5748
rect 416 -5916 424 -5748
rect 1140 -5748 1192 -5736
rect 1140 -5916 1150 -5748
rect 1150 -5916 1184 -5748
rect 1184 -5916 1192 -5748
rect 632 -6124 640 -5956
rect 640 -6124 674 -5956
rect 674 -6124 684 -5956
rect 632 -6136 684 -6124
rect 1400 -6124 1408 -5956
rect 1408 -6124 1442 -5956
rect 1442 -6124 1452 -5956
rect 1400 -6136 1452 -6124
rect 1656 -5748 1708 -5736
rect 1656 -5916 1666 -5748
rect 1666 -5916 1700 -5748
rect 1700 -5916 1708 -5748
rect 1916 -6124 1924 -5956
rect 1924 -6124 1958 -5956
rect 1958 -6124 1968 -5956
rect 1916 -6136 1968 -6124
rect 2172 -5748 2224 -5736
rect 2172 -5916 2182 -5748
rect 2182 -5916 2216 -5748
rect 2216 -5916 2224 -5748
rect 2940 -5748 2992 -5736
rect 2940 -5916 2950 -5748
rect 2950 -5916 2984 -5748
rect 2984 -5916 2992 -5748
rect 2432 -6124 2440 -5956
rect 2440 -6124 2474 -5956
rect 2474 -6124 2484 -5956
rect 2432 -6136 2484 -6124
rect 3200 -6124 3208 -5956
rect 3208 -6124 3242 -5956
rect 3242 -6124 3252 -5956
rect 3200 -6136 3252 -6124
rect 3456 -5748 3508 -5736
rect 3456 -5916 3466 -5748
rect 3466 -5916 3500 -5748
rect 3500 -5916 3508 -5748
rect 3716 -6124 3724 -5956
rect 3724 -6124 3758 -5956
rect 3758 -6124 3768 -5956
rect 3716 -6136 3768 -6124
rect 3972 -5748 4024 -5736
rect 3972 -5916 3982 -5748
rect 3982 -5916 4016 -5748
rect 4016 -5916 4024 -5748
rect 4232 -6124 4240 -5956
rect 4240 -6124 4274 -5956
rect 4274 -6124 4284 -5956
rect 4232 -6136 4284 -6124
rect -2460 -6366 -2408 -6352
rect -2460 -6532 -2450 -6366
rect -2450 -6532 -2416 -6366
rect -2416 -6532 -2408 -6366
rect -2200 -6742 -2192 -6572
rect -2192 -6742 -2158 -6572
rect -2158 -6742 -2148 -6572
rect -2200 -6752 -2148 -6742
rect -1944 -6366 -1892 -6352
rect -1944 -6532 -1934 -6366
rect -1934 -6532 -1900 -6366
rect -1900 -6532 -1892 -6366
rect -1684 -6742 -1676 -6572
rect -1676 -6742 -1642 -6572
rect -1642 -6742 -1632 -6572
rect -1684 -6752 -1632 -6742
rect -1428 -6366 -1376 -6352
rect -1428 -6532 -1418 -6366
rect -1418 -6532 -1384 -6366
rect -1384 -6532 -1376 -6366
rect -660 -6366 -608 -6352
rect -660 -6532 -650 -6366
rect -650 -6532 -616 -6366
rect -616 -6532 -608 -6366
rect -1168 -6742 -1160 -6572
rect -1160 -6742 -1126 -6572
rect -1126 -6742 -1116 -6572
rect -1168 -6752 -1116 -6742
rect -400 -6742 -392 -6572
rect -392 -6742 -358 -6572
rect -358 -6742 -348 -6572
rect -400 -6752 -348 -6742
rect -144 -6366 -92 -6352
rect -144 -6532 -134 -6366
rect -134 -6532 -100 -6366
rect -100 -6532 -92 -6366
rect 116 -6742 124 -6572
rect 124 -6742 158 -6572
rect 158 -6742 168 -6572
rect 116 -6752 168 -6742
rect 372 -6366 424 -6352
rect 372 -6532 382 -6366
rect 382 -6532 416 -6366
rect 416 -6532 424 -6366
rect 1140 -6366 1192 -6352
rect 1140 -6532 1150 -6366
rect 1150 -6532 1184 -6366
rect 1184 -6532 1192 -6366
rect 632 -6742 640 -6572
rect 640 -6742 674 -6572
rect 674 -6742 684 -6572
rect 632 -6752 684 -6742
rect 1400 -6742 1408 -6572
rect 1408 -6742 1442 -6572
rect 1442 -6742 1452 -6572
rect 1400 -6752 1452 -6742
rect 1656 -6366 1708 -6352
rect 1656 -6532 1666 -6366
rect 1666 -6532 1700 -6366
rect 1700 -6532 1708 -6366
rect 1916 -6742 1924 -6572
rect 1924 -6742 1958 -6572
rect 1958 -6742 1968 -6572
rect 1916 -6752 1968 -6742
rect 2172 -6366 2224 -6352
rect 2172 -6532 2182 -6366
rect 2182 -6532 2216 -6366
rect 2216 -6532 2224 -6366
rect 2940 -6366 2992 -6352
rect 2940 -6532 2950 -6366
rect 2950 -6532 2984 -6366
rect 2984 -6532 2992 -6366
rect 2432 -6742 2440 -6572
rect 2440 -6742 2474 -6572
rect 2474 -6742 2484 -6572
rect 2432 -6752 2484 -6742
rect 3200 -6742 3208 -6572
rect 3208 -6742 3242 -6572
rect 3242 -6742 3252 -6572
rect 3200 -6752 3252 -6742
rect 3456 -6366 3508 -6352
rect 3456 -6532 3466 -6366
rect 3466 -6532 3500 -6366
rect 3500 -6532 3508 -6366
rect 3716 -6742 3724 -6572
rect 3724 -6742 3758 -6572
rect 3758 -6742 3768 -6572
rect 3716 -6752 3768 -6742
rect 3972 -6366 4024 -6352
rect 3972 -6532 3982 -6366
rect 3982 -6532 4016 -6366
rect 4016 -6532 4024 -6366
rect 4232 -6742 4240 -6572
rect 4240 -6742 4274 -6572
rect 4274 -6742 4284 -6572
rect 4232 -6752 4284 -6742
rect -2460 -6984 -2408 -6972
rect -2460 -7152 -2450 -6984
rect -2450 -7152 -2416 -6984
rect -2416 -7152 -2408 -6984
rect -2200 -7360 -2192 -7192
rect -2192 -7360 -2158 -7192
rect -2158 -7360 -2148 -7192
rect -2200 -7372 -2148 -7360
rect -1944 -6984 -1892 -6972
rect -1944 -7152 -1934 -6984
rect -1934 -7152 -1900 -6984
rect -1900 -7152 -1892 -6984
rect -1684 -7360 -1676 -7192
rect -1676 -7360 -1642 -7192
rect -1642 -7360 -1632 -7192
rect -1684 -7372 -1632 -7360
rect -1428 -6984 -1376 -6972
rect -1428 -7152 -1418 -6984
rect -1418 -7152 -1384 -6984
rect -1384 -7152 -1376 -6984
rect -660 -6984 -608 -6972
rect -660 -7152 -650 -6984
rect -650 -7152 -616 -6984
rect -616 -7152 -608 -6984
rect -1168 -7360 -1160 -7192
rect -1160 -7360 -1126 -7192
rect -1126 -7360 -1116 -7192
rect -1168 -7372 -1116 -7360
rect -400 -7360 -392 -7192
rect -392 -7360 -358 -7192
rect -358 -7360 -348 -7192
rect -400 -7372 -348 -7360
rect -144 -6984 -92 -6972
rect -144 -7152 -134 -6984
rect -134 -7152 -100 -6984
rect -100 -7152 -92 -6984
rect 116 -7360 124 -7192
rect 124 -7360 158 -7192
rect 158 -7360 168 -7192
rect 116 -7372 168 -7360
rect 372 -6984 424 -6972
rect 372 -7152 382 -6984
rect 382 -7152 416 -6984
rect 416 -7152 424 -6984
rect 1140 -6984 1192 -6972
rect 1140 -7152 1150 -6984
rect 1150 -7152 1184 -6984
rect 1184 -7152 1192 -6984
rect 632 -7360 640 -7192
rect 640 -7360 674 -7192
rect 674 -7360 684 -7192
rect 632 -7372 684 -7360
rect 1400 -7360 1408 -7192
rect 1408 -7360 1442 -7192
rect 1442 -7360 1452 -7192
rect 1400 -7372 1452 -7360
rect 1656 -6984 1708 -6972
rect 1656 -7152 1666 -6984
rect 1666 -7152 1700 -6984
rect 1700 -7152 1708 -6984
rect 1916 -7360 1924 -7192
rect 1924 -7360 1958 -7192
rect 1958 -7360 1968 -7192
rect 1916 -7372 1968 -7360
rect 2172 -6984 2224 -6972
rect 2172 -7152 2182 -6984
rect 2182 -7152 2216 -6984
rect 2216 -7152 2224 -6984
rect 2940 -6984 2992 -6972
rect 2940 -7152 2950 -6984
rect 2950 -7152 2984 -6984
rect 2984 -7152 2992 -6984
rect 2432 -7360 2440 -7192
rect 2440 -7360 2474 -7192
rect 2474 -7360 2484 -7192
rect 2432 -7372 2484 -7360
rect 3200 -7360 3208 -7192
rect 3208 -7360 3242 -7192
rect 3242 -7360 3252 -7192
rect 3200 -7372 3252 -7360
rect 3456 -6984 3508 -6972
rect 3456 -7152 3466 -6984
rect 3466 -7152 3500 -6984
rect 3500 -7152 3508 -6984
rect 3716 -7360 3724 -7192
rect 3724 -7360 3758 -7192
rect 3758 -7360 3768 -7192
rect 3716 -7372 3768 -7360
rect 3972 -6984 4024 -6972
rect 3972 -7152 3982 -6984
rect 3982 -7152 4016 -6984
rect 4016 -7152 4024 -6984
rect 4232 -7360 4240 -7192
rect 4240 -7360 4274 -7192
rect 4274 -7360 4284 -7192
rect 4232 -7372 4284 -7360
rect -2460 -7602 -2408 -7588
rect -2460 -7768 -2450 -7602
rect -2450 -7768 -2416 -7602
rect -2416 -7768 -2408 -7602
rect -2200 -7978 -2192 -7808
rect -2192 -7978 -2158 -7808
rect -2158 -7978 -2148 -7808
rect -2200 -7988 -2148 -7978
rect -1944 -7602 -1892 -7588
rect -1944 -7768 -1934 -7602
rect -1934 -7768 -1900 -7602
rect -1900 -7768 -1892 -7602
rect -1684 -7978 -1676 -7808
rect -1676 -7978 -1642 -7808
rect -1642 -7978 -1632 -7808
rect -1684 -7988 -1632 -7978
rect -1428 -7602 -1376 -7588
rect -1428 -7768 -1418 -7602
rect -1418 -7768 -1384 -7602
rect -1384 -7768 -1376 -7602
rect -660 -7602 -608 -7588
rect -660 -7768 -650 -7602
rect -650 -7768 -616 -7602
rect -616 -7768 -608 -7602
rect -1168 -7978 -1160 -7808
rect -1160 -7978 -1126 -7808
rect -1126 -7978 -1116 -7808
rect -1168 -7988 -1116 -7978
rect -980 -8160 -800 -7960
rect -400 -7978 -392 -7808
rect -392 -7978 -358 -7808
rect -358 -7978 -348 -7808
rect -400 -7988 -348 -7978
rect -144 -7602 -92 -7588
rect -144 -7768 -134 -7602
rect -134 -7768 -100 -7602
rect -100 -7768 -92 -7602
rect 116 -7978 124 -7808
rect 124 -7978 158 -7808
rect 158 -7978 168 -7808
rect 116 -7988 168 -7978
rect 372 -7602 424 -7588
rect 372 -7768 382 -7602
rect 382 -7768 416 -7602
rect 416 -7768 424 -7602
rect 1140 -7602 1192 -7588
rect 1140 -7768 1150 -7602
rect 1150 -7768 1184 -7602
rect 1184 -7768 1192 -7602
rect 632 -7978 640 -7808
rect 640 -7978 674 -7808
rect 674 -7978 684 -7808
rect 632 -7988 684 -7978
rect 1400 -7978 1408 -7808
rect 1408 -7978 1442 -7808
rect 1442 -7978 1452 -7808
rect 1400 -7988 1452 -7978
rect 1656 -7602 1708 -7588
rect 1656 -7768 1666 -7602
rect 1666 -7768 1700 -7602
rect 1700 -7768 1708 -7602
rect 1916 -7978 1924 -7808
rect 1924 -7978 1958 -7808
rect 1958 -7978 1968 -7808
rect 1916 -7988 1968 -7978
rect 2172 -7602 2224 -7588
rect 2172 -7768 2182 -7602
rect 2182 -7768 2216 -7602
rect 2216 -7768 2224 -7602
rect 2940 -7602 2992 -7588
rect 2940 -7768 2950 -7602
rect 2950 -7768 2984 -7602
rect 2984 -7768 2992 -7602
rect 2432 -7978 2440 -7808
rect 2440 -7978 2474 -7808
rect 2474 -7978 2484 -7808
rect 2432 -7988 2484 -7978
rect 3200 -7978 3208 -7808
rect 3208 -7978 3242 -7808
rect 3242 -7978 3252 -7808
rect 3200 -7988 3252 -7978
rect 3456 -7602 3508 -7588
rect 3456 -7768 3466 -7602
rect 3466 -7768 3500 -7602
rect 3500 -7768 3508 -7602
rect 3716 -7978 3724 -7808
rect 3724 -7978 3758 -7808
rect 3758 -7978 3768 -7808
rect 3716 -7988 3768 -7978
rect 3972 -7602 4024 -7588
rect 3972 -7768 3982 -7602
rect 3982 -7768 4016 -7602
rect 4016 -7768 4024 -7602
rect 4232 -7978 4240 -7808
rect 4240 -7978 4274 -7808
rect 4274 -7978 4284 -7808
rect 4232 -7988 4284 -7978
rect -5444 -9416 -4636 -8610
<< metal2 >>
rect 3420 2580 3600 2590
rect 3420 2370 3600 2380
rect 2532 2136 4524 2152
rect -76 2122 492 2124
rect -80 2112 2096 2122
rect 2532 2056 3536 2136
rect 2532 1880 2536 2056
rect 2592 1880 2728 2056
rect 2536 1866 2592 1876
rect 2784 1880 2920 2056
rect 2728 1866 2784 1876
rect 2976 1880 3112 2056
rect 2920 1866 2976 1876
rect 3168 1880 3304 2056
rect 3112 1866 3168 1876
rect 3360 1880 3496 2056
rect 4512 1892 4524 2136
rect 6084 2064 6956 2074
rect 3304 1866 3360 1876
rect 3552 1880 3688 1892
rect 3496 1866 3552 1876
rect 3744 1880 3880 1892
rect 3688 1866 3744 1876
rect 3936 1880 4072 1892
rect 3880 1866 3936 1876
rect 4128 1880 4264 1892
rect 4072 1866 4128 1876
rect 4320 1880 4524 1892
rect 5032 2036 6084 2048
rect 4264 1866 4320 1876
rect 5032 1856 5036 2036
rect 5092 1856 5228 2036
rect 5036 1842 5092 1852
rect 5284 1856 5420 2036
rect 5228 1842 5284 1852
rect 5476 1856 5612 2036
rect 5420 1842 5476 1852
rect 5668 1856 5804 2036
rect 5612 1842 5668 1852
rect 5860 1856 5996 2036
rect 5804 1842 5860 1852
rect 6052 1864 6084 2036
rect 6052 1856 6188 1864
rect 6084 1854 6188 1856
rect 5996 1842 6052 1852
rect 6244 1854 6380 1864
rect 6188 1842 6244 1852
rect 6436 1854 6572 1864
rect 6380 1842 6436 1852
rect 6628 1854 6764 1864
rect 6572 1842 6628 1852
rect 6820 1854 6956 1864
rect 6764 1842 6820 1852
rect 2440 1834 2496 1842
rect 2632 1834 2688 1842
rect 2824 1834 2880 1842
rect 3016 1834 3072 1842
rect 3208 1834 3264 1842
rect 3400 1834 3456 1842
rect -80 1666 2096 1676
rect 2436 1832 3456 1834
rect 2436 1824 2440 1832
rect 2496 1824 2632 1832
rect 2688 1824 2824 1832
rect 2880 1824 3016 1832
rect 3072 1824 3208 1832
rect 3264 1824 3400 1832
rect 3592 1832 3648 1842
rect -76 1664 492 1666
rect 3456 1652 3592 1828
rect 3784 1832 3840 1842
rect 3648 1652 3784 1828
rect 3976 1832 4032 1842
rect 3840 1652 3976 1828
rect 4168 1832 4224 1842
rect 4032 1652 4168 1828
rect 4360 1832 4416 1842
rect 4224 1652 4360 1828
rect 4416 1652 4428 1828
rect 4940 1816 4996 1826
rect 3412 1568 4428 1652
rect 4932 1804 4940 1814
rect 5132 1816 5188 1826
rect 4996 1804 5132 1814
rect 5324 1816 5380 1826
rect 5188 1804 5324 1814
rect 5516 1816 5572 1826
rect 5380 1804 5516 1814
rect 5708 1816 5764 1826
rect 5572 1804 5708 1814
rect 5900 1816 5956 1826
rect 5764 1804 5900 1814
rect 6092 1816 6148 1826
rect 5956 1632 6092 1812
rect 6284 1816 6340 1826
rect 6148 1632 6284 1812
rect 6476 1816 6532 1826
rect 6340 1632 6476 1812
rect 6668 1816 6724 1826
rect 6532 1632 6668 1812
rect 6860 1816 6916 1826
rect 6724 1632 6860 1812
rect 5916 1620 6916 1632
rect 4932 1606 5916 1616
rect 2436 1556 4428 1568
rect 2524 1504 4516 1520
rect 2524 1424 3536 1504
rect 2524 1248 2536 1424
rect 2592 1248 2728 1424
rect 2536 1234 2592 1244
rect 2784 1248 2920 1424
rect 2728 1234 2784 1244
rect 2976 1248 3112 1424
rect 2920 1234 2976 1244
rect 3168 1248 3304 1424
rect 3112 1234 3168 1244
rect 3360 1248 3496 1424
rect 4512 1260 4516 1504
rect 6088 1448 6960 1458
rect 3304 1234 3360 1244
rect 3552 1248 3688 1260
rect 3496 1234 3552 1244
rect 3744 1248 3880 1260
rect 3688 1234 3744 1244
rect 3936 1248 4072 1260
rect 3880 1234 3936 1244
rect 4128 1248 4264 1260
rect 4072 1234 4128 1244
rect 4320 1248 4516 1260
rect 5032 1420 6088 1432
rect 4264 1234 4320 1244
rect 5032 1240 5036 1420
rect 5092 1240 5228 1420
rect 5036 1226 5092 1236
rect 5284 1240 5420 1420
rect 5228 1226 5284 1236
rect 5476 1240 5612 1420
rect 5420 1226 5476 1236
rect 5668 1240 5804 1420
rect 5612 1226 5668 1236
rect 5860 1240 5996 1420
rect 5804 1226 5860 1236
rect 6052 1248 6088 1420
rect 6052 1240 6188 1248
rect 6088 1238 6188 1240
rect 5996 1226 6052 1236
rect 6244 1238 6380 1248
rect 6188 1226 6244 1236
rect 6436 1238 6572 1248
rect 6380 1226 6436 1236
rect 6628 1238 6764 1248
rect 6572 1226 6628 1236
rect 6820 1238 6960 1248
rect 6764 1226 6820 1236
rect 2440 1202 2496 1210
rect 2632 1202 2688 1210
rect 2824 1202 2880 1210
rect 3016 1202 3072 1210
rect 3208 1202 3264 1210
rect 3400 1202 3456 1210
rect 2436 1200 3456 1202
rect 2436 1192 2440 1200
rect 2496 1192 2632 1200
rect 2688 1192 2824 1200
rect 2880 1192 3016 1200
rect 3072 1192 3208 1200
rect 3264 1192 3400 1200
rect 3592 1200 3648 1210
rect -5490 864 1760 1040
rect 3456 1020 3592 1196
rect 3784 1200 3840 1210
rect 3648 1020 3784 1196
rect 3976 1200 4032 1210
rect 3840 1020 3976 1196
rect 4168 1200 4224 1210
rect 4032 1020 4168 1196
rect 4360 1200 4416 1210
rect 4224 1020 4360 1196
rect 4940 1200 4996 1210
rect 4416 1020 4428 1196
rect 3412 932 4428 1020
rect 4936 1184 4940 1196
rect 5132 1200 5188 1210
rect 4996 1184 5132 1196
rect 5324 1200 5380 1210
rect 5188 1184 5324 1196
rect 5516 1200 5572 1210
rect 5380 1184 5516 1196
rect 5708 1200 5764 1210
rect 5572 1184 5708 1196
rect 5900 1200 5956 1210
rect 5764 1184 5900 1196
rect 6092 1200 6148 1210
rect 5956 1016 6092 1196
rect 6284 1200 6340 1210
rect 6148 1016 6284 1196
rect 6476 1200 6532 1210
rect 6340 1016 6476 1196
rect 6668 1200 6724 1210
rect 6532 1016 6668 1196
rect 6860 1200 6916 1210
rect 6724 1016 6860 1196
rect 5920 1004 6916 1016
rect 4936 986 5920 996
rect 2436 924 4428 932
rect 2436 922 3412 924
rect -5490 448 300 864
rect 6088 832 6960 842
rect 5032 800 6088 812
rect 5032 620 5036 800
rect 5092 620 5228 800
rect 5036 606 5092 616
rect 5284 620 5420 800
rect 5228 606 5284 616
rect 5476 620 5612 800
rect 5420 606 5476 616
rect 5668 620 5804 800
rect 5612 606 5668 616
rect 5860 620 5996 800
rect 5804 606 5860 616
rect 6052 632 6088 800
rect 6052 620 6188 632
rect 5996 606 6052 616
rect 6244 620 6380 632
rect 6188 606 6244 616
rect 6436 620 6572 632
rect 6380 606 6436 616
rect 6628 620 6764 632
rect 6572 606 6628 616
rect 6820 622 6960 632
rect 6820 620 6824 622
rect 6764 606 6820 616
rect 4940 580 4996 590
rect 4932 568 4940 578
rect 5132 580 5188 590
rect 4996 568 5132 578
rect 5324 580 5380 590
rect 5188 568 5324 578
rect 5516 580 5572 590
rect 5380 568 5516 578
rect 5708 580 5764 590
rect 5572 568 5708 578
rect 5900 580 5956 590
rect 5764 568 5900 578
rect 6092 580 6148 590
rect -5490 330 1760 448
rect 2532 556 4524 568
rect 2532 472 3548 556
rect 2144 420 2380 430
rect -5490 -110 90 330
rect 2140 152 2144 162
rect 2532 296 2536 472
rect 2592 296 2728 472
rect 2536 282 2592 292
rect 2784 296 2920 472
rect 2728 282 2784 292
rect 2976 296 3112 472
rect 2920 282 2976 292
rect 3168 296 3304 472
rect 3112 282 3168 292
rect 3360 296 3496 472
rect 5956 396 6092 576
rect 6284 580 6340 590
rect 6148 396 6284 576
rect 6476 580 6532 590
rect 6340 396 6476 576
rect 6668 580 6724 590
rect 6532 396 6668 576
rect 6860 580 6916 590
rect 6724 396 6860 576
rect 5916 384 6916 396
rect 4932 370 5916 380
rect 3304 282 3360 292
rect 3552 296 3688 308
rect 3496 282 3552 292
rect 3744 296 3880 308
rect 3688 282 3744 292
rect 3936 296 4072 308
rect 3880 282 3936 292
rect 4128 296 4264 308
rect 4072 282 4128 292
rect 4320 296 4524 308
rect 4264 282 4320 292
rect 2440 254 2496 258
rect 2632 254 2688 258
rect 2824 254 2880 258
rect 3016 254 3072 258
rect 3208 254 3264 258
rect 3400 254 3456 258
rect 2428 248 3456 254
rect 2428 244 2440 248
rect 2496 244 2632 248
rect 2688 244 2824 248
rect 2880 244 3016 248
rect 3072 244 3208 248
rect 3264 244 3400 248
rect 3592 248 3648 258
rect 290 130 1930 140
rect 212 28 290 44
rect 1930 28 2004 44
rect 212 -148 216 28
rect 272 -100 290 28
rect 1930 -100 1944 28
rect 272 -148 408 -100
rect 216 -162 272 -152
rect 464 -148 600 -100
rect 408 -162 464 -152
rect 656 -148 792 -100
rect 600 -162 656 -152
rect 848 -148 984 -100
rect 792 -162 848 -152
rect 1040 -148 1176 -100
rect 984 -162 1040 -152
rect 1232 -148 1368 -100
rect 1176 -162 1232 -152
rect 1424 -148 1560 -100
rect 1368 -162 1424 -152
rect 1616 -148 1752 -100
rect 1560 -162 1616 -152
rect 1808 -148 1944 -100
rect 1752 -162 1808 -152
rect 2000 -148 2004 28
rect 2380 -4 2428 244
rect 3456 68 3592 244
rect 3784 248 3840 258
rect 3648 68 3784 244
rect 3976 248 4032 258
rect 3840 68 3976 244
rect 4168 248 4224 258
rect 4032 68 4168 244
rect 4360 248 4416 258
rect 4224 68 4360 244
rect 6088 212 6960 222
rect 3404 -4 4416 68
rect 5032 184 6088 196
rect 5032 4 5036 184
rect 2380 -16 4416 -4
rect 5092 4 5228 184
rect 5036 -10 5092 0
rect 5284 4 5420 184
rect 5228 -10 5284 0
rect 5476 4 5612 184
rect 5420 -10 5476 0
rect 5668 4 5804 184
rect 5612 -10 5668 0
rect 5860 4 5996 184
rect 5804 -10 5860 0
rect 6052 12 6088 184
rect 6052 4 6188 12
rect 6088 2 6188 4
rect 5996 -10 6052 0
rect 6244 2 6380 12
rect 6188 -10 6244 0
rect 6436 2 6572 12
rect 6380 -10 6436 0
rect 6628 2 6764 12
rect 6572 -10 6628 0
rect 6820 2 6960 12
rect 6764 -10 6820 0
rect 2380 -120 2500 -16
rect 4940 -36 4996 -26
rect 4928 -48 4940 -38
rect 5132 -36 5188 -26
rect 4996 -48 5132 -38
rect 5324 -36 5380 -26
rect 5188 -48 5324 -38
rect 5516 -36 5572 -26
rect 5380 -48 5516 -38
rect 5708 -36 5764 -26
rect 5572 -48 5708 -38
rect 5900 -36 5956 -26
rect 5764 -48 5900 -38
rect 6092 -36 6148 -26
rect 2140 -130 2500 -120
rect 1944 -162 2000 -152
rect 120 -196 176 -186
rect -232 -376 120 -200
rect 312 -196 368 -186
rect 176 -376 312 -200
rect 504 -196 560 -186
rect 368 -376 504 -200
rect 696 -196 752 -186
rect 560 -376 696 -200
rect 888 -196 944 -186
rect 752 -376 888 -200
rect 1080 -196 1136 -186
rect 944 -376 1080 -200
rect 1272 -196 1328 -186
rect 1136 -376 1272 -200
rect 1464 -196 1520 -186
rect 1328 -376 1464 -200
rect 1656 -196 1712 -186
rect 1520 -376 1656 -200
rect 1848 -196 1904 -186
rect 1712 -376 1848 -200
rect 2040 -196 2096 -186
rect 1904 -376 2040 -200
rect 2096 -376 2244 -200
rect -232 -392 2244 -376
rect -232 -802 164 -392
rect 290 -490 1930 -480
rect 212 -588 290 -572
rect 1930 -588 2004 -572
rect 212 -764 216 -588
rect 272 -720 290 -588
rect 1930 -720 1944 -588
rect 272 -764 408 -720
rect 216 -778 272 -768
rect 464 -764 600 -720
rect 408 -778 464 -768
rect 656 -764 792 -720
rect 600 -778 656 -768
rect 848 -764 984 -720
rect 792 -778 848 -768
rect 1040 -764 1176 -720
rect 984 -778 1040 -768
rect 1232 -764 1368 -720
rect 1176 -778 1232 -768
rect 1424 -764 1560 -720
rect 1368 -778 1424 -768
rect 1616 -764 1752 -720
rect 1560 -778 1616 -768
rect 1808 -764 1944 -720
rect 1752 -778 1808 -768
rect 2000 -764 2004 -588
rect 1944 -778 2000 -768
rect 2044 -802 2244 -392
rect 2292 -370 2500 -130
rect 2532 -64 4524 -52
rect 2532 -148 3548 -64
rect 2532 -324 2536 -148
rect 2592 -324 2728 -148
rect 2536 -338 2592 -328
rect 2784 -324 2920 -148
rect 2728 -338 2784 -328
rect 2976 -324 3112 -148
rect 2920 -338 2976 -328
rect 3168 -324 3304 -148
rect 3112 -338 3168 -328
rect 3360 -324 3496 -148
rect 5956 -220 6092 -40
rect 6284 -36 6340 -26
rect 6148 -220 6284 -40
rect 6476 -36 6532 -26
rect 6340 -220 6476 -40
rect 6668 -36 6724 -26
rect 6532 -220 6668 -40
rect 6860 -36 6916 -26
rect 6724 -220 6860 -40
rect 5912 -232 6916 -220
rect 4928 -246 5912 -236
rect 3304 -338 3360 -328
rect 3552 -324 3688 -312
rect 3496 -338 3552 -328
rect 3744 -324 3880 -312
rect 3688 -338 3744 -328
rect 3936 -324 4072 -312
rect 3880 -338 3936 -328
rect 4128 -324 4264 -312
rect 4072 -338 4128 -328
rect 4320 -324 4524 -312
rect 4264 -338 4320 -328
rect 2632 -370 2688 -362
rect 2824 -370 2880 -362
rect 3016 -370 3072 -362
rect 3208 -370 3264 -362
rect 3400 -370 3456 -362
rect 2292 -372 3456 -370
rect 3592 -372 3648 -362
rect 3784 -372 3840 -362
rect 3976 -372 4032 -362
rect 4168 -372 4224 -362
rect 4360 -372 4416 -362
rect 2292 -380 2440 -372
rect 2496 -380 2632 -372
rect 2688 -380 2824 -372
rect 2880 -380 3016 -372
rect 3072 -380 3208 -372
rect 3264 -380 3400 -372
rect 2292 -628 2428 -380
rect 3456 -552 3592 -372
rect 3648 -552 3784 -372
rect 3840 -552 3976 -372
rect 4032 -552 4168 -372
rect 4224 -552 4360 -372
rect 4416 -552 4420 -372
rect 6088 -408 6960 -398
rect 3404 -628 4420 -552
rect 5032 -436 6088 -424
rect 5032 -616 5036 -436
rect 2292 -644 4420 -628
rect 5092 -616 5228 -436
rect 5036 -630 5092 -620
rect 5284 -616 5420 -436
rect 5228 -630 5284 -620
rect 5476 -616 5612 -436
rect 5420 -630 5476 -620
rect 5668 -616 5804 -436
rect 5612 -630 5668 -620
rect 5860 -616 5996 -436
rect 5804 -630 5860 -620
rect 6052 -608 6088 -436
rect 6052 -616 6188 -608
rect 6088 -618 6188 -616
rect 5996 -630 6052 -620
rect 6244 -618 6380 -608
rect 6188 -630 6244 -620
rect 6436 -618 6572 -608
rect 6380 -630 6436 -620
rect 6628 -618 6764 -608
rect 6572 -630 6628 -620
rect 6820 -618 6960 -608
rect 6764 -630 6820 -620
rect -232 -812 176 -802
rect -232 -992 120 -812
rect 312 -812 368 -802
rect 176 -992 312 -816
rect 504 -812 560 -802
rect 368 -992 504 -816
rect 696 -812 752 -802
rect 560 -992 696 -816
rect 888 -812 944 -802
rect 752 -992 888 -816
rect 1080 -812 1136 -802
rect 944 -992 1080 -816
rect 1272 -812 1328 -802
rect 1136 -992 1272 -816
rect 1464 -812 1520 -802
rect 1328 -992 1464 -816
rect 1656 -812 1712 -802
rect 1520 -992 1656 -816
rect 1848 -812 1904 -802
rect 1712 -992 1848 -816
rect 2040 -812 2244 -802
rect 1904 -992 2040 -816
rect 2096 -832 2244 -812
rect 2460 -756 2688 -644
rect 4940 -656 4996 -646
rect 4936 -662 4940 -660
rect 4932 -672 4940 -662
rect 5132 -656 5188 -646
rect 4996 -672 5132 -660
rect 5324 -656 5380 -646
rect 5188 -672 5324 -660
rect 5516 -656 5572 -646
rect 5380 -672 5516 -660
rect 5708 -656 5764 -646
rect 5572 -672 5708 -660
rect 5900 -656 5956 -646
rect 5764 -672 5900 -660
rect 6092 -656 6148 -646
rect 2096 -992 2352 -832
rect -232 -1008 2352 -992
rect -232 -1422 164 -1008
rect 290 -1110 1930 -1100
rect 212 -1208 290 -1192
rect 1930 -1208 2004 -1192
rect 212 -1384 216 -1208
rect 272 -1340 290 -1208
rect 1930 -1340 1944 -1208
rect 272 -1384 408 -1340
rect 216 -1398 272 -1388
rect 464 -1384 600 -1340
rect 408 -1398 464 -1388
rect 656 -1384 792 -1340
rect 600 -1398 656 -1388
rect 848 -1384 984 -1340
rect 792 -1398 848 -1388
rect 1040 -1384 1176 -1340
rect 984 -1398 1040 -1388
rect 1232 -1384 1368 -1340
rect 1176 -1398 1232 -1388
rect 1424 -1384 1560 -1340
rect 1368 -1398 1424 -1388
rect 1616 -1384 1752 -1340
rect 1560 -1398 1616 -1388
rect 1808 -1384 1944 -1340
rect 1752 -1398 1808 -1388
rect 2000 -1384 2004 -1208
rect 2044 -1300 2352 -1008
rect 2460 -1038 2688 -1028
rect 3708 -716 4400 -706
rect 5956 -840 6092 -660
rect 6284 -656 6340 -646
rect 6148 -840 6284 -660
rect 6476 -656 6532 -646
rect 6340 -840 6476 -660
rect 6668 -656 6724 -646
rect 6532 -840 6668 -660
rect 6860 -656 6916 -646
rect 6724 -840 6860 -660
rect 5916 -852 6916 -840
rect 4932 -870 5916 -860
rect 6088 -1024 6960 -1014
rect 3708 -1238 4400 -1228
rect 5032 -1052 6088 -1040
rect 5032 -1232 5036 -1052
rect 5092 -1232 5228 -1052
rect 5036 -1246 5092 -1236
rect 5284 -1232 5420 -1052
rect 5228 -1246 5284 -1236
rect 5476 -1232 5612 -1052
rect 5420 -1246 5476 -1236
rect 5668 -1232 5804 -1052
rect 5612 -1246 5668 -1236
rect 5860 -1232 5996 -1052
rect 5804 -1246 5860 -1236
rect 6052 -1224 6088 -1052
rect 6052 -1232 6188 -1224
rect 6088 -1234 6188 -1232
rect 5996 -1246 6052 -1236
rect 6244 -1234 6380 -1224
rect 6188 -1246 6244 -1236
rect 6436 -1234 6572 -1224
rect 6380 -1246 6436 -1236
rect 6628 -1234 6764 -1224
rect 6572 -1246 6628 -1236
rect 6820 -1234 6960 -1224
rect 6764 -1246 6820 -1236
rect 4940 -1272 4996 -1262
rect 4932 -1284 4940 -1274
rect 5132 -1272 5188 -1262
rect 4996 -1284 5132 -1274
rect 5324 -1272 5380 -1262
rect 5188 -1284 5324 -1274
rect 5516 -1272 5572 -1262
rect 5380 -1284 5516 -1274
rect 5708 -1272 5764 -1262
rect 5572 -1284 5708 -1274
rect 5900 -1272 5956 -1262
rect 5764 -1284 5900 -1274
rect 6092 -1272 6148 -1262
rect 4324 -1300 4852 -1290
rect 1944 -1398 2000 -1388
rect 2044 -1422 4324 -1300
rect -232 -1432 176 -1422
rect -232 -1436 120 -1432
rect -1416 -1612 120 -1436
rect 312 -1432 368 -1422
rect 176 -1612 312 -1436
rect 504 -1432 560 -1422
rect 368 -1612 504 -1436
rect 696 -1432 752 -1422
rect 560 -1612 696 -1436
rect 888 -1432 944 -1422
rect 752 -1612 888 -1436
rect 1080 -1432 1136 -1422
rect 944 -1612 1080 -1436
rect 1272 -1432 1328 -1422
rect 1136 -1612 1272 -1436
rect 1464 -1432 1520 -1422
rect 1328 -1612 1464 -1436
rect 1656 -1432 1712 -1422
rect 1520 -1612 1656 -1436
rect 1848 -1432 1904 -1422
rect 1712 -1612 1848 -1436
rect 2040 -1432 4324 -1422
rect 1904 -1612 2040 -1436
rect 2096 -1612 4324 -1432
rect -1416 -1628 4324 -1612
rect 5956 -1456 6092 -1276
rect 6284 -1272 6340 -1262
rect 6148 -1456 6284 -1276
rect 6476 -1272 6532 -1262
rect 6340 -1456 6476 -1276
rect 6668 -1272 6724 -1262
rect 6532 -1456 6668 -1276
rect 6860 -1272 6916 -1262
rect 6724 -1456 6860 -1276
rect 5916 -1468 6916 -1456
rect 4932 -1482 5916 -1472
rect -1416 -1638 4852 -1628
rect -1416 -1746 4528 -1638
rect 6088 -1640 6960 -1630
rect 5032 -1672 6088 -1660
rect -1416 -1756 4780 -1746
rect -1416 -1792 4284 -1756
rect -1416 -1884 -1104 -1792
rect 384 -1884 696 -1792
rect 2184 -1884 4284 -1792
rect -1416 -2072 4284 -1884
rect 5032 -1852 5036 -1672
rect 5092 -1852 5228 -1672
rect 5036 -1866 5092 -1856
rect 5284 -1852 5420 -1672
rect 5228 -1866 5284 -1856
rect 5476 -1852 5612 -1672
rect 5420 -1866 5476 -1856
rect 5668 -1852 5804 -1672
rect 5612 -1866 5668 -1856
rect 5860 -1852 5996 -1672
rect 5804 -1866 5860 -1856
rect 6052 -1840 6088 -1672
rect 6052 -1852 6188 -1840
rect 5996 -1866 6052 -1856
rect 6244 -1852 6380 -1840
rect 6188 -1866 6244 -1856
rect 6436 -1852 6572 -1840
rect 6380 -1866 6436 -1856
rect 6628 -1852 6764 -1840
rect 6572 -1866 6628 -1856
rect 6820 -1850 6960 -1840
rect 6820 -1852 6824 -1850
rect 6764 -1866 6820 -1856
rect 4940 -1892 4996 -1882
rect 4936 -1898 4940 -1896
rect -1416 -2082 4780 -2072
rect 4928 -1908 4940 -1898
rect 5132 -1892 5188 -1882
rect 4996 -1908 5132 -1896
rect 5324 -1892 5380 -1882
rect 5188 -1908 5324 -1896
rect 5516 -1892 5572 -1882
rect 5380 -1908 5516 -1896
rect 5708 -1892 5764 -1882
rect 5572 -1908 5708 -1896
rect 5900 -1892 5956 -1882
rect 5764 -1908 5900 -1896
rect 6092 -1892 6148 -1882
rect 5956 -2076 6092 -1896
rect 6284 -1892 6340 -1882
rect 6148 -2076 6284 -1896
rect 6476 -1892 6532 -1882
rect 6340 -2076 6476 -1896
rect 6668 -1892 6724 -1882
rect 6532 -2076 6668 -1896
rect 6860 -1892 6916 -1882
rect 6724 -2076 6860 -1896
rect -1416 -2120 4296 -2082
rect 5912 -2088 6916 -2076
rect 4928 -2106 5912 -2096
rect -1416 -2128 696 -2120
rect -2364 -2344 -1544 -2340
rect -1416 -2344 -1104 -2128
rect -2364 -2352 -1104 -2344
rect -2312 -2532 -2172 -2352
rect -2120 -2532 -1980 -2352
rect -1928 -2532 -1788 -2352
rect -1736 -2532 -1596 -2352
rect -1544 -2532 -1104 -2352
rect -2364 -2542 -2312 -2532
rect -2172 -2542 -2120 -2532
rect -1980 -2542 -1928 -2532
rect -1788 -2542 -1736 -2532
rect -1596 -2542 -1544 -2532
rect -2460 -2574 -2408 -2566
rect -2268 -2574 -2216 -2566
rect -2076 -2574 -2024 -2566
rect -1884 -2574 -1832 -2566
rect -2464 -2576 -1832 -2574
rect -1692 -2576 -1640 -2566
rect -1500 -2576 -1448 -2566
rect -2464 -2584 -2460 -2576
rect -2408 -2584 -2268 -2576
rect -2216 -2584 -2076 -2576
rect -2024 -2584 -1884 -2576
rect -1832 -2756 -1692 -2576
rect -1640 -2756 -1500 -2576
rect -1860 -2764 -1448 -2756
rect -1860 -2766 -1832 -2764
rect -1692 -2766 -1640 -2764
rect -1500 -2766 -1448 -2764
rect -2464 -2778 -1860 -2768
rect -2364 -2960 -1544 -2956
rect -1416 -2960 -1104 -2532
rect -564 -2344 256 -2340
rect 384 -2344 696 -2128
rect 2184 -2144 4296 -2120
rect 4412 -2144 4696 -2138
rect 2184 -2148 4696 -2144
rect 2184 -2176 4412 -2148
rect -564 -2352 696 -2344
rect -512 -2532 -372 -2352
rect -320 -2532 -180 -2352
rect -128 -2532 12 -2352
rect 64 -2532 204 -2352
rect 256 -2532 696 -2352
rect -564 -2542 -512 -2532
rect -372 -2542 -320 -2532
rect -180 -2542 -128 -2532
rect 12 -2542 64 -2532
rect 204 -2542 256 -2532
rect -660 -2574 -608 -2566
rect -468 -2574 -416 -2566
rect -276 -2574 -224 -2566
rect -84 -2574 -32 -2566
rect -664 -2576 -32 -2574
rect 108 -2576 160 -2566
rect 300 -2576 352 -2566
rect -664 -2584 -660 -2576
rect -608 -2584 -468 -2576
rect -416 -2584 -276 -2576
rect -224 -2584 -84 -2576
rect -32 -2756 108 -2576
rect 160 -2756 300 -2576
rect -60 -2764 352 -2756
rect -60 -2766 -32 -2764
rect 108 -2766 160 -2764
rect 300 -2766 352 -2764
rect -664 -2778 -60 -2768
rect -2364 -2968 -1104 -2960
rect -3080 -3136 -2648 -3126
rect -3484 -3412 -3080 -3402
rect -2312 -3148 -2172 -2968
rect -2120 -3148 -1980 -2968
rect -1928 -3148 -1788 -2968
rect -1736 -3148 -1596 -2968
rect -1544 -3148 -1104 -2968
rect -2364 -3158 -2312 -3148
rect -2172 -3158 -2120 -3148
rect -1980 -3158 -1928 -3148
rect -1788 -3158 -1736 -3148
rect -1596 -3158 -1544 -3148
rect -2460 -3190 -2408 -3182
rect -2268 -3190 -2216 -3182
rect -2076 -3190 -2024 -3182
rect -1884 -3190 -1832 -3182
rect -2464 -3192 -1832 -3190
rect -1692 -3192 -1640 -3182
rect -1500 -3192 -1448 -3182
rect -2464 -3200 -2460 -3192
rect -2408 -3200 -2268 -3192
rect -2216 -3200 -2076 -3192
rect -2024 -3200 -1884 -3192
rect -1832 -3372 -1692 -3192
rect -1640 -3372 -1500 -3192
rect -1860 -3380 -1448 -3372
rect -1860 -3382 -1832 -3380
rect -1692 -3382 -1640 -3380
rect -1500 -3382 -1448 -3380
rect -2464 -3394 -1860 -3384
rect -2364 -3584 -2312 -3578
rect -2172 -3584 -2120 -3578
rect -1980 -3584 -1928 -3578
rect -1788 -3584 -1736 -3578
rect -1596 -3584 -1544 -3578
rect -1416 -3584 -1104 -3148
rect -564 -2960 256 -2956
rect 384 -2960 696 -2532
rect 1236 -2344 2056 -2340
rect 2184 -2344 2496 -2176
rect 1236 -2352 2496 -2344
rect 1288 -2532 1428 -2352
rect 1480 -2532 1620 -2352
rect 1672 -2532 1812 -2352
rect 1864 -2532 2004 -2352
rect 2056 -2532 2496 -2352
rect 1236 -2542 1288 -2532
rect 1428 -2542 1480 -2532
rect 1620 -2542 1672 -2532
rect 1812 -2542 1864 -2532
rect 2004 -2542 2056 -2532
rect 1140 -2574 1192 -2566
rect 1332 -2574 1384 -2566
rect 1524 -2574 1576 -2566
rect 1716 -2574 1768 -2566
rect 1136 -2576 1768 -2574
rect 1908 -2576 1960 -2566
rect 2100 -2576 2152 -2566
rect 1136 -2584 1140 -2576
rect 1192 -2584 1332 -2576
rect 1384 -2584 1524 -2576
rect 1576 -2584 1716 -2576
rect 1768 -2756 1908 -2576
rect 1960 -2756 2100 -2576
rect 1740 -2764 2152 -2756
rect 1740 -2766 1768 -2764
rect 1908 -2766 1960 -2764
rect 2100 -2766 2152 -2764
rect 1136 -2778 1740 -2768
rect -564 -2968 696 -2960
rect -512 -3148 -372 -2968
rect -320 -3148 -180 -2968
rect -128 -3148 12 -2968
rect 64 -3148 204 -2968
rect 256 -3148 696 -2968
rect -564 -3158 -512 -3148
rect -372 -3158 -320 -3148
rect -180 -3158 -128 -3148
rect 12 -3158 64 -3148
rect 204 -3158 256 -3148
rect -660 -3190 -608 -3182
rect -468 -3190 -416 -3182
rect -276 -3190 -224 -3182
rect -84 -3190 -32 -3182
rect -664 -3192 -32 -3190
rect 108 -3192 160 -3182
rect 300 -3192 352 -3182
rect -664 -3200 -660 -3192
rect -608 -3200 -468 -3192
rect -416 -3200 -276 -3192
rect -224 -3200 -84 -3192
rect -32 -3372 108 -3192
rect 160 -3372 300 -3192
rect -60 -3380 352 -3372
rect -60 -3382 -32 -3380
rect 108 -3382 160 -3380
rect 300 -3382 352 -3380
rect -664 -3394 -60 -3384
rect -2364 -3588 -1104 -3584
rect -2312 -3768 -2172 -3588
rect -2120 -3768 -1980 -3588
rect -1928 -3768 -1788 -3588
rect -1736 -3768 -1596 -3588
rect -1544 -3768 -1104 -3588
rect -2364 -3772 -1104 -3768
rect -564 -3584 -512 -3578
rect -372 -3584 -320 -3578
rect -180 -3584 -128 -3578
rect 12 -3584 64 -3578
rect 204 -3584 256 -3578
rect 384 -3584 696 -3148
rect 1236 -2960 2056 -2956
rect 2184 -2960 2496 -2532
rect 3036 -2344 3856 -2340
rect 3984 -2344 4412 -2176
rect 3036 -2352 4412 -2344
rect 3088 -2532 3228 -2352
rect 3280 -2532 3420 -2352
rect 3472 -2532 3612 -2352
rect 3664 -2532 3804 -2352
rect 3856 -2532 4412 -2352
rect 3036 -2542 3088 -2532
rect 3228 -2542 3280 -2532
rect 3420 -2542 3472 -2532
rect 3612 -2542 3664 -2532
rect 3804 -2542 3856 -2532
rect 2940 -2574 2992 -2566
rect 3132 -2574 3184 -2566
rect 3324 -2574 3376 -2566
rect 3516 -2574 3568 -2566
rect 2936 -2576 3568 -2574
rect 3708 -2576 3760 -2566
rect 3900 -2576 3952 -2566
rect 2936 -2584 2940 -2576
rect 2992 -2584 3132 -2576
rect 3184 -2584 3324 -2576
rect 3376 -2584 3516 -2576
rect 3568 -2756 3708 -2576
rect 3760 -2756 3900 -2576
rect 3540 -2764 3952 -2756
rect 3540 -2766 3568 -2764
rect 3708 -2766 3760 -2764
rect 3900 -2766 3952 -2764
rect 3984 -2644 4412 -2532
rect 2936 -2778 3540 -2768
rect 1236 -2968 2496 -2960
rect 1288 -3148 1428 -2968
rect 1480 -3148 1620 -2968
rect 1672 -3148 1812 -2968
rect 1864 -3148 2004 -2968
rect 2056 -3148 2496 -2968
rect 1236 -3158 1288 -3148
rect 1428 -3158 1480 -3148
rect 1620 -3158 1672 -3148
rect 1812 -3158 1864 -3148
rect 2004 -3158 2056 -3148
rect 1140 -3190 1192 -3182
rect 1332 -3190 1384 -3182
rect 1524 -3190 1576 -3182
rect 1716 -3190 1768 -3182
rect 1136 -3192 1768 -3190
rect 1908 -3192 1960 -3182
rect 2100 -3192 2152 -3182
rect 1136 -3200 1140 -3192
rect 1192 -3200 1332 -3192
rect 1384 -3200 1524 -3192
rect 1576 -3200 1716 -3192
rect 1768 -3372 1908 -3192
rect 1960 -3372 2100 -3192
rect 1740 -3380 2152 -3372
rect 1740 -3382 1768 -3380
rect 1908 -3382 1960 -3380
rect 2100 -3382 2152 -3380
rect 1136 -3394 1740 -3384
rect -564 -3588 696 -3584
rect -512 -3768 -372 -3588
rect -320 -3768 -180 -3588
rect -128 -3768 12 -3588
rect 64 -3768 204 -3588
rect 256 -3768 696 -3588
rect -564 -3772 696 -3768
rect 1236 -3584 1288 -3578
rect 1428 -3584 1480 -3578
rect 1620 -3584 1672 -3578
rect 1812 -3584 1864 -3578
rect 2004 -3584 2056 -3578
rect 2184 -3584 2496 -3148
rect 3036 -2960 3856 -2956
rect 3984 -2960 4296 -2644
rect 6084 -2260 6956 -2250
rect 5032 -2288 6084 -2276
rect 5032 -2468 5036 -2288
rect 5092 -2468 5228 -2288
rect 5036 -2482 5092 -2472
rect 5284 -2468 5420 -2288
rect 5228 -2482 5284 -2472
rect 5476 -2468 5612 -2288
rect 5420 -2482 5476 -2472
rect 5668 -2468 5804 -2288
rect 5612 -2482 5668 -2472
rect 5860 -2468 5996 -2288
rect 5804 -2482 5860 -2472
rect 6052 -2460 6084 -2288
rect 6052 -2468 6188 -2460
rect 6084 -2470 6188 -2468
rect 5996 -2482 6052 -2472
rect 6244 -2470 6380 -2460
rect 6188 -2482 6244 -2472
rect 6436 -2470 6572 -2460
rect 6380 -2482 6436 -2472
rect 6628 -2470 6764 -2460
rect 6572 -2482 6628 -2472
rect 6820 -2470 6956 -2460
rect 6764 -2482 6820 -2472
rect 4940 -2508 4996 -2498
rect 4412 -2658 4696 -2648
rect 4928 -2520 4940 -2510
rect 5132 -2508 5188 -2498
rect 4996 -2520 5132 -2510
rect 5324 -2508 5380 -2498
rect 5188 -2520 5324 -2510
rect 5516 -2508 5572 -2498
rect 5380 -2520 5516 -2510
rect 5708 -2508 5764 -2498
rect 5572 -2520 5708 -2510
rect 5900 -2508 5956 -2498
rect 5764 -2520 5900 -2510
rect 6092 -2508 6148 -2498
rect 5956 -2692 6092 -2512
rect 6284 -2508 6340 -2498
rect 6148 -2692 6284 -2512
rect 6476 -2508 6532 -2498
rect 6340 -2692 6476 -2512
rect 6668 -2508 6724 -2498
rect 6532 -2692 6668 -2512
rect 6860 -2508 6916 -2498
rect 6724 -2692 6860 -2512
rect 5912 -2704 6916 -2692
rect 4928 -2718 5912 -2708
rect 6084 -2880 6956 -2870
rect 3036 -2968 4296 -2960
rect 3088 -3148 3228 -2968
rect 3280 -3148 3420 -2968
rect 3472 -3148 3612 -2968
rect 3664 -3148 3804 -2968
rect 3856 -3148 4296 -2968
rect 5032 -2908 6084 -2896
rect 5032 -3088 5036 -2908
rect 5092 -3088 5228 -2908
rect 5036 -3102 5092 -3092
rect 5284 -3088 5420 -2908
rect 5228 -3102 5284 -3092
rect 5476 -3088 5612 -2908
rect 5420 -3102 5476 -3092
rect 5668 -3088 5804 -2908
rect 5612 -3102 5668 -3092
rect 5860 -3088 5996 -2908
rect 5804 -3102 5860 -3092
rect 6052 -3080 6084 -2908
rect 6052 -3088 6188 -3080
rect 6084 -3090 6188 -3088
rect 5996 -3102 6052 -3092
rect 6244 -3090 6380 -3080
rect 6188 -3102 6244 -3092
rect 6436 -3090 6572 -3080
rect 6380 -3102 6436 -3092
rect 6628 -3090 6764 -3080
rect 6572 -3102 6628 -3092
rect 6820 -3090 6956 -3080
rect 6764 -3102 6820 -3092
rect 4940 -3128 4996 -3118
rect 4936 -3134 4940 -3132
rect 3036 -3158 3088 -3148
rect 3228 -3158 3280 -3148
rect 3420 -3158 3472 -3148
rect 3612 -3158 3664 -3148
rect 3804 -3158 3856 -3148
rect 2940 -3190 2992 -3182
rect 3132 -3190 3184 -3182
rect 3324 -3190 3376 -3182
rect 3516 -3190 3568 -3182
rect 2936 -3192 3568 -3190
rect 3708 -3192 3760 -3182
rect 3900 -3192 3952 -3182
rect 2936 -3200 2940 -3192
rect 2992 -3200 3132 -3192
rect 3184 -3200 3324 -3192
rect 3376 -3200 3516 -3192
rect 3568 -3372 3708 -3192
rect 3760 -3372 3900 -3192
rect 3540 -3380 3952 -3372
rect 3540 -3382 3568 -3380
rect 3708 -3382 3760 -3380
rect 3900 -3382 3952 -3380
rect 2936 -3394 3540 -3384
rect 1236 -3588 2496 -3584
rect 1288 -3768 1428 -3588
rect 1480 -3768 1620 -3588
rect 1672 -3768 1812 -3588
rect 1864 -3768 2004 -3588
rect 2056 -3768 2496 -3588
rect 1236 -3772 2496 -3768
rect 3036 -3584 3088 -3578
rect 3228 -3584 3280 -3578
rect 3420 -3584 3472 -3578
rect 3612 -3584 3664 -3578
rect 3804 -3584 3856 -3578
rect 3984 -3584 4296 -3148
rect 4928 -3144 4940 -3134
rect 5132 -3128 5188 -3118
rect 4996 -3144 5132 -3132
rect 5324 -3128 5380 -3118
rect 5188 -3144 5324 -3132
rect 5516 -3128 5572 -3118
rect 5380 -3144 5516 -3132
rect 5708 -3128 5764 -3118
rect 5572 -3144 5708 -3132
rect 5900 -3128 5956 -3118
rect 5764 -3144 5900 -3132
rect 6092 -3128 6148 -3118
rect 5956 -3312 6092 -3132
rect 6284 -3128 6340 -3118
rect 6148 -3312 6284 -3132
rect 6476 -3128 6532 -3118
rect 6340 -3312 6476 -3132
rect 6668 -3128 6724 -3118
rect 6532 -3312 6668 -3132
rect 6860 -3128 6916 -3118
rect 6724 -3312 6860 -3132
rect 5912 -3324 6916 -3312
rect 4928 -3342 5912 -3332
rect 3036 -3588 4296 -3584
rect 3088 -3768 3228 -3588
rect 3280 -3768 3420 -3588
rect 3472 -3768 3612 -3588
rect 3664 -3768 3804 -3588
rect 3856 -3768 4296 -3588
rect 3036 -3772 4296 -3768
rect -2364 -3778 -2312 -3772
rect -2172 -3778 -2120 -3772
rect -1980 -3778 -1928 -3772
rect -1788 -3778 -1736 -3772
rect -1596 -3778 -1544 -3772
rect -564 -3778 -512 -3772
rect -372 -3778 -320 -3772
rect -180 -3778 -128 -3772
rect 12 -3778 64 -3772
rect 204 -3778 256 -3772
rect 1236 -3778 1288 -3772
rect 1428 -3778 1480 -3772
rect 1620 -3778 1672 -3772
rect 1812 -3778 1864 -3772
rect 2004 -3778 2056 -3772
rect 3036 -3778 3088 -3772
rect 3228 -3778 3280 -3772
rect 3420 -3778 3472 -3772
rect 3612 -3778 3664 -3772
rect 3804 -3778 3856 -3772
rect -2460 -3810 -2408 -3802
rect -2268 -3810 -2216 -3802
rect -2076 -3810 -2024 -3802
rect -1884 -3810 -1832 -3802
rect -3484 -3828 -3080 -3824
rect -3484 -3834 -2648 -3828
rect -3080 -3838 -2648 -3834
rect -2468 -3812 -1832 -3810
rect -1692 -3812 -1640 -3802
rect -1500 -3812 -1448 -3802
rect -660 -3810 -608 -3802
rect -468 -3810 -416 -3802
rect -276 -3810 -224 -3802
rect -84 -3810 -32 -3802
rect -2468 -3820 -2460 -3812
rect -2408 -3820 -2268 -3812
rect -2216 -3820 -2076 -3812
rect -2024 -3820 -1884 -3812
rect -1832 -3992 -1692 -3812
rect -1640 -3992 -1500 -3812
rect -1864 -4000 -1448 -3992
rect -1864 -4002 -1832 -4000
rect -1692 -4002 -1640 -4000
rect -1500 -4002 -1448 -4000
rect -668 -3812 -32 -3810
rect 108 -3812 160 -3802
rect 300 -3812 352 -3802
rect 1140 -3810 1192 -3802
rect 1332 -3810 1384 -3802
rect 1524 -3810 1576 -3802
rect 1716 -3810 1768 -3802
rect -668 -3820 -660 -3812
rect -608 -3820 -468 -3812
rect -416 -3820 -276 -3812
rect -224 -3820 -84 -3812
rect -32 -3992 108 -3812
rect 160 -3992 300 -3812
rect -2468 -4014 -1864 -4004
rect -64 -4000 352 -3992
rect -64 -4002 -32 -4000
rect 108 -4002 160 -4000
rect 300 -4002 352 -4000
rect 1132 -3812 1768 -3810
rect 1908 -3812 1960 -3802
rect 2100 -3812 2152 -3802
rect 2940 -3810 2992 -3802
rect 3132 -3810 3184 -3802
rect 3324 -3810 3376 -3802
rect 3516 -3810 3568 -3802
rect 1132 -3820 1140 -3812
rect 1192 -3820 1332 -3812
rect 1384 -3820 1524 -3812
rect 1576 -3820 1716 -3812
rect 1768 -3992 1908 -3812
rect 1960 -3992 2100 -3812
rect -668 -4014 -64 -4004
rect 1736 -4000 2152 -3992
rect 1736 -4002 1768 -4000
rect 1908 -4002 1960 -4000
rect 2100 -4002 2152 -4000
rect 2932 -3812 3568 -3810
rect 3708 -3812 3760 -3802
rect 3900 -3812 3952 -3802
rect 2932 -3820 2940 -3812
rect 2992 -3820 3132 -3812
rect 3184 -3820 3324 -3812
rect 3376 -3820 3516 -3812
rect 3568 -3992 3708 -3812
rect 3760 -3992 3900 -3812
rect 1132 -4014 1736 -4004
rect 3536 -4000 3952 -3992
rect 3536 -4002 3568 -4000
rect 3708 -4002 3760 -4000
rect 3900 -4002 3952 -4000
rect 2932 -4014 3536 -4004
rect -2460 -4488 -1860 -4478
rect -1440 -4488 4036 -4464
rect -1860 -4500 -660 -4488
rect -60 -4500 1140 -4488
rect 1740 -4500 2940 -4488
rect 3540 -4500 4036 -4488
rect -1860 -4672 -1428 -4500
rect -2408 -4680 -1944 -4672
rect -1892 -4680 -1428 -4672
rect -1376 -4680 -660 -4500
rect -60 -4672 372 -4500
rect -608 -4680 -144 -4672
rect -92 -4680 372 -4672
rect 424 -4680 1140 -4500
rect 1740 -4672 2172 -4500
rect 1192 -4680 1656 -4672
rect 1708 -4680 2172 -4672
rect 2224 -4680 2940 -4500
rect 3540 -4672 3972 -4500
rect 2992 -4680 3456 -4672
rect 3508 -4680 3972 -4672
rect 4024 -4680 4036 -4500
rect -2460 -4682 -1860 -4680
rect -2460 -4690 -2408 -4682
rect -1944 -4690 -1892 -4682
rect -1428 -4690 -1376 -4680
rect -660 -4682 -60 -4680
rect -660 -4690 -608 -4682
rect -144 -4690 -92 -4682
rect 372 -4690 424 -4680
rect 1140 -4682 1740 -4680
rect 1140 -4690 1192 -4682
rect 1656 -4690 1708 -4682
rect 2172 -4690 2224 -4680
rect 2940 -4682 3540 -4680
rect 2940 -4690 2992 -4682
rect 3456 -4690 3508 -4682
rect 3972 -4690 4024 -4680
rect -2200 -4720 -2148 -4710
rect -1684 -4718 -1632 -4710
rect -1168 -4718 -1116 -4710
rect -1716 -4720 -1116 -4718
rect -2148 -4728 -1684 -4720
rect -1632 -4728 -1168 -4720
rect -2148 -4900 -1716 -4728
rect -2200 -4912 -1716 -4900
rect -400 -4720 -348 -4710
rect 116 -4718 168 -4710
rect 632 -4718 684 -4710
rect 84 -4720 684 -4718
rect -348 -4728 116 -4720
rect 168 -4728 632 -4720
rect -348 -4900 84 -4728
rect -400 -4912 84 -4900
rect 1400 -4720 1452 -4710
rect 1916 -4718 1968 -4710
rect 2432 -4718 2484 -4710
rect 1884 -4720 2484 -4718
rect 1452 -4728 1916 -4720
rect 1968 -4728 2432 -4720
rect 1452 -4900 1884 -4728
rect 1400 -4912 1884 -4900
rect 3200 -4720 3252 -4710
rect 3716 -4718 3768 -4710
rect 4232 -4718 4284 -4710
rect 3684 -4720 4284 -4718
rect 3252 -4728 3716 -4720
rect 3768 -4728 4232 -4720
rect 3252 -4900 3684 -4728
rect 3200 -4912 3684 -4900
rect -1716 -4922 -1116 -4912
rect 84 -4922 684 -4912
rect 1884 -4922 2484 -4912
rect 3684 -4922 4284 -4912
rect -2460 -5104 -1860 -5094
rect -660 -5104 -60 -5094
rect 1140 -5104 1740 -5094
rect 2940 -5104 3540 -5094
rect -1860 -5116 -1376 -5104
rect -1860 -5288 -1428 -5116
rect -2408 -5296 -1944 -5288
rect -1892 -5296 -1428 -5288
rect -2460 -5298 -1860 -5296
rect -2460 -5306 -2408 -5298
rect -1944 -5306 -1892 -5298
rect -1428 -5306 -1376 -5296
rect -60 -5116 424 -5104
rect -60 -5288 372 -5116
rect -608 -5296 -144 -5288
rect -92 -5296 372 -5288
rect -660 -5298 -60 -5296
rect -660 -5306 -608 -5298
rect -144 -5306 -92 -5298
rect 372 -5306 424 -5296
rect 1740 -5116 2224 -5104
rect 1740 -5288 2172 -5116
rect 1192 -5296 1656 -5288
rect 1708 -5296 2172 -5288
rect 1140 -5298 1740 -5296
rect 1140 -5306 1192 -5298
rect 1656 -5306 1708 -5298
rect 2172 -5306 2224 -5296
rect 3540 -5116 4024 -5104
rect 3540 -5288 3972 -5116
rect 2992 -5296 3456 -5288
rect 3508 -5296 3972 -5288
rect 2940 -5298 3540 -5296
rect 2940 -5306 2992 -5298
rect 3456 -5306 3508 -5298
rect 3972 -5306 4024 -5296
rect -2200 -5336 -2148 -5326
rect -1684 -5334 -1632 -5326
rect -1168 -5334 -1116 -5326
rect -1716 -5336 -1116 -5334
rect -2148 -5344 -1684 -5336
rect -1632 -5344 -1168 -5336
rect -2148 -5516 -1716 -5344
rect -2200 -5528 -1716 -5516
rect -400 -5336 -348 -5326
rect 116 -5334 168 -5326
rect 632 -5334 684 -5326
rect 84 -5336 684 -5334
rect -348 -5344 116 -5336
rect 168 -5344 632 -5336
rect -348 -5516 84 -5344
rect -400 -5528 84 -5516
rect 1400 -5336 1452 -5326
rect 1916 -5334 1968 -5326
rect 2432 -5334 2484 -5326
rect 1884 -5336 2484 -5334
rect 1452 -5344 1916 -5336
rect 1968 -5344 2432 -5336
rect 1452 -5516 1884 -5344
rect 1400 -5528 1884 -5516
rect 3200 -5336 3252 -5326
rect 3716 -5334 3768 -5326
rect 4232 -5334 4284 -5326
rect 3684 -5336 4284 -5334
rect 3252 -5344 3716 -5336
rect 3768 -5344 4232 -5336
rect 3252 -5516 3684 -5344
rect 3200 -5528 3684 -5516
rect -1716 -5538 -1116 -5528
rect 84 -5538 684 -5528
rect 1884 -5538 2484 -5528
rect 3684 -5538 4284 -5528
rect -2460 -5724 -1860 -5714
rect -660 -5724 -60 -5714
rect 1140 -5724 1740 -5714
rect 2940 -5724 3540 -5714
rect -1860 -5736 -1376 -5724
rect -1860 -5908 -1428 -5736
rect -2408 -5916 -1944 -5908
rect -1892 -5916 -1428 -5908
rect -2460 -5918 -1860 -5916
rect -2460 -5926 -2408 -5918
rect -1944 -5926 -1892 -5918
rect -1428 -5926 -1376 -5916
rect -60 -5736 424 -5724
rect -60 -5908 372 -5736
rect -608 -5916 -144 -5908
rect -92 -5916 372 -5908
rect -660 -5918 -60 -5916
rect -660 -5926 -608 -5918
rect -144 -5926 -92 -5918
rect 372 -5926 424 -5916
rect 1740 -5736 2224 -5724
rect 1740 -5908 2172 -5736
rect 1192 -5916 1656 -5908
rect 1708 -5916 2172 -5908
rect 1140 -5918 1740 -5916
rect 1140 -5926 1192 -5918
rect 1656 -5926 1708 -5918
rect 2172 -5926 2224 -5916
rect 3540 -5736 4024 -5724
rect 3540 -5908 3972 -5736
rect 2992 -5916 3456 -5908
rect 3508 -5916 3972 -5908
rect 2940 -5918 3540 -5916
rect 2940 -5926 2992 -5918
rect 3456 -5926 3508 -5918
rect 3972 -5926 4024 -5916
rect -2200 -5956 -2148 -5946
rect -1684 -5954 -1632 -5946
rect -1168 -5954 -1116 -5946
rect -1716 -5956 -1116 -5954
rect -2148 -5964 -1684 -5956
rect -1632 -5964 -1168 -5956
rect -2148 -6136 -1716 -5964
rect -2200 -6148 -1716 -6136
rect -400 -5956 -348 -5946
rect 116 -5954 168 -5946
rect 632 -5954 684 -5946
rect 84 -5956 684 -5954
rect -348 -5964 116 -5956
rect 168 -5964 632 -5956
rect -348 -6136 84 -5964
rect -400 -6148 84 -6136
rect 1400 -5956 1452 -5946
rect 1916 -5954 1968 -5946
rect 2432 -5954 2484 -5946
rect 1884 -5956 2484 -5954
rect 1452 -5964 1916 -5956
rect 1968 -5964 2432 -5956
rect 1452 -6136 1884 -5964
rect 1400 -6148 1884 -6136
rect 3200 -5956 3252 -5946
rect 3716 -5954 3768 -5946
rect 4232 -5954 4284 -5946
rect 3684 -5956 4284 -5954
rect 3252 -5964 3716 -5956
rect 3768 -5964 4232 -5956
rect 3252 -6136 3684 -5964
rect 3200 -6148 3684 -6136
rect -1716 -6158 -1116 -6148
rect 84 -6158 684 -6148
rect 1884 -6158 2484 -6148
rect 3684 -6158 4284 -6148
rect -2460 -6340 -1860 -6330
rect -660 -6340 -60 -6330
rect 1140 -6340 1740 -6330
rect 2940 -6340 3540 -6330
rect -1860 -6352 -1376 -6340
rect -1860 -6524 -1428 -6352
rect -2408 -6532 -1944 -6524
rect -1892 -6532 -1428 -6524
rect -2460 -6534 -1860 -6532
rect -2460 -6542 -2408 -6534
rect -1944 -6542 -1892 -6534
rect -1428 -6542 -1376 -6532
rect -60 -6352 424 -6340
rect -60 -6524 372 -6352
rect -608 -6532 -144 -6524
rect -92 -6532 372 -6524
rect -660 -6534 -60 -6532
rect -660 -6542 -608 -6534
rect -144 -6542 -92 -6534
rect 372 -6542 424 -6532
rect 1740 -6352 2224 -6340
rect 1740 -6524 2172 -6352
rect 1192 -6532 1656 -6524
rect 1708 -6532 2172 -6524
rect 1140 -6534 1740 -6532
rect 1140 -6542 1192 -6534
rect 1656 -6542 1708 -6534
rect 2172 -6542 2224 -6532
rect 3540 -6352 4024 -6340
rect 3540 -6524 3972 -6352
rect 2992 -6532 3456 -6524
rect 3508 -6532 3972 -6524
rect 2940 -6534 3540 -6532
rect 2940 -6542 2992 -6534
rect 3456 -6542 3508 -6534
rect 3972 -6542 4024 -6532
rect -2200 -6572 -2148 -6562
rect -1684 -6570 -1632 -6562
rect -1168 -6570 -1116 -6562
rect -1716 -6572 -1116 -6570
rect -2148 -6580 -1684 -6572
rect -1632 -6580 -1168 -6572
rect -2148 -6752 -1716 -6580
rect -2200 -6764 -1716 -6752
rect -400 -6572 -348 -6562
rect 116 -6570 168 -6562
rect 632 -6570 684 -6562
rect 84 -6572 684 -6570
rect -348 -6580 116 -6572
rect 168 -6580 632 -6572
rect -348 -6752 84 -6580
rect -400 -6764 84 -6752
rect 1400 -6572 1452 -6562
rect 1916 -6570 1968 -6562
rect 2432 -6570 2484 -6562
rect 1884 -6572 2484 -6570
rect 1452 -6580 1916 -6572
rect 1968 -6580 2432 -6572
rect 1452 -6752 1884 -6580
rect 1400 -6764 1884 -6752
rect 3200 -6572 3252 -6562
rect 3716 -6570 3768 -6562
rect 4232 -6570 4284 -6562
rect 3684 -6572 4284 -6570
rect 3252 -6580 3716 -6572
rect 3768 -6580 4232 -6572
rect 3252 -6752 3684 -6580
rect 3200 -6764 3684 -6752
rect -1716 -6774 -1116 -6764
rect 84 -6774 684 -6764
rect 1884 -6774 2484 -6764
rect 3684 -6774 4284 -6764
rect -2460 -6960 -1860 -6950
rect -660 -6960 -60 -6950
rect 1140 -6960 1740 -6950
rect 2940 -6960 3540 -6950
rect -1860 -6972 -1376 -6960
rect -1860 -7144 -1428 -6972
rect -2408 -7152 -1944 -7144
rect -1892 -7152 -1428 -7144
rect -2460 -7154 -1860 -7152
rect -2460 -7162 -2408 -7154
rect -1944 -7162 -1892 -7154
rect -1428 -7162 -1376 -7152
rect -60 -6972 424 -6960
rect -60 -7144 372 -6972
rect -608 -7152 -144 -7144
rect -92 -7152 372 -7144
rect -660 -7154 -60 -7152
rect -660 -7162 -608 -7154
rect -144 -7162 -92 -7154
rect 372 -7162 424 -7152
rect 1740 -6972 2224 -6960
rect 1740 -7144 2172 -6972
rect 1192 -7152 1656 -7144
rect 1708 -7152 2172 -7144
rect 1140 -7154 1740 -7152
rect 1140 -7162 1192 -7154
rect 1656 -7162 1708 -7154
rect 2172 -7162 2224 -7152
rect 3540 -6972 4024 -6960
rect 3540 -7144 3972 -6972
rect 2992 -7152 3456 -7144
rect 3508 -7152 3972 -7144
rect 2940 -7154 3540 -7152
rect 2940 -7162 2992 -7154
rect 3456 -7162 3508 -7154
rect 3972 -7162 4024 -7152
rect -2200 -7192 -2148 -7182
rect -1684 -7190 -1632 -7182
rect -1168 -7190 -1116 -7182
rect -1716 -7192 -1116 -7190
rect -2148 -7200 -1684 -7192
rect -1632 -7200 -1168 -7192
rect -2148 -7372 -1716 -7200
rect -2200 -7384 -1716 -7372
rect -400 -7192 -348 -7182
rect 116 -7190 168 -7182
rect 632 -7190 684 -7182
rect 84 -7192 684 -7190
rect -348 -7200 116 -7192
rect 168 -7200 632 -7192
rect -348 -7372 84 -7200
rect -400 -7384 84 -7372
rect 1400 -7192 1452 -7182
rect 1916 -7190 1968 -7182
rect 2432 -7190 2484 -7182
rect 1884 -7192 2484 -7190
rect 1452 -7200 1916 -7192
rect 1968 -7200 2432 -7192
rect 1452 -7372 1884 -7200
rect 1400 -7384 1884 -7372
rect 3200 -7192 3252 -7182
rect 3716 -7190 3768 -7182
rect 4232 -7190 4284 -7182
rect 3684 -7192 4284 -7190
rect 3252 -7200 3716 -7192
rect 3768 -7200 4232 -7192
rect 3252 -7372 3684 -7200
rect 3200 -7384 3684 -7372
rect -1716 -7394 -1116 -7384
rect 84 -7394 684 -7384
rect 1884 -7394 2484 -7384
rect 3684 -7394 4284 -7384
rect -2460 -7576 -1860 -7566
rect -660 -7576 -60 -7566
rect 1140 -7576 1740 -7566
rect 2940 -7576 3540 -7566
rect -1860 -7588 -1376 -7576
rect -1860 -7760 -1428 -7588
rect -2408 -7768 -1944 -7760
rect -1892 -7768 -1428 -7760
rect -2460 -7770 -1860 -7768
rect -2460 -7778 -2408 -7770
rect -1944 -7778 -1892 -7770
rect -1428 -7778 -1376 -7768
rect -60 -7588 424 -7576
rect -60 -7760 372 -7588
rect -608 -7768 -144 -7760
rect -92 -7768 372 -7760
rect -660 -7770 -60 -7768
rect -660 -7778 -608 -7770
rect -144 -7778 -92 -7770
rect 372 -7778 424 -7768
rect 1740 -7588 2224 -7576
rect 1740 -7760 2172 -7588
rect 1192 -7768 1656 -7760
rect 1708 -7768 2172 -7760
rect 1140 -7770 1740 -7768
rect 1140 -7778 1192 -7770
rect 1656 -7778 1708 -7770
rect 2172 -7778 2224 -7768
rect 3540 -7588 4024 -7576
rect 3540 -7760 3972 -7588
rect 2992 -7768 3456 -7760
rect 3508 -7768 3972 -7760
rect 2940 -7770 3540 -7768
rect 2940 -7778 2992 -7770
rect 3456 -7778 3508 -7770
rect 3972 -7778 4024 -7768
rect -2200 -7808 -2148 -7798
rect -1684 -7806 -1632 -7798
rect -1168 -7806 -1116 -7798
rect -1716 -7808 -1116 -7806
rect -2148 -7816 -1684 -7808
rect -1632 -7816 -1168 -7808
rect -2148 -7988 -1716 -7816
rect -400 -7808 -348 -7798
rect 116 -7806 168 -7798
rect 632 -7806 684 -7798
rect 84 -7808 684 -7806
rect -2200 -8000 -1716 -7988
rect -1716 -8010 -1116 -8000
rect -980 -7960 -800 -7950
rect -348 -7816 116 -7808
rect 168 -7816 632 -7808
rect -348 -7988 84 -7816
rect -400 -8000 84 -7988
rect 1400 -7808 1452 -7798
rect 1916 -7806 1968 -7798
rect 2432 -7806 2484 -7798
rect 1884 -7808 2484 -7806
rect 1452 -7816 1916 -7808
rect 1968 -7816 2432 -7808
rect 1452 -7988 1884 -7816
rect 1400 -8000 1884 -7988
rect 3200 -7808 3252 -7798
rect 3716 -7806 3768 -7798
rect 4232 -7806 4284 -7798
rect 3684 -7808 4284 -7806
rect 3252 -7816 3716 -7808
rect 3768 -7816 4232 -7808
rect 3252 -7988 3684 -7816
rect 3200 -8000 3684 -7988
rect 84 -8010 684 -8000
rect 1884 -8010 2484 -8000
rect 3684 -8010 4284 -8000
rect -980 -8170 -800 -8160
rect -5444 -8610 -4636 -8600
rect -5444 -9426 -4636 -9416
<< via2 >>
rect 3420 2380 3600 2580
rect -80 1676 2096 2112
rect 3536 2056 4512 2136
rect 3536 1892 3552 2056
rect 3552 1892 3688 2056
rect 3688 1892 3744 2056
rect 3744 1892 3880 2056
rect 3880 1892 3936 2056
rect 3936 1892 4072 2056
rect 4072 1892 4128 2056
rect 4128 1892 4264 2056
rect 4264 1892 4320 2056
rect 4320 1892 4512 2056
rect 6084 2036 6956 2064
rect 6084 1864 6188 2036
rect 6188 1864 6244 2036
rect 6244 1864 6380 2036
rect 6380 1864 6436 2036
rect 6436 1864 6572 2036
rect 6572 1864 6628 2036
rect 6628 1864 6764 2036
rect 6764 1864 6820 2036
rect 6820 1864 6956 2036
rect 2436 1652 2440 1824
rect 2440 1652 2496 1824
rect 2496 1652 2632 1824
rect 2632 1652 2688 1824
rect 2688 1652 2824 1824
rect 2824 1652 2880 1824
rect 2880 1652 3016 1824
rect 3016 1652 3072 1824
rect 3072 1652 3208 1824
rect 3208 1652 3264 1824
rect 3264 1652 3400 1824
rect 3400 1652 3412 1824
rect 2436 1568 3412 1652
rect 4932 1632 4940 1804
rect 4940 1632 4996 1804
rect 4996 1632 5132 1804
rect 5132 1632 5188 1804
rect 5188 1632 5324 1804
rect 5324 1632 5380 1804
rect 5380 1632 5516 1804
rect 5516 1632 5572 1804
rect 5572 1632 5708 1804
rect 5708 1632 5764 1804
rect 5764 1632 5900 1804
rect 5900 1632 5916 1804
rect 4932 1616 5916 1632
rect 3536 1424 4512 1504
rect 3536 1260 3552 1424
rect 3552 1260 3688 1424
rect 3688 1260 3744 1424
rect 3744 1260 3880 1424
rect 3880 1260 3936 1424
rect 3936 1260 4072 1424
rect 4072 1260 4128 1424
rect 4128 1260 4264 1424
rect 4264 1260 4320 1424
rect 4320 1260 4512 1424
rect 6088 1420 6960 1448
rect 6088 1248 6188 1420
rect 6188 1248 6244 1420
rect 6244 1248 6380 1420
rect 6380 1248 6436 1420
rect 6436 1248 6572 1420
rect 6572 1248 6628 1420
rect 6628 1248 6764 1420
rect 6764 1248 6820 1420
rect 6820 1248 6960 1420
rect 2436 1020 2440 1192
rect 2440 1020 2496 1192
rect 2496 1020 2632 1192
rect 2632 1020 2688 1192
rect 2688 1020 2824 1192
rect 2824 1020 2880 1192
rect 2880 1020 3016 1192
rect 3016 1020 3072 1192
rect 3072 1020 3208 1192
rect 3208 1020 3264 1192
rect 3264 1020 3400 1192
rect 3400 1020 3412 1192
rect 2436 932 3412 1020
rect 4936 1016 4940 1184
rect 4940 1016 4996 1184
rect 4996 1016 5132 1184
rect 5132 1016 5188 1184
rect 5188 1016 5324 1184
rect 5324 1016 5380 1184
rect 5380 1016 5516 1184
rect 5516 1016 5572 1184
rect 5572 1016 5708 1184
rect 5708 1016 5764 1184
rect 5764 1016 5900 1184
rect 5900 1016 5920 1184
rect 4936 996 5920 1016
rect 300 448 1760 864
rect 6088 800 6960 832
rect 6088 632 6188 800
rect 6188 632 6244 800
rect 6244 632 6380 800
rect 6380 632 6436 800
rect 6436 632 6572 800
rect 6572 632 6628 800
rect 6628 632 6764 800
rect 6764 632 6820 800
rect 6820 632 6960 800
rect 3548 472 4524 556
rect 3548 308 3552 472
rect 3552 308 3688 472
rect 3688 308 3744 472
rect 3744 308 3880 472
rect 3880 308 3936 472
rect 3936 308 4072 472
rect 4072 308 4128 472
rect 4128 308 4264 472
rect 4264 308 4320 472
rect 4320 308 4524 472
rect 4932 396 4940 568
rect 4940 396 4996 568
rect 4996 396 5132 568
rect 5132 396 5188 568
rect 5188 396 5324 568
rect 5324 396 5380 568
rect 5380 396 5516 568
rect 5516 396 5572 568
rect 5572 396 5708 568
rect 5708 396 5764 568
rect 5764 396 5900 568
rect 5900 396 5916 568
rect 4932 380 5916 396
rect 290 28 1930 130
rect 290 -100 408 28
rect 408 -100 464 28
rect 464 -100 600 28
rect 600 -100 656 28
rect 656 -100 792 28
rect 792 -100 848 28
rect 848 -100 984 28
rect 984 -100 1040 28
rect 1040 -100 1176 28
rect 1176 -100 1232 28
rect 1232 -100 1368 28
rect 1368 -100 1424 28
rect 1424 -100 1560 28
rect 1560 -100 1616 28
rect 1616 -100 1752 28
rect 1752 -100 1808 28
rect 1808 -100 1930 28
rect 2428 68 2440 244
rect 2440 68 2496 244
rect 2496 68 2632 244
rect 2632 68 2688 244
rect 2688 68 2824 244
rect 2824 68 2880 244
rect 2880 68 3016 244
rect 3016 68 3072 244
rect 3072 68 3208 244
rect 3208 68 3264 244
rect 3264 68 3400 244
rect 3400 68 3404 244
rect 2428 -4 3404 68
rect 6088 184 6960 212
rect 6088 12 6188 184
rect 6188 12 6244 184
rect 6244 12 6380 184
rect 6380 12 6436 184
rect 6436 12 6572 184
rect 6572 12 6628 184
rect 6628 12 6764 184
rect 6764 12 6820 184
rect 6820 12 6960 184
rect 290 -588 1930 -490
rect 290 -720 408 -588
rect 408 -720 464 -588
rect 464 -720 600 -588
rect 600 -720 656 -588
rect 656 -720 792 -588
rect 792 -720 848 -588
rect 848 -720 984 -588
rect 984 -720 1040 -588
rect 1040 -720 1176 -588
rect 1176 -720 1232 -588
rect 1232 -720 1368 -588
rect 1368 -720 1424 -588
rect 1424 -720 1560 -588
rect 1560 -720 1616 -588
rect 1616 -720 1752 -588
rect 1752 -720 1808 -588
rect 1808 -720 1930 -588
rect 3548 -148 4524 -64
rect 3548 -312 3552 -148
rect 3552 -312 3688 -148
rect 3688 -312 3744 -148
rect 3744 -312 3880 -148
rect 3880 -312 3936 -148
rect 3936 -312 4072 -148
rect 4072 -312 4128 -148
rect 4128 -312 4264 -148
rect 4264 -312 4320 -148
rect 4320 -312 4524 -148
rect 4928 -220 4940 -48
rect 4940 -220 4996 -48
rect 4996 -220 5132 -48
rect 5132 -220 5188 -48
rect 5188 -220 5324 -48
rect 5324 -220 5380 -48
rect 5380 -220 5516 -48
rect 5516 -220 5572 -48
rect 5572 -220 5708 -48
rect 5708 -220 5764 -48
rect 5764 -220 5900 -48
rect 5900 -220 5912 -48
rect 4928 -236 5912 -220
rect 2428 -552 2440 -380
rect 2440 -552 2496 -380
rect 2496 -552 2632 -380
rect 2632 -552 2688 -380
rect 2688 -552 2824 -380
rect 2824 -552 2880 -380
rect 2880 -552 3016 -380
rect 3016 -552 3072 -380
rect 3072 -552 3208 -380
rect 3208 -552 3264 -380
rect 3264 -552 3400 -380
rect 3400 -552 3404 -380
rect 2428 -628 3404 -552
rect 6088 -436 6960 -408
rect 6088 -608 6188 -436
rect 6188 -608 6244 -436
rect 6244 -608 6380 -436
rect 6380 -608 6436 -436
rect 6436 -608 6572 -436
rect 6572 -608 6628 -436
rect 6628 -608 6764 -436
rect 6764 -608 6820 -436
rect 6820 -608 6960 -436
rect 290 -1208 1930 -1110
rect 290 -1340 408 -1208
rect 408 -1340 464 -1208
rect 464 -1340 600 -1208
rect 600 -1340 656 -1208
rect 656 -1340 792 -1208
rect 792 -1340 848 -1208
rect 848 -1340 984 -1208
rect 984 -1340 1040 -1208
rect 1040 -1340 1176 -1208
rect 1176 -1340 1232 -1208
rect 1232 -1340 1368 -1208
rect 1368 -1340 1424 -1208
rect 1424 -1340 1560 -1208
rect 1560 -1340 1616 -1208
rect 1616 -1340 1752 -1208
rect 1752 -1340 1808 -1208
rect 1808 -1340 1930 -1208
rect 3708 -1228 4400 -716
rect 4932 -840 4940 -672
rect 4940 -840 4996 -672
rect 4996 -840 5132 -672
rect 5132 -840 5188 -672
rect 5188 -840 5324 -672
rect 5324 -840 5380 -672
rect 5380 -840 5516 -672
rect 5516 -840 5572 -672
rect 5572 -840 5708 -672
rect 5708 -840 5764 -672
rect 5764 -840 5900 -672
rect 5900 -840 5916 -672
rect 4932 -860 5916 -840
rect 6088 -1052 6960 -1024
rect 6088 -1224 6188 -1052
rect 6188 -1224 6244 -1052
rect 6244 -1224 6380 -1052
rect 6380 -1224 6436 -1052
rect 6436 -1224 6572 -1052
rect 6572 -1224 6628 -1052
rect 6628 -1224 6764 -1052
rect 6764 -1224 6820 -1052
rect 6820 -1224 6960 -1052
rect 4932 -1456 4940 -1284
rect 4940 -1456 4996 -1284
rect 4996 -1456 5132 -1284
rect 5132 -1456 5188 -1284
rect 5188 -1456 5324 -1284
rect 5324 -1456 5380 -1284
rect 5380 -1456 5516 -1284
rect 5516 -1456 5572 -1284
rect 5572 -1456 5708 -1284
rect 5708 -1456 5764 -1284
rect 5764 -1456 5900 -1284
rect 5900 -1456 5916 -1284
rect 4932 -1472 5916 -1456
rect 6088 -1672 6960 -1640
rect 6088 -1840 6188 -1672
rect 6188 -1840 6244 -1672
rect 6244 -1840 6380 -1672
rect 6380 -1840 6436 -1672
rect 6436 -1840 6572 -1672
rect 6572 -1840 6628 -1672
rect 6628 -1840 6764 -1672
rect 6764 -1840 6820 -1672
rect 6820 -1840 6960 -1672
rect 4928 -2076 4940 -1908
rect 4940 -2076 4996 -1908
rect 4996 -2076 5132 -1908
rect 5132 -2076 5188 -1908
rect 5188 -2076 5324 -1908
rect 5324 -2076 5380 -1908
rect 5380 -2076 5516 -1908
rect 5516 -2076 5572 -1908
rect 5572 -2076 5708 -1908
rect 5708 -2076 5764 -1908
rect 5764 -2076 5900 -1908
rect 5900 -2076 5912 -1908
rect 4928 -2096 5912 -2076
rect -2464 -2756 -2460 -2584
rect -2460 -2756 -2408 -2584
rect -2408 -2756 -2268 -2584
rect -2268 -2756 -2216 -2584
rect -2216 -2756 -2076 -2584
rect -2076 -2756 -2024 -2584
rect -2024 -2756 -1884 -2584
rect -1884 -2756 -1860 -2584
rect -2464 -2768 -1860 -2756
rect -664 -2756 -660 -2584
rect -660 -2756 -608 -2584
rect -608 -2756 -468 -2584
rect -468 -2756 -416 -2584
rect -416 -2756 -276 -2584
rect -276 -2756 -224 -2584
rect -224 -2756 -84 -2584
rect -84 -2756 -60 -2584
rect -664 -2768 -60 -2756
rect -2464 -3372 -2460 -3200
rect -2460 -3372 -2408 -3200
rect -2408 -3372 -2268 -3200
rect -2268 -3372 -2216 -3200
rect -2216 -3372 -2076 -3200
rect -2076 -3372 -2024 -3200
rect -2024 -3372 -1884 -3200
rect -1884 -3372 -1860 -3200
rect -2464 -3384 -1860 -3372
rect -3484 -3824 -3080 -3412
rect -3080 -3824 -2708 -3412
rect 1136 -2756 1140 -2584
rect 1140 -2756 1192 -2584
rect 1192 -2756 1332 -2584
rect 1332 -2756 1384 -2584
rect 1384 -2756 1524 -2584
rect 1524 -2756 1576 -2584
rect 1576 -2756 1716 -2584
rect 1716 -2756 1740 -2584
rect 1136 -2768 1740 -2756
rect -664 -3372 -660 -3200
rect -660 -3372 -608 -3200
rect -608 -3372 -468 -3200
rect -468 -3372 -416 -3200
rect -416 -3372 -276 -3200
rect -276 -3372 -224 -3200
rect -224 -3372 -84 -3200
rect -84 -3372 -60 -3200
rect -664 -3384 -60 -3372
rect 2936 -2756 2940 -2584
rect 2940 -2756 2992 -2584
rect 2992 -2756 3132 -2584
rect 3132 -2756 3184 -2584
rect 3184 -2756 3324 -2584
rect 3324 -2756 3376 -2584
rect 3376 -2756 3516 -2584
rect 3516 -2756 3540 -2584
rect 2936 -2768 3540 -2756
rect 1136 -3372 1140 -3200
rect 1140 -3372 1192 -3200
rect 1192 -3372 1332 -3200
rect 1332 -3372 1384 -3200
rect 1384 -3372 1524 -3200
rect 1524 -3372 1576 -3200
rect 1576 -3372 1716 -3200
rect 1716 -3372 1740 -3200
rect 1136 -3384 1740 -3372
rect 6084 -2288 6956 -2260
rect 6084 -2460 6188 -2288
rect 6188 -2460 6244 -2288
rect 6244 -2460 6380 -2288
rect 6380 -2460 6436 -2288
rect 6436 -2460 6572 -2288
rect 6572 -2460 6628 -2288
rect 6628 -2460 6764 -2288
rect 6764 -2460 6820 -2288
rect 6820 -2460 6956 -2288
rect 4928 -2692 4940 -2520
rect 4940 -2692 4996 -2520
rect 4996 -2692 5132 -2520
rect 5132 -2692 5188 -2520
rect 5188 -2692 5324 -2520
rect 5324 -2692 5380 -2520
rect 5380 -2692 5516 -2520
rect 5516 -2692 5572 -2520
rect 5572 -2692 5708 -2520
rect 5708 -2692 5764 -2520
rect 5764 -2692 5900 -2520
rect 5900 -2692 5912 -2520
rect 4928 -2708 5912 -2692
rect 6084 -2908 6956 -2880
rect 6084 -3080 6188 -2908
rect 6188 -3080 6244 -2908
rect 6244 -3080 6380 -2908
rect 6380 -3080 6436 -2908
rect 6436 -3080 6572 -2908
rect 6572 -3080 6628 -2908
rect 6628 -3080 6764 -2908
rect 6764 -3080 6820 -2908
rect 6820 -3080 6956 -2908
rect 2936 -3372 2940 -3200
rect 2940 -3372 2992 -3200
rect 2992 -3372 3132 -3200
rect 3132 -3372 3184 -3200
rect 3184 -3372 3324 -3200
rect 3324 -3372 3376 -3200
rect 3376 -3372 3516 -3200
rect 3516 -3372 3540 -3200
rect 2936 -3384 3540 -3372
rect 4928 -3312 4940 -3144
rect 4940 -3312 4996 -3144
rect 4996 -3312 5132 -3144
rect 5132 -3312 5188 -3144
rect 5188 -3312 5324 -3144
rect 5324 -3312 5380 -3144
rect 5380 -3312 5516 -3144
rect 5516 -3312 5572 -3144
rect 5572 -3312 5708 -3144
rect 5708 -3312 5764 -3144
rect 5764 -3312 5900 -3144
rect 5900 -3312 5912 -3144
rect 4928 -3332 5912 -3312
rect -2468 -3992 -2460 -3820
rect -2460 -3992 -2408 -3820
rect -2408 -3992 -2268 -3820
rect -2268 -3992 -2216 -3820
rect -2216 -3992 -2076 -3820
rect -2076 -3992 -2024 -3820
rect -2024 -3992 -1884 -3820
rect -1884 -3992 -1864 -3820
rect -2468 -4004 -1864 -3992
rect -668 -3992 -660 -3820
rect -660 -3992 -608 -3820
rect -608 -3992 -468 -3820
rect -468 -3992 -416 -3820
rect -416 -3992 -276 -3820
rect -276 -3992 -224 -3820
rect -224 -3992 -84 -3820
rect -84 -3992 -64 -3820
rect -668 -4004 -64 -3992
rect 1132 -3992 1140 -3820
rect 1140 -3992 1192 -3820
rect 1192 -3992 1332 -3820
rect 1332 -3992 1384 -3820
rect 1384 -3992 1524 -3820
rect 1524 -3992 1576 -3820
rect 1576 -3992 1716 -3820
rect 1716 -3992 1736 -3820
rect 1132 -4004 1736 -3992
rect 2932 -3992 2940 -3820
rect 2940 -3992 2992 -3820
rect 2992 -3992 3132 -3820
rect 3132 -3992 3184 -3820
rect 3184 -3992 3324 -3820
rect 3324 -3992 3376 -3820
rect 3376 -3992 3516 -3820
rect 3516 -3992 3536 -3820
rect 2932 -4004 3536 -3992
rect -2460 -4500 -1860 -4488
rect -660 -4500 -60 -4488
rect 1140 -4500 1740 -4488
rect 2940 -4500 3540 -4488
rect -2460 -4672 -2408 -4500
rect -2408 -4672 -1944 -4500
rect -1944 -4672 -1892 -4500
rect -1892 -4672 -1860 -4500
rect -660 -4672 -608 -4500
rect -608 -4672 -144 -4500
rect -144 -4672 -92 -4500
rect -92 -4672 -60 -4500
rect 1140 -4672 1192 -4500
rect 1192 -4672 1656 -4500
rect 1656 -4672 1708 -4500
rect 1708 -4672 1740 -4500
rect 2940 -4672 2992 -4500
rect 2992 -4672 3456 -4500
rect 3456 -4672 3508 -4500
rect 3508 -4672 3540 -4500
rect -1716 -4900 -1684 -4728
rect -1684 -4900 -1632 -4728
rect -1632 -4900 -1168 -4728
rect -1168 -4900 -1116 -4728
rect -1716 -4912 -1116 -4900
rect 84 -4900 116 -4728
rect 116 -4900 168 -4728
rect 168 -4900 632 -4728
rect 632 -4900 684 -4728
rect 84 -4912 684 -4900
rect 1884 -4900 1916 -4728
rect 1916 -4900 1968 -4728
rect 1968 -4900 2432 -4728
rect 2432 -4900 2484 -4728
rect 1884 -4912 2484 -4900
rect 3684 -4900 3716 -4728
rect 3716 -4900 3768 -4728
rect 3768 -4900 4232 -4728
rect 4232 -4900 4284 -4728
rect 3684 -4912 4284 -4900
rect -2460 -5116 -1860 -5104
rect -2460 -5288 -2408 -5116
rect -2408 -5288 -1944 -5116
rect -1944 -5288 -1892 -5116
rect -1892 -5288 -1860 -5116
rect -660 -5116 -60 -5104
rect -660 -5288 -608 -5116
rect -608 -5288 -144 -5116
rect -144 -5288 -92 -5116
rect -92 -5288 -60 -5116
rect 1140 -5116 1740 -5104
rect 1140 -5288 1192 -5116
rect 1192 -5288 1656 -5116
rect 1656 -5288 1708 -5116
rect 1708 -5288 1740 -5116
rect 2940 -5116 3540 -5104
rect 2940 -5288 2992 -5116
rect 2992 -5288 3456 -5116
rect 3456 -5288 3508 -5116
rect 3508 -5288 3540 -5116
rect -1716 -5516 -1684 -5344
rect -1684 -5516 -1632 -5344
rect -1632 -5516 -1168 -5344
rect -1168 -5516 -1116 -5344
rect -1716 -5528 -1116 -5516
rect 84 -5516 116 -5344
rect 116 -5516 168 -5344
rect 168 -5516 632 -5344
rect 632 -5516 684 -5344
rect 84 -5528 684 -5516
rect 1884 -5516 1916 -5344
rect 1916 -5516 1968 -5344
rect 1968 -5516 2432 -5344
rect 2432 -5516 2484 -5344
rect 1884 -5528 2484 -5516
rect 3684 -5516 3716 -5344
rect 3716 -5516 3768 -5344
rect 3768 -5516 4232 -5344
rect 4232 -5516 4284 -5344
rect 3684 -5528 4284 -5516
rect -2460 -5736 -1860 -5724
rect -2460 -5908 -2408 -5736
rect -2408 -5908 -1944 -5736
rect -1944 -5908 -1892 -5736
rect -1892 -5908 -1860 -5736
rect -660 -5736 -60 -5724
rect -660 -5908 -608 -5736
rect -608 -5908 -144 -5736
rect -144 -5908 -92 -5736
rect -92 -5908 -60 -5736
rect 1140 -5736 1740 -5724
rect 1140 -5908 1192 -5736
rect 1192 -5908 1656 -5736
rect 1656 -5908 1708 -5736
rect 1708 -5908 1740 -5736
rect 2940 -5736 3540 -5724
rect 2940 -5908 2992 -5736
rect 2992 -5908 3456 -5736
rect 3456 -5908 3508 -5736
rect 3508 -5908 3540 -5736
rect -1716 -6136 -1684 -5964
rect -1684 -6136 -1632 -5964
rect -1632 -6136 -1168 -5964
rect -1168 -6136 -1116 -5964
rect -1716 -6148 -1116 -6136
rect 84 -6136 116 -5964
rect 116 -6136 168 -5964
rect 168 -6136 632 -5964
rect 632 -6136 684 -5964
rect 84 -6148 684 -6136
rect 1884 -6136 1916 -5964
rect 1916 -6136 1968 -5964
rect 1968 -6136 2432 -5964
rect 2432 -6136 2484 -5964
rect 1884 -6148 2484 -6136
rect 3684 -6136 3716 -5964
rect 3716 -6136 3768 -5964
rect 3768 -6136 4232 -5964
rect 4232 -6136 4284 -5964
rect 3684 -6148 4284 -6136
rect -2460 -6352 -1860 -6340
rect -2460 -6524 -2408 -6352
rect -2408 -6524 -1944 -6352
rect -1944 -6524 -1892 -6352
rect -1892 -6524 -1860 -6352
rect -660 -6352 -60 -6340
rect -660 -6524 -608 -6352
rect -608 -6524 -144 -6352
rect -144 -6524 -92 -6352
rect -92 -6524 -60 -6352
rect 1140 -6352 1740 -6340
rect 1140 -6524 1192 -6352
rect 1192 -6524 1656 -6352
rect 1656 -6524 1708 -6352
rect 1708 -6524 1740 -6352
rect 2940 -6352 3540 -6340
rect 2940 -6524 2992 -6352
rect 2992 -6524 3456 -6352
rect 3456 -6524 3508 -6352
rect 3508 -6524 3540 -6352
rect -1716 -6752 -1684 -6580
rect -1684 -6752 -1632 -6580
rect -1632 -6752 -1168 -6580
rect -1168 -6752 -1116 -6580
rect -1716 -6764 -1116 -6752
rect 84 -6752 116 -6580
rect 116 -6752 168 -6580
rect 168 -6752 632 -6580
rect 632 -6752 684 -6580
rect 84 -6764 684 -6752
rect 1884 -6752 1916 -6580
rect 1916 -6752 1968 -6580
rect 1968 -6752 2432 -6580
rect 2432 -6752 2484 -6580
rect 1884 -6764 2484 -6752
rect 3684 -6752 3716 -6580
rect 3716 -6752 3768 -6580
rect 3768 -6752 4232 -6580
rect 4232 -6752 4284 -6580
rect 3684 -6764 4284 -6752
rect -2460 -6972 -1860 -6960
rect -2460 -7144 -2408 -6972
rect -2408 -7144 -1944 -6972
rect -1944 -7144 -1892 -6972
rect -1892 -7144 -1860 -6972
rect -660 -6972 -60 -6960
rect -660 -7144 -608 -6972
rect -608 -7144 -144 -6972
rect -144 -7144 -92 -6972
rect -92 -7144 -60 -6972
rect 1140 -6972 1740 -6960
rect 1140 -7144 1192 -6972
rect 1192 -7144 1656 -6972
rect 1656 -7144 1708 -6972
rect 1708 -7144 1740 -6972
rect 2940 -6972 3540 -6960
rect 2940 -7144 2992 -6972
rect 2992 -7144 3456 -6972
rect 3456 -7144 3508 -6972
rect 3508 -7144 3540 -6972
rect -1716 -7372 -1684 -7200
rect -1684 -7372 -1632 -7200
rect -1632 -7372 -1168 -7200
rect -1168 -7372 -1116 -7200
rect -1716 -7384 -1116 -7372
rect 84 -7372 116 -7200
rect 116 -7372 168 -7200
rect 168 -7372 632 -7200
rect 632 -7372 684 -7200
rect 84 -7384 684 -7372
rect 1884 -7372 1916 -7200
rect 1916 -7372 1968 -7200
rect 1968 -7372 2432 -7200
rect 2432 -7372 2484 -7200
rect 1884 -7384 2484 -7372
rect 3684 -7372 3716 -7200
rect 3716 -7372 3768 -7200
rect 3768 -7372 4232 -7200
rect 4232 -7372 4284 -7200
rect 3684 -7384 4284 -7372
rect -2460 -7588 -1860 -7576
rect -2460 -7760 -2408 -7588
rect -2408 -7760 -1944 -7588
rect -1944 -7760 -1892 -7588
rect -1892 -7760 -1860 -7588
rect -660 -7588 -60 -7576
rect -660 -7760 -608 -7588
rect -608 -7760 -144 -7588
rect -144 -7760 -92 -7588
rect -92 -7760 -60 -7588
rect 1140 -7588 1740 -7576
rect 1140 -7760 1192 -7588
rect 1192 -7760 1656 -7588
rect 1656 -7760 1708 -7588
rect 1708 -7760 1740 -7588
rect 2940 -7588 3540 -7576
rect 2940 -7760 2992 -7588
rect 2992 -7760 3456 -7588
rect 3456 -7760 3508 -7588
rect 3508 -7760 3540 -7588
rect -1716 -7988 -1684 -7816
rect -1684 -7988 -1632 -7816
rect -1632 -7988 -1168 -7816
rect -1168 -7988 -1116 -7816
rect -1716 -8000 -1116 -7988
rect -980 -8160 -800 -7960
rect 84 -7988 116 -7816
rect 116 -7988 168 -7816
rect 168 -7988 632 -7816
rect 632 -7988 684 -7816
rect 84 -8000 684 -7988
rect 1884 -7988 1916 -7816
rect 1916 -7988 1968 -7816
rect 1968 -7988 2432 -7816
rect 2432 -7988 2484 -7816
rect 1884 -8000 2484 -7988
rect 3684 -7988 3716 -7816
rect 3716 -7988 3768 -7816
rect 3768 -7988 4232 -7816
rect 4232 -7988 4284 -7816
rect 3684 -8000 4284 -7988
rect -5444 -9416 -4636 -8610
<< metal3 >>
rect -4448 2580 4644 3244
rect -4448 2496 3420 2580
rect -4536 2476 3420 2496
rect -4536 2412 -4508 2476
rect -484 2412 3420 2476
rect -4536 2380 3420 2412
rect 3600 2380 4644 2580
rect -4536 2136 4644 2380
rect -4536 2112 3536 2136
rect -4536 1932 -80 2112
rect -4536 -1876 -456 1932
rect -90 1676 -80 1932
rect 2096 1932 3536 2112
rect 2096 1676 2106 1932
rect 3526 1892 3536 1932
rect 4512 1932 4644 2136
rect 6074 2064 6966 2069
rect 4512 1892 4552 1932
rect 3526 1887 4552 1892
rect 2426 1828 3422 1829
rect -90 1671 2106 1676
rect 2416 1824 3422 1828
rect -80 1668 2096 1671
rect 2416 1568 2436 1824
rect 3412 1568 3422 1824
rect 2416 1563 3422 1568
rect 2416 1197 3412 1563
rect 3536 1509 4552 1887
rect 6074 1864 6084 2064
rect 6956 1864 6966 2064
rect 6074 1859 6966 1864
rect 4924 1809 5924 1812
rect 4922 1804 5926 1809
rect 4922 1616 4932 1804
rect 5916 1616 5926 1804
rect 4922 1611 5926 1616
rect 3526 1504 4552 1509
rect 3526 1260 3536 1504
rect 4512 1260 4552 1504
rect 3526 1255 4552 1260
rect 3536 1248 4552 1255
rect 2416 1192 3422 1197
rect 2416 932 2436 1192
rect 3412 932 3422 1192
rect 2416 927 3422 932
rect 4924 1189 5924 1611
rect 6084 1453 6960 1859
rect 6078 1448 6970 1453
rect 6078 1248 6088 1448
rect 6960 1248 6970 1448
rect 6078 1243 6970 1248
rect 4924 1184 5930 1189
rect 4924 996 4936 1184
rect 5920 996 5930 1184
rect 4924 991 5930 996
rect 292 869 1768 872
rect 290 864 1770 869
rect 290 448 300 864
rect 1760 448 1770 864
rect 290 443 1770 448
rect 292 280 1768 443
rect 290 135 1770 280
rect 2416 249 3412 927
rect 4924 573 5924 991
rect 6084 837 6960 1243
rect 6078 832 6970 837
rect 6078 632 6088 832
rect 6960 632 6970 832
rect 6078 627 6970 632
rect 4922 568 5926 573
rect 3538 556 4534 561
rect 3538 308 3548 556
rect 4524 492 4534 556
rect 4922 492 4932 568
rect 4524 380 4932 492
rect 5916 380 5926 568
rect 4524 375 5926 380
rect 4524 308 5924 375
rect 3538 303 5924 308
rect 2416 244 3414 249
rect 280 130 1940 135
rect 280 -100 290 130
rect 1930 -100 1940 130
rect 280 -105 1940 -100
rect 2416 -4 2428 244
rect 3404 -4 3414 244
rect 2416 -9 3414 -4
rect 290 -485 1770 -105
rect 2416 -375 3412 -9
rect 3548 -48 5924 303
rect 6084 217 6960 627
rect 6078 212 6970 217
rect 6078 12 6088 212
rect 6960 12 6970 212
rect 6078 7 6970 12
rect 3548 -59 4928 -48
rect 3538 -64 4928 -59
rect 3538 -312 3548 -64
rect 4524 -236 4928 -64
rect 5912 -236 5924 -48
rect 4524 -312 5924 -236
rect 3538 -317 5924 -312
rect 3548 -324 5924 -317
rect 2416 -380 3414 -375
rect 280 -490 1940 -485
rect 280 -720 290 -490
rect 1930 -720 1940 -490
rect 2416 -572 2428 -380
rect 2418 -628 2428 -572
rect 3404 -628 3414 -380
rect 2418 -633 3414 -628
rect 4924 -667 5924 -324
rect 6084 -403 6960 7
rect 6078 -408 6970 -403
rect 6078 -608 6088 -408
rect 6960 -608 6970 -408
rect 6078 -613 6970 -608
rect 4922 -672 5926 -667
rect 3708 -711 4716 -676
rect 280 -725 1940 -720
rect 3698 -716 4716 -711
rect 290 -1105 1770 -725
rect 280 -1110 1940 -1105
rect 280 -1340 290 -1110
rect 1930 -1340 1940 -1110
rect 3698 -1228 3708 -716
rect 4400 -1228 4716 -716
rect 4922 -860 4932 -672
rect 5916 -860 5926 -672
rect 4922 -865 5926 -860
rect 3698 -1233 4716 -1228
rect 280 -1345 1940 -1340
rect 290 -1390 1770 -1345
rect -2464 -2579 -1860 -2576
rect -664 -2579 -60 -2576
rect 1136 -2579 1740 -2576
rect 2936 -2579 3540 -2576
rect -2474 -2584 -1850 -2579
rect -2474 -2768 -2464 -2584
rect -1860 -2768 -1850 -2584
rect -2474 -2773 -1850 -2768
rect -674 -2584 -50 -2579
rect -674 -2768 -664 -2584
rect -60 -2768 -50 -2584
rect -674 -2773 -50 -2768
rect 1126 -2584 1750 -2579
rect 1126 -2768 1136 -2584
rect 1740 -2768 1750 -2584
rect 1126 -2773 1750 -2768
rect 2926 -2584 3550 -2579
rect 2926 -2768 2936 -2584
rect 3540 -2768 3550 -2584
rect 2926 -2773 3550 -2768
rect -2464 -3195 -1860 -2773
rect -664 -3195 -60 -2773
rect 1136 -3195 1740 -2773
rect 2936 -3195 3540 -2773
rect -2474 -3200 -1850 -3195
rect -2474 -3384 -2464 -3200
rect -1860 -3384 -1850 -3200
rect -2474 -3389 -1850 -3384
rect -674 -3200 -50 -3195
rect -674 -3384 -664 -3200
rect -60 -3384 -50 -3200
rect -674 -3389 -50 -3384
rect 1126 -3200 1750 -3195
rect 1126 -3384 1136 -3200
rect 1740 -3384 1750 -3200
rect 1126 -3389 1750 -3384
rect 2926 -3200 3550 -3195
rect 2926 -3384 2936 -3200
rect 3540 -3384 3550 -3200
rect 2926 -3389 3550 -3384
rect -3494 -3412 -2698 -3407
rect -3494 -3824 -3484 -3412
rect -2708 -3824 -2698 -3412
rect -2464 -3815 -1860 -3389
rect -664 -3815 -60 -3389
rect 1136 -3815 1740 -3389
rect 2936 -3815 3540 -3389
rect 3708 -3772 4716 -1233
rect 4924 -1279 5924 -865
rect 6084 -1019 6960 -613
rect 6078 -1024 6970 -1019
rect 6078 -1224 6088 -1024
rect 6960 -1224 6970 -1024
rect 6078 -1229 6970 -1224
rect 4922 -1284 5926 -1279
rect 4922 -1472 4932 -1284
rect 5916 -1472 5926 -1284
rect 4922 -1477 5926 -1472
rect 4924 -1903 5924 -1477
rect 6084 -1635 6960 -1229
rect 6078 -1640 6970 -1635
rect 6078 -1840 6088 -1640
rect 6960 -1840 6970 -1640
rect 6078 -1845 6970 -1840
rect 4918 -1908 5924 -1903
rect 4918 -2096 4928 -1908
rect 5912 -2096 5924 -1908
rect 4918 -2101 5924 -2096
rect 4924 -2515 5924 -2101
rect 6084 -2208 6960 -1845
rect 6084 -2255 6096 -2208
rect 6074 -2260 6096 -2255
rect 6940 -2255 6960 -2208
rect 6940 -2260 6966 -2255
rect 6074 -2460 6084 -2260
rect 6956 -2460 6966 -2260
rect 6074 -2465 6096 -2460
rect 4918 -2520 5924 -2515
rect 4918 -2708 4928 -2520
rect 5912 -2708 5924 -2520
rect 4918 -2713 5924 -2708
rect 4924 -3139 5924 -2713
rect 6084 -2875 6096 -2465
rect 6074 -2880 6096 -2875
rect 6940 -2465 6966 -2460
rect 6940 -2875 6960 -2465
rect 6940 -2880 6966 -2875
rect 6074 -3080 6084 -2880
rect 6956 -3080 6966 -2880
rect 6074 -3085 6966 -3080
rect 6084 -3088 6960 -3085
rect 4918 -3144 5924 -3139
rect 4918 -3332 4928 -3144
rect 5912 -3324 5924 -3144
rect 5912 -3332 5922 -3324
rect 4918 -3337 5922 -3332
rect -3494 -3829 -2698 -3824
rect -2478 -3820 -1854 -3815
rect -3480 -4100 -2704 -3829
rect -2478 -4004 -2468 -3820
rect -1864 -4004 -1854 -3820
rect -2478 -4009 -1854 -4004
rect -678 -3820 -54 -3815
rect -678 -4004 -668 -3820
rect -64 -4004 -54 -3820
rect -678 -4009 -54 -4004
rect 1122 -3820 1746 -3815
rect 1122 -4004 1132 -3820
rect 1736 -4004 1746 -3820
rect 1122 -4009 1746 -4004
rect 2922 -3820 3546 -3815
rect 2922 -4004 2932 -3820
rect 3536 -4004 3546 -3820
rect 2922 -4009 3546 -4004
rect -6076 -4128 -2704 -4100
rect -6076 -8152 -2788 -4128
rect -2724 -8152 -2704 -4128
rect -2464 -4483 -1860 -4009
rect -664 -4483 -60 -4009
rect 1136 -4483 1740 -4009
rect 2936 -4483 3540 -4009
rect 3708 -4120 4720 -3772
rect 3708 -4148 7876 -4120
rect 3708 -4176 7792 -4148
rect -2470 -4488 -1850 -4483
rect -2470 -4672 -2460 -4488
rect -1860 -4672 -1850 -4488
rect -2470 -4677 -1850 -4672
rect -670 -4488 -50 -4483
rect -670 -4672 -660 -4488
rect -60 -4672 -50 -4488
rect -670 -4677 -50 -4672
rect 1130 -4488 1750 -4483
rect 1130 -4672 1140 -4488
rect 1740 -4672 1750 -4488
rect 1130 -4677 1750 -4672
rect 2930 -4488 3550 -4483
rect 3712 -4488 7792 -4176
rect 2930 -4672 2940 -4488
rect 3540 -4672 3550 -4488
rect 2930 -4677 3550 -4672
rect -2464 -5099 -1860 -4677
rect -1726 -4728 -1106 -4723
rect -1726 -4912 -1716 -4728
rect -1116 -4912 -1106 -4728
rect -1726 -4917 -1106 -4912
rect -2470 -5104 -1850 -5099
rect -2470 -5288 -2460 -5104
rect -1860 -5288 -1850 -5104
rect -2470 -5293 -1850 -5288
rect -2464 -5719 -1860 -5293
rect -1716 -5339 -1116 -4917
rect -664 -5099 -60 -4677
rect 74 -4728 694 -4723
rect 74 -4912 84 -4728
rect 684 -4912 694 -4728
rect 74 -4917 694 -4912
rect -670 -5104 -50 -5099
rect -670 -5288 -660 -5104
rect -60 -5288 -50 -5104
rect -670 -5293 -50 -5288
rect -1726 -5344 -1106 -5339
rect -1726 -5528 -1716 -5344
rect -1116 -5528 -1106 -5344
rect -1726 -5533 -1106 -5528
rect -2470 -5724 -1850 -5719
rect -2470 -5908 -2460 -5724
rect -1860 -5908 -1850 -5724
rect -2470 -5913 -1850 -5908
rect -2464 -6335 -1860 -5913
rect -1716 -5959 -1116 -5533
rect -664 -5719 -60 -5293
rect 84 -5339 684 -4917
rect 1136 -5099 1740 -4677
rect 1874 -4728 2494 -4723
rect 1874 -4912 1884 -4728
rect 2484 -4912 2494 -4728
rect 1874 -4917 2494 -4912
rect 1130 -5104 1750 -5099
rect 1130 -5288 1140 -5104
rect 1740 -5288 1750 -5104
rect 1130 -5293 1750 -5288
rect 74 -5344 694 -5339
rect 74 -5528 84 -5344
rect 684 -5528 694 -5344
rect 74 -5533 694 -5528
rect -670 -5724 -50 -5719
rect -670 -5908 -660 -5724
rect -60 -5908 -50 -5724
rect -670 -5913 -50 -5908
rect -1726 -5964 -1106 -5959
rect -1726 -6148 -1716 -5964
rect -1116 -6148 -1106 -5964
rect -1726 -6153 -1106 -6148
rect -2470 -6340 -1850 -6335
rect -2470 -6524 -2460 -6340
rect -1860 -6524 -1850 -6340
rect -2470 -6529 -1850 -6524
rect -2464 -6955 -1860 -6529
rect -1716 -6575 -1116 -6153
rect -664 -6335 -60 -5913
rect 84 -5959 684 -5533
rect 1136 -5719 1740 -5293
rect 1884 -5339 2484 -4917
rect 2936 -5099 3540 -4677
rect 3674 -4728 4294 -4723
rect 3674 -4912 3684 -4728
rect 4284 -4912 4294 -4728
rect 3674 -4917 4294 -4912
rect 2930 -5104 3550 -5099
rect 2930 -5288 2940 -5104
rect 3540 -5288 3550 -5104
rect 2930 -5293 3550 -5288
rect 1874 -5344 2494 -5339
rect 1874 -5528 1884 -5344
rect 2484 -5528 2494 -5344
rect 1874 -5533 2494 -5528
rect 1130 -5724 1750 -5719
rect 1130 -5908 1140 -5724
rect 1740 -5908 1750 -5724
rect 1130 -5913 1750 -5908
rect 74 -5964 694 -5959
rect 74 -6148 84 -5964
rect 684 -6148 694 -5964
rect 74 -6153 694 -6148
rect -670 -6340 -50 -6335
rect -670 -6524 -660 -6340
rect -60 -6524 -50 -6340
rect -670 -6529 -50 -6524
rect -1726 -6580 -1106 -6575
rect -1726 -6764 -1716 -6580
rect -1116 -6764 -1106 -6580
rect -1726 -6769 -1106 -6764
rect -2470 -6960 -1850 -6955
rect -2470 -7144 -2460 -6960
rect -1860 -7144 -1850 -6960
rect -2470 -7149 -1850 -7144
rect -2464 -7571 -1860 -7149
rect -1716 -7195 -1116 -6769
rect -664 -6955 -60 -6529
rect 84 -6575 684 -6153
rect 1136 -6335 1740 -5913
rect 1884 -5959 2484 -5533
rect 2936 -5719 3540 -5293
rect 3684 -5339 4284 -4917
rect 3674 -5344 4294 -5339
rect 3674 -5528 3684 -5344
rect 4284 -5528 4294 -5344
rect 3674 -5533 4294 -5528
rect 2930 -5724 3550 -5719
rect 2930 -5908 2940 -5724
rect 3540 -5908 3550 -5724
rect 2930 -5913 3550 -5908
rect 1874 -5964 2494 -5959
rect 1874 -6148 1884 -5964
rect 2484 -6148 2494 -5964
rect 1874 -6153 2494 -6148
rect 1130 -6340 1750 -6335
rect 1130 -6524 1140 -6340
rect 1740 -6524 1750 -6340
rect 1130 -6529 1750 -6524
rect 74 -6580 694 -6575
rect 74 -6764 84 -6580
rect 684 -6764 694 -6580
rect 74 -6769 694 -6764
rect -670 -6960 -50 -6955
rect -670 -7144 -660 -6960
rect -60 -7144 -50 -6960
rect -670 -7149 -50 -7144
rect -1726 -7200 -1106 -7195
rect -1726 -7384 -1716 -7200
rect -1116 -7384 -1106 -7200
rect -1726 -7389 -1106 -7384
rect -1716 -7548 -1116 -7389
rect -2470 -7576 -1850 -7571
rect -2470 -7760 -2460 -7576
rect -1860 -7760 -1850 -7576
rect -2470 -7765 -1850 -7760
rect -2464 -7784 -1860 -7765
rect -1716 -7811 -1700 -7548
rect -1726 -7816 -1700 -7811
rect -1128 -7811 -1116 -7548
rect -664 -7571 -60 -7149
rect 84 -7195 684 -6769
rect 1136 -6955 1740 -6529
rect 1884 -6575 2484 -6153
rect 2936 -6335 3540 -5913
rect 3684 -5959 4284 -5533
rect 3674 -5964 4294 -5959
rect 3674 -6148 3684 -5964
rect 4284 -6148 4294 -5964
rect 3674 -6153 4294 -6148
rect 2930 -6340 3550 -6335
rect 2930 -6524 2940 -6340
rect 3540 -6524 3550 -6340
rect 2930 -6529 3550 -6524
rect 1874 -6580 2494 -6575
rect 1874 -6764 1884 -6580
rect 2484 -6764 2494 -6580
rect 1874 -6769 2494 -6764
rect 1130 -6960 1750 -6955
rect 1130 -7144 1140 -6960
rect 1740 -7144 1750 -6960
rect 1130 -7149 1750 -7144
rect 74 -7200 694 -7195
rect 74 -7384 84 -7200
rect 684 -7384 694 -7200
rect 74 -7389 694 -7384
rect 84 -7548 684 -7389
rect -670 -7576 -50 -7571
rect -670 -7760 -660 -7576
rect -60 -7760 -50 -7576
rect -670 -7765 -50 -7760
rect -664 -7784 -60 -7765
rect 84 -7811 100 -7548
rect -1128 -7816 -1106 -7811
rect -1726 -8000 -1716 -7816
rect -1116 -8000 -1106 -7816
rect 74 -7816 100 -7811
rect 672 -7811 684 -7548
rect 1136 -7571 1740 -7149
rect 1884 -7195 2484 -6769
rect 2936 -6955 3540 -6529
rect 3684 -6575 4284 -6153
rect 3674 -6580 4294 -6575
rect 3674 -6764 3684 -6580
rect 4284 -6764 4294 -6580
rect 3674 -6769 4294 -6764
rect 2930 -6960 3550 -6955
rect 2930 -7144 2940 -6960
rect 3540 -7144 3550 -6960
rect 2930 -7149 3550 -7144
rect 1874 -7200 2494 -7195
rect 1874 -7384 1884 -7200
rect 2484 -7384 2494 -7200
rect 1874 -7389 2494 -7384
rect 1884 -7552 2484 -7389
rect 1130 -7576 1750 -7571
rect 1130 -7760 1140 -7576
rect 1740 -7760 1750 -7576
rect 1130 -7765 1750 -7760
rect 1136 -7784 1740 -7765
rect 1884 -7811 1896 -7552
rect 672 -7816 694 -7811
rect -1726 -8005 -1106 -8000
rect -990 -7960 -790 -7955
rect -6076 -8180 -2704 -8152
rect -990 -8160 -980 -7960
rect -800 -8160 -790 -7960
rect 74 -8000 84 -7816
rect 684 -8000 694 -7816
rect 74 -8005 694 -8000
rect 1874 -7816 1896 -7811
rect 2468 -7811 2484 -7552
rect 2936 -7571 3540 -7149
rect 3684 -7195 4284 -6769
rect 3674 -7200 4294 -7195
rect 3674 -7384 3684 -7200
rect 4284 -7384 4294 -7200
rect 3674 -7389 4294 -7384
rect 3684 -7552 4284 -7389
rect 2930 -7576 3550 -7571
rect 2930 -7760 2940 -7576
rect 3540 -7760 3550 -7576
rect 2930 -7765 3550 -7760
rect 2936 -7784 3540 -7765
rect 3684 -7811 3696 -7552
rect 2468 -7816 2494 -7811
rect 1874 -8000 1884 -7816
rect 2484 -8000 2494 -7816
rect 1874 -8005 2494 -8000
rect 3674 -7816 3696 -7811
rect 4268 -7811 4284 -7552
rect 4268 -7816 4294 -7811
rect 3674 -8000 3684 -7816
rect 4284 -8000 4294 -7816
rect 3674 -8005 4294 -8000
rect -990 -8165 -790 -8160
rect 4504 -8172 7792 -4488
rect 7856 -8172 7876 -4148
rect 4504 -8200 7876 -8172
rect -5454 -8610 -4626 -8605
rect -5454 -9416 -5444 -8610
rect -4636 -9416 -4626 -8610
rect -5454 -9421 -4626 -9416
<< via3 >>
rect -4508 2412 -484 2476
rect 6096 -2260 6940 -2208
rect 6096 -2460 6940 -2260
rect 6096 -2880 6940 -2460
rect 6096 -3068 6940 -2880
rect -2788 -8152 -2724 -4128
rect -1700 -7816 -1128 -7548
rect -1700 -7988 -1128 -7816
rect 100 -7816 672 -7548
rect -980 -8160 -800 -7960
rect 100 -7988 672 -7816
rect 1896 -7816 2468 -7552
rect 1896 -7992 2468 -7816
rect 3696 -7816 4268 -7552
rect 3696 -7992 4268 -7816
rect 7792 -8172 7856 -4148
rect -5444 -9416 -4636 -8610
<< mimcap >>
rect -4496 2124 -496 2164
rect -4496 -1796 -4456 2124
rect -536 -1796 -496 2124
rect -4496 -1836 -496 -1796
rect -6036 -4180 -3036 -4140
rect -6036 -8100 -5996 -4180
rect -3076 -8100 -3036 -4180
rect -6036 -8140 -3036 -8100
rect 4544 -4200 7544 -4160
rect 4544 -8120 4584 -4200
rect 7504 -8120 7544 -4200
rect 4544 -8160 7544 -8120
<< mimcapcontact >>
rect -4456 -1796 -536 2124
rect -5996 -8100 -3076 -4180
rect 4584 -8120 7504 -4200
<< metal4 >>
rect -4524 2476 -468 2492
rect -4524 2412 -4508 2476
rect -484 2412 -468 2476
rect -4524 2396 -468 2412
rect -4457 2124 -535 2125
rect -4457 -548 -4456 2124
rect -4780 -1796 -4456 -548
rect -536 -1796 -535 2124
rect -4780 -1797 -535 -1796
rect -4780 -4179 -3108 -1797
rect 6084 -2208 6960 -2192
rect 6084 -3068 6096 -2208
rect 6940 -3068 6960 -2208
rect -2804 -4128 -2708 -4112
rect -5997 -4180 -3075 -4179
rect -5997 -8100 -5996 -4180
rect -3076 -8100 -3075 -4180
rect -5997 -8101 -3075 -8100
rect -4780 -8324 -3108 -8101
rect -2804 -8152 -2788 -4128
rect -2724 -8152 -2708 -4128
rect 6084 -4199 6960 -3068
rect 7776 -4148 7872 -4132
rect 4583 -4200 7505 -4199
rect -2804 -8168 -2708 -8152
rect -1716 -7548 -1116 -7540
rect -1716 -7988 -1700 -7548
rect -1128 -7900 -1116 -7548
rect 84 -7548 684 -7540
rect -1128 -7960 -740 -7900
rect -1128 -7988 -980 -7960
rect -1716 -8160 -980 -7988
rect -800 -8160 -740 -7960
rect -1716 -8324 -740 -8160
rect 84 -7988 100 -7548
rect 672 -7988 684 -7548
rect 84 -8324 684 -7988
rect 1884 -7552 2484 -7540
rect 1884 -7992 1896 -7552
rect 2468 -7992 2484 -7552
rect 1884 -8324 2484 -7992
rect 3684 -7552 4284 -7544
rect 3684 -7992 3696 -7552
rect 4268 -7992 4284 -7552
rect 3684 -8324 4284 -7992
rect 4583 -8120 4584 -4200
rect 7504 -8120 7505 -4200
rect 4583 -8121 7505 -8120
rect 5040 -8324 6416 -8121
rect 7776 -8172 7792 -4148
rect 7856 -8172 7872 -4148
rect 7776 -8188 7872 -8172
rect -5692 -8332 7964 -8324
rect -5708 -8610 7964 -8332
rect -5708 -9416 -5444 -8610
rect -4636 -9132 7964 -8610
rect -4636 -9416 7956 -9132
rect -5708 -9628 7956 -9416
<< res1p41 >>
rect -76 876 210 1680
rect 302 876 588 1680
rect 680 876 966 1680
rect 1058 876 1344 1680
rect 1436 876 1722 1680
rect 1814 876 2100 1680
<< labels >>
rlabel metal3 -4130 2670 -3760 3010 1 VP
port 1 n
rlabel metal2 -5350 60 -4820 790 1 Out_2
port 2 n
rlabel metal2 2930 -1900 3400 -1490 1 Input
port 3 n
rlabel metal3 2560 700 2730 780 1 V_Bias1
port 5 n
rlabel metal4 -4390 -9320 -4050 -8750 1 VN
port 6 n
rlabel metal1 -3014 -2800 -2722 -2328 1 V_Bias1
port 5 n
rlabel metal3 4432 -3892 4656 -3608 1 V_Bias2
port 4 n
<< end >>
