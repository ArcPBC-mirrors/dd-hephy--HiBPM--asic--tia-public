magic
tech sky130A
magscale 1 2
timestamp 1684492973
<< dnwell >>
rect 1320 6260 4020 9160
rect 15720 6260 18420 9160
<< nwell >>
rect 6340 25196 8254 27306
rect 8560 25196 10474 27306
rect 10740 25196 12654 27306
rect 12920 25196 14834 27306
rect 15120 25196 17034 27306
rect 6340 23736 8114 25196
rect 8560 23736 10334 25196
rect 10740 23736 12514 25196
rect 12920 23736 14694 25196
rect 15120 23736 16894 25196
rect 18820 23242 19458 25232
rect 18160 23240 19458 23242
rect 18160 22404 19454 23240
rect 1240 8954 4100 9240
rect 4976 9028 7230 10502
rect 1240 6466 1526 8954
rect 3814 6466 4100 8954
rect 1240 6180 4100 6466
rect 15640 8954 18500 9240
rect 19376 9028 21630 10502
rect 15640 6466 15926 8954
rect 18214 6466 18500 8954
rect 15640 6180 18500 6466
<< pwell >>
rect 6460 21576 7754 23632
rect 8180 21576 9474 23632
rect 18160 23256 18774 25252
rect 6460 17576 8084 21486
rect 8180 17576 9804 21486
rect 18160 20936 19454 22374
rect 10020 19116 11026 19936
rect 10020 17576 11314 19014
rect 18160 18216 19784 20890
rect 2436 9288 4940 11284
rect -10200 6388 -8906 8444
rect -8880 6388 -8260 8380
rect 1540 6480 3794 8940
rect 4976 7468 7230 8906
rect -10200 4308 -8906 6364
rect -10200 308 -8576 4218
rect 76 4028 1370 6084
rect 1876 4028 3170 6084
rect 3676 4028 4970 6084
rect 5476 4028 6770 6084
rect 7476 4708 9730 10472
rect 16836 9288 19340 11284
rect 15940 6480 18194 8940
rect 19376 7468 21630 8906
rect 14476 4028 15770 6084
rect 16276 4028 17570 6084
rect 18076 4028 19370 6084
rect 19876 4028 21170 6084
rect 21876 4708 24130 10472
rect 76 28 1700 3938
rect 1876 28 3500 3938
rect 3676 28 5300 3938
rect 5476 28 7100 3938
rect 14476 28 16100 3938
rect 16276 28 17900 3938
rect 18076 28 19700 3938
rect 19876 28 21500 3938
<< pmos >>
rect 6536 26687 6636 27087
rect 6694 26687 6794 27087
rect 6852 26687 6952 27087
rect 7010 26687 7110 27087
rect 7168 26687 7268 27087
rect 7326 26687 7426 27087
rect 7484 26687 7584 27087
rect 7642 26687 7742 27087
rect 7800 26687 7900 27087
rect 7958 26687 8058 27087
rect 6536 26051 6636 26451
rect 6694 26051 6794 26451
rect 6852 26051 6952 26451
rect 7010 26051 7110 26451
rect 7168 26051 7268 26451
rect 7326 26051 7426 26451
rect 7484 26051 7584 26451
rect 7642 26051 7742 26451
rect 7800 26051 7900 26451
rect 7958 26051 8058 26451
rect 6536 25415 6636 25815
rect 6694 25415 6794 25815
rect 6852 25415 6952 25815
rect 7010 25415 7110 25815
rect 7168 25415 7268 25815
rect 7326 25415 7426 25815
rect 7484 25415 7584 25815
rect 7642 25415 7742 25815
rect 7800 25415 7900 25815
rect 7958 25415 8058 25815
rect 8756 26687 8856 27087
rect 8914 26687 9014 27087
rect 9072 26687 9172 27087
rect 9230 26687 9330 27087
rect 9388 26687 9488 27087
rect 9546 26687 9646 27087
rect 9704 26687 9804 27087
rect 9862 26687 9962 27087
rect 10020 26687 10120 27087
rect 10178 26687 10278 27087
rect 8756 26051 8856 26451
rect 8914 26051 9014 26451
rect 9072 26051 9172 26451
rect 9230 26051 9330 26451
rect 9388 26051 9488 26451
rect 9546 26051 9646 26451
rect 9704 26051 9804 26451
rect 9862 26051 9962 26451
rect 10020 26051 10120 26451
rect 10178 26051 10278 26451
rect 8756 25415 8856 25815
rect 8914 25415 9014 25815
rect 9072 25415 9172 25815
rect 9230 25415 9330 25815
rect 9388 25415 9488 25815
rect 9546 25415 9646 25815
rect 9704 25415 9804 25815
rect 9862 25415 9962 25815
rect 10020 25415 10120 25815
rect 10178 25415 10278 25815
rect 10936 26687 11036 27087
rect 11094 26687 11194 27087
rect 11252 26687 11352 27087
rect 11410 26687 11510 27087
rect 11568 26687 11668 27087
rect 11726 26687 11826 27087
rect 11884 26687 11984 27087
rect 12042 26687 12142 27087
rect 12200 26687 12300 27087
rect 12358 26687 12458 27087
rect 10936 26051 11036 26451
rect 11094 26051 11194 26451
rect 11252 26051 11352 26451
rect 11410 26051 11510 26451
rect 11568 26051 11668 26451
rect 11726 26051 11826 26451
rect 11884 26051 11984 26451
rect 12042 26051 12142 26451
rect 12200 26051 12300 26451
rect 12358 26051 12458 26451
rect 10936 25415 11036 25815
rect 11094 25415 11194 25815
rect 11252 25415 11352 25815
rect 11410 25415 11510 25815
rect 11568 25415 11668 25815
rect 11726 25415 11826 25815
rect 11884 25415 11984 25815
rect 12042 25415 12142 25815
rect 12200 25415 12300 25815
rect 12358 25415 12458 25815
rect 13116 26687 13216 27087
rect 13274 26687 13374 27087
rect 13432 26687 13532 27087
rect 13590 26687 13690 27087
rect 13748 26687 13848 27087
rect 13906 26687 14006 27087
rect 14064 26687 14164 27087
rect 14222 26687 14322 27087
rect 14380 26687 14480 27087
rect 14538 26687 14638 27087
rect 13116 26051 13216 26451
rect 13274 26051 13374 26451
rect 13432 26051 13532 26451
rect 13590 26051 13690 26451
rect 13748 26051 13848 26451
rect 13906 26051 14006 26451
rect 14064 26051 14164 26451
rect 14222 26051 14322 26451
rect 14380 26051 14480 26451
rect 14538 26051 14638 26451
rect 13116 25415 13216 25815
rect 13274 25415 13374 25815
rect 13432 25415 13532 25815
rect 13590 25415 13690 25815
rect 13748 25415 13848 25815
rect 13906 25415 14006 25815
rect 14064 25415 14164 25815
rect 14222 25415 14322 25815
rect 14380 25415 14480 25815
rect 14538 25415 14638 25815
rect 15316 26687 15416 27087
rect 15474 26687 15574 27087
rect 15632 26687 15732 27087
rect 15790 26687 15890 27087
rect 15948 26687 16048 27087
rect 16106 26687 16206 27087
rect 16264 26687 16364 27087
rect 16422 26687 16522 27087
rect 16580 26687 16680 27087
rect 16738 26687 16838 27087
rect 15316 26051 15416 26451
rect 15474 26051 15574 26451
rect 15632 26051 15732 26451
rect 15790 26051 15890 26451
rect 15948 26051 16048 26451
rect 16106 26051 16206 26451
rect 16264 26051 16364 26451
rect 16422 26051 16522 26451
rect 16580 26051 16680 26451
rect 16738 26051 16838 26451
rect 15316 25415 15416 25815
rect 15474 25415 15574 25815
rect 15632 25415 15732 25815
rect 15790 25415 15890 25815
rect 15948 25415 16048 25815
rect 16106 25415 16206 25815
rect 16264 25415 16364 25815
rect 16422 25415 16522 25815
rect 16580 25415 16680 25815
rect 16738 25415 16838 25815
rect 6540 24591 6570 24991
rect 6636 24591 6666 24991
rect 6732 24591 6762 24991
rect 6828 24591 6858 24991
rect 6924 24591 6954 24991
rect 7020 24591 7050 24991
rect 7116 24591 7146 24991
rect 7212 24591 7242 24991
rect 7308 24591 7338 24991
rect 7404 24591 7434 24991
rect 7500 24591 7530 24991
rect 7596 24591 7626 24991
rect 7692 24591 7722 24991
rect 7788 24591 7818 24991
rect 7884 24591 7914 24991
rect 6540 23955 6570 24355
rect 6636 23955 6666 24355
rect 6732 23955 6762 24355
rect 6828 23955 6858 24355
rect 6924 23955 6954 24355
rect 7020 23955 7050 24355
rect 7116 23955 7146 24355
rect 7212 23955 7242 24355
rect 7308 23955 7338 24355
rect 7404 23955 7434 24355
rect 7500 23955 7530 24355
rect 7596 23955 7626 24355
rect 7692 23955 7722 24355
rect 7788 23955 7818 24355
rect 7884 23955 7914 24355
rect 8760 24591 8790 24991
rect 8856 24591 8886 24991
rect 8952 24591 8982 24991
rect 9048 24591 9078 24991
rect 9144 24591 9174 24991
rect 9240 24591 9270 24991
rect 9336 24591 9366 24991
rect 9432 24591 9462 24991
rect 9528 24591 9558 24991
rect 9624 24591 9654 24991
rect 9720 24591 9750 24991
rect 9816 24591 9846 24991
rect 9912 24591 9942 24991
rect 10008 24591 10038 24991
rect 10104 24591 10134 24991
rect 8760 23955 8790 24355
rect 8856 23955 8886 24355
rect 8952 23955 8982 24355
rect 9048 23955 9078 24355
rect 9144 23955 9174 24355
rect 9240 23955 9270 24355
rect 9336 23955 9366 24355
rect 9432 23955 9462 24355
rect 9528 23955 9558 24355
rect 9624 23955 9654 24355
rect 9720 23955 9750 24355
rect 9816 23955 9846 24355
rect 9912 23955 9942 24355
rect 10008 23955 10038 24355
rect 10104 23955 10134 24355
rect 10940 24591 10970 24991
rect 11036 24591 11066 24991
rect 11132 24591 11162 24991
rect 11228 24591 11258 24991
rect 11324 24591 11354 24991
rect 11420 24591 11450 24991
rect 11516 24591 11546 24991
rect 11612 24591 11642 24991
rect 11708 24591 11738 24991
rect 11804 24591 11834 24991
rect 11900 24591 11930 24991
rect 11996 24591 12026 24991
rect 12092 24591 12122 24991
rect 12188 24591 12218 24991
rect 12284 24591 12314 24991
rect 10940 23955 10970 24355
rect 11036 23955 11066 24355
rect 11132 23955 11162 24355
rect 11228 23955 11258 24355
rect 11324 23955 11354 24355
rect 11420 23955 11450 24355
rect 11516 23955 11546 24355
rect 11612 23955 11642 24355
rect 11708 23955 11738 24355
rect 11804 23955 11834 24355
rect 11900 23955 11930 24355
rect 11996 23955 12026 24355
rect 12092 23955 12122 24355
rect 12188 23955 12218 24355
rect 12284 23955 12314 24355
rect 13120 24591 13150 24991
rect 13216 24591 13246 24991
rect 13312 24591 13342 24991
rect 13408 24591 13438 24991
rect 13504 24591 13534 24991
rect 13600 24591 13630 24991
rect 13696 24591 13726 24991
rect 13792 24591 13822 24991
rect 13888 24591 13918 24991
rect 13984 24591 14014 24991
rect 14080 24591 14110 24991
rect 14176 24591 14206 24991
rect 14272 24591 14302 24991
rect 14368 24591 14398 24991
rect 14464 24591 14494 24991
rect 13120 23955 13150 24355
rect 13216 23955 13246 24355
rect 13312 23955 13342 24355
rect 13408 23955 13438 24355
rect 13504 23955 13534 24355
rect 13600 23955 13630 24355
rect 13696 23955 13726 24355
rect 13792 23955 13822 24355
rect 13888 23955 13918 24355
rect 13984 23955 14014 24355
rect 14080 23955 14110 24355
rect 14176 23955 14206 24355
rect 14272 23955 14302 24355
rect 14368 23955 14398 24355
rect 14464 23955 14494 24355
rect 15320 24591 15350 24991
rect 15416 24591 15446 24991
rect 15512 24591 15542 24991
rect 15608 24591 15638 24991
rect 15704 24591 15734 24991
rect 15800 24591 15830 24991
rect 15896 24591 15926 24991
rect 15992 24591 16022 24991
rect 16088 24591 16118 24991
rect 16184 24591 16214 24991
rect 16280 24591 16310 24991
rect 16376 24591 16406 24991
rect 16472 24591 16502 24991
rect 16568 24591 16598 24991
rect 16664 24591 16694 24991
rect 15320 23955 15350 24355
rect 15416 23955 15446 24355
rect 15512 23955 15542 24355
rect 15608 23955 15638 24355
rect 15704 23955 15734 24355
rect 15800 23955 15830 24355
rect 15896 23955 15926 24355
rect 15992 23955 16022 24355
rect 16088 23955 16118 24355
rect 16184 23955 16214 24355
rect 16280 23955 16310 24355
rect 16376 23955 16406 24355
rect 16472 23955 16502 24355
rect 16568 23955 16598 24355
rect 16664 23955 16694 24355
rect 19039 23436 19239 25036
rect 18360 22623 18390 23023
rect 18456 22623 18486 23023
rect 18552 22623 18582 23023
rect 18648 22623 18678 23023
rect 18744 22623 18774 23023
rect 18840 22623 18870 23023
rect 18936 22623 18966 23023
rect 19032 22623 19062 23023
rect 19128 22623 19158 23023
rect 19224 22623 19254 23023
rect 5176 9883 5206 10283
rect 5272 9883 5302 10283
rect 5368 9883 5398 10283
rect 5464 9883 5494 10283
rect 5560 9883 5590 10283
rect 5656 9883 5686 10283
rect 5752 9883 5782 10283
rect 5848 9883 5878 10283
rect 5944 9883 5974 10283
rect 6040 9883 6070 10283
rect 6136 9883 6166 10283
rect 6232 9883 6262 10283
rect 6328 9883 6358 10283
rect 6424 9883 6454 10283
rect 6520 9883 6550 10283
rect 6616 9883 6646 10283
rect 6712 9883 6742 10283
rect 6808 9883 6838 10283
rect 6904 9883 6934 10283
rect 7000 9883 7030 10283
rect 5176 9247 5206 9647
rect 5272 9247 5302 9647
rect 5368 9247 5398 9647
rect 5464 9247 5494 9647
rect 5560 9247 5590 9647
rect 5656 9247 5686 9647
rect 5752 9247 5782 9647
rect 5848 9247 5878 9647
rect 5944 9247 5974 9647
rect 6040 9247 6070 9647
rect 6136 9247 6166 9647
rect 6232 9247 6262 9647
rect 6328 9247 6358 9647
rect 6424 9247 6454 9647
rect 6520 9247 6550 9647
rect 6616 9247 6646 9647
rect 6712 9247 6742 9647
rect 6808 9247 6838 9647
rect 6904 9247 6934 9647
rect 7000 9247 7030 9647
rect 19576 9883 19606 10283
rect 19672 9883 19702 10283
rect 19768 9883 19798 10283
rect 19864 9883 19894 10283
rect 19960 9883 19990 10283
rect 20056 9883 20086 10283
rect 20152 9883 20182 10283
rect 20248 9883 20278 10283
rect 20344 9883 20374 10283
rect 20440 9883 20470 10283
rect 20536 9883 20566 10283
rect 20632 9883 20662 10283
rect 20728 9883 20758 10283
rect 20824 9883 20854 10283
rect 20920 9883 20950 10283
rect 21016 9883 21046 10283
rect 21112 9883 21142 10283
rect 21208 9883 21238 10283
rect 21304 9883 21334 10283
rect 21400 9883 21430 10283
rect 19576 9247 19606 9647
rect 19672 9247 19702 9647
rect 19768 9247 19798 9647
rect 19864 9247 19894 9647
rect 19960 9247 19990 9647
rect 20056 9247 20086 9647
rect 20152 9247 20182 9647
rect 20248 9247 20278 9647
rect 20344 9247 20374 9647
rect 20440 9247 20470 9647
rect 20536 9247 20566 9647
rect 20632 9247 20662 9647
rect 20728 9247 20758 9647
rect 20824 9247 20854 9647
rect 20920 9247 20950 9647
rect 21016 9247 21046 9647
rect 21112 9247 21142 9647
rect 21208 9247 21238 9647
rect 21304 9247 21334 9647
rect 21400 9247 21430 9647
<< nmoslvt >>
rect 6660 23022 6690 23422
rect 6756 23022 6786 23422
rect 6852 23022 6882 23422
rect 6948 23022 6978 23422
rect 7044 23022 7074 23422
rect 7140 23022 7170 23422
rect 7236 23022 7266 23422
rect 7332 23022 7362 23422
rect 7428 23022 7458 23422
rect 7524 23022 7554 23422
rect 6660 22404 6690 22804
rect 6756 22404 6786 22804
rect 6852 22404 6882 22804
rect 6948 22404 6978 22804
rect 7044 22404 7074 22804
rect 7140 22404 7170 22804
rect 7236 22404 7266 22804
rect 7332 22404 7362 22804
rect 7428 22404 7458 22804
rect 7524 22404 7554 22804
rect 6660 21786 6690 22186
rect 6756 21786 6786 22186
rect 6852 21786 6882 22186
rect 6948 21786 6978 22186
rect 7044 21786 7074 22186
rect 7140 21786 7170 22186
rect 7236 21786 7266 22186
rect 7332 21786 7362 22186
rect 7428 21786 7458 22186
rect 7524 21786 7554 22186
rect 8380 23022 8410 23422
rect 8476 23022 8506 23422
rect 8572 23022 8602 23422
rect 8668 23022 8698 23422
rect 8764 23022 8794 23422
rect 8860 23022 8890 23422
rect 8956 23022 8986 23422
rect 9052 23022 9082 23422
rect 9148 23022 9178 23422
rect 9244 23022 9274 23422
rect 8380 22404 8410 22804
rect 8476 22404 8506 22804
rect 8572 22404 8602 22804
rect 8668 22404 8698 22804
rect 8764 22404 8794 22804
rect 8860 22404 8890 22804
rect 8956 22404 8986 22804
rect 9052 22404 9082 22804
rect 9148 22404 9178 22804
rect 9244 22404 9274 22804
rect 8380 21786 8410 22186
rect 8476 21786 8506 22186
rect 8572 21786 8602 22186
rect 8668 21786 8698 22186
rect 8764 21786 8794 22186
rect 8860 21786 8890 22186
rect 8956 21786 8986 22186
rect 9052 21786 9082 22186
rect 9148 21786 9178 22186
rect 9244 21786 9274 22186
rect 6656 20876 6856 21276
rect 6914 20876 7114 21276
rect 7172 20876 7372 21276
rect 7430 20876 7630 21276
rect 7688 20876 7888 21276
rect 6656 20258 6856 20658
rect 6914 20258 7114 20658
rect 7172 20258 7372 20658
rect 7430 20258 7630 20658
rect 7688 20258 7888 20658
rect 6656 19640 6856 20040
rect 6914 19640 7114 20040
rect 7172 19640 7372 20040
rect 7430 19640 7630 20040
rect 7688 19640 7888 20040
rect 6656 19022 6856 19422
rect 6914 19022 7114 19422
rect 7172 19022 7372 19422
rect 7430 19022 7630 19422
rect 7688 19022 7888 19422
rect 6656 18404 6856 18804
rect 6914 18404 7114 18804
rect 7172 18404 7372 18804
rect 7430 18404 7630 18804
rect 7688 18404 7888 18804
rect 6656 17786 6856 18186
rect 6914 17786 7114 18186
rect 7172 17786 7372 18186
rect 7430 17786 7630 18186
rect 7688 17786 7888 18186
rect 8376 20876 8576 21276
rect 8634 20876 8834 21276
rect 8892 20876 9092 21276
rect 9150 20876 9350 21276
rect 9408 20876 9608 21276
rect 8376 20258 8576 20658
rect 8634 20258 8834 20658
rect 8892 20258 9092 20658
rect 9150 20258 9350 20658
rect 9408 20258 9608 20658
rect 8376 19640 8576 20040
rect 8634 19640 8834 20040
rect 8892 19640 9092 20040
rect 9150 19640 9350 20040
rect 9408 19640 9608 20040
rect 8376 19022 8576 19422
rect 8634 19022 8834 19422
rect 8892 19022 9092 19422
rect 9150 19022 9350 19422
rect 9408 19022 9608 19422
rect 8376 18404 8576 18804
rect 8634 18404 8834 18804
rect 8892 18404 9092 18804
rect 9150 18404 9350 18804
rect 9408 18404 9608 18804
rect 8376 17786 8576 18186
rect 8634 17786 8834 18186
rect 8892 17786 9092 18186
rect 9150 17786 9350 18186
rect 9408 17786 9608 18186
rect 18360 21764 18390 22164
rect 18456 21764 18486 22164
rect 18552 21764 18582 22164
rect 18648 21764 18678 22164
rect 18744 21764 18774 22164
rect 18840 21764 18870 22164
rect 18936 21764 18966 22164
rect 19032 21764 19062 22164
rect 19128 21764 19158 22164
rect 19224 21764 19254 22164
rect 18360 21146 18390 21546
rect 18456 21146 18486 21546
rect 18552 21146 18582 21546
rect 18648 21146 18678 21546
rect 18744 21146 18774 21546
rect 18840 21146 18870 21546
rect 18936 21146 18966 21546
rect 19032 21146 19062 21546
rect 19128 21146 19158 21546
rect 19224 21146 19254 21546
rect 10220 19326 10250 19726
rect 10316 19326 10346 19726
rect 10412 19326 10442 19726
rect 10508 19326 10538 19726
rect 10604 19326 10634 19726
rect 10700 19326 10730 19726
rect 10796 19326 10826 19726
rect 10220 18404 10250 18804
rect 10316 18404 10346 18804
rect 10412 18404 10442 18804
rect 10508 18404 10538 18804
rect 10604 18404 10634 18804
rect 10700 18404 10730 18804
rect 10796 18404 10826 18804
rect 10892 18404 10922 18804
rect 10988 18404 11018 18804
rect 11084 18404 11114 18804
rect 10220 17786 10250 18186
rect 10316 17786 10346 18186
rect 10412 17786 10442 18186
rect 10508 17786 10538 18186
rect 10604 17786 10634 18186
rect 10700 17786 10730 18186
rect 10796 17786 10826 18186
rect 10892 17786 10922 18186
rect 10988 17786 11018 18186
rect 11084 17786 11114 18186
rect 18356 20280 18556 20680
rect 18614 20280 18814 20680
rect 18872 20280 19072 20680
rect 19130 20280 19330 20680
rect 19388 20280 19588 20680
rect 18356 19662 18556 20062
rect 18614 19662 18814 20062
rect 18872 19662 19072 20062
rect 19130 19662 19330 20062
rect 19388 19662 19588 20062
rect 18356 19044 18556 19444
rect 18614 19044 18814 19444
rect 18872 19044 19072 19444
rect 19130 19044 19330 19444
rect 19388 19044 19588 19444
rect 18356 18426 18556 18826
rect 18614 18426 18814 18826
rect 18872 18426 19072 18826
rect 19130 18426 19330 18826
rect 19388 18426 19588 18826
rect -10000 7834 -9970 8234
rect -9904 7834 -9874 8234
rect -9808 7834 -9778 8234
rect -9712 7834 -9682 8234
rect -9616 7834 -9586 8234
rect -9520 7834 -9490 8234
rect -9424 7834 -9394 8234
rect -9328 7834 -9298 8234
rect -9232 7834 -9202 8234
rect -9136 7834 -9106 8234
rect -10000 7216 -9970 7616
rect -9904 7216 -9874 7616
rect -9808 7216 -9778 7616
rect -9712 7216 -9682 7616
rect -9616 7216 -9586 7616
rect -9520 7216 -9490 7616
rect -9424 7216 -9394 7616
rect -9328 7216 -9298 7616
rect -9232 7216 -9202 7616
rect -9136 7216 -9106 7616
rect -10000 6598 -9970 6998
rect -9904 6598 -9874 6998
rect -9808 6598 -9778 6998
rect -9712 6598 -9682 6998
rect -9616 6598 -9586 6998
rect -9520 6598 -9490 6998
rect -9424 6598 -9394 6998
rect -9328 6598 -9298 6998
rect -9232 6598 -9202 6998
rect -9136 6598 -9106 6998
rect -8670 6584 -8470 8184
rect -10000 5754 -9970 6154
rect -9904 5754 -9874 6154
rect -9808 5754 -9778 6154
rect -9712 5754 -9682 6154
rect -9616 5754 -9586 6154
rect -9520 5754 -9490 6154
rect -9424 5754 -9394 6154
rect -9328 5754 -9298 6154
rect -9232 5754 -9202 6154
rect -9136 5754 -9106 6154
rect -10000 5136 -9970 5536
rect -9904 5136 -9874 5536
rect -9808 5136 -9778 5536
rect -9712 5136 -9682 5536
rect -9616 5136 -9586 5536
rect -9520 5136 -9490 5536
rect -9424 5136 -9394 5536
rect -9328 5136 -9298 5536
rect -9232 5136 -9202 5536
rect -9136 5136 -9106 5536
rect -10000 4518 -9970 4918
rect -9904 4518 -9874 4918
rect -9808 4518 -9778 4918
rect -9712 4518 -9682 4918
rect -9616 4518 -9586 4918
rect -9520 4518 -9490 4918
rect -9424 4518 -9394 4918
rect -9328 4518 -9298 4918
rect -9232 4518 -9202 4918
rect -9136 4518 -9106 4918
rect 1740 8330 1770 8730
rect 1836 8330 1866 8730
rect 1932 8330 1962 8730
rect 2028 8330 2058 8730
rect 2124 8330 2154 8730
rect 2220 8330 2250 8730
rect 2316 8330 2346 8730
rect 2412 8330 2442 8730
rect 2508 8330 2538 8730
rect 2604 8330 2634 8730
rect 2700 8330 2730 8730
rect 2796 8330 2826 8730
rect 2892 8330 2922 8730
rect 2988 8330 3018 8730
rect 3084 8330 3114 8730
rect 3180 8330 3210 8730
rect 3276 8330 3306 8730
rect 3372 8330 3402 8730
rect 3468 8330 3498 8730
rect 3564 8330 3594 8730
rect 1740 7510 1770 7910
rect 1836 7510 1866 7910
rect 1932 7510 1962 7910
rect 2028 7510 2058 7910
rect 2124 7510 2154 7910
rect 2220 7510 2250 7910
rect 2316 7510 2346 7910
rect 2412 7510 2442 7910
rect 2508 7510 2538 7910
rect 2604 7510 2634 7910
rect 2700 7510 2730 7910
rect 2796 7510 2826 7910
rect 2892 7510 2922 7910
rect 2988 7510 3018 7910
rect 3084 7510 3114 7910
rect 3180 7510 3210 7910
rect 3276 7510 3306 7910
rect 3372 7510 3402 7910
rect 3468 7510 3498 7910
rect 3564 7510 3594 7910
rect 1740 6690 1770 7090
rect 1836 6690 1866 7090
rect 1932 6690 1962 7090
rect 2028 6690 2058 7090
rect 2124 6690 2154 7090
rect 2220 6690 2250 7090
rect 2316 6690 2346 7090
rect 2412 6690 2442 7090
rect 2508 6690 2538 7090
rect 2604 6690 2634 7090
rect 2700 6690 2730 7090
rect 2796 6690 2826 7090
rect 2892 6690 2922 7090
rect 2988 6690 3018 7090
rect 3084 6690 3114 7090
rect 3180 6690 3210 7090
rect 3276 6690 3306 7090
rect 3372 6690 3402 7090
rect 3468 6690 3498 7090
rect 3564 6690 3594 7090
rect 5176 8296 5206 8696
rect 5272 8296 5302 8696
rect 5368 8296 5398 8696
rect 5464 8296 5494 8696
rect 5560 8296 5590 8696
rect 5656 8296 5686 8696
rect 5752 8296 5782 8696
rect 5848 8296 5878 8696
rect 5944 8296 5974 8696
rect 6040 8296 6070 8696
rect 6136 8296 6166 8696
rect 6232 8296 6262 8696
rect 6328 8296 6358 8696
rect 6424 8296 6454 8696
rect 6520 8296 6550 8696
rect 6616 8296 6646 8696
rect 6712 8296 6742 8696
rect 6808 8296 6838 8696
rect 6904 8296 6934 8696
rect 7000 8296 7030 8696
rect 5176 7678 5206 8078
rect 5272 7678 5302 8078
rect 5368 7678 5398 8078
rect 5464 7678 5494 8078
rect 5560 7678 5590 8078
rect 5656 7678 5686 8078
rect 5752 7678 5782 8078
rect 5848 7678 5878 8078
rect 5944 7678 5974 8078
rect 6040 7678 6070 8078
rect 6136 7678 6166 8078
rect 6232 7678 6262 8078
rect 6328 7678 6358 8078
rect 6424 7678 6454 8078
rect 6520 7678 6550 8078
rect 6616 7678 6646 8078
rect 6712 7678 6742 8078
rect 6808 7678 6838 8078
rect 6904 7678 6934 8078
rect 7000 7678 7030 8078
rect -10004 3608 -9804 4008
rect -9746 3608 -9546 4008
rect -9488 3608 -9288 4008
rect -9230 3608 -9030 4008
rect -8972 3608 -8772 4008
rect -10004 2990 -9804 3390
rect -9746 2990 -9546 3390
rect -9488 2990 -9288 3390
rect -9230 2990 -9030 3390
rect -8972 2990 -8772 3390
rect -10004 2372 -9804 2772
rect -9746 2372 -9546 2772
rect -9488 2372 -9288 2772
rect -9230 2372 -9030 2772
rect -8972 2372 -8772 2772
rect -10004 1754 -9804 2154
rect -9746 1754 -9546 2154
rect -9488 1754 -9288 2154
rect -9230 1754 -9030 2154
rect -8972 1754 -8772 2154
rect -10004 1136 -9804 1536
rect -9746 1136 -9546 1536
rect -9488 1136 -9288 1536
rect -9230 1136 -9030 1536
rect -8972 1136 -8772 1536
rect -10004 518 -9804 918
rect -9746 518 -9546 918
rect -9488 518 -9288 918
rect -9230 518 -9030 918
rect -8972 518 -8772 918
rect 276 5474 306 5874
rect 372 5474 402 5874
rect 468 5474 498 5874
rect 564 5474 594 5874
rect 660 5474 690 5874
rect 756 5474 786 5874
rect 852 5474 882 5874
rect 948 5474 978 5874
rect 1044 5474 1074 5874
rect 1140 5474 1170 5874
rect 276 4856 306 5256
rect 372 4856 402 5256
rect 468 4856 498 5256
rect 564 4856 594 5256
rect 660 4856 690 5256
rect 756 4856 786 5256
rect 852 4856 882 5256
rect 948 4856 978 5256
rect 1044 4856 1074 5256
rect 1140 4856 1170 5256
rect 276 4238 306 4638
rect 372 4238 402 4638
rect 468 4238 498 4638
rect 564 4238 594 4638
rect 660 4238 690 4638
rect 756 4238 786 4638
rect 852 4238 882 4638
rect 948 4238 978 4638
rect 1044 4238 1074 4638
rect 1140 4238 1170 4638
rect 2076 5474 2106 5874
rect 2172 5474 2202 5874
rect 2268 5474 2298 5874
rect 2364 5474 2394 5874
rect 2460 5474 2490 5874
rect 2556 5474 2586 5874
rect 2652 5474 2682 5874
rect 2748 5474 2778 5874
rect 2844 5474 2874 5874
rect 2940 5474 2970 5874
rect 2076 4856 2106 5256
rect 2172 4856 2202 5256
rect 2268 4856 2298 5256
rect 2364 4856 2394 5256
rect 2460 4856 2490 5256
rect 2556 4856 2586 5256
rect 2652 4856 2682 5256
rect 2748 4856 2778 5256
rect 2844 4856 2874 5256
rect 2940 4856 2970 5256
rect 2076 4238 2106 4638
rect 2172 4238 2202 4638
rect 2268 4238 2298 4638
rect 2364 4238 2394 4638
rect 2460 4238 2490 4638
rect 2556 4238 2586 4638
rect 2652 4238 2682 4638
rect 2748 4238 2778 4638
rect 2844 4238 2874 4638
rect 2940 4238 2970 4638
rect 3876 5474 3906 5874
rect 3972 5474 4002 5874
rect 4068 5474 4098 5874
rect 4164 5474 4194 5874
rect 4260 5474 4290 5874
rect 4356 5474 4386 5874
rect 4452 5474 4482 5874
rect 4548 5474 4578 5874
rect 4644 5474 4674 5874
rect 4740 5474 4770 5874
rect 3876 4856 3906 5256
rect 3972 4856 4002 5256
rect 4068 4856 4098 5256
rect 4164 4856 4194 5256
rect 4260 4856 4290 5256
rect 4356 4856 4386 5256
rect 4452 4856 4482 5256
rect 4548 4856 4578 5256
rect 4644 4856 4674 5256
rect 4740 4856 4770 5256
rect 3876 4238 3906 4638
rect 3972 4238 4002 4638
rect 4068 4238 4098 4638
rect 4164 4238 4194 4638
rect 4260 4238 4290 4638
rect 4356 4238 4386 4638
rect 4452 4238 4482 4638
rect 4548 4238 4578 4638
rect 4644 4238 4674 4638
rect 4740 4238 4770 4638
rect 5676 5474 5706 5874
rect 5772 5474 5802 5874
rect 5868 5474 5898 5874
rect 5964 5474 5994 5874
rect 6060 5474 6090 5874
rect 6156 5474 6186 5874
rect 6252 5474 6282 5874
rect 6348 5474 6378 5874
rect 6444 5474 6474 5874
rect 6540 5474 6570 5874
rect 5676 4856 5706 5256
rect 5772 4856 5802 5256
rect 5868 4856 5898 5256
rect 5964 4856 5994 5256
rect 6060 4856 6090 5256
rect 6156 4856 6186 5256
rect 6252 4856 6282 5256
rect 6348 4856 6378 5256
rect 6444 4856 6474 5256
rect 6540 4856 6570 5256
rect 5676 4238 5706 4638
rect 5772 4238 5802 4638
rect 5868 4238 5898 4638
rect 5964 4238 5994 4638
rect 6060 4238 6090 4638
rect 6156 4238 6186 4638
rect 6252 4238 6282 4638
rect 6348 4238 6378 4638
rect 6444 4238 6474 4638
rect 6540 4238 6570 4638
rect 7676 9862 7706 10262
rect 7772 9862 7802 10262
rect 7868 9862 7898 10262
rect 7964 9862 7994 10262
rect 8060 9862 8090 10262
rect 8156 9862 8186 10262
rect 8252 9862 8282 10262
rect 8348 9862 8378 10262
rect 8444 9862 8474 10262
rect 8540 9862 8570 10262
rect 8636 9862 8666 10262
rect 8732 9862 8762 10262
rect 8828 9862 8858 10262
rect 8924 9862 8954 10262
rect 9020 9862 9050 10262
rect 9116 9862 9146 10262
rect 9212 9862 9242 10262
rect 9308 9862 9338 10262
rect 9404 9862 9434 10262
rect 9500 9862 9530 10262
rect 7676 9244 7706 9644
rect 7772 9244 7802 9644
rect 7868 9244 7898 9644
rect 7964 9244 7994 9644
rect 8060 9244 8090 9644
rect 8156 9244 8186 9644
rect 8252 9244 8282 9644
rect 8348 9244 8378 9644
rect 8444 9244 8474 9644
rect 8540 9244 8570 9644
rect 8636 9244 8666 9644
rect 8732 9244 8762 9644
rect 8828 9244 8858 9644
rect 8924 9244 8954 9644
rect 9020 9244 9050 9644
rect 9116 9244 9146 9644
rect 9212 9244 9242 9644
rect 9308 9244 9338 9644
rect 9404 9244 9434 9644
rect 9500 9244 9530 9644
rect 7676 8626 7706 9026
rect 7772 8626 7802 9026
rect 7868 8626 7898 9026
rect 7964 8626 7994 9026
rect 8060 8626 8090 9026
rect 8156 8626 8186 9026
rect 8252 8626 8282 9026
rect 8348 8626 8378 9026
rect 8444 8626 8474 9026
rect 8540 8626 8570 9026
rect 8636 8626 8666 9026
rect 8732 8626 8762 9026
rect 8828 8626 8858 9026
rect 8924 8626 8954 9026
rect 9020 8626 9050 9026
rect 9116 8626 9146 9026
rect 9212 8626 9242 9026
rect 9308 8626 9338 9026
rect 9404 8626 9434 9026
rect 9500 8626 9530 9026
rect 7676 8008 7706 8408
rect 7772 8008 7802 8408
rect 7868 8008 7898 8408
rect 7964 8008 7994 8408
rect 8060 8008 8090 8408
rect 8156 8008 8186 8408
rect 8252 8008 8282 8408
rect 8348 8008 8378 8408
rect 8444 8008 8474 8408
rect 8540 8008 8570 8408
rect 8636 8008 8666 8408
rect 8732 8008 8762 8408
rect 8828 8008 8858 8408
rect 8924 8008 8954 8408
rect 9020 8008 9050 8408
rect 9116 8008 9146 8408
rect 9212 8008 9242 8408
rect 9308 8008 9338 8408
rect 9404 8008 9434 8408
rect 9500 8008 9530 8408
rect 7676 7390 7706 7790
rect 7772 7390 7802 7790
rect 7868 7390 7898 7790
rect 7964 7390 7994 7790
rect 8060 7390 8090 7790
rect 8156 7390 8186 7790
rect 8252 7390 8282 7790
rect 8348 7390 8378 7790
rect 8444 7390 8474 7790
rect 8540 7390 8570 7790
rect 8636 7390 8666 7790
rect 8732 7390 8762 7790
rect 8828 7390 8858 7790
rect 8924 7390 8954 7790
rect 9020 7390 9050 7790
rect 9116 7390 9146 7790
rect 9212 7390 9242 7790
rect 9308 7390 9338 7790
rect 9404 7390 9434 7790
rect 9500 7390 9530 7790
rect 7676 6772 7706 7172
rect 7772 6772 7802 7172
rect 7868 6772 7898 7172
rect 7964 6772 7994 7172
rect 8060 6772 8090 7172
rect 8156 6772 8186 7172
rect 8252 6772 8282 7172
rect 8348 6772 8378 7172
rect 8444 6772 8474 7172
rect 8540 6772 8570 7172
rect 8636 6772 8666 7172
rect 8732 6772 8762 7172
rect 8828 6772 8858 7172
rect 8924 6772 8954 7172
rect 9020 6772 9050 7172
rect 9116 6772 9146 7172
rect 9212 6772 9242 7172
rect 9308 6772 9338 7172
rect 9404 6772 9434 7172
rect 9500 6772 9530 7172
rect 7676 6154 7706 6554
rect 7772 6154 7802 6554
rect 7868 6154 7898 6554
rect 7964 6154 7994 6554
rect 8060 6154 8090 6554
rect 8156 6154 8186 6554
rect 8252 6154 8282 6554
rect 8348 6154 8378 6554
rect 8444 6154 8474 6554
rect 8540 6154 8570 6554
rect 8636 6154 8666 6554
rect 8732 6154 8762 6554
rect 8828 6154 8858 6554
rect 8924 6154 8954 6554
rect 9020 6154 9050 6554
rect 9116 6154 9146 6554
rect 9212 6154 9242 6554
rect 9308 6154 9338 6554
rect 9404 6154 9434 6554
rect 9500 6154 9530 6554
rect 7676 5536 7706 5936
rect 7772 5536 7802 5936
rect 7868 5536 7898 5936
rect 7964 5536 7994 5936
rect 8060 5536 8090 5936
rect 8156 5536 8186 5936
rect 8252 5536 8282 5936
rect 8348 5536 8378 5936
rect 8444 5536 8474 5936
rect 8540 5536 8570 5936
rect 8636 5536 8666 5936
rect 8732 5536 8762 5936
rect 8828 5536 8858 5936
rect 8924 5536 8954 5936
rect 9020 5536 9050 5936
rect 9116 5536 9146 5936
rect 9212 5536 9242 5936
rect 9308 5536 9338 5936
rect 9404 5536 9434 5936
rect 9500 5536 9530 5936
rect 7676 4918 7706 5318
rect 7772 4918 7802 5318
rect 7868 4918 7898 5318
rect 7964 4918 7994 5318
rect 8060 4918 8090 5318
rect 8156 4918 8186 5318
rect 8252 4918 8282 5318
rect 8348 4918 8378 5318
rect 8444 4918 8474 5318
rect 8540 4918 8570 5318
rect 8636 4918 8666 5318
rect 8732 4918 8762 5318
rect 8828 4918 8858 5318
rect 8924 4918 8954 5318
rect 9020 4918 9050 5318
rect 9116 4918 9146 5318
rect 9212 4918 9242 5318
rect 9308 4918 9338 5318
rect 9404 4918 9434 5318
rect 9500 4918 9530 5318
rect 16140 8330 16170 8730
rect 16236 8330 16266 8730
rect 16332 8330 16362 8730
rect 16428 8330 16458 8730
rect 16524 8330 16554 8730
rect 16620 8330 16650 8730
rect 16716 8330 16746 8730
rect 16812 8330 16842 8730
rect 16908 8330 16938 8730
rect 17004 8330 17034 8730
rect 17100 8330 17130 8730
rect 17196 8330 17226 8730
rect 17292 8330 17322 8730
rect 17388 8330 17418 8730
rect 17484 8330 17514 8730
rect 17580 8330 17610 8730
rect 17676 8330 17706 8730
rect 17772 8330 17802 8730
rect 17868 8330 17898 8730
rect 17964 8330 17994 8730
rect 16140 7510 16170 7910
rect 16236 7510 16266 7910
rect 16332 7510 16362 7910
rect 16428 7510 16458 7910
rect 16524 7510 16554 7910
rect 16620 7510 16650 7910
rect 16716 7510 16746 7910
rect 16812 7510 16842 7910
rect 16908 7510 16938 7910
rect 17004 7510 17034 7910
rect 17100 7510 17130 7910
rect 17196 7510 17226 7910
rect 17292 7510 17322 7910
rect 17388 7510 17418 7910
rect 17484 7510 17514 7910
rect 17580 7510 17610 7910
rect 17676 7510 17706 7910
rect 17772 7510 17802 7910
rect 17868 7510 17898 7910
rect 17964 7510 17994 7910
rect 16140 6690 16170 7090
rect 16236 6690 16266 7090
rect 16332 6690 16362 7090
rect 16428 6690 16458 7090
rect 16524 6690 16554 7090
rect 16620 6690 16650 7090
rect 16716 6690 16746 7090
rect 16812 6690 16842 7090
rect 16908 6690 16938 7090
rect 17004 6690 17034 7090
rect 17100 6690 17130 7090
rect 17196 6690 17226 7090
rect 17292 6690 17322 7090
rect 17388 6690 17418 7090
rect 17484 6690 17514 7090
rect 17580 6690 17610 7090
rect 17676 6690 17706 7090
rect 17772 6690 17802 7090
rect 17868 6690 17898 7090
rect 17964 6690 17994 7090
rect 19576 8296 19606 8696
rect 19672 8296 19702 8696
rect 19768 8296 19798 8696
rect 19864 8296 19894 8696
rect 19960 8296 19990 8696
rect 20056 8296 20086 8696
rect 20152 8296 20182 8696
rect 20248 8296 20278 8696
rect 20344 8296 20374 8696
rect 20440 8296 20470 8696
rect 20536 8296 20566 8696
rect 20632 8296 20662 8696
rect 20728 8296 20758 8696
rect 20824 8296 20854 8696
rect 20920 8296 20950 8696
rect 21016 8296 21046 8696
rect 21112 8296 21142 8696
rect 21208 8296 21238 8696
rect 21304 8296 21334 8696
rect 21400 8296 21430 8696
rect 19576 7678 19606 8078
rect 19672 7678 19702 8078
rect 19768 7678 19798 8078
rect 19864 7678 19894 8078
rect 19960 7678 19990 8078
rect 20056 7678 20086 8078
rect 20152 7678 20182 8078
rect 20248 7678 20278 8078
rect 20344 7678 20374 8078
rect 20440 7678 20470 8078
rect 20536 7678 20566 8078
rect 20632 7678 20662 8078
rect 20728 7678 20758 8078
rect 20824 7678 20854 8078
rect 20920 7678 20950 8078
rect 21016 7678 21046 8078
rect 21112 7678 21142 8078
rect 21208 7678 21238 8078
rect 21304 7678 21334 8078
rect 21400 7678 21430 8078
rect 14676 5474 14706 5874
rect 14772 5474 14802 5874
rect 14868 5474 14898 5874
rect 14964 5474 14994 5874
rect 15060 5474 15090 5874
rect 15156 5474 15186 5874
rect 15252 5474 15282 5874
rect 15348 5474 15378 5874
rect 15444 5474 15474 5874
rect 15540 5474 15570 5874
rect 14676 4856 14706 5256
rect 14772 4856 14802 5256
rect 14868 4856 14898 5256
rect 14964 4856 14994 5256
rect 15060 4856 15090 5256
rect 15156 4856 15186 5256
rect 15252 4856 15282 5256
rect 15348 4856 15378 5256
rect 15444 4856 15474 5256
rect 15540 4856 15570 5256
rect 14676 4238 14706 4638
rect 14772 4238 14802 4638
rect 14868 4238 14898 4638
rect 14964 4238 14994 4638
rect 15060 4238 15090 4638
rect 15156 4238 15186 4638
rect 15252 4238 15282 4638
rect 15348 4238 15378 4638
rect 15444 4238 15474 4638
rect 15540 4238 15570 4638
rect 16476 5474 16506 5874
rect 16572 5474 16602 5874
rect 16668 5474 16698 5874
rect 16764 5474 16794 5874
rect 16860 5474 16890 5874
rect 16956 5474 16986 5874
rect 17052 5474 17082 5874
rect 17148 5474 17178 5874
rect 17244 5474 17274 5874
rect 17340 5474 17370 5874
rect 16476 4856 16506 5256
rect 16572 4856 16602 5256
rect 16668 4856 16698 5256
rect 16764 4856 16794 5256
rect 16860 4856 16890 5256
rect 16956 4856 16986 5256
rect 17052 4856 17082 5256
rect 17148 4856 17178 5256
rect 17244 4856 17274 5256
rect 17340 4856 17370 5256
rect 16476 4238 16506 4638
rect 16572 4238 16602 4638
rect 16668 4238 16698 4638
rect 16764 4238 16794 4638
rect 16860 4238 16890 4638
rect 16956 4238 16986 4638
rect 17052 4238 17082 4638
rect 17148 4238 17178 4638
rect 17244 4238 17274 4638
rect 17340 4238 17370 4638
rect 18276 5474 18306 5874
rect 18372 5474 18402 5874
rect 18468 5474 18498 5874
rect 18564 5474 18594 5874
rect 18660 5474 18690 5874
rect 18756 5474 18786 5874
rect 18852 5474 18882 5874
rect 18948 5474 18978 5874
rect 19044 5474 19074 5874
rect 19140 5474 19170 5874
rect 18276 4856 18306 5256
rect 18372 4856 18402 5256
rect 18468 4856 18498 5256
rect 18564 4856 18594 5256
rect 18660 4856 18690 5256
rect 18756 4856 18786 5256
rect 18852 4856 18882 5256
rect 18948 4856 18978 5256
rect 19044 4856 19074 5256
rect 19140 4856 19170 5256
rect 18276 4238 18306 4638
rect 18372 4238 18402 4638
rect 18468 4238 18498 4638
rect 18564 4238 18594 4638
rect 18660 4238 18690 4638
rect 18756 4238 18786 4638
rect 18852 4238 18882 4638
rect 18948 4238 18978 4638
rect 19044 4238 19074 4638
rect 19140 4238 19170 4638
rect 20076 5474 20106 5874
rect 20172 5474 20202 5874
rect 20268 5474 20298 5874
rect 20364 5474 20394 5874
rect 20460 5474 20490 5874
rect 20556 5474 20586 5874
rect 20652 5474 20682 5874
rect 20748 5474 20778 5874
rect 20844 5474 20874 5874
rect 20940 5474 20970 5874
rect 20076 4856 20106 5256
rect 20172 4856 20202 5256
rect 20268 4856 20298 5256
rect 20364 4856 20394 5256
rect 20460 4856 20490 5256
rect 20556 4856 20586 5256
rect 20652 4856 20682 5256
rect 20748 4856 20778 5256
rect 20844 4856 20874 5256
rect 20940 4856 20970 5256
rect 20076 4238 20106 4638
rect 20172 4238 20202 4638
rect 20268 4238 20298 4638
rect 20364 4238 20394 4638
rect 20460 4238 20490 4638
rect 20556 4238 20586 4638
rect 20652 4238 20682 4638
rect 20748 4238 20778 4638
rect 20844 4238 20874 4638
rect 20940 4238 20970 4638
rect 22076 9862 22106 10262
rect 22172 9862 22202 10262
rect 22268 9862 22298 10262
rect 22364 9862 22394 10262
rect 22460 9862 22490 10262
rect 22556 9862 22586 10262
rect 22652 9862 22682 10262
rect 22748 9862 22778 10262
rect 22844 9862 22874 10262
rect 22940 9862 22970 10262
rect 23036 9862 23066 10262
rect 23132 9862 23162 10262
rect 23228 9862 23258 10262
rect 23324 9862 23354 10262
rect 23420 9862 23450 10262
rect 23516 9862 23546 10262
rect 23612 9862 23642 10262
rect 23708 9862 23738 10262
rect 23804 9862 23834 10262
rect 23900 9862 23930 10262
rect 22076 9244 22106 9644
rect 22172 9244 22202 9644
rect 22268 9244 22298 9644
rect 22364 9244 22394 9644
rect 22460 9244 22490 9644
rect 22556 9244 22586 9644
rect 22652 9244 22682 9644
rect 22748 9244 22778 9644
rect 22844 9244 22874 9644
rect 22940 9244 22970 9644
rect 23036 9244 23066 9644
rect 23132 9244 23162 9644
rect 23228 9244 23258 9644
rect 23324 9244 23354 9644
rect 23420 9244 23450 9644
rect 23516 9244 23546 9644
rect 23612 9244 23642 9644
rect 23708 9244 23738 9644
rect 23804 9244 23834 9644
rect 23900 9244 23930 9644
rect 22076 8626 22106 9026
rect 22172 8626 22202 9026
rect 22268 8626 22298 9026
rect 22364 8626 22394 9026
rect 22460 8626 22490 9026
rect 22556 8626 22586 9026
rect 22652 8626 22682 9026
rect 22748 8626 22778 9026
rect 22844 8626 22874 9026
rect 22940 8626 22970 9026
rect 23036 8626 23066 9026
rect 23132 8626 23162 9026
rect 23228 8626 23258 9026
rect 23324 8626 23354 9026
rect 23420 8626 23450 9026
rect 23516 8626 23546 9026
rect 23612 8626 23642 9026
rect 23708 8626 23738 9026
rect 23804 8626 23834 9026
rect 23900 8626 23930 9026
rect 22076 8008 22106 8408
rect 22172 8008 22202 8408
rect 22268 8008 22298 8408
rect 22364 8008 22394 8408
rect 22460 8008 22490 8408
rect 22556 8008 22586 8408
rect 22652 8008 22682 8408
rect 22748 8008 22778 8408
rect 22844 8008 22874 8408
rect 22940 8008 22970 8408
rect 23036 8008 23066 8408
rect 23132 8008 23162 8408
rect 23228 8008 23258 8408
rect 23324 8008 23354 8408
rect 23420 8008 23450 8408
rect 23516 8008 23546 8408
rect 23612 8008 23642 8408
rect 23708 8008 23738 8408
rect 23804 8008 23834 8408
rect 23900 8008 23930 8408
rect 22076 7390 22106 7790
rect 22172 7390 22202 7790
rect 22268 7390 22298 7790
rect 22364 7390 22394 7790
rect 22460 7390 22490 7790
rect 22556 7390 22586 7790
rect 22652 7390 22682 7790
rect 22748 7390 22778 7790
rect 22844 7390 22874 7790
rect 22940 7390 22970 7790
rect 23036 7390 23066 7790
rect 23132 7390 23162 7790
rect 23228 7390 23258 7790
rect 23324 7390 23354 7790
rect 23420 7390 23450 7790
rect 23516 7390 23546 7790
rect 23612 7390 23642 7790
rect 23708 7390 23738 7790
rect 23804 7390 23834 7790
rect 23900 7390 23930 7790
rect 22076 6772 22106 7172
rect 22172 6772 22202 7172
rect 22268 6772 22298 7172
rect 22364 6772 22394 7172
rect 22460 6772 22490 7172
rect 22556 6772 22586 7172
rect 22652 6772 22682 7172
rect 22748 6772 22778 7172
rect 22844 6772 22874 7172
rect 22940 6772 22970 7172
rect 23036 6772 23066 7172
rect 23132 6772 23162 7172
rect 23228 6772 23258 7172
rect 23324 6772 23354 7172
rect 23420 6772 23450 7172
rect 23516 6772 23546 7172
rect 23612 6772 23642 7172
rect 23708 6772 23738 7172
rect 23804 6772 23834 7172
rect 23900 6772 23930 7172
rect 22076 6154 22106 6554
rect 22172 6154 22202 6554
rect 22268 6154 22298 6554
rect 22364 6154 22394 6554
rect 22460 6154 22490 6554
rect 22556 6154 22586 6554
rect 22652 6154 22682 6554
rect 22748 6154 22778 6554
rect 22844 6154 22874 6554
rect 22940 6154 22970 6554
rect 23036 6154 23066 6554
rect 23132 6154 23162 6554
rect 23228 6154 23258 6554
rect 23324 6154 23354 6554
rect 23420 6154 23450 6554
rect 23516 6154 23546 6554
rect 23612 6154 23642 6554
rect 23708 6154 23738 6554
rect 23804 6154 23834 6554
rect 23900 6154 23930 6554
rect 22076 5536 22106 5936
rect 22172 5536 22202 5936
rect 22268 5536 22298 5936
rect 22364 5536 22394 5936
rect 22460 5536 22490 5936
rect 22556 5536 22586 5936
rect 22652 5536 22682 5936
rect 22748 5536 22778 5936
rect 22844 5536 22874 5936
rect 22940 5536 22970 5936
rect 23036 5536 23066 5936
rect 23132 5536 23162 5936
rect 23228 5536 23258 5936
rect 23324 5536 23354 5936
rect 23420 5536 23450 5936
rect 23516 5536 23546 5936
rect 23612 5536 23642 5936
rect 23708 5536 23738 5936
rect 23804 5536 23834 5936
rect 23900 5536 23930 5936
rect 22076 4918 22106 5318
rect 22172 4918 22202 5318
rect 22268 4918 22298 5318
rect 22364 4918 22394 5318
rect 22460 4918 22490 5318
rect 22556 4918 22586 5318
rect 22652 4918 22682 5318
rect 22748 4918 22778 5318
rect 22844 4918 22874 5318
rect 22940 4918 22970 5318
rect 23036 4918 23066 5318
rect 23132 4918 23162 5318
rect 23228 4918 23258 5318
rect 23324 4918 23354 5318
rect 23420 4918 23450 5318
rect 23516 4918 23546 5318
rect 23612 4918 23642 5318
rect 23708 4918 23738 5318
rect 23804 4918 23834 5318
rect 23900 4918 23930 5318
rect 272 3328 472 3728
rect 530 3328 730 3728
rect 788 3328 988 3728
rect 1046 3328 1246 3728
rect 1304 3328 1504 3728
rect 272 2710 472 3110
rect 530 2710 730 3110
rect 788 2710 988 3110
rect 1046 2710 1246 3110
rect 1304 2710 1504 3110
rect 272 2092 472 2492
rect 530 2092 730 2492
rect 788 2092 988 2492
rect 1046 2092 1246 2492
rect 1304 2092 1504 2492
rect 272 1474 472 1874
rect 530 1474 730 1874
rect 788 1474 988 1874
rect 1046 1474 1246 1874
rect 1304 1474 1504 1874
rect 272 856 472 1256
rect 530 856 730 1256
rect 788 856 988 1256
rect 1046 856 1246 1256
rect 1304 856 1504 1256
rect 272 238 472 638
rect 530 238 730 638
rect 788 238 988 638
rect 1046 238 1246 638
rect 1304 238 1504 638
rect 2072 3328 2272 3728
rect 2330 3328 2530 3728
rect 2588 3328 2788 3728
rect 2846 3328 3046 3728
rect 3104 3328 3304 3728
rect 2072 2710 2272 3110
rect 2330 2710 2530 3110
rect 2588 2710 2788 3110
rect 2846 2710 3046 3110
rect 3104 2710 3304 3110
rect 2072 2092 2272 2492
rect 2330 2092 2530 2492
rect 2588 2092 2788 2492
rect 2846 2092 3046 2492
rect 3104 2092 3304 2492
rect 2072 1474 2272 1874
rect 2330 1474 2530 1874
rect 2588 1474 2788 1874
rect 2846 1474 3046 1874
rect 3104 1474 3304 1874
rect 2072 856 2272 1256
rect 2330 856 2530 1256
rect 2588 856 2788 1256
rect 2846 856 3046 1256
rect 3104 856 3304 1256
rect 2072 238 2272 638
rect 2330 238 2530 638
rect 2588 238 2788 638
rect 2846 238 3046 638
rect 3104 238 3304 638
rect 3872 3328 4072 3728
rect 4130 3328 4330 3728
rect 4388 3328 4588 3728
rect 4646 3328 4846 3728
rect 4904 3328 5104 3728
rect 3872 2710 4072 3110
rect 4130 2710 4330 3110
rect 4388 2710 4588 3110
rect 4646 2710 4846 3110
rect 4904 2710 5104 3110
rect 3872 2092 4072 2492
rect 4130 2092 4330 2492
rect 4388 2092 4588 2492
rect 4646 2092 4846 2492
rect 4904 2092 5104 2492
rect 3872 1474 4072 1874
rect 4130 1474 4330 1874
rect 4388 1474 4588 1874
rect 4646 1474 4846 1874
rect 4904 1474 5104 1874
rect 3872 856 4072 1256
rect 4130 856 4330 1256
rect 4388 856 4588 1256
rect 4646 856 4846 1256
rect 4904 856 5104 1256
rect 3872 238 4072 638
rect 4130 238 4330 638
rect 4388 238 4588 638
rect 4646 238 4846 638
rect 4904 238 5104 638
rect 5672 3328 5872 3728
rect 5930 3328 6130 3728
rect 6188 3328 6388 3728
rect 6446 3328 6646 3728
rect 6704 3328 6904 3728
rect 5672 2710 5872 3110
rect 5930 2710 6130 3110
rect 6188 2710 6388 3110
rect 6446 2710 6646 3110
rect 6704 2710 6904 3110
rect 5672 2092 5872 2492
rect 5930 2092 6130 2492
rect 6188 2092 6388 2492
rect 6446 2092 6646 2492
rect 6704 2092 6904 2492
rect 5672 1474 5872 1874
rect 5930 1474 6130 1874
rect 6188 1474 6388 1874
rect 6446 1474 6646 1874
rect 6704 1474 6904 1874
rect 5672 856 5872 1256
rect 5930 856 6130 1256
rect 6188 856 6388 1256
rect 6446 856 6646 1256
rect 6704 856 6904 1256
rect 5672 238 5872 638
rect 5930 238 6130 638
rect 6188 238 6388 638
rect 6446 238 6646 638
rect 6704 238 6904 638
rect 14672 3328 14872 3728
rect 14930 3328 15130 3728
rect 15188 3328 15388 3728
rect 15446 3328 15646 3728
rect 15704 3328 15904 3728
rect 14672 2710 14872 3110
rect 14930 2710 15130 3110
rect 15188 2710 15388 3110
rect 15446 2710 15646 3110
rect 15704 2710 15904 3110
rect 14672 2092 14872 2492
rect 14930 2092 15130 2492
rect 15188 2092 15388 2492
rect 15446 2092 15646 2492
rect 15704 2092 15904 2492
rect 14672 1474 14872 1874
rect 14930 1474 15130 1874
rect 15188 1474 15388 1874
rect 15446 1474 15646 1874
rect 15704 1474 15904 1874
rect 14672 856 14872 1256
rect 14930 856 15130 1256
rect 15188 856 15388 1256
rect 15446 856 15646 1256
rect 15704 856 15904 1256
rect 14672 238 14872 638
rect 14930 238 15130 638
rect 15188 238 15388 638
rect 15446 238 15646 638
rect 15704 238 15904 638
rect 16472 3328 16672 3728
rect 16730 3328 16930 3728
rect 16988 3328 17188 3728
rect 17246 3328 17446 3728
rect 17504 3328 17704 3728
rect 16472 2710 16672 3110
rect 16730 2710 16930 3110
rect 16988 2710 17188 3110
rect 17246 2710 17446 3110
rect 17504 2710 17704 3110
rect 16472 2092 16672 2492
rect 16730 2092 16930 2492
rect 16988 2092 17188 2492
rect 17246 2092 17446 2492
rect 17504 2092 17704 2492
rect 16472 1474 16672 1874
rect 16730 1474 16930 1874
rect 16988 1474 17188 1874
rect 17246 1474 17446 1874
rect 17504 1474 17704 1874
rect 16472 856 16672 1256
rect 16730 856 16930 1256
rect 16988 856 17188 1256
rect 17246 856 17446 1256
rect 17504 856 17704 1256
rect 16472 238 16672 638
rect 16730 238 16930 638
rect 16988 238 17188 638
rect 17246 238 17446 638
rect 17504 238 17704 638
rect 18272 3328 18472 3728
rect 18530 3328 18730 3728
rect 18788 3328 18988 3728
rect 19046 3328 19246 3728
rect 19304 3328 19504 3728
rect 18272 2710 18472 3110
rect 18530 2710 18730 3110
rect 18788 2710 18988 3110
rect 19046 2710 19246 3110
rect 19304 2710 19504 3110
rect 18272 2092 18472 2492
rect 18530 2092 18730 2492
rect 18788 2092 18988 2492
rect 19046 2092 19246 2492
rect 19304 2092 19504 2492
rect 18272 1474 18472 1874
rect 18530 1474 18730 1874
rect 18788 1474 18988 1874
rect 19046 1474 19246 1874
rect 19304 1474 19504 1874
rect 18272 856 18472 1256
rect 18530 856 18730 1256
rect 18788 856 18988 1256
rect 19046 856 19246 1256
rect 19304 856 19504 1256
rect 18272 238 18472 638
rect 18530 238 18730 638
rect 18788 238 18988 638
rect 19046 238 19246 638
rect 19304 238 19504 638
rect 20072 3328 20272 3728
rect 20330 3328 20530 3728
rect 20588 3328 20788 3728
rect 20846 3328 21046 3728
rect 21104 3328 21304 3728
rect 20072 2710 20272 3110
rect 20330 2710 20530 3110
rect 20588 2710 20788 3110
rect 20846 2710 21046 3110
rect 21104 2710 21304 3110
rect 20072 2092 20272 2492
rect 20330 2092 20530 2492
rect 20588 2092 20788 2492
rect 20846 2092 21046 2492
rect 21104 2092 21304 2492
rect 20072 1474 20272 1874
rect 20330 1474 20530 1874
rect 20588 1474 20788 1874
rect 20846 1474 21046 1874
rect 21104 1474 21304 1874
rect 20072 856 20272 1256
rect 20330 856 20530 1256
rect 20588 856 20788 1256
rect 20846 856 21046 1256
rect 21104 856 21304 1256
rect 20072 238 20272 638
rect 20330 238 20530 638
rect 20588 238 20788 638
rect 20846 238 21046 638
rect 21104 238 21304 638
<< ndiff >>
rect 6598 23410 6660 23422
rect 6598 23034 6610 23410
rect 6644 23034 6660 23410
rect 6598 23022 6660 23034
rect 6690 23410 6756 23422
rect 6690 23034 6706 23410
rect 6740 23034 6756 23410
rect 6690 23022 6756 23034
rect 6786 23410 6852 23422
rect 6786 23034 6802 23410
rect 6836 23034 6852 23410
rect 6786 23022 6852 23034
rect 6882 23410 6948 23422
rect 6882 23034 6898 23410
rect 6932 23034 6948 23410
rect 6882 23022 6948 23034
rect 6978 23410 7044 23422
rect 6978 23034 6994 23410
rect 7028 23034 7044 23410
rect 6978 23022 7044 23034
rect 7074 23410 7140 23422
rect 7074 23034 7090 23410
rect 7124 23034 7140 23410
rect 7074 23022 7140 23034
rect 7170 23410 7236 23422
rect 7170 23034 7186 23410
rect 7220 23034 7236 23410
rect 7170 23022 7236 23034
rect 7266 23410 7332 23422
rect 7266 23034 7282 23410
rect 7316 23034 7332 23410
rect 7266 23022 7332 23034
rect 7362 23410 7428 23422
rect 7362 23034 7378 23410
rect 7412 23034 7428 23410
rect 7362 23022 7428 23034
rect 7458 23410 7524 23422
rect 7458 23034 7474 23410
rect 7508 23034 7524 23410
rect 7458 23022 7524 23034
rect 7554 23410 7616 23422
rect 7554 23034 7570 23410
rect 7604 23034 7616 23410
rect 7554 23022 7616 23034
rect 6598 22792 6660 22804
rect 6598 22416 6610 22792
rect 6644 22416 6660 22792
rect 6598 22404 6660 22416
rect 6690 22792 6756 22804
rect 6690 22416 6706 22792
rect 6740 22416 6756 22792
rect 6690 22404 6756 22416
rect 6786 22792 6852 22804
rect 6786 22416 6802 22792
rect 6836 22416 6852 22792
rect 6786 22404 6852 22416
rect 6882 22792 6948 22804
rect 6882 22416 6898 22792
rect 6932 22416 6948 22792
rect 6882 22404 6948 22416
rect 6978 22792 7044 22804
rect 6978 22416 6994 22792
rect 7028 22416 7044 22792
rect 6978 22404 7044 22416
rect 7074 22792 7140 22804
rect 7074 22416 7090 22792
rect 7124 22416 7140 22792
rect 7074 22404 7140 22416
rect 7170 22792 7236 22804
rect 7170 22416 7186 22792
rect 7220 22416 7236 22792
rect 7170 22404 7236 22416
rect 7266 22792 7332 22804
rect 7266 22416 7282 22792
rect 7316 22416 7332 22792
rect 7266 22404 7332 22416
rect 7362 22792 7428 22804
rect 7362 22416 7378 22792
rect 7412 22416 7428 22792
rect 7362 22404 7428 22416
rect 7458 22792 7524 22804
rect 7458 22416 7474 22792
rect 7508 22416 7524 22792
rect 7458 22404 7524 22416
rect 7554 22792 7616 22804
rect 7554 22416 7570 22792
rect 7604 22416 7616 22792
rect 7554 22404 7616 22416
rect 6598 22174 6660 22186
rect 6598 21798 6610 22174
rect 6644 21798 6660 22174
rect 6598 21786 6660 21798
rect 6690 22174 6756 22186
rect 6690 21798 6706 22174
rect 6740 21798 6756 22174
rect 6690 21786 6756 21798
rect 6786 22174 6852 22186
rect 6786 21798 6802 22174
rect 6836 21798 6852 22174
rect 6786 21786 6852 21798
rect 6882 22174 6948 22186
rect 6882 21798 6898 22174
rect 6932 21798 6948 22174
rect 6882 21786 6948 21798
rect 6978 22174 7044 22186
rect 6978 21798 6994 22174
rect 7028 21798 7044 22174
rect 6978 21786 7044 21798
rect 7074 22174 7140 22186
rect 7074 21798 7090 22174
rect 7124 21798 7140 22174
rect 7074 21786 7140 21798
rect 7170 22174 7236 22186
rect 7170 21798 7186 22174
rect 7220 21798 7236 22174
rect 7170 21786 7236 21798
rect 7266 22174 7332 22186
rect 7266 21798 7282 22174
rect 7316 21798 7332 22174
rect 7266 21786 7332 21798
rect 7362 22174 7428 22186
rect 7362 21798 7378 22174
rect 7412 21798 7428 22174
rect 7362 21786 7428 21798
rect 7458 22174 7524 22186
rect 7458 21798 7474 22174
rect 7508 21798 7524 22174
rect 7458 21786 7524 21798
rect 7554 22174 7616 22186
rect 7554 21798 7570 22174
rect 7604 21798 7616 22174
rect 7554 21786 7616 21798
rect 8318 23410 8380 23422
rect 8318 23034 8330 23410
rect 8364 23034 8380 23410
rect 8318 23022 8380 23034
rect 8410 23410 8476 23422
rect 8410 23034 8426 23410
rect 8460 23034 8476 23410
rect 8410 23022 8476 23034
rect 8506 23410 8572 23422
rect 8506 23034 8522 23410
rect 8556 23034 8572 23410
rect 8506 23022 8572 23034
rect 8602 23410 8668 23422
rect 8602 23034 8618 23410
rect 8652 23034 8668 23410
rect 8602 23022 8668 23034
rect 8698 23410 8764 23422
rect 8698 23034 8714 23410
rect 8748 23034 8764 23410
rect 8698 23022 8764 23034
rect 8794 23410 8860 23422
rect 8794 23034 8810 23410
rect 8844 23034 8860 23410
rect 8794 23022 8860 23034
rect 8890 23410 8956 23422
rect 8890 23034 8906 23410
rect 8940 23034 8956 23410
rect 8890 23022 8956 23034
rect 8986 23410 9052 23422
rect 8986 23034 9002 23410
rect 9036 23034 9052 23410
rect 8986 23022 9052 23034
rect 9082 23410 9148 23422
rect 9082 23034 9098 23410
rect 9132 23034 9148 23410
rect 9082 23022 9148 23034
rect 9178 23410 9244 23422
rect 9178 23034 9194 23410
rect 9228 23034 9244 23410
rect 9178 23022 9244 23034
rect 9274 23410 9336 23422
rect 9274 23034 9290 23410
rect 9324 23034 9336 23410
rect 9274 23022 9336 23034
rect 8318 22792 8380 22804
rect 8318 22416 8330 22792
rect 8364 22416 8380 22792
rect 8318 22404 8380 22416
rect 8410 22792 8476 22804
rect 8410 22416 8426 22792
rect 8460 22416 8476 22792
rect 8410 22404 8476 22416
rect 8506 22792 8572 22804
rect 8506 22416 8522 22792
rect 8556 22416 8572 22792
rect 8506 22404 8572 22416
rect 8602 22792 8668 22804
rect 8602 22416 8618 22792
rect 8652 22416 8668 22792
rect 8602 22404 8668 22416
rect 8698 22792 8764 22804
rect 8698 22416 8714 22792
rect 8748 22416 8764 22792
rect 8698 22404 8764 22416
rect 8794 22792 8860 22804
rect 8794 22416 8810 22792
rect 8844 22416 8860 22792
rect 8794 22404 8860 22416
rect 8890 22792 8956 22804
rect 8890 22416 8906 22792
rect 8940 22416 8956 22792
rect 8890 22404 8956 22416
rect 8986 22792 9052 22804
rect 8986 22416 9002 22792
rect 9036 22416 9052 22792
rect 8986 22404 9052 22416
rect 9082 22792 9148 22804
rect 9082 22416 9098 22792
rect 9132 22416 9148 22792
rect 9082 22404 9148 22416
rect 9178 22792 9244 22804
rect 9178 22416 9194 22792
rect 9228 22416 9244 22792
rect 9178 22404 9244 22416
rect 9274 22792 9336 22804
rect 9274 22416 9290 22792
rect 9324 22416 9336 22792
rect 9274 22404 9336 22416
rect 8318 22174 8380 22186
rect 8318 21798 8330 22174
rect 8364 21798 8380 22174
rect 8318 21786 8380 21798
rect 8410 22174 8476 22186
rect 8410 21798 8426 22174
rect 8460 21798 8476 22174
rect 8410 21786 8476 21798
rect 8506 22174 8572 22186
rect 8506 21798 8522 22174
rect 8556 21798 8572 22174
rect 8506 21786 8572 21798
rect 8602 22174 8668 22186
rect 8602 21798 8618 22174
rect 8652 21798 8668 22174
rect 8602 21786 8668 21798
rect 8698 22174 8764 22186
rect 8698 21798 8714 22174
rect 8748 21798 8764 22174
rect 8698 21786 8764 21798
rect 8794 22174 8860 22186
rect 8794 21798 8810 22174
rect 8844 21798 8860 22174
rect 8794 21786 8860 21798
rect 8890 22174 8956 22186
rect 8890 21798 8906 22174
rect 8940 21798 8956 22174
rect 8890 21786 8956 21798
rect 8986 22174 9052 22186
rect 8986 21798 9002 22174
rect 9036 21798 9052 22174
rect 8986 21786 9052 21798
rect 9082 22174 9148 22186
rect 9082 21798 9098 22174
rect 9132 21798 9148 22174
rect 9082 21786 9148 21798
rect 9178 22174 9244 22186
rect 9178 21798 9194 22174
rect 9228 21798 9244 22174
rect 9178 21786 9244 21798
rect 9274 22174 9336 22186
rect 9274 21798 9290 22174
rect 9324 21798 9336 22174
rect 9274 21786 9336 21798
rect 6598 21264 6656 21276
rect 6598 20888 6610 21264
rect 6644 20888 6656 21264
rect 6598 20876 6656 20888
rect 6856 21264 6914 21276
rect 6856 20888 6868 21264
rect 6902 20888 6914 21264
rect 6856 20876 6914 20888
rect 7114 21264 7172 21276
rect 7114 20888 7126 21264
rect 7160 20888 7172 21264
rect 7114 20876 7172 20888
rect 7372 21264 7430 21276
rect 7372 20888 7384 21264
rect 7418 20888 7430 21264
rect 7372 20876 7430 20888
rect 7630 21264 7688 21276
rect 7630 20888 7642 21264
rect 7676 20888 7688 21264
rect 7630 20876 7688 20888
rect 7888 21264 7946 21276
rect 7888 20888 7900 21264
rect 7934 20888 7946 21264
rect 7888 20876 7946 20888
rect 6598 20646 6656 20658
rect 6598 20270 6610 20646
rect 6644 20270 6656 20646
rect 6598 20258 6656 20270
rect 6856 20646 6914 20658
rect 6856 20270 6868 20646
rect 6902 20270 6914 20646
rect 6856 20258 6914 20270
rect 7114 20646 7172 20658
rect 7114 20270 7126 20646
rect 7160 20270 7172 20646
rect 7114 20258 7172 20270
rect 7372 20646 7430 20658
rect 7372 20270 7384 20646
rect 7418 20270 7430 20646
rect 7372 20258 7430 20270
rect 7630 20646 7688 20658
rect 7630 20270 7642 20646
rect 7676 20270 7688 20646
rect 7630 20258 7688 20270
rect 7888 20646 7946 20658
rect 7888 20270 7900 20646
rect 7934 20270 7946 20646
rect 7888 20258 7946 20270
rect 6598 20028 6656 20040
rect 6598 19652 6610 20028
rect 6644 19652 6656 20028
rect 6598 19640 6656 19652
rect 6856 20028 6914 20040
rect 6856 19652 6868 20028
rect 6902 19652 6914 20028
rect 6856 19640 6914 19652
rect 7114 20028 7172 20040
rect 7114 19652 7126 20028
rect 7160 19652 7172 20028
rect 7114 19640 7172 19652
rect 7372 20028 7430 20040
rect 7372 19652 7384 20028
rect 7418 19652 7430 20028
rect 7372 19640 7430 19652
rect 7630 20028 7688 20040
rect 7630 19652 7642 20028
rect 7676 19652 7688 20028
rect 7630 19640 7688 19652
rect 7888 20028 7946 20040
rect 7888 19652 7900 20028
rect 7934 19652 7946 20028
rect 7888 19640 7946 19652
rect 6598 19410 6656 19422
rect 6598 19034 6610 19410
rect 6644 19034 6656 19410
rect 6598 19022 6656 19034
rect 6856 19410 6914 19422
rect 6856 19034 6868 19410
rect 6902 19034 6914 19410
rect 6856 19022 6914 19034
rect 7114 19410 7172 19422
rect 7114 19034 7126 19410
rect 7160 19034 7172 19410
rect 7114 19022 7172 19034
rect 7372 19410 7430 19422
rect 7372 19034 7384 19410
rect 7418 19034 7430 19410
rect 7372 19022 7430 19034
rect 7630 19410 7688 19422
rect 7630 19034 7642 19410
rect 7676 19034 7688 19410
rect 7630 19022 7688 19034
rect 7888 19410 7946 19422
rect 7888 19034 7900 19410
rect 7934 19034 7946 19410
rect 7888 19022 7946 19034
rect 6598 18792 6656 18804
rect 6598 18416 6610 18792
rect 6644 18416 6656 18792
rect 6598 18404 6656 18416
rect 6856 18792 6914 18804
rect 6856 18416 6868 18792
rect 6902 18416 6914 18792
rect 6856 18404 6914 18416
rect 7114 18792 7172 18804
rect 7114 18416 7126 18792
rect 7160 18416 7172 18792
rect 7114 18404 7172 18416
rect 7372 18792 7430 18804
rect 7372 18416 7384 18792
rect 7418 18416 7430 18792
rect 7372 18404 7430 18416
rect 7630 18792 7688 18804
rect 7630 18416 7642 18792
rect 7676 18416 7688 18792
rect 7630 18404 7688 18416
rect 7888 18792 7946 18804
rect 7888 18416 7900 18792
rect 7934 18416 7946 18792
rect 7888 18404 7946 18416
rect 6598 18174 6656 18186
rect 6598 17798 6610 18174
rect 6644 17798 6656 18174
rect 6598 17786 6656 17798
rect 6856 18174 6914 18186
rect 6856 17798 6868 18174
rect 6902 17798 6914 18174
rect 6856 17786 6914 17798
rect 7114 18174 7172 18186
rect 7114 17798 7126 18174
rect 7160 17798 7172 18174
rect 7114 17786 7172 17798
rect 7372 18174 7430 18186
rect 7372 17798 7384 18174
rect 7418 17798 7430 18174
rect 7372 17786 7430 17798
rect 7630 18174 7688 18186
rect 7630 17798 7642 18174
rect 7676 17798 7688 18174
rect 7630 17786 7688 17798
rect 7888 18174 7946 18186
rect 7888 17798 7900 18174
rect 7934 17798 7946 18174
rect 7888 17786 7946 17798
rect 8318 21264 8376 21276
rect 8318 20888 8330 21264
rect 8364 20888 8376 21264
rect 8318 20876 8376 20888
rect 8576 21264 8634 21276
rect 8576 20888 8588 21264
rect 8622 20888 8634 21264
rect 8576 20876 8634 20888
rect 8834 21264 8892 21276
rect 8834 20888 8846 21264
rect 8880 20888 8892 21264
rect 8834 20876 8892 20888
rect 9092 21264 9150 21276
rect 9092 20888 9104 21264
rect 9138 20888 9150 21264
rect 9092 20876 9150 20888
rect 9350 21264 9408 21276
rect 9350 20888 9362 21264
rect 9396 20888 9408 21264
rect 9350 20876 9408 20888
rect 9608 21264 9666 21276
rect 9608 20888 9620 21264
rect 9654 20888 9666 21264
rect 9608 20876 9666 20888
rect 8318 20646 8376 20658
rect 8318 20270 8330 20646
rect 8364 20270 8376 20646
rect 8318 20258 8376 20270
rect 8576 20646 8634 20658
rect 8576 20270 8588 20646
rect 8622 20270 8634 20646
rect 8576 20258 8634 20270
rect 8834 20646 8892 20658
rect 8834 20270 8846 20646
rect 8880 20270 8892 20646
rect 8834 20258 8892 20270
rect 9092 20646 9150 20658
rect 9092 20270 9104 20646
rect 9138 20270 9150 20646
rect 9092 20258 9150 20270
rect 9350 20646 9408 20658
rect 9350 20270 9362 20646
rect 9396 20270 9408 20646
rect 9350 20258 9408 20270
rect 9608 20646 9666 20658
rect 9608 20270 9620 20646
rect 9654 20270 9666 20646
rect 9608 20258 9666 20270
rect 8318 20028 8376 20040
rect 8318 19652 8330 20028
rect 8364 19652 8376 20028
rect 8318 19640 8376 19652
rect 8576 20028 8634 20040
rect 8576 19652 8588 20028
rect 8622 19652 8634 20028
rect 8576 19640 8634 19652
rect 8834 20028 8892 20040
rect 8834 19652 8846 20028
rect 8880 19652 8892 20028
rect 8834 19640 8892 19652
rect 9092 20028 9150 20040
rect 9092 19652 9104 20028
rect 9138 19652 9150 20028
rect 9092 19640 9150 19652
rect 9350 20028 9408 20040
rect 9350 19652 9362 20028
rect 9396 19652 9408 20028
rect 9350 19640 9408 19652
rect 9608 20028 9666 20040
rect 9608 19652 9620 20028
rect 9654 19652 9666 20028
rect 9608 19640 9666 19652
rect 8318 19410 8376 19422
rect 8318 19034 8330 19410
rect 8364 19034 8376 19410
rect 8318 19022 8376 19034
rect 8576 19410 8634 19422
rect 8576 19034 8588 19410
rect 8622 19034 8634 19410
rect 8576 19022 8634 19034
rect 8834 19410 8892 19422
rect 8834 19034 8846 19410
rect 8880 19034 8892 19410
rect 8834 19022 8892 19034
rect 9092 19410 9150 19422
rect 9092 19034 9104 19410
rect 9138 19034 9150 19410
rect 9092 19022 9150 19034
rect 9350 19410 9408 19422
rect 9350 19034 9362 19410
rect 9396 19034 9408 19410
rect 9350 19022 9408 19034
rect 9608 19410 9666 19422
rect 9608 19034 9620 19410
rect 9654 19034 9666 19410
rect 9608 19022 9666 19034
rect 8318 18792 8376 18804
rect 8318 18416 8330 18792
rect 8364 18416 8376 18792
rect 8318 18404 8376 18416
rect 8576 18792 8634 18804
rect 8576 18416 8588 18792
rect 8622 18416 8634 18792
rect 8576 18404 8634 18416
rect 8834 18792 8892 18804
rect 8834 18416 8846 18792
rect 8880 18416 8892 18792
rect 8834 18404 8892 18416
rect 9092 18792 9150 18804
rect 9092 18416 9104 18792
rect 9138 18416 9150 18792
rect 9092 18404 9150 18416
rect 9350 18792 9408 18804
rect 9350 18416 9362 18792
rect 9396 18416 9408 18792
rect 9350 18404 9408 18416
rect 9608 18792 9666 18804
rect 9608 18416 9620 18792
rect 9654 18416 9666 18792
rect 9608 18404 9666 18416
rect 8318 18174 8376 18186
rect 8318 17798 8330 18174
rect 8364 17798 8376 18174
rect 8318 17786 8376 17798
rect 8576 18174 8634 18186
rect 8576 17798 8588 18174
rect 8622 17798 8634 18174
rect 8576 17786 8634 17798
rect 8834 18174 8892 18186
rect 8834 17798 8846 18174
rect 8880 17798 8892 18174
rect 8834 17786 8892 17798
rect 9092 18174 9150 18186
rect 9092 17798 9104 18174
rect 9138 17798 9150 18174
rect 9092 17786 9150 17798
rect 9350 18174 9408 18186
rect 9350 17798 9362 18174
rect 9396 17798 9408 18174
rect 9350 17786 9408 17798
rect 9608 18174 9666 18186
rect 9608 17798 9620 18174
rect 9654 17798 9666 18174
rect 9608 17786 9666 17798
rect 18298 22152 18360 22164
rect 18298 21776 18310 22152
rect 18344 21776 18360 22152
rect 18298 21764 18360 21776
rect 18390 22152 18456 22164
rect 18390 21776 18406 22152
rect 18440 21776 18456 22152
rect 18390 21764 18456 21776
rect 18486 22152 18552 22164
rect 18486 21776 18502 22152
rect 18536 21776 18552 22152
rect 18486 21764 18552 21776
rect 18582 22152 18648 22164
rect 18582 21776 18598 22152
rect 18632 21776 18648 22152
rect 18582 21764 18648 21776
rect 18678 22152 18744 22164
rect 18678 21776 18694 22152
rect 18728 21776 18744 22152
rect 18678 21764 18744 21776
rect 18774 22152 18840 22164
rect 18774 21776 18790 22152
rect 18824 21776 18840 22152
rect 18774 21764 18840 21776
rect 18870 22152 18936 22164
rect 18870 21776 18886 22152
rect 18920 21776 18936 22152
rect 18870 21764 18936 21776
rect 18966 22152 19032 22164
rect 18966 21776 18982 22152
rect 19016 21776 19032 22152
rect 18966 21764 19032 21776
rect 19062 22152 19128 22164
rect 19062 21776 19078 22152
rect 19112 21776 19128 22152
rect 19062 21764 19128 21776
rect 19158 22152 19224 22164
rect 19158 21776 19174 22152
rect 19208 21776 19224 22152
rect 19158 21764 19224 21776
rect 19254 22152 19316 22164
rect 19254 21776 19270 22152
rect 19304 21776 19316 22152
rect 19254 21764 19316 21776
rect 18298 21534 18360 21546
rect 18298 21158 18310 21534
rect 18344 21158 18360 21534
rect 18298 21146 18360 21158
rect 18390 21534 18456 21546
rect 18390 21158 18406 21534
rect 18440 21158 18456 21534
rect 18390 21146 18456 21158
rect 18486 21534 18552 21546
rect 18486 21158 18502 21534
rect 18536 21158 18552 21534
rect 18486 21146 18552 21158
rect 18582 21534 18648 21546
rect 18582 21158 18598 21534
rect 18632 21158 18648 21534
rect 18582 21146 18648 21158
rect 18678 21534 18744 21546
rect 18678 21158 18694 21534
rect 18728 21158 18744 21534
rect 18678 21146 18744 21158
rect 18774 21534 18840 21546
rect 18774 21158 18790 21534
rect 18824 21158 18840 21534
rect 18774 21146 18840 21158
rect 18870 21534 18936 21546
rect 18870 21158 18886 21534
rect 18920 21158 18936 21534
rect 18870 21146 18936 21158
rect 18966 21534 19032 21546
rect 18966 21158 18982 21534
rect 19016 21158 19032 21534
rect 18966 21146 19032 21158
rect 19062 21534 19128 21546
rect 19062 21158 19078 21534
rect 19112 21158 19128 21534
rect 19062 21146 19128 21158
rect 19158 21534 19224 21546
rect 19158 21158 19174 21534
rect 19208 21158 19224 21534
rect 19158 21146 19224 21158
rect 19254 21534 19316 21546
rect 19254 21158 19270 21534
rect 19304 21158 19316 21534
rect 19254 21146 19316 21158
rect 10158 19714 10220 19726
rect 10158 19338 10170 19714
rect 10204 19338 10220 19714
rect 10158 19326 10220 19338
rect 10250 19714 10316 19726
rect 10250 19338 10266 19714
rect 10300 19338 10316 19714
rect 10250 19326 10316 19338
rect 10346 19714 10412 19726
rect 10346 19338 10362 19714
rect 10396 19338 10412 19714
rect 10346 19326 10412 19338
rect 10442 19714 10508 19726
rect 10442 19338 10458 19714
rect 10492 19338 10508 19714
rect 10442 19326 10508 19338
rect 10538 19714 10604 19726
rect 10538 19338 10554 19714
rect 10588 19338 10604 19714
rect 10538 19326 10604 19338
rect 10634 19714 10700 19726
rect 10634 19338 10650 19714
rect 10684 19338 10700 19714
rect 10634 19326 10700 19338
rect 10730 19714 10796 19726
rect 10730 19338 10746 19714
rect 10780 19338 10796 19714
rect 10730 19326 10796 19338
rect 10826 19714 10888 19726
rect 10826 19338 10842 19714
rect 10876 19338 10888 19714
rect 10826 19326 10888 19338
rect 10158 18792 10220 18804
rect 10158 18416 10170 18792
rect 10204 18416 10220 18792
rect 10158 18404 10220 18416
rect 10250 18792 10316 18804
rect 10250 18416 10266 18792
rect 10300 18416 10316 18792
rect 10250 18404 10316 18416
rect 10346 18792 10412 18804
rect 10346 18416 10362 18792
rect 10396 18416 10412 18792
rect 10346 18404 10412 18416
rect 10442 18792 10508 18804
rect 10442 18416 10458 18792
rect 10492 18416 10508 18792
rect 10442 18404 10508 18416
rect 10538 18792 10604 18804
rect 10538 18416 10554 18792
rect 10588 18416 10604 18792
rect 10538 18404 10604 18416
rect 10634 18792 10700 18804
rect 10634 18416 10650 18792
rect 10684 18416 10700 18792
rect 10634 18404 10700 18416
rect 10730 18792 10796 18804
rect 10730 18416 10746 18792
rect 10780 18416 10796 18792
rect 10730 18404 10796 18416
rect 10826 18792 10892 18804
rect 10826 18416 10842 18792
rect 10876 18416 10892 18792
rect 10826 18404 10892 18416
rect 10922 18792 10988 18804
rect 10922 18416 10938 18792
rect 10972 18416 10988 18792
rect 10922 18404 10988 18416
rect 11018 18792 11084 18804
rect 11018 18416 11034 18792
rect 11068 18416 11084 18792
rect 11018 18404 11084 18416
rect 11114 18792 11176 18804
rect 11114 18416 11130 18792
rect 11164 18416 11176 18792
rect 11114 18404 11176 18416
rect 10158 18174 10220 18186
rect 10158 17798 10170 18174
rect 10204 17798 10220 18174
rect 10158 17786 10220 17798
rect 10250 18174 10316 18186
rect 10250 17798 10266 18174
rect 10300 17798 10316 18174
rect 10250 17786 10316 17798
rect 10346 18174 10412 18186
rect 10346 17798 10362 18174
rect 10396 17798 10412 18174
rect 10346 17786 10412 17798
rect 10442 18174 10508 18186
rect 10442 17798 10458 18174
rect 10492 17798 10508 18174
rect 10442 17786 10508 17798
rect 10538 18174 10604 18186
rect 10538 17798 10554 18174
rect 10588 17798 10604 18174
rect 10538 17786 10604 17798
rect 10634 18174 10700 18186
rect 10634 17798 10650 18174
rect 10684 17798 10700 18174
rect 10634 17786 10700 17798
rect 10730 18174 10796 18186
rect 10730 17798 10746 18174
rect 10780 17798 10796 18174
rect 10730 17786 10796 17798
rect 10826 18174 10892 18186
rect 10826 17798 10842 18174
rect 10876 17798 10892 18174
rect 10826 17786 10892 17798
rect 10922 18174 10988 18186
rect 10922 17798 10938 18174
rect 10972 17798 10988 18174
rect 10922 17786 10988 17798
rect 11018 18174 11084 18186
rect 11018 17798 11034 18174
rect 11068 17798 11084 18174
rect 11018 17786 11084 17798
rect 11114 18174 11176 18186
rect 11114 17798 11130 18174
rect 11164 17798 11176 18174
rect 11114 17786 11176 17798
rect 18298 20668 18356 20680
rect 18298 20292 18310 20668
rect 18344 20292 18356 20668
rect 18298 20280 18356 20292
rect 18556 20668 18614 20680
rect 18556 20292 18568 20668
rect 18602 20292 18614 20668
rect 18556 20280 18614 20292
rect 18814 20668 18872 20680
rect 18814 20292 18826 20668
rect 18860 20292 18872 20668
rect 18814 20280 18872 20292
rect 19072 20668 19130 20680
rect 19072 20292 19084 20668
rect 19118 20292 19130 20668
rect 19072 20280 19130 20292
rect 19330 20668 19388 20680
rect 19330 20292 19342 20668
rect 19376 20292 19388 20668
rect 19330 20280 19388 20292
rect 19588 20668 19646 20680
rect 19588 20292 19600 20668
rect 19634 20292 19646 20668
rect 19588 20280 19646 20292
rect 18298 20050 18356 20062
rect 18298 19674 18310 20050
rect 18344 19674 18356 20050
rect 18298 19662 18356 19674
rect 18556 20050 18614 20062
rect 18556 19674 18568 20050
rect 18602 19674 18614 20050
rect 18556 19662 18614 19674
rect 18814 20050 18872 20062
rect 18814 19674 18826 20050
rect 18860 19674 18872 20050
rect 18814 19662 18872 19674
rect 19072 20050 19130 20062
rect 19072 19674 19084 20050
rect 19118 19674 19130 20050
rect 19072 19662 19130 19674
rect 19330 20050 19388 20062
rect 19330 19674 19342 20050
rect 19376 19674 19388 20050
rect 19330 19662 19388 19674
rect 19588 20050 19646 20062
rect 19588 19674 19600 20050
rect 19634 19674 19646 20050
rect 19588 19662 19646 19674
rect 18298 19432 18356 19444
rect 18298 19056 18310 19432
rect 18344 19056 18356 19432
rect 18298 19044 18356 19056
rect 18556 19432 18614 19444
rect 18556 19056 18568 19432
rect 18602 19056 18614 19432
rect 18556 19044 18614 19056
rect 18814 19432 18872 19444
rect 18814 19056 18826 19432
rect 18860 19056 18872 19432
rect 18814 19044 18872 19056
rect 19072 19432 19130 19444
rect 19072 19056 19084 19432
rect 19118 19056 19130 19432
rect 19072 19044 19130 19056
rect 19330 19432 19388 19444
rect 19330 19056 19342 19432
rect 19376 19056 19388 19432
rect 19330 19044 19388 19056
rect 19588 19432 19646 19444
rect 19588 19056 19600 19432
rect 19634 19056 19646 19432
rect 19588 19044 19646 19056
rect 18298 18814 18356 18826
rect 18298 18438 18310 18814
rect 18344 18438 18356 18814
rect 18298 18426 18356 18438
rect 18556 18814 18614 18826
rect 18556 18438 18568 18814
rect 18602 18438 18614 18814
rect 18556 18426 18614 18438
rect 18814 18814 18872 18826
rect 18814 18438 18826 18814
rect 18860 18438 18872 18814
rect 18814 18426 18872 18438
rect 19072 18814 19130 18826
rect 19072 18438 19084 18814
rect 19118 18438 19130 18814
rect 19072 18426 19130 18438
rect 19330 18814 19388 18826
rect 19330 18438 19342 18814
rect 19376 18438 19388 18814
rect 19330 18426 19388 18438
rect 19588 18814 19646 18826
rect 19588 18438 19600 18814
rect 19634 18438 19646 18814
rect 19588 18426 19646 18438
rect -10062 8222 -10000 8234
rect -10062 7846 -10050 8222
rect -10016 7846 -10000 8222
rect -10062 7834 -10000 7846
rect -9970 8222 -9904 8234
rect -9970 7846 -9954 8222
rect -9920 7846 -9904 8222
rect -9970 7834 -9904 7846
rect -9874 8222 -9808 8234
rect -9874 7846 -9858 8222
rect -9824 7846 -9808 8222
rect -9874 7834 -9808 7846
rect -9778 8222 -9712 8234
rect -9778 7846 -9762 8222
rect -9728 7846 -9712 8222
rect -9778 7834 -9712 7846
rect -9682 8222 -9616 8234
rect -9682 7846 -9666 8222
rect -9632 7846 -9616 8222
rect -9682 7834 -9616 7846
rect -9586 8222 -9520 8234
rect -9586 7846 -9570 8222
rect -9536 7846 -9520 8222
rect -9586 7834 -9520 7846
rect -9490 8222 -9424 8234
rect -9490 7846 -9474 8222
rect -9440 7846 -9424 8222
rect -9490 7834 -9424 7846
rect -9394 8222 -9328 8234
rect -9394 7846 -9378 8222
rect -9344 7846 -9328 8222
rect -9394 7834 -9328 7846
rect -9298 8222 -9232 8234
rect -9298 7846 -9282 8222
rect -9248 7846 -9232 8222
rect -9298 7834 -9232 7846
rect -9202 8222 -9136 8234
rect -9202 7846 -9186 8222
rect -9152 7846 -9136 8222
rect -9202 7834 -9136 7846
rect -9106 8222 -9044 8234
rect -9106 7846 -9090 8222
rect -9056 7846 -9044 8222
rect -9106 7834 -9044 7846
rect -10062 7604 -10000 7616
rect -10062 7228 -10050 7604
rect -10016 7228 -10000 7604
rect -10062 7216 -10000 7228
rect -9970 7604 -9904 7616
rect -9970 7228 -9954 7604
rect -9920 7228 -9904 7604
rect -9970 7216 -9904 7228
rect -9874 7604 -9808 7616
rect -9874 7228 -9858 7604
rect -9824 7228 -9808 7604
rect -9874 7216 -9808 7228
rect -9778 7604 -9712 7616
rect -9778 7228 -9762 7604
rect -9728 7228 -9712 7604
rect -9778 7216 -9712 7228
rect -9682 7604 -9616 7616
rect -9682 7228 -9666 7604
rect -9632 7228 -9616 7604
rect -9682 7216 -9616 7228
rect -9586 7604 -9520 7616
rect -9586 7228 -9570 7604
rect -9536 7228 -9520 7604
rect -9586 7216 -9520 7228
rect -9490 7604 -9424 7616
rect -9490 7228 -9474 7604
rect -9440 7228 -9424 7604
rect -9490 7216 -9424 7228
rect -9394 7604 -9328 7616
rect -9394 7228 -9378 7604
rect -9344 7228 -9328 7604
rect -9394 7216 -9328 7228
rect -9298 7604 -9232 7616
rect -9298 7228 -9282 7604
rect -9248 7228 -9232 7604
rect -9298 7216 -9232 7228
rect -9202 7604 -9136 7616
rect -9202 7228 -9186 7604
rect -9152 7228 -9136 7604
rect -9202 7216 -9136 7228
rect -9106 7604 -9044 7616
rect -9106 7228 -9090 7604
rect -9056 7228 -9044 7604
rect -9106 7216 -9044 7228
rect -10062 6986 -10000 6998
rect -10062 6610 -10050 6986
rect -10016 6610 -10000 6986
rect -10062 6598 -10000 6610
rect -9970 6986 -9904 6998
rect -9970 6610 -9954 6986
rect -9920 6610 -9904 6986
rect -9970 6598 -9904 6610
rect -9874 6986 -9808 6998
rect -9874 6610 -9858 6986
rect -9824 6610 -9808 6986
rect -9874 6598 -9808 6610
rect -9778 6986 -9712 6998
rect -9778 6610 -9762 6986
rect -9728 6610 -9712 6986
rect -9778 6598 -9712 6610
rect -9682 6986 -9616 6998
rect -9682 6610 -9666 6986
rect -9632 6610 -9616 6986
rect -9682 6598 -9616 6610
rect -9586 6986 -9520 6998
rect -9586 6610 -9570 6986
rect -9536 6610 -9520 6986
rect -9586 6598 -9520 6610
rect -9490 6986 -9424 6998
rect -9490 6610 -9474 6986
rect -9440 6610 -9424 6986
rect -9490 6598 -9424 6610
rect -9394 6986 -9328 6998
rect -9394 6610 -9378 6986
rect -9344 6610 -9328 6986
rect -9394 6598 -9328 6610
rect -9298 6986 -9232 6998
rect -9298 6610 -9282 6986
rect -9248 6610 -9232 6986
rect -9298 6598 -9232 6610
rect -9202 6986 -9136 6998
rect -9202 6610 -9186 6986
rect -9152 6610 -9136 6986
rect -9202 6598 -9136 6610
rect -9106 6986 -9044 6998
rect -9106 6610 -9090 6986
rect -9056 6610 -9044 6986
rect -9106 6598 -9044 6610
rect -8670 8230 -8470 8242
rect -8670 8196 -8658 8230
rect -8482 8196 -8470 8230
rect -8670 8184 -8470 8196
rect -8670 6572 -8470 6584
rect -8670 6538 -8658 6572
rect -8482 6538 -8470 6572
rect -8670 6526 -8470 6538
rect -10062 6142 -10000 6154
rect -10062 5766 -10050 6142
rect -10016 5766 -10000 6142
rect -10062 5754 -10000 5766
rect -9970 6142 -9904 6154
rect -9970 5766 -9954 6142
rect -9920 5766 -9904 6142
rect -9970 5754 -9904 5766
rect -9874 6142 -9808 6154
rect -9874 5766 -9858 6142
rect -9824 5766 -9808 6142
rect -9874 5754 -9808 5766
rect -9778 6142 -9712 6154
rect -9778 5766 -9762 6142
rect -9728 5766 -9712 6142
rect -9778 5754 -9712 5766
rect -9682 6142 -9616 6154
rect -9682 5766 -9666 6142
rect -9632 5766 -9616 6142
rect -9682 5754 -9616 5766
rect -9586 6142 -9520 6154
rect -9586 5766 -9570 6142
rect -9536 5766 -9520 6142
rect -9586 5754 -9520 5766
rect -9490 6142 -9424 6154
rect -9490 5766 -9474 6142
rect -9440 5766 -9424 6142
rect -9490 5754 -9424 5766
rect -9394 6142 -9328 6154
rect -9394 5766 -9378 6142
rect -9344 5766 -9328 6142
rect -9394 5754 -9328 5766
rect -9298 6142 -9232 6154
rect -9298 5766 -9282 6142
rect -9248 5766 -9232 6142
rect -9298 5754 -9232 5766
rect -9202 6142 -9136 6154
rect -9202 5766 -9186 6142
rect -9152 5766 -9136 6142
rect -9202 5754 -9136 5766
rect -9106 6142 -9044 6154
rect -9106 5766 -9090 6142
rect -9056 5766 -9044 6142
rect -9106 5754 -9044 5766
rect -10062 5524 -10000 5536
rect -10062 5148 -10050 5524
rect -10016 5148 -10000 5524
rect -10062 5136 -10000 5148
rect -9970 5524 -9904 5536
rect -9970 5148 -9954 5524
rect -9920 5148 -9904 5524
rect -9970 5136 -9904 5148
rect -9874 5524 -9808 5536
rect -9874 5148 -9858 5524
rect -9824 5148 -9808 5524
rect -9874 5136 -9808 5148
rect -9778 5524 -9712 5536
rect -9778 5148 -9762 5524
rect -9728 5148 -9712 5524
rect -9778 5136 -9712 5148
rect -9682 5524 -9616 5536
rect -9682 5148 -9666 5524
rect -9632 5148 -9616 5524
rect -9682 5136 -9616 5148
rect -9586 5524 -9520 5536
rect -9586 5148 -9570 5524
rect -9536 5148 -9520 5524
rect -9586 5136 -9520 5148
rect -9490 5524 -9424 5536
rect -9490 5148 -9474 5524
rect -9440 5148 -9424 5524
rect -9490 5136 -9424 5148
rect -9394 5524 -9328 5536
rect -9394 5148 -9378 5524
rect -9344 5148 -9328 5524
rect -9394 5136 -9328 5148
rect -9298 5524 -9232 5536
rect -9298 5148 -9282 5524
rect -9248 5148 -9232 5524
rect -9298 5136 -9232 5148
rect -9202 5524 -9136 5536
rect -9202 5148 -9186 5524
rect -9152 5148 -9136 5524
rect -9202 5136 -9136 5148
rect -9106 5524 -9044 5536
rect -9106 5148 -9090 5524
rect -9056 5148 -9044 5524
rect -9106 5136 -9044 5148
rect -10062 4906 -10000 4918
rect -10062 4530 -10050 4906
rect -10016 4530 -10000 4906
rect -10062 4518 -10000 4530
rect -9970 4906 -9904 4918
rect -9970 4530 -9954 4906
rect -9920 4530 -9904 4906
rect -9970 4518 -9904 4530
rect -9874 4906 -9808 4918
rect -9874 4530 -9858 4906
rect -9824 4530 -9808 4906
rect -9874 4518 -9808 4530
rect -9778 4906 -9712 4918
rect -9778 4530 -9762 4906
rect -9728 4530 -9712 4906
rect -9778 4518 -9712 4530
rect -9682 4906 -9616 4918
rect -9682 4530 -9666 4906
rect -9632 4530 -9616 4906
rect -9682 4518 -9616 4530
rect -9586 4906 -9520 4918
rect -9586 4530 -9570 4906
rect -9536 4530 -9520 4906
rect -9586 4518 -9520 4530
rect -9490 4906 -9424 4918
rect -9490 4530 -9474 4906
rect -9440 4530 -9424 4906
rect -9490 4518 -9424 4530
rect -9394 4906 -9328 4918
rect -9394 4530 -9378 4906
rect -9344 4530 -9328 4906
rect -9394 4518 -9328 4530
rect -9298 4906 -9232 4918
rect -9298 4530 -9282 4906
rect -9248 4530 -9232 4906
rect -9298 4518 -9232 4530
rect -9202 4906 -9136 4918
rect -9202 4530 -9186 4906
rect -9152 4530 -9136 4906
rect -9202 4518 -9136 4530
rect -9106 4906 -9044 4918
rect -9106 4530 -9090 4906
rect -9056 4530 -9044 4906
rect -9106 4518 -9044 4530
rect 1678 8718 1740 8730
rect 1678 8342 1690 8718
rect 1724 8342 1740 8718
rect 1678 8330 1740 8342
rect 1770 8718 1836 8730
rect 1770 8342 1786 8718
rect 1820 8342 1836 8718
rect 1770 8330 1836 8342
rect 1866 8718 1932 8730
rect 1866 8342 1882 8718
rect 1916 8342 1932 8718
rect 1866 8330 1932 8342
rect 1962 8718 2028 8730
rect 1962 8342 1978 8718
rect 2012 8342 2028 8718
rect 1962 8330 2028 8342
rect 2058 8718 2124 8730
rect 2058 8342 2074 8718
rect 2108 8342 2124 8718
rect 2058 8330 2124 8342
rect 2154 8718 2220 8730
rect 2154 8342 2170 8718
rect 2204 8342 2220 8718
rect 2154 8330 2220 8342
rect 2250 8718 2316 8730
rect 2250 8342 2266 8718
rect 2300 8342 2316 8718
rect 2250 8330 2316 8342
rect 2346 8718 2412 8730
rect 2346 8342 2362 8718
rect 2396 8342 2412 8718
rect 2346 8330 2412 8342
rect 2442 8718 2508 8730
rect 2442 8342 2458 8718
rect 2492 8342 2508 8718
rect 2442 8330 2508 8342
rect 2538 8718 2604 8730
rect 2538 8342 2554 8718
rect 2588 8342 2604 8718
rect 2538 8330 2604 8342
rect 2634 8718 2700 8730
rect 2634 8342 2650 8718
rect 2684 8342 2700 8718
rect 2634 8330 2700 8342
rect 2730 8718 2796 8730
rect 2730 8342 2746 8718
rect 2780 8342 2796 8718
rect 2730 8330 2796 8342
rect 2826 8718 2892 8730
rect 2826 8342 2842 8718
rect 2876 8342 2892 8718
rect 2826 8330 2892 8342
rect 2922 8718 2988 8730
rect 2922 8342 2938 8718
rect 2972 8342 2988 8718
rect 2922 8330 2988 8342
rect 3018 8718 3084 8730
rect 3018 8342 3034 8718
rect 3068 8342 3084 8718
rect 3018 8330 3084 8342
rect 3114 8718 3180 8730
rect 3114 8342 3130 8718
rect 3164 8342 3180 8718
rect 3114 8330 3180 8342
rect 3210 8718 3276 8730
rect 3210 8342 3226 8718
rect 3260 8342 3276 8718
rect 3210 8330 3276 8342
rect 3306 8718 3372 8730
rect 3306 8342 3322 8718
rect 3356 8342 3372 8718
rect 3306 8330 3372 8342
rect 3402 8718 3468 8730
rect 3402 8342 3418 8718
rect 3452 8342 3468 8718
rect 3402 8330 3468 8342
rect 3498 8718 3564 8730
rect 3498 8342 3514 8718
rect 3548 8342 3564 8718
rect 3498 8330 3564 8342
rect 3594 8718 3656 8730
rect 3594 8342 3610 8718
rect 3644 8342 3656 8718
rect 3594 8330 3656 8342
rect 1678 7898 1740 7910
rect 1678 7522 1690 7898
rect 1724 7522 1740 7898
rect 1678 7510 1740 7522
rect 1770 7898 1836 7910
rect 1770 7522 1786 7898
rect 1820 7522 1836 7898
rect 1770 7510 1836 7522
rect 1866 7898 1932 7910
rect 1866 7522 1882 7898
rect 1916 7522 1932 7898
rect 1866 7510 1932 7522
rect 1962 7898 2028 7910
rect 1962 7522 1978 7898
rect 2012 7522 2028 7898
rect 1962 7510 2028 7522
rect 2058 7898 2124 7910
rect 2058 7522 2074 7898
rect 2108 7522 2124 7898
rect 2058 7510 2124 7522
rect 2154 7898 2220 7910
rect 2154 7522 2170 7898
rect 2204 7522 2220 7898
rect 2154 7510 2220 7522
rect 2250 7898 2316 7910
rect 2250 7522 2266 7898
rect 2300 7522 2316 7898
rect 2250 7510 2316 7522
rect 2346 7898 2412 7910
rect 2346 7522 2362 7898
rect 2396 7522 2412 7898
rect 2346 7510 2412 7522
rect 2442 7898 2508 7910
rect 2442 7522 2458 7898
rect 2492 7522 2508 7898
rect 2442 7510 2508 7522
rect 2538 7898 2604 7910
rect 2538 7522 2554 7898
rect 2588 7522 2604 7898
rect 2538 7510 2604 7522
rect 2634 7898 2700 7910
rect 2634 7522 2650 7898
rect 2684 7522 2700 7898
rect 2634 7510 2700 7522
rect 2730 7898 2796 7910
rect 2730 7522 2746 7898
rect 2780 7522 2796 7898
rect 2730 7510 2796 7522
rect 2826 7898 2892 7910
rect 2826 7522 2842 7898
rect 2876 7522 2892 7898
rect 2826 7510 2892 7522
rect 2922 7898 2988 7910
rect 2922 7522 2938 7898
rect 2972 7522 2988 7898
rect 2922 7510 2988 7522
rect 3018 7898 3084 7910
rect 3018 7522 3034 7898
rect 3068 7522 3084 7898
rect 3018 7510 3084 7522
rect 3114 7898 3180 7910
rect 3114 7522 3130 7898
rect 3164 7522 3180 7898
rect 3114 7510 3180 7522
rect 3210 7898 3276 7910
rect 3210 7522 3226 7898
rect 3260 7522 3276 7898
rect 3210 7510 3276 7522
rect 3306 7898 3372 7910
rect 3306 7522 3322 7898
rect 3356 7522 3372 7898
rect 3306 7510 3372 7522
rect 3402 7898 3468 7910
rect 3402 7522 3418 7898
rect 3452 7522 3468 7898
rect 3402 7510 3468 7522
rect 3498 7898 3564 7910
rect 3498 7522 3514 7898
rect 3548 7522 3564 7898
rect 3498 7510 3564 7522
rect 3594 7898 3656 7910
rect 3594 7522 3610 7898
rect 3644 7522 3656 7898
rect 3594 7510 3656 7522
rect 1678 7078 1740 7090
rect 1678 6702 1690 7078
rect 1724 6702 1740 7078
rect 1678 6690 1740 6702
rect 1770 7078 1836 7090
rect 1770 6702 1786 7078
rect 1820 6702 1836 7078
rect 1770 6690 1836 6702
rect 1866 7078 1932 7090
rect 1866 6702 1882 7078
rect 1916 6702 1932 7078
rect 1866 6690 1932 6702
rect 1962 7078 2028 7090
rect 1962 6702 1978 7078
rect 2012 6702 2028 7078
rect 1962 6690 2028 6702
rect 2058 7078 2124 7090
rect 2058 6702 2074 7078
rect 2108 6702 2124 7078
rect 2058 6690 2124 6702
rect 2154 7078 2220 7090
rect 2154 6702 2170 7078
rect 2204 6702 2220 7078
rect 2154 6690 2220 6702
rect 2250 7078 2316 7090
rect 2250 6702 2266 7078
rect 2300 6702 2316 7078
rect 2250 6690 2316 6702
rect 2346 7078 2412 7090
rect 2346 6702 2362 7078
rect 2396 6702 2412 7078
rect 2346 6690 2412 6702
rect 2442 7078 2508 7090
rect 2442 6702 2458 7078
rect 2492 6702 2508 7078
rect 2442 6690 2508 6702
rect 2538 7078 2604 7090
rect 2538 6702 2554 7078
rect 2588 6702 2604 7078
rect 2538 6690 2604 6702
rect 2634 7078 2700 7090
rect 2634 6702 2650 7078
rect 2684 6702 2700 7078
rect 2634 6690 2700 6702
rect 2730 7078 2796 7090
rect 2730 6702 2746 7078
rect 2780 6702 2796 7078
rect 2730 6690 2796 6702
rect 2826 7078 2892 7090
rect 2826 6702 2842 7078
rect 2876 6702 2892 7078
rect 2826 6690 2892 6702
rect 2922 7078 2988 7090
rect 2922 6702 2938 7078
rect 2972 6702 2988 7078
rect 2922 6690 2988 6702
rect 3018 7078 3084 7090
rect 3018 6702 3034 7078
rect 3068 6702 3084 7078
rect 3018 6690 3084 6702
rect 3114 7078 3180 7090
rect 3114 6702 3130 7078
rect 3164 6702 3180 7078
rect 3114 6690 3180 6702
rect 3210 7078 3276 7090
rect 3210 6702 3226 7078
rect 3260 6702 3276 7078
rect 3210 6690 3276 6702
rect 3306 7078 3372 7090
rect 3306 6702 3322 7078
rect 3356 6702 3372 7078
rect 3306 6690 3372 6702
rect 3402 7078 3468 7090
rect 3402 6702 3418 7078
rect 3452 6702 3468 7078
rect 3402 6690 3468 6702
rect 3498 7078 3564 7090
rect 3498 6702 3514 7078
rect 3548 6702 3564 7078
rect 3498 6690 3564 6702
rect 3594 7078 3656 7090
rect 3594 6702 3610 7078
rect 3644 6702 3656 7078
rect 3594 6690 3656 6702
rect 5114 8684 5176 8696
rect 5114 8308 5126 8684
rect 5160 8308 5176 8684
rect 5114 8296 5176 8308
rect 5206 8684 5272 8696
rect 5206 8308 5222 8684
rect 5256 8308 5272 8684
rect 5206 8296 5272 8308
rect 5302 8684 5368 8696
rect 5302 8308 5318 8684
rect 5352 8308 5368 8684
rect 5302 8296 5368 8308
rect 5398 8684 5464 8696
rect 5398 8308 5414 8684
rect 5448 8308 5464 8684
rect 5398 8296 5464 8308
rect 5494 8684 5560 8696
rect 5494 8308 5510 8684
rect 5544 8308 5560 8684
rect 5494 8296 5560 8308
rect 5590 8684 5656 8696
rect 5590 8308 5606 8684
rect 5640 8308 5656 8684
rect 5590 8296 5656 8308
rect 5686 8684 5752 8696
rect 5686 8308 5702 8684
rect 5736 8308 5752 8684
rect 5686 8296 5752 8308
rect 5782 8684 5848 8696
rect 5782 8308 5798 8684
rect 5832 8308 5848 8684
rect 5782 8296 5848 8308
rect 5878 8684 5944 8696
rect 5878 8308 5894 8684
rect 5928 8308 5944 8684
rect 5878 8296 5944 8308
rect 5974 8684 6040 8696
rect 5974 8308 5990 8684
rect 6024 8308 6040 8684
rect 5974 8296 6040 8308
rect 6070 8684 6136 8696
rect 6070 8308 6086 8684
rect 6120 8308 6136 8684
rect 6070 8296 6136 8308
rect 6166 8684 6232 8696
rect 6166 8308 6182 8684
rect 6216 8308 6232 8684
rect 6166 8296 6232 8308
rect 6262 8684 6328 8696
rect 6262 8308 6278 8684
rect 6312 8308 6328 8684
rect 6262 8296 6328 8308
rect 6358 8684 6424 8696
rect 6358 8308 6374 8684
rect 6408 8308 6424 8684
rect 6358 8296 6424 8308
rect 6454 8684 6520 8696
rect 6454 8308 6470 8684
rect 6504 8308 6520 8684
rect 6454 8296 6520 8308
rect 6550 8684 6616 8696
rect 6550 8308 6566 8684
rect 6600 8308 6616 8684
rect 6550 8296 6616 8308
rect 6646 8684 6712 8696
rect 6646 8308 6662 8684
rect 6696 8308 6712 8684
rect 6646 8296 6712 8308
rect 6742 8684 6808 8696
rect 6742 8308 6758 8684
rect 6792 8308 6808 8684
rect 6742 8296 6808 8308
rect 6838 8684 6904 8696
rect 6838 8308 6854 8684
rect 6888 8308 6904 8684
rect 6838 8296 6904 8308
rect 6934 8684 7000 8696
rect 6934 8308 6950 8684
rect 6984 8308 7000 8684
rect 6934 8296 7000 8308
rect 7030 8684 7092 8696
rect 7030 8308 7046 8684
rect 7080 8308 7092 8684
rect 7030 8296 7092 8308
rect 5114 8066 5176 8078
rect 5114 7690 5126 8066
rect 5160 7690 5176 8066
rect 5114 7678 5176 7690
rect 5206 8066 5272 8078
rect 5206 7690 5222 8066
rect 5256 7690 5272 8066
rect 5206 7678 5272 7690
rect 5302 8066 5368 8078
rect 5302 7690 5318 8066
rect 5352 7690 5368 8066
rect 5302 7678 5368 7690
rect 5398 8066 5464 8078
rect 5398 7690 5414 8066
rect 5448 7690 5464 8066
rect 5398 7678 5464 7690
rect 5494 8066 5560 8078
rect 5494 7690 5510 8066
rect 5544 7690 5560 8066
rect 5494 7678 5560 7690
rect 5590 8066 5656 8078
rect 5590 7690 5606 8066
rect 5640 7690 5656 8066
rect 5590 7678 5656 7690
rect 5686 8066 5752 8078
rect 5686 7690 5702 8066
rect 5736 7690 5752 8066
rect 5686 7678 5752 7690
rect 5782 8066 5848 8078
rect 5782 7690 5798 8066
rect 5832 7690 5848 8066
rect 5782 7678 5848 7690
rect 5878 8066 5944 8078
rect 5878 7690 5894 8066
rect 5928 7690 5944 8066
rect 5878 7678 5944 7690
rect 5974 8066 6040 8078
rect 5974 7690 5990 8066
rect 6024 7690 6040 8066
rect 5974 7678 6040 7690
rect 6070 8066 6136 8078
rect 6070 7690 6086 8066
rect 6120 7690 6136 8066
rect 6070 7678 6136 7690
rect 6166 8066 6232 8078
rect 6166 7690 6182 8066
rect 6216 7690 6232 8066
rect 6166 7678 6232 7690
rect 6262 8066 6328 8078
rect 6262 7690 6278 8066
rect 6312 7690 6328 8066
rect 6262 7678 6328 7690
rect 6358 8066 6424 8078
rect 6358 7690 6374 8066
rect 6408 7690 6424 8066
rect 6358 7678 6424 7690
rect 6454 8066 6520 8078
rect 6454 7690 6470 8066
rect 6504 7690 6520 8066
rect 6454 7678 6520 7690
rect 6550 8066 6616 8078
rect 6550 7690 6566 8066
rect 6600 7690 6616 8066
rect 6550 7678 6616 7690
rect 6646 8066 6712 8078
rect 6646 7690 6662 8066
rect 6696 7690 6712 8066
rect 6646 7678 6712 7690
rect 6742 8066 6808 8078
rect 6742 7690 6758 8066
rect 6792 7690 6808 8066
rect 6742 7678 6808 7690
rect 6838 8066 6904 8078
rect 6838 7690 6854 8066
rect 6888 7690 6904 8066
rect 6838 7678 6904 7690
rect 6934 8066 7000 8078
rect 6934 7690 6950 8066
rect 6984 7690 7000 8066
rect 6934 7678 7000 7690
rect 7030 8066 7092 8078
rect 7030 7690 7046 8066
rect 7080 7690 7092 8066
rect 7030 7678 7092 7690
rect -10062 3996 -10004 4008
rect -10062 3620 -10050 3996
rect -10016 3620 -10004 3996
rect -10062 3608 -10004 3620
rect -9804 3996 -9746 4008
rect -9804 3620 -9792 3996
rect -9758 3620 -9746 3996
rect -9804 3608 -9746 3620
rect -9546 3996 -9488 4008
rect -9546 3620 -9534 3996
rect -9500 3620 -9488 3996
rect -9546 3608 -9488 3620
rect -9288 3996 -9230 4008
rect -9288 3620 -9276 3996
rect -9242 3620 -9230 3996
rect -9288 3608 -9230 3620
rect -9030 3996 -8972 4008
rect -9030 3620 -9018 3996
rect -8984 3620 -8972 3996
rect -9030 3608 -8972 3620
rect -8772 3996 -8714 4008
rect -8772 3620 -8760 3996
rect -8726 3620 -8714 3996
rect -8772 3608 -8714 3620
rect -10062 3378 -10004 3390
rect -10062 3002 -10050 3378
rect -10016 3002 -10004 3378
rect -10062 2990 -10004 3002
rect -9804 3378 -9746 3390
rect -9804 3002 -9792 3378
rect -9758 3002 -9746 3378
rect -9804 2990 -9746 3002
rect -9546 3378 -9488 3390
rect -9546 3002 -9534 3378
rect -9500 3002 -9488 3378
rect -9546 2990 -9488 3002
rect -9288 3378 -9230 3390
rect -9288 3002 -9276 3378
rect -9242 3002 -9230 3378
rect -9288 2990 -9230 3002
rect -9030 3378 -8972 3390
rect -9030 3002 -9018 3378
rect -8984 3002 -8972 3378
rect -9030 2990 -8972 3002
rect -8772 3378 -8714 3390
rect -8772 3002 -8760 3378
rect -8726 3002 -8714 3378
rect -8772 2990 -8714 3002
rect -10062 2760 -10004 2772
rect -10062 2384 -10050 2760
rect -10016 2384 -10004 2760
rect -10062 2372 -10004 2384
rect -9804 2760 -9746 2772
rect -9804 2384 -9792 2760
rect -9758 2384 -9746 2760
rect -9804 2372 -9746 2384
rect -9546 2760 -9488 2772
rect -9546 2384 -9534 2760
rect -9500 2384 -9488 2760
rect -9546 2372 -9488 2384
rect -9288 2760 -9230 2772
rect -9288 2384 -9276 2760
rect -9242 2384 -9230 2760
rect -9288 2372 -9230 2384
rect -9030 2760 -8972 2772
rect -9030 2384 -9018 2760
rect -8984 2384 -8972 2760
rect -9030 2372 -8972 2384
rect -8772 2760 -8714 2772
rect -8772 2384 -8760 2760
rect -8726 2384 -8714 2760
rect -8772 2372 -8714 2384
rect -10062 2142 -10004 2154
rect -10062 1766 -10050 2142
rect -10016 1766 -10004 2142
rect -10062 1754 -10004 1766
rect -9804 2142 -9746 2154
rect -9804 1766 -9792 2142
rect -9758 1766 -9746 2142
rect -9804 1754 -9746 1766
rect -9546 2142 -9488 2154
rect -9546 1766 -9534 2142
rect -9500 1766 -9488 2142
rect -9546 1754 -9488 1766
rect -9288 2142 -9230 2154
rect -9288 1766 -9276 2142
rect -9242 1766 -9230 2142
rect -9288 1754 -9230 1766
rect -9030 2142 -8972 2154
rect -9030 1766 -9018 2142
rect -8984 1766 -8972 2142
rect -9030 1754 -8972 1766
rect -8772 2142 -8714 2154
rect -8772 1766 -8760 2142
rect -8726 1766 -8714 2142
rect -8772 1754 -8714 1766
rect -10062 1524 -10004 1536
rect -10062 1148 -10050 1524
rect -10016 1148 -10004 1524
rect -10062 1136 -10004 1148
rect -9804 1524 -9746 1536
rect -9804 1148 -9792 1524
rect -9758 1148 -9746 1524
rect -9804 1136 -9746 1148
rect -9546 1524 -9488 1536
rect -9546 1148 -9534 1524
rect -9500 1148 -9488 1524
rect -9546 1136 -9488 1148
rect -9288 1524 -9230 1536
rect -9288 1148 -9276 1524
rect -9242 1148 -9230 1524
rect -9288 1136 -9230 1148
rect -9030 1524 -8972 1536
rect -9030 1148 -9018 1524
rect -8984 1148 -8972 1524
rect -9030 1136 -8972 1148
rect -8772 1524 -8714 1536
rect -8772 1148 -8760 1524
rect -8726 1148 -8714 1524
rect -8772 1136 -8714 1148
rect -10062 906 -10004 918
rect -10062 530 -10050 906
rect -10016 530 -10004 906
rect -10062 518 -10004 530
rect -9804 906 -9746 918
rect -9804 530 -9792 906
rect -9758 530 -9746 906
rect -9804 518 -9746 530
rect -9546 906 -9488 918
rect -9546 530 -9534 906
rect -9500 530 -9488 906
rect -9546 518 -9488 530
rect -9288 906 -9230 918
rect -9288 530 -9276 906
rect -9242 530 -9230 906
rect -9288 518 -9230 530
rect -9030 906 -8972 918
rect -9030 530 -9018 906
rect -8984 530 -8972 906
rect -9030 518 -8972 530
rect -8772 906 -8714 918
rect -8772 530 -8760 906
rect -8726 530 -8714 906
rect -8772 518 -8714 530
rect 214 5862 276 5874
rect 214 5486 226 5862
rect 260 5486 276 5862
rect 214 5474 276 5486
rect 306 5862 372 5874
rect 306 5486 322 5862
rect 356 5486 372 5862
rect 306 5474 372 5486
rect 402 5862 468 5874
rect 402 5486 418 5862
rect 452 5486 468 5862
rect 402 5474 468 5486
rect 498 5862 564 5874
rect 498 5486 514 5862
rect 548 5486 564 5862
rect 498 5474 564 5486
rect 594 5862 660 5874
rect 594 5486 610 5862
rect 644 5486 660 5862
rect 594 5474 660 5486
rect 690 5862 756 5874
rect 690 5486 706 5862
rect 740 5486 756 5862
rect 690 5474 756 5486
rect 786 5862 852 5874
rect 786 5486 802 5862
rect 836 5486 852 5862
rect 786 5474 852 5486
rect 882 5862 948 5874
rect 882 5486 898 5862
rect 932 5486 948 5862
rect 882 5474 948 5486
rect 978 5862 1044 5874
rect 978 5486 994 5862
rect 1028 5486 1044 5862
rect 978 5474 1044 5486
rect 1074 5862 1140 5874
rect 1074 5486 1090 5862
rect 1124 5486 1140 5862
rect 1074 5474 1140 5486
rect 1170 5862 1232 5874
rect 1170 5486 1186 5862
rect 1220 5486 1232 5862
rect 1170 5474 1232 5486
rect 214 5244 276 5256
rect 214 4868 226 5244
rect 260 4868 276 5244
rect 214 4856 276 4868
rect 306 5244 372 5256
rect 306 4868 322 5244
rect 356 4868 372 5244
rect 306 4856 372 4868
rect 402 5244 468 5256
rect 402 4868 418 5244
rect 452 4868 468 5244
rect 402 4856 468 4868
rect 498 5244 564 5256
rect 498 4868 514 5244
rect 548 4868 564 5244
rect 498 4856 564 4868
rect 594 5244 660 5256
rect 594 4868 610 5244
rect 644 4868 660 5244
rect 594 4856 660 4868
rect 690 5244 756 5256
rect 690 4868 706 5244
rect 740 4868 756 5244
rect 690 4856 756 4868
rect 786 5244 852 5256
rect 786 4868 802 5244
rect 836 4868 852 5244
rect 786 4856 852 4868
rect 882 5244 948 5256
rect 882 4868 898 5244
rect 932 4868 948 5244
rect 882 4856 948 4868
rect 978 5244 1044 5256
rect 978 4868 994 5244
rect 1028 4868 1044 5244
rect 978 4856 1044 4868
rect 1074 5244 1140 5256
rect 1074 4868 1090 5244
rect 1124 4868 1140 5244
rect 1074 4856 1140 4868
rect 1170 5244 1232 5256
rect 1170 4868 1186 5244
rect 1220 4868 1232 5244
rect 1170 4856 1232 4868
rect 214 4626 276 4638
rect 214 4250 226 4626
rect 260 4250 276 4626
rect 214 4238 276 4250
rect 306 4626 372 4638
rect 306 4250 322 4626
rect 356 4250 372 4626
rect 306 4238 372 4250
rect 402 4626 468 4638
rect 402 4250 418 4626
rect 452 4250 468 4626
rect 402 4238 468 4250
rect 498 4626 564 4638
rect 498 4250 514 4626
rect 548 4250 564 4626
rect 498 4238 564 4250
rect 594 4626 660 4638
rect 594 4250 610 4626
rect 644 4250 660 4626
rect 594 4238 660 4250
rect 690 4626 756 4638
rect 690 4250 706 4626
rect 740 4250 756 4626
rect 690 4238 756 4250
rect 786 4626 852 4638
rect 786 4250 802 4626
rect 836 4250 852 4626
rect 786 4238 852 4250
rect 882 4626 948 4638
rect 882 4250 898 4626
rect 932 4250 948 4626
rect 882 4238 948 4250
rect 978 4626 1044 4638
rect 978 4250 994 4626
rect 1028 4250 1044 4626
rect 978 4238 1044 4250
rect 1074 4626 1140 4638
rect 1074 4250 1090 4626
rect 1124 4250 1140 4626
rect 1074 4238 1140 4250
rect 1170 4626 1232 4638
rect 1170 4250 1186 4626
rect 1220 4250 1232 4626
rect 1170 4238 1232 4250
rect 2014 5862 2076 5874
rect 2014 5486 2026 5862
rect 2060 5486 2076 5862
rect 2014 5474 2076 5486
rect 2106 5862 2172 5874
rect 2106 5486 2122 5862
rect 2156 5486 2172 5862
rect 2106 5474 2172 5486
rect 2202 5862 2268 5874
rect 2202 5486 2218 5862
rect 2252 5486 2268 5862
rect 2202 5474 2268 5486
rect 2298 5862 2364 5874
rect 2298 5486 2314 5862
rect 2348 5486 2364 5862
rect 2298 5474 2364 5486
rect 2394 5862 2460 5874
rect 2394 5486 2410 5862
rect 2444 5486 2460 5862
rect 2394 5474 2460 5486
rect 2490 5862 2556 5874
rect 2490 5486 2506 5862
rect 2540 5486 2556 5862
rect 2490 5474 2556 5486
rect 2586 5862 2652 5874
rect 2586 5486 2602 5862
rect 2636 5486 2652 5862
rect 2586 5474 2652 5486
rect 2682 5862 2748 5874
rect 2682 5486 2698 5862
rect 2732 5486 2748 5862
rect 2682 5474 2748 5486
rect 2778 5862 2844 5874
rect 2778 5486 2794 5862
rect 2828 5486 2844 5862
rect 2778 5474 2844 5486
rect 2874 5862 2940 5874
rect 2874 5486 2890 5862
rect 2924 5486 2940 5862
rect 2874 5474 2940 5486
rect 2970 5862 3032 5874
rect 2970 5486 2986 5862
rect 3020 5486 3032 5862
rect 2970 5474 3032 5486
rect 2014 5244 2076 5256
rect 2014 4868 2026 5244
rect 2060 4868 2076 5244
rect 2014 4856 2076 4868
rect 2106 5244 2172 5256
rect 2106 4868 2122 5244
rect 2156 4868 2172 5244
rect 2106 4856 2172 4868
rect 2202 5244 2268 5256
rect 2202 4868 2218 5244
rect 2252 4868 2268 5244
rect 2202 4856 2268 4868
rect 2298 5244 2364 5256
rect 2298 4868 2314 5244
rect 2348 4868 2364 5244
rect 2298 4856 2364 4868
rect 2394 5244 2460 5256
rect 2394 4868 2410 5244
rect 2444 4868 2460 5244
rect 2394 4856 2460 4868
rect 2490 5244 2556 5256
rect 2490 4868 2506 5244
rect 2540 4868 2556 5244
rect 2490 4856 2556 4868
rect 2586 5244 2652 5256
rect 2586 4868 2602 5244
rect 2636 4868 2652 5244
rect 2586 4856 2652 4868
rect 2682 5244 2748 5256
rect 2682 4868 2698 5244
rect 2732 4868 2748 5244
rect 2682 4856 2748 4868
rect 2778 5244 2844 5256
rect 2778 4868 2794 5244
rect 2828 4868 2844 5244
rect 2778 4856 2844 4868
rect 2874 5244 2940 5256
rect 2874 4868 2890 5244
rect 2924 4868 2940 5244
rect 2874 4856 2940 4868
rect 2970 5244 3032 5256
rect 2970 4868 2986 5244
rect 3020 4868 3032 5244
rect 2970 4856 3032 4868
rect 2014 4626 2076 4638
rect 2014 4250 2026 4626
rect 2060 4250 2076 4626
rect 2014 4238 2076 4250
rect 2106 4626 2172 4638
rect 2106 4250 2122 4626
rect 2156 4250 2172 4626
rect 2106 4238 2172 4250
rect 2202 4626 2268 4638
rect 2202 4250 2218 4626
rect 2252 4250 2268 4626
rect 2202 4238 2268 4250
rect 2298 4626 2364 4638
rect 2298 4250 2314 4626
rect 2348 4250 2364 4626
rect 2298 4238 2364 4250
rect 2394 4626 2460 4638
rect 2394 4250 2410 4626
rect 2444 4250 2460 4626
rect 2394 4238 2460 4250
rect 2490 4626 2556 4638
rect 2490 4250 2506 4626
rect 2540 4250 2556 4626
rect 2490 4238 2556 4250
rect 2586 4626 2652 4638
rect 2586 4250 2602 4626
rect 2636 4250 2652 4626
rect 2586 4238 2652 4250
rect 2682 4626 2748 4638
rect 2682 4250 2698 4626
rect 2732 4250 2748 4626
rect 2682 4238 2748 4250
rect 2778 4626 2844 4638
rect 2778 4250 2794 4626
rect 2828 4250 2844 4626
rect 2778 4238 2844 4250
rect 2874 4626 2940 4638
rect 2874 4250 2890 4626
rect 2924 4250 2940 4626
rect 2874 4238 2940 4250
rect 2970 4626 3032 4638
rect 2970 4250 2986 4626
rect 3020 4250 3032 4626
rect 2970 4238 3032 4250
rect 3814 5862 3876 5874
rect 3814 5486 3826 5862
rect 3860 5486 3876 5862
rect 3814 5474 3876 5486
rect 3906 5862 3972 5874
rect 3906 5486 3922 5862
rect 3956 5486 3972 5862
rect 3906 5474 3972 5486
rect 4002 5862 4068 5874
rect 4002 5486 4018 5862
rect 4052 5486 4068 5862
rect 4002 5474 4068 5486
rect 4098 5862 4164 5874
rect 4098 5486 4114 5862
rect 4148 5486 4164 5862
rect 4098 5474 4164 5486
rect 4194 5862 4260 5874
rect 4194 5486 4210 5862
rect 4244 5486 4260 5862
rect 4194 5474 4260 5486
rect 4290 5862 4356 5874
rect 4290 5486 4306 5862
rect 4340 5486 4356 5862
rect 4290 5474 4356 5486
rect 4386 5862 4452 5874
rect 4386 5486 4402 5862
rect 4436 5486 4452 5862
rect 4386 5474 4452 5486
rect 4482 5862 4548 5874
rect 4482 5486 4498 5862
rect 4532 5486 4548 5862
rect 4482 5474 4548 5486
rect 4578 5862 4644 5874
rect 4578 5486 4594 5862
rect 4628 5486 4644 5862
rect 4578 5474 4644 5486
rect 4674 5862 4740 5874
rect 4674 5486 4690 5862
rect 4724 5486 4740 5862
rect 4674 5474 4740 5486
rect 4770 5862 4832 5874
rect 4770 5486 4786 5862
rect 4820 5486 4832 5862
rect 4770 5474 4832 5486
rect 3814 5244 3876 5256
rect 3814 4868 3826 5244
rect 3860 4868 3876 5244
rect 3814 4856 3876 4868
rect 3906 5244 3972 5256
rect 3906 4868 3922 5244
rect 3956 4868 3972 5244
rect 3906 4856 3972 4868
rect 4002 5244 4068 5256
rect 4002 4868 4018 5244
rect 4052 4868 4068 5244
rect 4002 4856 4068 4868
rect 4098 5244 4164 5256
rect 4098 4868 4114 5244
rect 4148 4868 4164 5244
rect 4098 4856 4164 4868
rect 4194 5244 4260 5256
rect 4194 4868 4210 5244
rect 4244 4868 4260 5244
rect 4194 4856 4260 4868
rect 4290 5244 4356 5256
rect 4290 4868 4306 5244
rect 4340 4868 4356 5244
rect 4290 4856 4356 4868
rect 4386 5244 4452 5256
rect 4386 4868 4402 5244
rect 4436 4868 4452 5244
rect 4386 4856 4452 4868
rect 4482 5244 4548 5256
rect 4482 4868 4498 5244
rect 4532 4868 4548 5244
rect 4482 4856 4548 4868
rect 4578 5244 4644 5256
rect 4578 4868 4594 5244
rect 4628 4868 4644 5244
rect 4578 4856 4644 4868
rect 4674 5244 4740 5256
rect 4674 4868 4690 5244
rect 4724 4868 4740 5244
rect 4674 4856 4740 4868
rect 4770 5244 4832 5256
rect 4770 4868 4786 5244
rect 4820 4868 4832 5244
rect 4770 4856 4832 4868
rect 3814 4626 3876 4638
rect 3814 4250 3826 4626
rect 3860 4250 3876 4626
rect 3814 4238 3876 4250
rect 3906 4626 3972 4638
rect 3906 4250 3922 4626
rect 3956 4250 3972 4626
rect 3906 4238 3972 4250
rect 4002 4626 4068 4638
rect 4002 4250 4018 4626
rect 4052 4250 4068 4626
rect 4002 4238 4068 4250
rect 4098 4626 4164 4638
rect 4098 4250 4114 4626
rect 4148 4250 4164 4626
rect 4098 4238 4164 4250
rect 4194 4626 4260 4638
rect 4194 4250 4210 4626
rect 4244 4250 4260 4626
rect 4194 4238 4260 4250
rect 4290 4626 4356 4638
rect 4290 4250 4306 4626
rect 4340 4250 4356 4626
rect 4290 4238 4356 4250
rect 4386 4626 4452 4638
rect 4386 4250 4402 4626
rect 4436 4250 4452 4626
rect 4386 4238 4452 4250
rect 4482 4626 4548 4638
rect 4482 4250 4498 4626
rect 4532 4250 4548 4626
rect 4482 4238 4548 4250
rect 4578 4626 4644 4638
rect 4578 4250 4594 4626
rect 4628 4250 4644 4626
rect 4578 4238 4644 4250
rect 4674 4626 4740 4638
rect 4674 4250 4690 4626
rect 4724 4250 4740 4626
rect 4674 4238 4740 4250
rect 4770 4626 4832 4638
rect 4770 4250 4786 4626
rect 4820 4250 4832 4626
rect 4770 4238 4832 4250
rect 5614 5862 5676 5874
rect 5614 5486 5626 5862
rect 5660 5486 5676 5862
rect 5614 5474 5676 5486
rect 5706 5862 5772 5874
rect 5706 5486 5722 5862
rect 5756 5486 5772 5862
rect 5706 5474 5772 5486
rect 5802 5862 5868 5874
rect 5802 5486 5818 5862
rect 5852 5486 5868 5862
rect 5802 5474 5868 5486
rect 5898 5862 5964 5874
rect 5898 5486 5914 5862
rect 5948 5486 5964 5862
rect 5898 5474 5964 5486
rect 5994 5862 6060 5874
rect 5994 5486 6010 5862
rect 6044 5486 6060 5862
rect 5994 5474 6060 5486
rect 6090 5862 6156 5874
rect 6090 5486 6106 5862
rect 6140 5486 6156 5862
rect 6090 5474 6156 5486
rect 6186 5862 6252 5874
rect 6186 5486 6202 5862
rect 6236 5486 6252 5862
rect 6186 5474 6252 5486
rect 6282 5862 6348 5874
rect 6282 5486 6298 5862
rect 6332 5486 6348 5862
rect 6282 5474 6348 5486
rect 6378 5862 6444 5874
rect 6378 5486 6394 5862
rect 6428 5486 6444 5862
rect 6378 5474 6444 5486
rect 6474 5862 6540 5874
rect 6474 5486 6490 5862
rect 6524 5486 6540 5862
rect 6474 5474 6540 5486
rect 6570 5862 6632 5874
rect 6570 5486 6586 5862
rect 6620 5486 6632 5862
rect 6570 5474 6632 5486
rect 5614 5244 5676 5256
rect 5614 4868 5626 5244
rect 5660 4868 5676 5244
rect 5614 4856 5676 4868
rect 5706 5244 5772 5256
rect 5706 4868 5722 5244
rect 5756 4868 5772 5244
rect 5706 4856 5772 4868
rect 5802 5244 5868 5256
rect 5802 4868 5818 5244
rect 5852 4868 5868 5244
rect 5802 4856 5868 4868
rect 5898 5244 5964 5256
rect 5898 4868 5914 5244
rect 5948 4868 5964 5244
rect 5898 4856 5964 4868
rect 5994 5244 6060 5256
rect 5994 4868 6010 5244
rect 6044 4868 6060 5244
rect 5994 4856 6060 4868
rect 6090 5244 6156 5256
rect 6090 4868 6106 5244
rect 6140 4868 6156 5244
rect 6090 4856 6156 4868
rect 6186 5244 6252 5256
rect 6186 4868 6202 5244
rect 6236 4868 6252 5244
rect 6186 4856 6252 4868
rect 6282 5244 6348 5256
rect 6282 4868 6298 5244
rect 6332 4868 6348 5244
rect 6282 4856 6348 4868
rect 6378 5244 6444 5256
rect 6378 4868 6394 5244
rect 6428 4868 6444 5244
rect 6378 4856 6444 4868
rect 6474 5244 6540 5256
rect 6474 4868 6490 5244
rect 6524 4868 6540 5244
rect 6474 4856 6540 4868
rect 6570 5244 6632 5256
rect 6570 4868 6586 5244
rect 6620 4868 6632 5244
rect 6570 4856 6632 4868
rect 5614 4626 5676 4638
rect 5614 4250 5626 4626
rect 5660 4250 5676 4626
rect 5614 4238 5676 4250
rect 5706 4626 5772 4638
rect 5706 4250 5722 4626
rect 5756 4250 5772 4626
rect 5706 4238 5772 4250
rect 5802 4626 5868 4638
rect 5802 4250 5818 4626
rect 5852 4250 5868 4626
rect 5802 4238 5868 4250
rect 5898 4626 5964 4638
rect 5898 4250 5914 4626
rect 5948 4250 5964 4626
rect 5898 4238 5964 4250
rect 5994 4626 6060 4638
rect 5994 4250 6010 4626
rect 6044 4250 6060 4626
rect 5994 4238 6060 4250
rect 6090 4626 6156 4638
rect 6090 4250 6106 4626
rect 6140 4250 6156 4626
rect 6090 4238 6156 4250
rect 6186 4626 6252 4638
rect 6186 4250 6202 4626
rect 6236 4250 6252 4626
rect 6186 4238 6252 4250
rect 6282 4626 6348 4638
rect 6282 4250 6298 4626
rect 6332 4250 6348 4626
rect 6282 4238 6348 4250
rect 6378 4626 6444 4638
rect 6378 4250 6394 4626
rect 6428 4250 6444 4626
rect 6378 4238 6444 4250
rect 6474 4626 6540 4638
rect 6474 4250 6490 4626
rect 6524 4250 6540 4626
rect 6474 4238 6540 4250
rect 6570 4626 6632 4638
rect 6570 4250 6586 4626
rect 6620 4250 6632 4626
rect 6570 4238 6632 4250
rect 7614 10250 7676 10262
rect 7614 9874 7626 10250
rect 7660 9874 7676 10250
rect 7614 9862 7676 9874
rect 7706 10250 7772 10262
rect 7706 9874 7722 10250
rect 7756 9874 7772 10250
rect 7706 9862 7772 9874
rect 7802 10250 7868 10262
rect 7802 9874 7818 10250
rect 7852 9874 7868 10250
rect 7802 9862 7868 9874
rect 7898 10250 7964 10262
rect 7898 9874 7914 10250
rect 7948 9874 7964 10250
rect 7898 9862 7964 9874
rect 7994 10250 8060 10262
rect 7994 9874 8010 10250
rect 8044 9874 8060 10250
rect 7994 9862 8060 9874
rect 8090 10250 8156 10262
rect 8090 9874 8106 10250
rect 8140 9874 8156 10250
rect 8090 9862 8156 9874
rect 8186 10250 8252 10262
rect 8186 9874 8202 10250
rect 8236 9874 8252 10250
rect 8186 9862 8252 9874
rect 8282 10250 8348 10262
rect 8282 9874 8298 10250
rect 8332 9874 8348 10250
rect 8282 9862 8348 9874
rect 8378 10250 8444 10262
rect 8378 9874 8394 10250
rect 8428 9874 8444 10250
rect 8378 9862 8444 9874
rect 8474 10250 8540 10262
rect 8474 9874 8490 10250
rect 8524 9874 8540 10250
rect 8474 9862 8540 9874
rect 8570 10250 8636 10262
rect 8570 9874 8586 10250
rect 8620 9874 8636 10250
rect 8570 9862 8636 9874
rect 8666 10250 8732 10262
rect 8666 9874 8682 10250
rect 8716 9874 8732 10250
rect 8666 9862 8732 9874
rect 8762 10250 8828 10262
rect 8762 9874 8778 10250
rect 8812 9874 8828 10250
rect 8762 9862 8828 9874
rect 8858 10250 8924 10262
rect 8858 9874 8874 10250
rect 8908 9874 8924 10250
rect 8858 9862 8924 9874
rect 8954 10250 9020 10262
rect 8954 9874 8970 10250
rect 9004 9874 9020 10250
rect 8954 9862 9020 9874
rect 9050 10250 9116 10262
rect 9050 9874 9066 10250
rect 9100 9874 9116 10250
rect 9050 9862 9116 9874
rect 9146 10250 9212 10262
rect 9146 9874 9162 10250
rect 9196 9874 9212 10250
rect 9146 9862 9212 9874
rect 9242 10250 9308 10262
rect 9242 9874 9258 10250
rect 9292 9874 9308 10250
rect 9242 9862 9308 9874
rect 9338 10250 9404 10262
rect 9338 9874 9354 10250
rect 9388 9874 9404 10250
rect 9338 9862 9404 9874
rect 9434 10250 9500 10262
rect 9434 9874 9450 10250
rect 9484 9874 9500 10250
rect 9434 9862 9500 9874
rect 9530 10250 9592 10262
rect 9530 9874 9546 10250
rect 9580 9874 9592 10250
rect 9530 9862 9592 9874
rect 7614 9632 7676 9644
rect 7614 9256 7626 9632
rect 7660 9256 7676 9632
rect 7614 9244 7676 9256
rect 7706 9632 7772 9644
rect 7706 9256 7722 9632
rect 7756 9256 7772 9632
rect 7706 9244 7772 9256
rect 7802 9632 7868 9644
rect 7802 9256 7818 9632
rect 7852 9256 7868 9632
rect 7802 9244 7868 9256
rect 7898 9632 7964 9644
rect 7898 9256 7914 9632
rect 7948 9256 7964 9632
rect 7898 9244 7964 9256
rect 7994 9632 8060 9644
rect 7994 9256 8010 9632
rect 8044 9256 8060 9632
rect 7994 9244 8060 9256
rect 8090 9632 8156 9644
rect 8090 9256 8106 9632
rect 8140 9256 8156 9632
rect 8090 9244 8156 9256
rect 8186 9632 8252 9644
rect 8186 9256 8202 9632
rect 8236 9256 8252 9632
rect 8186 9244 8252 9256
rect 8282 9632 8348 9644
rect 8282 9256 8298 9632
rect 8332 9256 8348 9632
rect 8282 9244 8348 9256
rect 8378 9632 8444 9644
rect 8378 9256 8394 9632
rect 8428 9256 8444 9632
rect 8378 9244 8444 9256
rect 8474 9632 8540 9644
rect 8474 9256 8490 9632
rect 8524 9256 8540 9632
rect 8474 9244 8540 9256
rect 8570 9632 8636 9644
rect 8570 9256 8586 9632
rect 8620 9256 8636 9632
rect 8570 9244 8636 9256
rect 8666 9632 8732 9644
rect 8666 9256 8682 9632
rect 8716 9256 8732 9632
rect 8666 9244 8732 9256
rect 8762 9632 8828 9644
rect 8762 9256 8778 9632
rect 8812 9256 8828 9632
rect 8762 9244 8828 9256
rect 8858 9632 8924 9644
rect 8858 9256 8874 9632
rect 8908 9256 8924 9632
rect 8858 9244 8924 9256
rect 8954 9632 9020 9644
rect 8954 9256 8970 9632
rect 9004 9256 9020 9632
rect 8954 9244 9020 9256
rect 9050 9632 9116 9644
rect 9050 9256 9066 9632
rect 9100 9256 9116 9632
rect 9050 9244 9116 9256
rect 9146 9632 9212 9644
rect 9146 9256 9162 9632
rect 9196 9256 9212 9632
rect 9146 9244 9212 9256
rect 9242 9632 9308 9644
rect 9242 9256 9258 9632
rect 9292 9256 9308 9632
rect 9242 9244 9308 9256
rect 9338 9632 9404 9644
rect 9338 9256 9354 9632
rect 9388 9256 9404 9632
rect 9338 9244 9404 9256
rect 9434 9632 9500 9644
rect 9434 9256 9450 9632
rect 9484 9256 9500 9632
rect 9434 9244 9500 9256
rect 9530 9632 9592 9644
rect 9530 9256 9546 9632
rect 9580 9256 9592 9632
rect 9530 9244 9592 9256
rect 7614 9014 7676 9026
rect 7614 8638 7626 9014
rect 7660 8638 7676 9014
rect 7614 8626 7676 8638
rect 7706 9014 7772 9026
rect 7706 8638 7722 9014
rect 7756 8638 7772 9014
rect 7706 8626 7772 8638
rect 7802 9014 7868 9026
rect 7802 8638 7818 9014
rect 7852 8638 7868 9014
rect 7802 8626 7868 8638
rect 7898 9014 7964 9026
rect 7898 8638 7914 9014
rect 7948 8638 7964 9014
rect 7898 8626 7964 8638
rect 7994 9014 8060 9026
rect 7994 8638 8010 9014
rect 8044 8638 8060 9014
rect 7994 8626 8060 8638
rect 8090 9014 8156 9026
rect 8090 8638 8106 9014
rect 8140 8638 8156 9014
rect 8090 8626 8156 8638
rect 8186 9014 8252 9026
rect 8186 8638 8202 9014
rect 8236 8638 8252 9014
rect 8186 8626 8252 8638
rect 8282 9014 8348 9026
rect 8282 8638 8298 9014
rect 8332 8638 8348 9014
rect 8282 8626 8348 8638
rect 8378 9014 8444 9026
rect 8378 8638 8394 9014
rect 8428 8638 8444 9014
rect 8378 8626 8444 8638
rect 8474 9014 8540 9026
rect 8474 8638 8490 9014
rect 8524 8638 8540 9014
rect 8474 8626 8540 8638
rect 8570 9014 8636 9026
rect 8570 8638 8586 9014
rect 8620 8638 8636 9014
rect 8570 8626 8636 8638
rect 8666 9014 8732 9026
rect 8666 8638 8682 9014
rect 8716 8638 8732 9014
rect 8666 8626 8732 8638
rect 8762 9014 8828 9026
rect 8762 8638 8778 9014
rect 8812 8638 8828 9014
rect 8762 8626 8828 8638
rect 8858 9014 8924 9026
rect 8858 8638 8874 9014
rect 8908 8638 8924 9014
rect 8858 8626 8924 8638
rect 8954 9014 9020 9026
rect 8954 8638 8970 9014
rect 9004 8638 9020 9014
rect 8954 8626 9020 8638
rect 9050 9014 9116 9026
rect 9050 8638 9066 9014
rect 9100 8638 9116 9014
rect 9050 8626 9116 8638
rect 9146 9014 9212 9026
rect 9146 8638 9162 9014
rect 9196 8638 9212 9014
rect 9146 8626 9212 8638
rect 9242 9014 9308 9026
rect 9242 8638 9258 9014
rect 9292 8638 9308 9014
rect 9242 8626 9308 8638
rect 9338 9014 9404 9026
rect 9338 8638 9354 9014
rect 9388 8638 9404 9014
rect 9338 8626 9404 8638
rect 9434 9014 9500 9026
rect 9434 8638 9450 9014
rect 9484 8638 9500 9014
rect 9434 8626 9500 8638
rect 9530 9014 9592 9026
rect 9530 8638 9546 9014
rect 9580 8638 9592 9014
rect 9530 8626 9592 8638
rect 7614 8396 7676 8408
rect 7614 8020 7626 8396
rect 7660 8020 7676 8396
rect 7614 8008 7676 8020
rect 7706 8396 7772 8408
rect 7706 8020 7722 8396
rect 7756 8020 7772 8396
rect 7706 8008 7772 8020
rect 7802 8396 7868 8408
rect 7802 8020 7818 8396
rect 7852 8020 7868 8396
rect 7802 8008 7868 8020
rect 7898 8396 7964 8408
rect 7898 8020 7914 8396
rect 7948 8020 7964 8396
rect 7898 8008 7964 8020
rect 7994 8396 8060 8408
rect 7994 8020 8010 8396
rect 8044 8020 8060 8396
rect 7994 8008 8060 8020
rect 8090 8396 8156 8408
rect 8090 8020 8106 8396
rect 8140 8020 8156 8396
rect 8090 8008 8156 8020
rect 8186 8396 8252 8408
rect 8186 8020 8202 8396
rect 8236 8020 8252 8396
rect 8186 8008 8252 8020
rect 8282 8396 8348 8408
rect 8282 8020 8298 8396
rect 8332 8020 8348 8396
rect 8282 8008 8348 8020
rect 8378 8396 8444 8408
rect 8378 8020 8394 8396
rect 8428 8020 8444 8396
rect 8378 8008 8444 8020
rect 8474 8396 8540 8408
rect 8474 8020 8490 8396
rect 8524 8020 8540 8396
rect 8474 8008 8540 8020
rect 8570 8396 8636 8408
rect 8570 8020 8586 8396
rect 8620 8020 8636 8396
rect 8570 8008 8636 8020
rect 8666 8396 8732 8408
rect 8666 8020 8682 8396
rect 8716 8020 8732 8396
rect 8666 8008 8732 8020
rect 8762 8396 8828 8408
rect 8762 8020 8778 8396
rect 8812 8020 8828 8396
rect 8762 8008 8828 8020
rect 8858 8396 8924 8408
rect 8858 8020 8874 8396
rect 8908 8020 8924 8396
rect 8858 8008 8924 8020
rect 8954 8396 9020 8408
rect 8954 8020 8970 8396
rect 9004 8020 9020 8396
rect 8954 8008 9020 8020
rect 9050 8396 9116 8408
rect 9050 8020 9066 8396
rect 9100 8020 9116 8396
rect 9050 8008 9116 8020
rect 9146 8396 9212 8408
rect 9146 8020 9162 8396
rect 9196 8020 9212 8396
rect 9146 8008 9212 8020
rect 9242 8396 9308 8408
rect 9242 8020 9258 8396
rect 9292 8020 9308 8396
rect 9242 8008 9308 8020
rect 9338 8396 9404 8408
rect 9338 8020 9354 8396
rect 9388 8020 9404 8396
rect 9338 8008 9404 8020
rect 9434 8396 9500 8408
rect 9434 8020 9450 8396
rect 9484 8020 9500 8396
rect 9434 8008 9500 8020
rect 9530 8396 9592 8408
rect 9530 8020 9546 8396
rect 9580 8020 9592 8396
rect 9530 8008 9592 8020
rect 7614 7778 7676 7790
rect 7614 7402 7626 7778
rect 7660 7402 7676 7778
rect 7614 7390 7676 7402
rect 7706 7778 7772 7790
rect 7706 7402 7722 7778
rect 7756 7402 7772 7778
rect 7706 7390 7772 7402
rect 7802 7778 7868 7790
rect 7802 7402 7818 7778
rect 7852 7402 7868 7778
rect 7802 7390 7868 7402
rect 7898 7778 7964 7790
rect 7898 7402 7914 7778
rect 7948 7402 7964 7778
rect 7898 7390 7964 7402
rect 7994 7778 8060 7790
rect 7994 7402 8010 7778
rect 8044 7402 8060 7778
rect 7994 7390 8060 7402
rect 8090 7778 8156 7790
rect 8090 7402 8106 7778
rect 8140 7402 8156 7778
rect 8090 7390 8156 7402
rect 8186 7778 8252 7790
rect 8186 7402 8202 7778
rect 8236 7402 8252 7778
rect 8186 7390 8252 7402
rect 8282 7778 8348 7790
rect 8282 7402 8298 7778
rect 8332 7402 8348 7778
rect 8282 7390 8348 7402
rect 8378 7778 8444 7790
rect 8378 7402 8394 7778
rect 8428 7402 8444 7778
rect 8378 7390 8444 7402
rect 8474 7778 8540 7790
rect 8474 7402 8490 7778
rect 8524 7402 8540 7778
rect 8474 7390 8540 7402
rect 8570 7778 8636 7790
rect 8570 7402 8586 7778
rect 8620 7402 8636 7778
rect 8570 7390 8636 7402
rect 8666 7778 8732 7790
rect 8666 7402 8682 7778
rect 8716 7402 8732 7778
rect 8666 7390 8732 7402
rect 8762 7778 8828 7790
rect 8762 7402 8778 7778
rect 8812 7402 8828 7778
rect 8762 7390 8828 7402
rect 8858 7778 8924 7790
rect 8858 7402 8874 7778
rect 8908 7402 8924 7778
rect 8858 7390 8924 7402
rect 8954 7778 9020 7790
rect 8954 7402 8970 7778
rect 9004 7402 9020 7778
rect 8954 7390 9020 7402
rect 9050 7778 9116 7790
rect 9050 7402 9066 7778
rect 9100 7402 9116 7778
rect 9050 7390 9116 7402
rect 9146 7778 9212 7790
rect 9146 7402 9162 7778
rect 9196 7402 9212 7778
rect 9146 7390 9212 7402
rect 9242 7778 9308 7790
rect 9242 7402 9258 7778
rect 9292 7402 9308 7778
rect 9242 7390 9308 7402
rect 9338 7778 9404 7790
rect 9338 7402 9354 7778
rect 9388 7402 9404 7778
rect 9338 7390 9404 7402
rect 9434 7778 9500 7790
rect 9434 7402 9450 7778
rect 9484 7402 9500 7778
rect 9434 7390 9500 7402
rect 9530 7778 9592 7790
rect 9530 7402 9546 7778
rect 9580 7402 9592 7778
rect 9530 7390 9592 7402
rect 7614 7160 7676 7172
rect 7614 6784 7626 7160
rect 7660 6784 7676 7160
rect 7614 6772 7676 6784
rect 7706 7160 7772 7172
rect 7706 6784 7722 7160
rect 7756 6784 7772 7160
rect 7706 6772 7772 6784
rect 7802 7160 7868 7172
rect 7802 6784 7818 7160
rect 7852 6784 7868 7160
rect 7802 6772 7868 6784
rect 7898 7160 7964 7172
rect 7898 6784 7914 7160
rect 7948 6784 7964 7160
rect 7898 6772 7964 6784
rect 7994 7160 8060 7172
rect 7994 6784 8010 7160
rect 8044 6784 8060 7160
rect 7994 6772 8060 6784
rect 8090 7160 8156 7172
rect 8090 6784 8106 7160
rect 8140 6784 8156 7160
rect 8090 6772 8156 6784
rect 8186 7160 8252 7172
rect 8186 6784 8202 7160
rect 8236 6784 8252 7160
rect 8186 6772 8252 6784
rect 8282 7160 8348 7172
rect 8282 6784 8298 7160
rect 8332 6784 8348 7160
rect 8282 6772 8348 6784
rect 8378 7160 8444 7172
rect 8378 6784 8394 7160
rect 8428 6784 8444 7160
rect 8378 6772 8444 6784
rect 8474 7160 8540 7172
rect 8474 6784 8490 7160
rect 8524 6784 8540 7160
rect 8474 6772 8540 6784
rect 8570 7160 8636 7172
rect 8570 6784 8586 7160
rect 8620 6784 8636 7160
rect 8570 6772 8636 6784
rect 8666 7160 8732 7172
rect 8666 6784 8682 7160
rect 8716 6784 8732 7160
rect 8666 6772 8732 6784
rect 8762 7160 8828 7172
rect 8762 6784 8778 7160
rect 8812 6784 8828 7160
rect 8762 6772 8828 6784
rect 8858 7160 8924 7172
rect 8858 6784 8874 7160
rect 8908 6784 8924 7160
rect 8858 6772 8924 6784
rect 8954 7160 9020 7172
rect 8954 6784 8970 7160
rect 9004 6784 9020 7160
rect 8954 6772 9020 6784
rect 9050 7160 9116 7172
rect 9050 6784 9066 7160
rect 9100 6784 9116 7160
rect 9050 6772 9116 6784
rect 9146 7160 9212 7172
rect 9146 6784 9162 7160
rect 9196 6784 9212 7160
rect 9146 6772 9212 6784
rect 9242 7160 9308 7172
rect 9242 6784 9258 7160
rect 9292 6784 9308 7160
rect 9242 6772 9308 6784
rect 9338 7160 9404 7172
rect 9338 6784 9354 7160
rect 9388 6784 9404 7160
rect 9338 6772 9404 6784
rect 9434 7160 9500 7172
rect 9434 6784 9450 7160
rect 9484 6784 9500 7160
rect 9434 6772 9500 6784
rect 9530 7160 9592 7172
rect 9530 6784 9546 7160
rect 9580 6784 9592 7160
rect 9530 6772 9592 6784
rect 7614 6542 7676 6554
rect 7614 6166 7626 6542
rect 7660 6166 7676 6542
rect 7614 6154 7676 6166
rect 7706 6542 7772 6554
rect 7706 6166 7722 6542
rect 7756 6166 7772 6542
rect 7706 6154 7772 6166
rect 7802 6542 7868 6554
rect 7802 6166 7818 6542
rect 7852 6166 7868 6542
rect 7802 6154 7868 6166
rect 7898 6542 7964 6554
rect 7898 6166 7914 6542
rect 7948 6166 7964 6542
rect 7898 6154 7964 6166
rect 7994 6542 8060 6554
rect 7994 6166 8010 6542
rect 8044 6166 8060 6542
rect 7994 6154 8060 6166
rect 8090 6542 8156 6554
rect 8090 6166 8106 6542
rect 8140 6166 8156 6542
rect 8090 6154 8156 6166
rect 8186 6542 8252 6554
rect 8186 6166 8202 6542
rect 8236 6166 8252 6542
rect 8186 6154 8252 6166
rect 8282 6542 8348 6554
rect 8282 6166 8298 6542
rect 8332 6166 8348 6542
rect 8282 6154 8348 6166
rect 8378 6542 8444 6554
rect 8378 6166 8394 6542
rect 8428 6166 8444 6542
rect 8378 6154 8444 6166
rect 8474 6542 8540 6554
rect 8474 6166 8490 6542
rect 8524 6166 8540 6542
rect 8474 6154 8540 6166
rect 8570 6542 8636 6554
rect 8570 6166 8586 6542
rect 8620 6166 8636 6542
rect 8570 6154 8636 6166
rect 8666 6542 8732 6554
rect 8666 6166 8682 6542
rect 8716 6166 8732 6542
rect 8666 6154 8732 6166
rect 8762 6542 8828 6554
rect 8762 6166 8778 6542
rect 8812 6166 8828 6542
rect 8762 6154 8828 6166
rect 8858 6542 8924 6554
rect 8858 6166 8874 6542
rect 8908 6166 8924 6542
rect 8858 6154 8924 6166
rect 8954 6542 9020 6554
rect 8954 6166 8970 6542
rect 9004 6166 9020 6542
rect 8954 6154 9020 6166
rect 9050 6542 9116 6554
rect 9050 6166 9066 6542
rect 9100 6166 9116 6542
rect 9050 6154 9116 6166
rect 9146 6542 9212 6554
rect 9146 6166 9162 6542
rect 9196 6166 9212 6542
rect 9146 6154 9212 6166
rect 9242 6542 9308 6554
rect 9242 6166 9258 6542
rect 9292 6166 9308 6542
rect 9242 6154 9308 6166
rect 9338 6542 9404 6554
rect 9338 6166 9354 6542
rect 9388 6166 9404 6542
rect 9338 6154 9404 6166
rect 9434 6542 9500 6554
rect 9434 6166 9450 6542
rect 9484 6166 9500 6542
rect 9434 6154 9500 6166
rect 9530 6542 9592 6554
rect 9530 6166 9546 6542
rect 9580 6166 9592 6542
rect 9530 6154 9592 6166
rect 7614 5924 7676 5936
rect 7614 5548 7626 5924
rect 7660 5548 7676 5924
rect 7614 5536 7676 5548
rect 7706 5924 7772 5936
rect 7706 5548 7722 5924
rect 7756 5548 7772 5924
rect 7706 5536 7772 5548
rect 7802 5924 7868 5936
rect 7802 5548 7818 5924
rect 7852 5548 7868 5924
rect 7802 5536 7868 5548
rect 7898 5924 7964 5936
rect 7898 5548 7914 5924
rect 7948 5548 7964 5924
rect 7898 5536 7964 5548
rect 7994 5924 8060 5936
rect 7994 5548 8010 5924
rect 8044 5548 8060 5924
rect 7994 5536 8060 5548
rect 8090 5924 8156 5936
rect 8090 5548 8106 5924
rect 8140 5548 8156 5924
rect 8090 5536 8156 5548
rect 8186 5924 8252 5936
rect 8186 5548 8202 5924
rect 8236 5548 8252 5924
rect 8186 5536 8252 5548
rect 8282 5924 8348 5936
rect 8282 5548 8298 5924
rect 8332 5548 8348 5924
rect 8282 5536 8348 5548
rect 8378 5924 8444 5936
rect 8378 5548 8394 5924
rect 8428 5548 8444 5924
rect 8378 5536 8444 5548
rect 8474 5924 8540 5936
rect 8474 5548 8490 5924
rect 8524 5548 8540 5924
rect 8474 5536 8540 5548
rect 8570 5924 8636 5936
rect 8570 5548 8586 5924
rect 8620 5548 8636 5924
rect 8570 5536 8636 5548
rect 8666 5924 8732 5936
rect 8666 5548 8682 5924
rect 8716 5548 8732 5924
rect 8666 5536 8732 5548
rect 8762 5924 8828 5936
rect 8762 5548 8778 5924
rect 8812 5548 8828 5924
rect 8762 5536 8828 5548
rect 8858 5924 8924 5936
rect 8858 5548 8874 5924
rect 8908 5548 8924 5924
rect 8858 5536 8924 5548
rect 8954 5924 9020 5936
rect 8954 5548 8970 5924
rect 9004 5548 9020 5924
rect 8954 5536 9020 5548
rect 9050 5924 9116 5936
rect 9050 5548 9066 5924
rect 9100 5548 9116 5924
rect 9050 5536 9116 5548
rect 9146 5924 9212 5936
rect 9146 5548 9162 5924
rect 9196 5548 9212 5924
rect 9146 5536 9212 5548
rect 9242 5924 9308 5936
rect 9242 5548 9258 5924
rect 9292 5548 9308 5924
rect 9242 5536 9308 5548
rect 9338 5924 9404 5936
rect 9338 5548 9354 5924
rect 9388 5548 9404 5924
rect 9338 5536 9404 5548
rect 9434 5924 9500 5936
rect 9434 5548 9450 5924
rect 9484 5548 9500 5924
rect 9434 5536 9500 5548
rect 9530 5924 9592 5936
rect 9530 5548 9546 5924
rect 9580 5548 9592 5924
rect 9530 5536 9592 5548
rect 7614 5306 7676 5318
rect 7614 4930 7626 5306
rect 7660 4930 7676 5306
rect 7614 4918 7676 4930
rect 7706 5306 7772 5318
rect 7706 4930 7722 5306
rect 7756 4930 7772 5306
rect 7706 4918 7772 4930
rect 7802 5306 7868 5318
rect 7802 4930 7818 5306
rect 7852 4930 7868 5306
rect 7802 4918 7868 4930
rect 7898 5306 7964 5318
rect 7898 4930 7914 5306
rect 7948 4930 7964 5306
rect 7898 4918 7964 4930
rect 7994 5306 8060 5318
rect 7994 4930 8010 5306
rect 8044 4930 8060 5306
rect 7994 4918 8060 4930
rect 8090 5306 8156 5318
rect 8090 4930 8106 5306
rect 8140 4930 8156 5306
rect 8090 4918 8156 4930
rect 8186 5306 8252 5318
rect 8186 4930 8202 5306
rect 8236 4930 8252 5306
rect 8186 4918 8252 4930
rect 8282 5306 8348 5318
rect 8282 4930 8298 5306
rect 8332 4930 8348 5306
rect 8282 4918 8348 4930
rect 8378 5306 8444 5318
rect 8378 4930 8394 5306
rect 8428 4930 8444 5306
rect 8378 4918 8444 4930
rect 8474 5306 8540 5318
rect 8474 4930 8490 5306
rect 8524 4930 8540 5306
rect 8474 4918 8540 4930
rect 8570 5306 8636 5318
rect 8570 4930 8586 5306
rect 8620 4930 8636 5306
rect 8570 4918 8636 4930
rect 8666 5306 8732 5318
rect 8666 4930 8682 5306
rect 8716 4930 8732 5306
rect 8666 4918 8732 4930
rect 8762 5306 8828 5318
rect 8762 4930 8778 5306
rect 8812 4930 8828 5306
rect 8762 4918 8828 4930
rect 8858 5306 8924 5318
rect 8858 4930 8874 5306
rect 8908 4930 8924 5306
rect 8858 4918 8924 4930
rect 8954 5306 9020 5318
rect 8954 4930 8970 5306
rect 9004 4930 9020 5306
rect 8954 4918 9020 4930
rect 9050 5306 9116 5318
rect 9050 4930 9066 5306
rect 9100 4930 9116 5306
rect 9050 4918 9116 4930
rect 9146 5306 9212 5318
rect 9146 4930 9162 5306
rect 9196 4930 9212 5306
rect 9146 4918 9212 4930
rect 9242 5306 9308 5318
rect 9242 4930 9258 5306
rect 9292 4930 9308 5306
rect 9242 4918 9308 4930
rect 9338 5306 9404 5318
rect 9338 4930 9354 5306
rect 9388 4930 9404 5306
rect 9338 4918 9404 4930
rect 9434 5306 9500 5318
rect 9434 4930 9450 5306
rect 9484 4930 9500 5306
rect 9434 4918 9500 4930
rect 9530 5306 9592 5318
rect 9530 4930 9546 5306
rect 9580 4930 9592 5306
rect 9530 4918 9592 4930
rect 16078 8718 16140 8730
rect 16078 8342 16090 8718
rect 16124 8342 16140 8718
rect 16078 8330 16140 8342
rect 16170 8718 16236 8730
rect 16170 8342 16186 8718
rect 16220 8342 16236 8718
rect 16170 8330 16236 8342
rect 16266 8718 16332 8730
rect 16266 8342 16282 8718
rect 16316 8342 16332 8718
rect 16266 8330 16332 8342
rect 16362 8718 16428 8730
rect 16362 8342 16378 8718
rect 16412 8342 16428 8718
rect 16362 8330 16428 8342
rect 16458 8718 16524 8730
rect 16458 8342 16474 8718
rect 16508 8342 16524 8718
rect 16458 8330 16524 8342
rect 16554 8718 16620 8730
rect 16554 8342 16570 8718
rect 16604 8342 16620 8718
rect 16554 8330 16620 8342
rect 16650 8718 16716 8730
rect 16650 8342 16666 8718
rect 16700 8342 16716 8718
rect 16650 8330 16716 8342
rect 16746 8718 16812 8730
rect 16746 8342 16762 8718
rect 16796 8342 16812 8718
rect 16746 8330 16812 8342
rect 16842 8718 16908 8730
rect 16842 8342 16858 8718
rect 16892 8342 16908 8718
rect 16842 8330 16908 8342
rect 16938 8718 17004 8730
rect 16938 8342 16954 8718
rect 16988 8342 17004 8718
rect 16938 8330 17004 8342
rect 17034 8718 17100 8730
rect 17034 8342 17050 8718
rect 17084 8342 17100 8718
rect 17034 8330 17100 8342
rect 17130 8718 17196 8730
rect 17130 8342 17146 8718
rect 17180 8342 17196 8718
rect 17130 8330 17196 8342
rect 17226 8718 17292 8730
rect 17226 8342 17242 8718
rect 17276 8342 17292 8718
rect 17226 8330 17292 8342
rect 17322 8718 17388 8730
rect 17322 8342 17338 8718
rect 17372 8342 17388 8718
rect 17322 8330 17388 8342
rect 17418 8718 17484 8730
rect 17418 8342 17434 8718
rect 17468 8342 17484 8718
rect 17418 8330 17484 8342
rect 17514 8718 17580 8730
rect 17514 8342 17530 8718
rect 17564 8342 17580 8718
rect 17514 8330 17580 8342
rect 17610 8718 17676 8730
rect 17610 8342 17626 8718
rect 17660 8342 17676 8718
rect 17610 8330 17676 8342
rect 17706 8718 17772 8730
rect 17706 8342 17722 8718
rect 17756 8342 17772 8718
rect 17706 8330 17772 8342
rect 17802 8718 17868 8730
rect 17802 8342 17818 8718
rect 17852 8342 17868 8718
rect 17802 8330 17868 8342
rect 17898 8718 17964 8730
rect 17898 8342 17914 8718
rect 17948 8342 17964 8718
rect 17898 8330 17964 8342
rect 17994 8718 18056 8730
rect 17994 8342 18010 8718
rect 18044 8342 18056 8718
rect 17994 8330 18056 8342
rect 16078 7898 16140 7910
rect 16078 7522 16090 7898
rect 16124 7522 16140 7898
rect 16078 7510 16140 7522
rect 16170 7898 16236 7910
rect 16170 7522 16186 7898
rect 16220 7522 16236 7898
rect 16170 7510 16236 7522
rect 16266 7898 16332 7910
rect 16266 7522 16282 7898
rect 16316 7522 16332 7898
rect 16266 7510 16332 7522
rect 16362 7898 16428 7910
rect 16362 7522 16378 7898
rect 16412 7522 16428 7898
rect 16362 7510 16428 7522
rect 16458 7898 16524 7910
rect 16458 7522 16474 7898
rect 16508 7522 16524 7898
rect 16458 7510 16524 7522
rect 16554 7898 16620 7910
rect 16554 7522 16570 7898
rect 16604 7522 16620 7898
rect 16554 7510 16620 7522
rect 16650 7898 16716 7910
rect 16650 7522 16666 7898
rect 16700 7522 16716 7898
rect 16650 7510 16716 7522
rect 16746 7898 16812 7910
rect 16746 7522 16762 7898
rect 16796 7522 16812 7898
rect 16746 7510 16812 7522
rect 16842 7898 16908 7910
rect 16842 7522 16858 7898
rect 16892 7522 16908 7898
rect 16842 7510 16908 7522
rect 16938 7898 17004 7910
rect 16938 7522 16954 7898
rect 16988 7522 17004 7898
rect 16938 7510 17004 7522
rect 17034 7898 17100 7910
rect 17034 7522 17050 7898
rect 17084 7522 17100 7898
rect 17034 7510 17100 7522
rect 17130 7898 17196 7910
rect 17130 7522 17146 7898
rect 17180 7522 17196 7898
rect 17130 7510 17196 7522
rect 17226 7898 17292 7910
rect 17226 7522 17242 7898
rect 17276 7522 17292 7898
rect 17226 7510 17292 7522
rect 17322 7898 17388 7910
rect 17322 7522 17338 7898
rect 17372 7522 17388 7898
rect 17322 7510 17388 7522
rect 17418 7898 17484 7910
rect 17418 7522 17434 7898
rect 17468 7522 17484 7898
rect 17418 7510 17484 7522
rect 17514 7898 17580 7910
rect 17514 7522 17530 7898
rect 17564 7522 17580 7898
rect 17514 7510 17580 7522
rect 17610 7898 17676 7910
rect 17610 7522 17626 7898
rect 17660 7522 17676 7898
rect 17610 7510 17676 7522
rect 17706 7898 17772 7910
rect 17706 7522 17722 7898
rect 17756 7522 17772 7898
rect 17706 7510 17772 7522
rect 17802 7898 17868 7910
rect 17802 7522 17818 7898
rect 17852 7522 17868 7898
rect 17802 7510 17868 7522
rect 17898 7898 17964 7910
rect 17898 7522 17914 7898
rect 17948 7522 17964 7898
rect 17898 7510 17964 7522
rect 17994 7898 18056 7910
rect 17994 7522 18010 7898
rect 18044 7522 18056 7898
rect 17994 7510 18056 7522
rect 16078 7078 16140 7090
rect 16078 6702 16090 7078
rect 16124 6702 16140 7078
rect 16078 6690 16140 6702
rect 16170 7078 16236 7090
rect 16170 6702 16186 7078
rect 16220 6702 16236 7078
rect 16170 6690 16236 6702
rect 16266 7078 16332 7090
rect 16266 6702 16282 7078
rect 16316 6702 16332 7078
rect 16266 6690 16332 6702
rect 16362 7078 16428 7090
rect 16362 6702 16378 7078
rect 16412 6702 16428 7078
rect 16362 6690 16428 6702
rect 16458 7078 16524 7090
rect 16458 6702 16474 7078
rect 16508 6702 16524 7078
rect 16458 6690 16524 6702
rect 16554 7078 16620 7090
rect 16554 6702 16570 7078
rect 16604 6702 16620 7078
rect 16554 6690 16620 6702
rect 16650 7078 16716 7090
rect 16650 6702 16666 7078
rect 16700 6702 16716 7078
rect 16650 6690 16716 6702
rect 16746 7078 16812 7090
rect 16746 6702 16762 7078
rect 16796 6702 16812 7078
rect 16746 6690 16812 6702
rect 16842 7078 16908 7090
rect 16842 6702 16858 7078
rect 16892 6702 16908 7078
rect 16842 6690 16908 6702
rect 16938 7078 17004 7090
rect 16938 6702 16954 7078
rect 16988 6702 17004 7078
rect 16938 6690 17004 6702
rect 17034 7078 17100 7090
rect 17034 6702 17050 7078
rect 17084 6702 17100 7078
rect 17034 6690 17100 6702
rect 17130 7078 17196 7090
rect 17130 6702 17146 7078
rect 17180 6702 17196 7078
rect 17130 6690 17196 6702
rect 17226 7078 17292 7090
rect 17226 6702 17242 7078
rect 17276 6702 17292 7078
rect 17226 6690 17292 6702
rect 17322 7078 17388 7090
rect 17322 6702 17338 7078
rect 17372 6702 17388 7078
rect 17322 6690 17388 6702
rect 17418 7078 17484 7090
rect 17418 6702 17434 7078
rect 17468 6702 17484 7078
rect 17418 6690 17484 6702
rect 17514 7078 17580 7090
rect 17514 6702 17530 7078
rect 17564 6702 17580 7078
rect 17514 6690 17580 6702
rect 17610 7078 17676 7090
rect 17610 6702 17626 7078
rect 17660 6702 17676 7078
rect 17610 6690 17676 6702
rect 17706 7078 17772 7090
rect 17706 6702 17722 7078
rect 17756 6702 17772 7078
rect 17706 6690 17772 6702
rect 17802 7078 17868 7090
rect 17802 6702 17818 7078
rect 17852 6702 17868 7078
rect 17802 6690 17868 6702
rect 17898 7078 17964 7090
rect 17898 6702 17914 7078
rect 17948 6702 17964 7078
rect 17898 6690 17964 6702
rect 17994 7078 18056 7090
rect 17994 6702 18010 7078
rect 18044 6702 18056 7078
rect 17994 6690 18056 6702
rect 19514 8684 19576 8696
rect 19514 8308 19526 8684
rect 19560 8308 19576 8684
rect 19514 8296 19576 8308
rect 19606 8684 19672 8696
rect 19606 8308 19622 8684
rect 19656 8308 19672 8684
rect 19606 8296 19672 8308
rect 19702 8684 19768 8696
rect 19702 8308 19718 8684
rect 19752 8308 19768 8684
rect 19702 8296 19768 8308
rect 19798 8684 19864 8696
rect 19798 8308 19814 8684
rect 19848 8308 19864 8684
rect 19798 8296 19864 8308
rect 19894 8684 19960 8696
rect 19894 8308 19910 8684
rect 19944 8308 19960 8684
rect 19894 8296 19960 8308
rect 19990 8684 20056 8696
rect 19990 8308 20006 8684
rect 20040 8308 20056 8684
rect 19990 8296 20056 8308
rect 20086 8684 20152 8696
rect 20086 8308 20102 8684
rect 20136 8308 20152 8684
rect 20086 8296 20152 8308
rect 20182 8684 20248 8696
rect 20182 8308 20198 8684
rect 20232 8308 20248 8684
rect 20182 8296 20248 8308
rect 20278 8684 20344 8696
rect 20278 8308 20294 8684
rect 20328 8308 20344 8684
rect 20278 8296 20344 8308
rect 20374 8684 20440 8696
rect 20374 8308 20390 8684
rect 20424 8308 20440 8684
rect 20374 8296 20440 8308
rect 20470 8684 20536 8696
rect 20470 8308 20486 8684
rect 20520 8308 20536 8684
rect 20470 8296 20536 8308
rect 20566 8684 20632 8696
rect 20566 8308 20582 8684
rect 20616 8308 20632 8684
rect 20566 8296 20632 8308
rect 20662 8684 20728 8696
rect 20662 8308 20678 8684
rect 20712 8308 20728 8684
rect 20662 8296 20728 8308
rect 20758 8684 20824 8696
rect 20758 8308 20774 8684
rect 20808 8308 20824 8684
rect 20758 8296 20824 8308
rect 20854 8684 20920 8696
rect 20854 8308 20870 8684
rect 20904 8308 20920 8684
rect 20854 8296 20920 8308
rect 20950 8684 21016 8696
rect 20950 8308 20966 8684
rect 21000 8308 21016 8684
rect 20950 8296 21016 8308
rect 21046 8684 21112 8696
rect 21046 8308 21062 8684
rect 21096 8308 21112 8684
rect 21046 8296 21112 8308
rect 21142 8684 21208 8696
rect 21142 8308 21158 8684
rect 21192 8308 21208 8684
rect 21142 8296 21208 8308
rect 21238 8684 21304 8696
rect 21238 8308 21254 8684
rect 21288 8308 21304 8684
rect 21238 8296 21304 8308
rect 21334 8684 21400 8696
rect 21334 8308 21350 8684
rect 21384 8308 21400 8684
rect 21334 8296 21400 8308
rect 21430 8684 21492 8696
rect 21430 8308 21446 8684
rect 21480 8308 21492 8684
rect 21430 8296 21492 8308
rect 19514 8066 19576 8078
rect 19514 7690 19526 8066
rect 19560 7690 19576 8066
rect 19514 7678 19576 7690
rect 19606 8066 19672 8078
rect 19606 7690 19622 8066
rect 19656 7690 19672 8066
rect 19606 7678 19672 7690
rect 19702 8066 19768 8078
rect 19702 7690 19718 8066
rect 19752 7690 19768 8066
rect 19702 7678 19768 7690
rect 19798 8066 19864 8078
rect 19798 7690 19814 8066
rect 19848 7690 19864 8066
rect 19798 7678 19864 7690
rect 19894 8066 19960 8078
rect 19894 7690 19910 8066
rect 19944 7690 19960 8066
rect 19894 7678 19960 7690
rect 19990 8066 20056 8078
rect 19990 7690 20006 8066
rect 20040 7690 20056 8066
rect 19990 7678 20056 7690
rect 20086 8066 20152 8078
rect 20086 7690 20102 8066
rect 20136 7690 20152 8066
rect 20086 7678 20152 7690
rect 20182 8066 20248 8078
rect 20182 7690 20198 8066
rect 20232 7690 20248 8066
rect 20182 7678 20248 7690
rect 20278 8066 20344 8078
rect 20278 7690 20294 8066
rect 20328 7690 20344 8066
rect 20278 7678 20344 7690
rect 20374 8066 20440 8078
rect 20374 7690 20390 8066
rect 20424 7690 20440 8066
rect 20374 7678 20440 7690
rect 20470 8066 20536 8078
rect 20470 7690 20486 8066
rect 20520 7690 20536 8066
rect 20470 7678 20536 7690
rect 20566 8066 20632 8078
rect 20566 7690 20582 8066
rect 20616 7690 20632 8066
rect 20566 7678 20632 7690
rect 20662 8066 20728 8078
rect 20662 7690 20678 8066
rect 20712 7690 20728 8066
rect 20662 7678 20728 7690
rect 20758 8066 20824 8078
rect 20758 7690 20774 8066
rect 20808 7690 20824 8066
rect 20758 7678 20824 7690
rect 20854 8066 20920 8078
rect 20854 7690 20870 8066
rect 20904 7690 20920 8066
rect 20854 7678 20920 7690
rect 20950 8066 21016 8078
rect 20950 7690 20966 8066
rect 21000 7690 21016 8066
rect 20950 7678 21016 7690
rect 21046 8066 21112 8078
rect 21046 7690 21062 8066
rect 21096 7690 21112 8066
rect 21046 7678 21112 7690
rect 21142 8066 21208 8078
rect 21142 7690 21158 8066
rect 21192 7690 21208 8066
rect 21142 7678 21208 7690
rect 21238 8066 21304 8078
rect 21238 7690 21254 8066
rect 21288 7690 21304 8066
rect 21238 7678 21304 7690
rect 21334 8066 21400 8078
rect 21334 7690 21350 8066
rect 21384 7690 21400 8066
rect 21334 7678 21400 7690
rect 21430 8066 21492 8078
rect 21430 7690 21446 8066
rect 21480 7690 21492 8066
rect 21430 7678 21492 7690
rect 14614 5862 14676 5874
rect 14614 5486 14626 5862
rect 14660 5486 14676 5862
rect 14614 5474 14676 5486
rect 14706 5862 14772 5874
rect 14706 5486 14722 5862
rect 14756 5486 14772 5862
rect 14706 5474 14772 5486
rect 14802 5862 14868 5874
rect 14802 5486 14818 5862
rect 14852 5486 14868 5862
rect 14802 5474 14868 5486
rect 14898 5862 14964 5874
rect 14898 5486 14914 5862
rect 14948 5486 14964 5862
rect 14898 5474 14964 5486
rect 14994 5862 15060 5874
rect 14994 5486 15010 5862
rect 15044 5486 15060 5862
rect 14994 5474 15060 5486
rect 15090 5862 15156 5874
rect 15090 5486 15106 5862
rect 15140 5486 15156 5862
rect 15090 5474 15156 5486
rect 15186 5862 15252 5874
rect 15186 5486 15202 5862
rect 15236 5486 15252 5862
rect 15186 5474 15252 5486
rect 15282 5862 15348 5874
rect 15282 5486 15298 5862
rect 15332 5486 15348 5862
rect 15282 5474 15348 5486
rect 15378 5862 15444 5874
rect 15378 5486 15394 5862
rect 15428 5486 15444 5862
rect 15378 5474 15444 5486
rect 15474 5862 15540 5874
rect 15474 5486 15490 5862
rect 15524 5486 15540 5862
rect 15474 5474 15540 5486
rect 15570 5862 15632 5874
rect 15570 5486 15586 5862
rect 15620 5486 15632 5862
rect 15570 5474 15632 5486
rect 14614 5244 14676 5256
rect 14614 4868 14626 5244
rect 14660 4868 14676 5244
rect 14614 4856 14676 4868
rect 14706 5244 14772 5256
rect 14706 4868 14722 5244
rect 14756 4868 14772 5244
rect 14706 4856 14772 4868
rect 14802 5244 14868 5256
rect 14802 4868 14818 5244
rect 14852 4868 14868 5244
rect 14802 4856 14868 4868
rect 14898 5244 14964 5256
rect 14898 4868 14914 5244
rect 14948 4868 14964 5244
rect 14898 4856 14964 4868
rect 14994 5244 15060 5256
rect 14994 4868 15010 5244
rect 15044 4868 15060 5244
rect 14994 4856 15060 4868
rect 15090 5244 15156 5256
rect 15090 4868 15106 5244
rect 15140 4868 15156 5244
rect 15090 4856 15156 4868
rect 15186 5244 15252 5256
rect 15186 4868 15202 5244
rect 15236 4868 15252 5244
rect 15186 4856 15252 4868
rect 15282 5244 15348 5256
rect 15282 4868 15298 5244
rect 15332 4868 15348 5244
rect 15282 4856 15348 4868
rect 15378 5244 15444 5256
rect 15378 4868 15394 5244
rect 15428 4868 15444 5244
rect 15378 4856 15444 4868
rect 15474 5244 15540 5256
rect 15474 4868 15490 5244
rect 15524 4868 15540 5244
rect 15474 4856 15540 4868
rect 15570 5244 15632 5256
rect 15570 4868 15586 5244
rect 15620 4868 15632 5244
rect 15570 4856 15632 4868
rect 14614 4626 14676 4638
rect 14614 4250 14626 4626
rect 14660 4250 14676 4626
rect 14614 4238 14676 4250
rect 14706 4626 14772 4638
rect 14706 4250 14722 4626
rect 14756 4250 14772 4626
rect 14706 4238 14772 4250
rect 14802 4626 14868 4638
rect 14802 4250 14818 4626
rect 14852 4250 14868 4626
rect 14802 4238 14868 4250
rect 14898 4626 14964 4638
rect 14898 4250 14914 4626
rect 14948 4250 14964 4626
rect 14898 4238 14964 4250
rect 14994 4626 15060 4638
rect 14994 4250 15010 4626
rect 15044 4250 15060 4626
rect 14994 4238 15060 4250
rect 15090 4626 15156 4638
rect 15090 4250 15106 4626
rect 15140 4250 15156 4626
rect 15090 4238 15156 4250
rect 15186 4626 15252 4638
rect 15186 4250 15202 4626
rect 15236 4250 15252 4626
rect 15186 4238 15252 4250
rect 15282 4626 15348 4638
rect 15282 4250 15298 4626
rect 15332 4250 15348 4626
rect 15282 4238 15348 4250
rect 15378 4626 15444 4638
rect 15378 4250 15394 4626
rect 15428 4250 15444 4626
rect 15378 4238 15444 4250
rect 15474 4626 15540 4638
rect 15474 4250 15490 4626
rect 15524 4250 15540 4626
rect 15474 4238 15540 4250
rect 15570 4626 15632 4638
rect 15570 4250 15586 4626
rect 15620 4250 15632 4626
rect 15570 4238 15632 4250
rect 16414 5862 16476 5874
rect 16414 5486 16426 5862
rect 16460 5486 16476 5862
rect 16414 5474 16476 5486
rect 16506 5862 16572 5874
rect 16506 5486 16522 5862
rect 16556 5486 16572 5862
rect 16506 5474 16572 5486
rect 16602 5862 16668 5874
rect 16602 5486 16618 5862
rect 16652 5486 16668 5862
rect 16602 5474 16668 5486
rect 16698 5862 16764 5874
rect 16698 5486 16714 5862
rect 16748 5486 16764 5862
rect 16698 5474 16764 5486
rect 16794 5862 16860 5874
rect 16794 5486 16810 5862
rect 16844 5486 16860 5862
rect 16794 5474 16860 5486
rect 16890 5862 16956 5874
rect 16890 5486 16906 5862
rect 16940 5486 16956 5862
rect 16890 5474 16956 5486
rect 16986 5862 17052 5874
rect 16986 5486 17002 5862
rect 17036 5486 17052 5862
rect 16986 5474 17052 5486
rect 17082 5862 17148 5874
rect 17082 5486 17098 5862
rect 17132 5486 17148 5862
rect 17082 5474 17148 5486
rect 17178 5862 17244 5874
rect 17178 5486 17194 5862
rect 17228 5486 17244 5862
rect 17178 5474 17244 5486
rect 17274 5862 17340 5874
rect 17274 5486 17290 5862
rect 17324 5486 17340 5862
rect 17274 5474 17340 5486
rect 17370 5862 17432 5874
rect 17370 5486 17386 5862
rect 17420 5486 17432 5862
rect 17370 5474 17432 5486
rect 16414 5244 16476 5256
rect 16414 4868 16426 5244
rect 16460 4868 16476 5244
rect 16414 4856 16476 4868
rect 16506 5244 16572 5256
rect 16506 4868 16522 5244
rect 16556 4868 16572 5244
rect 16506 4856 16572 4868
rect 16602 5244 16668 5256
rect 16602 4868 16618 5244
rect 16652 4868 16668 5244
rect 16602 4856 16668 4868
rect 16698 5244 16764 5256
rect 16698 4868 16714 5244
rect 16748 4868 16764 5244
rect 16698 4856 16764 4868
rect 16794 5244 16860 5256
rect 16794 4868 16810 5244
rect 16844 4868 16860 5244
rect 16794 4856 16860 4868
rect 16890 5244 16956 5256
rect 16890 4868 16906 5244
rect 16940 4868 16956 5244
rect 16890 4856 16956 4868
rect 16986 5244 17052 5256
rect 16986 4868 17002 5244
rect 17036 4868 17052 5244
rect 16986 4856 17052 4868
rect 17082 5244 17148 5256
rect 17082 4868 17098 5244
rect 17132 4868 17148 5244
rect 17082 4856 17148 4868
rect 17178 5244 17244 5256
rect 17178 4868 17194 5244
rect 17228 4868 17244 5244
rect 17178 4856 17244 4868
rect 17274 5244 17340 5256
rect 17274 4868 17290 5244
rect 17324 4868 17340 5244
rect 17274 4856 17340 4868
rect 17370 5244 17432 5256
rect 17370 4868 17386 5244
rect 17420 4868 17432 5244
rect 17370 4856 17432 4868
rect 16414 4626 16476 4638
rect 16414 4250 16426 4626
rect 16460 4250 16476 4626
rect 16414 4238 16476 4250
rect 16506 4626 16572 4638
rect 16506 4250 16522 4626
rect 16556 4250 16572 4626
rect 16506 4238 16572 4250
rect 16602 4626 16668 4638
rect 16602 4250 16618 4626
rect 16652 4250 16668 4626
rect 16602 4238 16668 4250
rect 16698 4626 16764 4638
rect 16698 4250 16714 4626
rect 16748 4250 16764 4626
rect 16698 4238 16764 4250
rect 16794 4626 16860 4638
rect 16794 4250 16810 4626
rect 16844 4250 16860 4626
rect 16794 4238 16860 4250
rect 16890 4626 16956 4638
rect 16890 4250 16906 4626
rect 16940 4250 16956 4626
rect 16890 4238 16956 4250
rect 16986 4626 17052 4638
rect 16986 4250 17002 4626
rect 17036 4250 17052 4626
rect 16986 4238 17052 4250
rect 17082 4626 17148 4638
rect 17082 4250 17098 4626
rect 17132 4250 17148 4626
rect 17082 4238 17148 4250
rect 17178 4626 17244 4638
rect 17178 4250 17194 4626
rect 17228 4250 17244 4626
rect 17178 4238 17244 4250
rect 17274 4626 17340 4638
rect 17274 4250 17290 4626
rect 17324 4250 17340 4626
rect 17274 4238 17340 4250
rect 17370 4626 17432 4638
rect 17370 4250 17386 4626
rect 17420 4250 17432 4626
rect 17370 4238 17432 4250
rect 18214 5862 18276 5874
rect 18214 5486 18226 5862
rect 18260 5486 18276 5862
rect 18214 5474 18276 5486
rect 18306 5862 18372 5874
rect 18306 5486 18322 5862
rect 18356 5486 18372 5862
rect 18306 5474 18372 5486
rect 18402 5862 18468 5874
rect 18402 5486 18418 5862
rect 18452 5486 18468 5862
rect 18402 5474 18468 5486
rect 18498 5862 18564 5874
rect 18498 5486 18514 5862
rect 18548 5486 18564 5862
rect 18498 5474 18564 5486
rect 18594 5862 18660 5874
rect 18594 5486 18610 5862
rect 18644 5486 18660 5862
rect 18594 5474 18660 5486
rect 18690 5862 18756 5874
rect 18690 5486 18706 5862
rect 18740 5486 18756 5862
rect 18690 5474 18756 5486
rect 18786 5862 18852 5874
rect 18786 5486 18802 5862
rect 18836 5486 18852 5862
rect 18786 5474 18852 5486
rect 18882 5862 18948 5874
rect 18882 5486 18898 5862
rect 18932 5486 18948 5862
rect 18882 5474 18948 5486
rect 18978 5862 19044 5874
rect 18978 5486 18994 5862
rect 19028 5486 19044 5862
rect 18978 5474 19044 5486
rect 19074 5862 19140 5874
rect 19074 5486 19090 5862
rect 19124 5486 19140 5862
rect 19074 5474 19140 5486
rect 19170 5862 19232 5874
rect 19170 5486 19186 5862
rect 19220 5486 19232 5862
rect 19170 5474 19232 5486
rect 18214 5244 18276 5256
rect 18214 4868 18226 5244
rect 18260 4868 18276 5244
rect 18214 4856 18276 4868
rect 18306 5244 18372 5256
rect 18306 4868 18322 5244
rect 18356 4868 18372 5244
rect 18306 4856 18372 4868
rect 18402 5244 18468 5256
rect 18402 4868 18418 5244
rect 18452 4868 18468 5244
rect 18402 4856 18468 4868
rect 18498 5244 18564 5256
rect 18498 4868 18514 5244
rect 18548 4868 18564 5244
rect 18498 4856 18564 4868
rect 18594 5244 18660 5256
rect 18594 4868 18610 5244
rect 18644 4868 18660 5244
rect 18594 4856 18660 4868
rect 18690 5244 18756 5256
rect 18690 4868 18706 5244
rect 18740 4868 18756 5244
rect 18690 4856 18756 4868
rect 18786 5244 18852 5256
rect 18786 4868 18802 5244
rect 18836 4868 18852 5244
rect 18786 4856 18852 4868
rect 18882 5244 18948 5256
rect 18882 4868 18898 5244
rect 18932 4868 18948 5244
rect 18882 4856 18948 4868
rect 18978 5244 19044 5256
rect 18978 4868 18994 5244
rect 19028 4868 19044 5244
rect 18978 4856 19044 4868
rect 19074 5244 19140 5256
rect 19074 4868 19090 5244
rect 19124 4868 19140 5244
rect 19074 4856 19140 4868
rect 19170 5244 19232 5256
rect 19170 4868 19186 5244
rect 19220 4868 19232 5244
rect 19170 4856 19232 4868
rect 18214 4626 18276 4638
rect 18214 4250 18226 4626
rect 18260 4250 18276 4626
rect 18214 4238 18276 4250
rect 18306 4626 18372 4638
rect 18306 4250 18322 4626
rect 18356 4250 18372 4626
rect 18306 4238 18372 4250
rect 18402 4626 18468 4638
rect 18402 4250 18418 4626
rect 18452 4250 18468 4626
rect 18402 4238 18468 4250
rect 18498 4626 18564 4638
rect 18498 4250 18514 4626
rect 18548 4250 18564 4626
rect 18498 4238 18564 4250
rect 18594 4626 18660 4638
rect 18594 4250 18610 4626
rect 18644 4250 18660 4626
rect 18594 4238 18660 4250
rect 18690 4626 18756 4638
rect 18690 4250 18706 4626
rect 18740 4250 18756 4626
rect 18690 4238 18756 4250
rect 18786 4626 18852 4638
rect 18786 4250 18802 4626
rect 18836 4250 18852 4626
rect 18786 4238 18852 4250
rect 18882 4626 18948 4638
rect 18882 4250 18898 4626
rect 18932 4250 18948 4626
rect 18882 4238 18948 4250
rect 18978 4626 19044 4638
rect 18978 4250 18994 4626
rect 19028 4250 19044 4626
rect 18978 4238 19044 4250
rect 19074 4626 19140 4638
rect 19074 4250 19090 4626
rect 19124 4250 19140 4626
rect 19074 4238 19140 4250
rect 19170 4626 19232 4638
rect 19170 4250 19186 4626
rect 19220 4250 19232 4626
rect 19170 4238 19232 4250
rect 20014 5862 20076 5874
rect 20014 5486 20026 5862
rect 20060 5486 20076 5862
rect 20014 5474 20076 5486
rect 20106 5862 20172 5874
rect 20106 5486 20122 5862
rect 20156 5486 20172 5862
rect 20106 5474 20172 5486
rect 20202 5862 20268 5874
rect 20202 5486 20218 5862
rect 20252 5486 20268 5862
rect 20202 5474 20268 5486
rect 20298 5862 20364 5874
rect 20298 5486 20314 5862
rect 20348 5486 20364 5862
rect 20298 5474 20364 5486
rect 20394 5862 20460 5874
rect 20394 5486 20410 5862
rect 20444 5486 20460 5862
rect 20394 5474 20460 5486
rect 20490 5862 20556 5874
rect 20490 5486 20506 5862
rect 20540 5486 20556 5862
rect 20490 5474 20556 5486
rect 20586 5862 20652 5874
rect 20586 5486 20602 5862
rect 20636 5486 20652 5862
rect 20586 5474 20652 5486
rect 20682 5862 20748 5874
rect 20682 5486 20698 5862
rect 20732 5486 20748 5862
rect 20682 5474 20748 5486
rect 20778 5862 20844 5874
rect 20778 5486 20794 5862
rect 20828 5486 20844 5862
rect 20778 5474 20844 5486
rect 20874 5862 20940 5874
rect 20874 5486 20890 5862
rect 20924 5486 20940 5862
rect 20874 5474 20940 5486
rect 20970 5862 21032 5874
rect 20970 5486 20986 5862
rect 21020 5486 21032 5862
rect 20970 5474 21032 5486
rect 20014 5244 20076 5256
rect 20014 4868 20026 5244
rect 20060 4868 20076 5244
rect 20014 4856 20076 4868
rect 20106 5244 20172 5256
rect 20106 4868 20122 5244
rect 20156 4868 20172 5244
rect 20106 4856 20172 4868
rect 20202 5244 20268 5256
rect 20202 4868 20218 5244
rect 20252 4868 20268 5244
rect 20202 4856 20268 4868
rect 20298 5244 20364 5256
rect 20298 4868 20314 5244
rect 20348 4868 20364 5244
rect 20298 4856 20364 4868
rect 20394 5244 20460 5256
rect 20394 4868 20410 5244
rect 20444 4868 20460 5244
rect 20394 4856 20460 4868
rect 20490 5244 20556 5256
rect 20490 4868 20506 5244
rect 20540 4868 20556 5244
rect 20490 4856 20556 4868
rect 20586 5244 20652 5256
rect 20586 4868 20602 5244
rect 20636 4868 20652 5244
rect 20586 4856 20652 4868
rect 20682 5244 20748 5256
rect 20682 4868 20698 5244
rect 20732 4868 20748 5244
rect 20682 4856 20748 4868
rect 20778 5244 20844 5256
rect 20778 4868 20794 5244
rect 20828 4868 20844 5244
rect 20778 4856 20844 4868
rect 20874 5244 20940 5256
rect 20874 4868 20890 5244
rect 20924 4868 20940 5244
rect 20874 4856 20940 4868
rect 20970 5244 21032 5256
rect 20970 4868 20986 5244
rect 21020 4868 21032 5244
rect 20970 4856 21032 4868
rect 20014 4626 20076 4638
rect 20014 4250 20026 4626
rect 20060 4250 20076 4626
rect 20014 4238 20076 4250
rect 20106 4626 20172 4638
rect 20106 4250 20122 4626
rect 20156 4250 20172 4626
rect 20106 4238 20172 4250
rect 20202 4626 20268 4638
rect 20202 4250 20218 4626
rect 20252 4250 20268 4626
rect 20202 4238 20268 4250
rect 20298 4626 20364 4638
rect 20298 4250 20314 4626
rect 20348 4250 20364 4626
rect 20298 4238 20364 4250
rect 20394 4626 20460 4638
rect 20394 4250 20410 4626
rect 20444 4250 20460 4626
rect 20394 4238 20460 4250
rect 20490 4626 20556 4638
rect 20490 4250 20506 4626
rect 20540 4250 20556 4626
rect 20490 4238 20556 4250
rect 20586 4626 20652 4638
rect 20586 4250 20602 4626
rect 20636 4250 20652 4626
rect 20586 4238 20652 4250
rect 20682 4626 20748 4638
rect 20682 4250 20698 4626
rect 20732 4250 20748 4626
rect 20682 4238 20748 4250
rect 20778 4626 20844 4638
rect 20778 4250 20794 4626
rect 20828 4250 20844 4626
rect 20778 4238 20844 4250
rect 20874 4626 20940 4638
rect 20874 4250 20890 4626
rect 20924 4250 20940 4626
rect 20874 4238 20940 4250
rect 20970 4626 21032 4638
rect 20970 4250 20986 4626
rect 21020 4250 21032 4626
rect 20970 4238 21032 4250
rect 22014 10250 22076 10262
rect 22014 9874 22026 10250
rect 22060 9874 22076 10250
rect 22014 9862 22076 9874
rect 22106 10250 22172 10262
rect 22106 9874 22122 10250
rect 22156 9874 22172 10250
rect 22106 9862 22172 9874
rect 22202 10250 22268 10262
rect 22202 9874 22218 10250
rect 22252 9874 22268 10250
rect 22202 9862 22268 9874
rect 22298 10250 22364 10262
rect 22298 9874 22314 10250
rect 22348 9874 22364 10250
rect 22298 9862 22364 9874
rect 22394 10250 22460 10262
rect 22394 9874 22410 10250
rect 22444 9874 22460 10250
rect 22394 9862 22460 9874
rect 22490 10250 22556 10262
rect 22490 9874 22506 10250
rect 22540 9874 22556 10250
rect 22490 9862 22556 9874
rect 22586 10250 22652 10262
rect 22586 9874 22602 10250
rect 22636 9874 22652 10250
rect 22586 9862 22652 9874
rect 22682 10250 22748 10262
rect 22682 9874 22698 10250
rect 22732 9874 22748 10250
rect 22682 9862 22748 9874
rect 22778 10250 22844 10262
rect 22778 9874 22794 10250
rect 22828 9874 22844 10250
rect 22778 9862 22844 9874
rect 22874 10250 22940 10262
rect 22874 9874 22890 10250
rect 22924 9874 22940 10250
rect 22874 9862 22940 9874
rect 22970 10250 23036 10262
rect 22970 9874 22986 10250
rect 23020 9874 23036 10250
rect 22970 9862 23036 9874
rect 23066 10250 23132 10262
rect 23066 9874 23082 10250
rect 23116 9874 23132 10250
rect 23066 9862 23132 9874
rect 23162 10250 23228 10262
rect 23162 9874 23178 10250
rect 23212 9874 23228 10250
rect 23162 9862 23228 9874
rect 23258 10250 23324 10262
rect 23258 9874 23274 10250
rect 23308 9874 23324 10250
rect 23258 9862 23324 9874
rect 23354 10250 23420 10262
rect 23354 9874 23370 10250
rect 23404 9874 23420 10250
rect 23354 9862 23420 9874
rect 23450 10250 23516 10262
rect 23450 9874 23466 10250
rect 23500 9874 23516 10250
rect 23450 9862 23516 9874
rect 23546 10250 23612 10262
rect 23546 9874 23562 10250
rect 23596 9874 23612 10250
rect 23546 9862 23612 9874
rect 23642 10250 23708 10262
rect 23642 9874 23658 10250
rect 23692 9874 23708 10250
rect 23642 9862 23708 9874
rect 23738 10250 23804 10262
rect 23738 9874 23754 10250
rect 23788 9874 23804 10250
rect 23738 9862 23804 9874
rect 23834 10250 23900 10262
rect 23834 9874 23850 10250
rect 23884 9874 23900 10250
rect 23834 9862 23900 9874
rect 23930 10250 23992 10262
rect 23930 9874 23946 10250
rect 23980 9874 23992 10250
rect 23930 9862 23992 9874
rect 22014 9632 22076 9644
rect 22014 9256 22026 9632
rect 22060 9256 22076 9632
rect 22014 9244 22076 9256
rect 22106 9632 22172 9644
rect 22106 9256 22122 9632
rect 22156 9256 22172 9632
rect 22106 9244 22172 9256
rect 22202 9632 22268 9644
rect 22202 9256 22218 9632
rect 22252 9256 22268 9632
rect 22202 9244 22268 9256
rect 22298 9632 22364 9644
rect 22298 9256 22314 9632
rect 22348 9256 22364 9632
rect 22298 9244 22364 9256
rect 22394 9632 22460 9644
rect 22394 9256 22410 9632
rect 22444 9256 22460 9632
rect 22394 9244 22460 9256
rect 22490 9632 22556 9644
rect 22490 9256 22506 9632
rect 22540 9256 22556 9632
rect 22490 9244 22556 9256
rect 22586 9632 22652 9644
rect 22586 9256 22602 9632
rect 22636 9256 22652 9632
rect 22586 9244 22652 9256
rect 22682 9632 22748 9644
rect 22682 9256 22698 9632
rect 22732 9256 22748 9632
rect 22682 9244 22748 9256
rect 22778 9632 22844 9644
rect 22778 9256 22794 9632
rect 22828 9256 22844 9632
rect 22778 9244 22844 9256
rect 22874 9632 22940 9644
rect 22874 9256 22890 9632
rect 22924 9256 22940 9632
rect 22874 9244 22940 9256
rect 22970 9632 23036 9644
rect 22970 9256 22986 9632
rect 23020 9256 23036 9632
rect 22970 9244 23036 9256
rect 23066 9632 23132 9644
rect 23066 9256 23082 9632
rect 23116 9256 23132 9632
rect 23066 9244 23132 9256
rect 23162 9632 23228 9644
rect 23162 9256 23178 9632
rect 23212 9256 23228 9632
rect 23162 9244 23228 9256
rect 23258 9632 23324 9644
rect 23258 9256 23274 9632
rect 23308 9256 23324 9632
rect 23258 9244 23324 9256
rect 23354 9632 23420 9644
rect 23354 9256 23370 9632
rect 23404 9256 23420 9632
rect 23354 9244 23420 9256
rect 23450 9632 23516 9644
rect 23450 9256 23466 9632
rect 23500 9256 23516 9632
rect 23450 9244 23516 9256
rect 23546 9632 23612 9644
rect 23546 9256 23562 9632
rect 23596 9256 23612 9632
rect 23546 9244 23612 9256
rect 23642 9632 23708 9644
rect 23642 9256 23658 9632
rect 23692 9256 23708 9632
rect 23642 9244 23708 9256
rect 23738 9632 23804 9644
rect 23738 9256 23754 9632
rect 23788 9256 23804 9632
rect 23738 9244 23804 9256
rect 23834 9632 23900 9644
rect 23834 9256 23850 9632
rect 23884 9256 23900 9632
rect 23834 9244 23900 9256
rect 23930 9632 23992 9644
rect 23930 9256 23946 9632
rect 23980 9256 23992 9632
rect 23930 9244 23992 9256
rect 22014 9014 22076 9026
rect 22014 8638 22026 9014
rect 22060 8638 22076 9014
rect 22014 8626 22076 8638
rect 22106 9014 22172 9026
rect 22106 8638 22122 9014
rect 22156 8638 22172 9014
rect 22106 8626 22172 8638
rect 22202 9014 22268 9026
rect 22202 8638 22218 9014
rect 22252 8638 22268 9014
rect 22202 8626 22268 8638
rect 22298 9014 22364 9026
rect 22298 8638 22314 9014
rect 22348 8638 22364 9014
rect 22298 8626 22364 8638
rect 22394 9014 22460 9026
rect 22394 8638 22410 9014
rect 22444 8638 22460 9014
rect 22394 8626 22460 8638
rect 22490 9014 22556 9026
rect 22490 8638 22506 9014
rect 22540 8638 22556 9014
rect 22490 8626 22556 8638
rect 22586 9014 22652 9026
rect 22586 8638 22602 9014
rect 22636 8638 22652 9014
rect 22586 8626 22652 8638
rect 22682 9014 22748 9026
rect 22682 8638 22698 9014
rect 22732 8638 22748 9014
rect 22682 8626 22748 8638
rect 22778 9014 22844 9026
rect 22778 8638 22794 9014
rect 22828 8638 22844 9014
rect 22778 8626 22844 8638
rect 22874 9014 22940 9026
rect 22874 8638 22890 9014
rect 22924 8638 22940 9014
rect 22874 8626 22940 8638
rect 22970 9014 23036 9026
rect 22970 8638 22986 9014
rect 23020 8638 23036 9014
rect 22970 8626 23036 8638
rect 23066 9014 23132 9026
rect 23066 8638 23082 9014
rect 23116 8638 23132 9014
rect 23066 8626 23132 8638
rect 23162 9014 23228 9026
rect 23162 8638 23178 9014
rect 23212 8638 23228 9014
rect 23162 8626 23228 8638
rect 23258 9014 23324 9026
rect 23258 8638 23274 9014
rect 23308 8638 23324 9014
rect 23258 8626 23324 8638
rect 23354 9014 23420 9026
rect 23354 8638 23370 9014
rect 23404 8638 23420 9014
rect 23354 8626 23420 8638
rect 23450 9014 23516 9026
rect 23450 8638 23466 9014
rect 23500 8638 23516 9014
rect 23450 8626 23516 8638
rect 23546 9014 23612 9026
rect 23546 8638 23562 9014
rect 23596 8638 23612 9014
rect 23546 8626 23612 8638
rect 23642 9014 23708 9026
rect 23642 8638 23658 9014
rect 23692 8638 23708 9014
rect 23642 8626 23708 8638
rect 23738 9014 23804 9026
rect 23738 8638 23754 9014
rect 23788 8638 23804 9014
rect 23738 8626 23804 8638
rect 23834 9014 23900 9026
rect 23834 8638 23850 9014
rect 23884 8638 23900 9014
rect 23834 8626 23900 8638
rect 23930 9014 23992 9026
rect 23930 8638 23946 9014
rect 23980 8638 23992 9014
rect 23930 8626 23992 8638
rect 22014 8396 22076 8408
rect 22014 8020 22026 8396
rect 22060 8020 22076 8396
rect 22014 8008 22076 8020
rect 22106 8396 22172 8408
rect 22106 8020 22122 8396
rect 22156 8020 22172 8396
rect 22106 8008 22172 8020
rect 22202 8396 22268 8408
rect 22202 8020 22218 8396
rect 22252 8020 22268 8396
rect 22202 8008 22268 8020
rect 22298 8396 22364 8408
rect 22298 8020 22314 8396
rect 22348 8020 22364 8396
rect 22298 8008 22364 8020
rect 22394 8396 22460 8408
rect 22394 8020 22410 8396
rect 22444 8020 22460 8396
rect 22394 8008 22460 8020
rect 22490 8396 22556 8408
rect 22490 8020 22506 8396
rect 22540 8020 22556 8396
rect 22490 8008 22556 8020
rect 22586 8396 22652 8408
rect 22586 8020 22602 8396
rect 22636 8020 22652 8396
rect 22586 8008 22652 8020
rect 22682 8396 22748 8408
rect 22682 8020 22698 8396
rect 22732 8020 22748 8396
rect 22682 8008 22748 8020
rect 22778 8396 22844 8408
rect 22778 8020 22794 8396
rect 22828 8020 22844 8396
rect 22778 8008 22844 8020
rect 22874 8396 22940 8408
rect 22874 8020 22890 8396
rect 22924 8020 22940 8396
rect 22874 8008 22940 8020
rect 22970 8396 23036 8408
rect 22970 8020 22986 8396
rect 23020 8020 23036 8396
rect 22970 8008 23036 8020
rect 23066 8396 23132 8408
rect 23066 8020 23082 8396
rect 23116 8020 23132 8396
rect 23066 8008 23132 8020
rect 23162 8396 23228 8408
rect 23162 8020 23178 8396
rect 23212 8020 23228 8396
rect 23162 8008 23228 8020
rect 23258 8396 23324 8408
rect 23258 8020 23274 8396
rect 23308 8020 23324 8396
rect 23258 8008 23324 8020
rect 23354 8396 23420 8408
rect 23354 8020 23370 8396
rect 23404 8020 23420 8396
rect 23354 8008 23420 8020
rect 23450 8396 23516 8408
rect 23450 8020 23466 8396
rect 23500 8020 23516 8396
rect 23450 8008 23516 8020
rect 23546 8396 23612 8408
rect 23546 8020 23562 8396
rect 23596 8020 23612 8396
rect 23546 8008 23612 8020
rect 23642 8396 23708 8408
rect 23642 8020 23658 8396
rect 23692 8020 23708 8396
rect 23642 8008 23708 8020
rect 23738 8396 23804 8408
rect 23738 8020 23754 8396
rect 23788 8020 23804 8396
rect 23738 8008 23804 8020
rect 23834 8396 23900 8408
rect 23834 8020 23850 8396
rect 23884 8020 23900 8396
rect 23834 8008 23900 8020
rect 23930 8396 23992 8408
rect 23930 8020 23946 8396
rect 23980 8020 23992 8396
rect 23930 8008 23992 8020
rect 22014 7778 22076 7790
rect 22014 7402 22026 7778
rect 22060 7402 22076 7778
rect 22014 7390 22076 7402
rect 22106 7778 22172 7790
rect 22106 7402 22122 7778
rect 22156 7402 22172 7778
rect 22106 7390 22172 7402
rect 22202 7778 22268 7790
rect 22202 7402 22218 7778
rect 22252 7402 22268 7778
rect 22202 7390 22268 7402
rect 22298 7778 22364 7790
rect 22298 7402 22314 7778
rect 22348 7402 22364 7778
rect 22298 7390 22364 7402
rect 22394 7778 22460 7790
rect 22394 7402 22410 7778
rect 22444 7402 22460 7778
rect 22394 7390 22460 7402
rect 22490 7778 22556 7790
rect 22490 7402 22506 7778
rect 22540 7402 22556 7778
rect 22490 7390 22556 7402
rect 22586 7778 22652 7790
rect 22586 7402 22602 7778
rect 22636 7402 22652 7778
rect 22586 7390 22652 7402
rect 22682 7778 22748 7790
rect 22682 7402 22698 7778
rect 22732 7402 22748 7778
rect 22682 7390 22748 7402
rect 22778 7778 22844 7790
rect 22778 7402 22794 7778
rect 22828 7402 22844 7778
rect 22778 7390 22844 7402
rect 22874 7778 22940 7790
rect 22874 7402 22890 7778
rect 22924 7402 22940 7778
rect 22874 7390 22940 7402
rect 22970 7778 23036 7790
rect 22970 7402 22986 7778
rect 23020 7402 23036 7778
rect 22970 7390 23036 7402
rect 23066 7778 23132 7790
rect 23066 7402 23082 7778
rect 23116 7402 23132 7778
rect 23066 7390 23132 7402
rect 23162 7778 23228 7790
rect 23162 7402 23178 7778
rect 23212 7402 23228 7778
rect 23162 7390 23228 7402
rect 23258 7778 23324 7790
rect 23258 7402 23274 7778
rect 23308 7402 23324 7778
rect 23258 7390 23324 7402
rect 23354 7778 23420 7790
rect 23354 7402 23370 7778
rect 23404 7402 23420 7778
rect 23354 7390 23420 7402
rect 23450 7778 23516 7790
rect 23450 7402 23466 7778
rect 23500 7402 23516 7778
rect 23450 7390 23516 7402
rect 23546 7778 23612 7790
rect 23546 7402 23562 7778
rect 23596 7402 23612 7778
rect 23546 7390 23612 7402
rect 23642 7778 23708 7790
rect 23642 7402 23658 7778
rect 23692 7402 23708 7778
rect 23642 7390 23708 7402
rect 23738 7778 23804 7790
rect 23738 7402 23754 7778
rect 23788 7402 23804 7778
rect 23738 7390 23804 7402
rect 23834 7778 23900 7790
rect 23834 7402 23850 7778
rect 23884 7402 23900 7778
rect 23834 7390 23900 7402
rect 23930 7778 23992 7790
rect 23930 7402 23946 7778
rect 23980 7402 23992 7778
rect 23930 7390 23992 7402
rect 22014 7160 22076 7172
rect 22014 6784 22026 7160
rect 22060 6784 22076 7160
rect 22014 6772 22076 6784
rect 22106 7160 22172 7172
rect 22106 6784 22122 7160
rect 22156 6784 22172 7160
rect 22106 6772 22172 6784
rect 22202 7160 22268 7172
rect 22202 6784 22218 7160
rect 22252 6784 22268 7160
rect 22202 6772 22268 6784
rect 22298 7160 22364 7172
rect 22298 6784 22314 7160
rect 22348 6784 22364 7160
rect 22298 6772 22364 6784
rect 22394 7160 22460 7172
rect 22394 6784 22410 7160
rect 22444 6784 22460 7160
rect 22394 6772 22460 6784
rect 22490 7160 22556 7172
rect 22490 6784 22506 7160
rect 22540 6784 22556 7160
rect 22490 6772 22556 6784
rect 22586 7160 22652 7172
rect 22586 6784 22602 7160
rect 22636 6784 22652 7160
rect 22586 6772 22652 6784
rect 22682 7160 22748 7172
rect 22682 6784 22698 7160
rect 22732 6784 22748 7160
rect 22682 6772 22748 6784
rect 22778 7160 22844 7172
rect 22778 6784 22794 7160
rect 22828 6784 22844 7160
rect 22778 6772 22844 6784
rect 22874 7160 22940 7172
rect 22874 6784 22890 7160
rect 22924 6784 22940 7160
rect 22874 6772 22940 6784
rect 22970 7160 23036 7172
rect 22970 6784 22986 7160
rect 23020 6784 23036 7160
rect 22970 6772 23036 6784
rect 23066 7160 23132 7172
rect 23066 6784 23082 7160
rect 23116 6784 23132 7160
rect 23066 6772 23132 6784
rect 23162 7160 23228 7172
rect 23162 6784 23178 7160
rect 23212 6784 23228 7160
rect 23162 6772 23228 6784
rect 23258 7160 23324 7172
rect 23258 6784 23274 7160
rect 23308 6784 23324 7160
rect 23258 6772 23324 6784
rect 23354 7160 23420 7172
rect 23354 6784 23370 7160
rect 23404 6784 23420 7160
rect 23354 6772 23420 6784
rect 23450 7160 23516 7172
rect 23450 6784 23466 7160
rect 23500 6784 23516 7160
rect 23450 6772 23516 6784
rect 23546 7160 23612 7172
rect 23546 6784 23562 7160
rect 23596 6784 23612 7160
rect 23546 6772 23612 6784
rect 23642 7160 23708 7172
rect 23642 6784 23658 7160
rect 23692 6784 23708 7160
rect 23642 6772 23708 6784
rect 23738 7160 23804 7172
rect 23738 6784 23754 7160
rect 23788 6784 23804 7160
rect 23738 6772 23804 6784
rect 23834 7160 23900 7172
rect 23834 6784 23850 7160
rect 23884 6784 23900 7160
rect 23834 6772 23900 6784
rect 23930 7160 23992 7172
rect 23930 6784 23946 7160
rect 23980 6784 23992 7160
rect 23930 6772 23992 6784
rect 22014 6542 22076 6554
rect 22014 6166 22026 6542
rect 22060 6166 22076 6542
rect 22014 6154 22076 6166
rect 22106 6542 22172 6554
rect 22106 6166 22122 6542
rect 22156 6166 22172 6542
rect 22106 6154 22172 6166
rect 22202 6542 22268 6554
rect 22202 6166 22218 6542
rect 22252 6166 22268 6542
rect 22202 6154 22268 6166
rect 22298 6542 22364 6554
rect 22298 6166 22314 6542
rect 22348 6166 22364 6542
rect 22298 6154 22364 6166
rect 22394 6542 22460 6554
rect 22394 6166 22410 6542
rect 22444 6166 22460 6542
rect 22394 6154 22460 6166
rect 22490 6542 22556 6554
rect 22490 6166 22506 6542
rect 22540 6166 22556 6542
rect 22490 6154 22556 6166
rect 22586 6542 22652 6554
rect 22586 6166 22602 6542
rect 22636 6166 22652 6542
rect 22586 6154 22652 6166
rect 22682 6542 22748 6554
rect 22682 6166 22698 6542
rect 22732 6166 22748 6542
rect 22682 6154 22748 6166
rect 22778 6542 22844 6554
rect 22778 6166 22794 6542
rect 22828 6166 22844 6542
rect 22778 6154 22844 6166
rect 22874 6542 22940 6554
rect 22874 6166 22890 6542
rect 22924 6166 22940 6542
rect 22874 6154 22940 6166
rect 22970 6542 23036 6554
rect 22970 6166 22986 6542
rect 23020 6166 23036 6542
rect 22970 6154 23036 6166
rect 23066 6542 23132 6554
rect 23066 6166 23082 6542
rect 23116 6166 23132 6542
rect 23066 6154 23132 6166
rect 23162 6542 23228 6554
rect 23162 6166 23178 6542
rect 23212 6166 23228 6542
rect 23162 6154 23228 6166
rect 23258 6542 23324 6554
rect 23258 6166 23274 6542
rect 23308 6166 23324 6542
rect 23258 6154 23324 6166
rect 23354 6542 23420 6554
rect 23354 6166 23370 6542
rect 23404 6166 23420 6542
rect 23354 6154 23420 6166
rect 23450 6542 23516 6554
rect 23450 6166 23466 6542
rect 23500 6166 23516 6542
rect 23450 6154 23516 6166
rect 23546 6542 23612 6554
rect 23546 6166 23562 6542
rect 23596 6166 23612 6542
rect 23546 6154 23612 6166
rect 23642 6542 23708 6554
rect 23642 6166 23658 6542
rect 23692 6166 23708 6542
rect 23642 6154 23708 6166
rect 23738 6542 23804 6554
rect 23738 6166 23754 6542
rect 23788 6166 23804 6542
rect 23738 6154 23804 6166
rect 23834 6542 23900 6554
rect 23834 6166 23850 6542
rect 23884 6166 23900 6542
rect 23834 6154 23900 6166
rect 23930 6542 23992 6554
rect 23930 6166 23946 6542
rect 23980 6166 23992 6542
rect 23930 6154 23992 6166
rect 22014 5924 22076 5936
rect 22014 5548 22026 5924
rect 22060 5548 22076 5924
rect 22014 5536 22076 5548
rect 22106 5924 22172 5936
rect 22106 5548 22122 5924
rect 22156 5548 22172 5924
rect 22106 5536 22172 5548
rect 22202 5924 22268 5936
rect 22202 5548 22218 5924
rect 22252 5548 22268 5924
rect 22202 5536 22268 5548
rect 22298 5924 22364 5936
rect 22298 5548 22314 5924
rect 22348 5548 22364 5924
rect 22298 5536 22364 5548
rect 22394 5924 22460 5936
rect 22394 5548 22410 5924
rect 22444 5548 22460 5924
rect 22394 5536 22460 5548
rect 22490 5924 22556 5936
rect 22490 5548 22506 5924
rect 22540 5548 22556 5924
rect 22490 5536 22556 5548
rect 22586 5924 22652 5936
rect 22586 5548 22602 5924
rect 22636 5548 22652 5924
rect 22586 5536 22652 5548
rect 22682 5924 22748 5936
rect 22682 5548 22698 5924
rect 22732 5548 22748 5924
rect 22682 5536 22748 5548
rect 22778 5924 22844 5936
rect 22778 5548 22794 5924
rect 22828 5548 22844 5924
rect 22778 5536 22844 5548
rect 22874 5924 22940 5936
rect 22874 5548 22890 5924
rect 22924 5548 22940 5924
rect 22874 5536 22940 5548
rect 22970 5924 23036 5936
rect 22970 5548 22986 5924
rect 23020 5548 23036 5924
rect 22970 5536 23036 5548
rect 23066 5924 23132 5936
rect 23066 5548 23082 5924
rect 23116 5548 23132 5924
rect 23066 5536 23132 5548
rect 23162 5924 23228 5936
rect 23162 5548 23178 5924
rect 23212 5548 23228 5924
rect 23162 5536 23228 5548
rect 23258 5924 23324 5936
rect 23258 5548 23274 5924
rect 23308 5548 23324 5924
rect 23258 5536 23324 5548
rect 23354 5924 23420 5936
rect 23354 5548 23370 5924
rect 23404 5548 23420 5924
rect 23354 5536 23420 5548
rect 23450 5924 23516 5936
rect 23450 5548 23466 5924
rect 23500 5548 23516 5924
rect 23450 5536 23516 5548
rect 23546 5924 23612 5936
rect 23546 5548 23562 5924
rect 23596 5548 23612 5924
rect 23546 5536 23612 5548
rect 23642 5924 23708 5936
rect 23642 5548 23658 5924
rect 23692 5548 23708 5924
rect 23642 5536 23708 5548
rect 23738 5924 23804 5936
rect 23738 5548 23754 5924
rect 23788 5548 23804 5924
rect 23738 5536 23804 5548
rect 23834 5924 23900 5936
rect 23834 5548 23850 5924
rect 23884 5548 23900 5924
rect 23834 5536 23900 5548
rect 23930 5924 23992 5936
rect 23930 5548 23946 5924
rect 23980 5548 23992 5924
rect 23930 5536 23992 5548
rect 22014 5306 22076 5318
rect 22014 4930 22026 5306
rect 22060 4930 22076 5306
rect 22014 4918 22076 4930
rect 22106 5306 22172 5318
rect 22106 4930 22122 5306
rect 22156 4930 22172 5306
rect 22106 4918 22172 4930
rect 22202 5306 22268 5318
rect 22202 4930 22218 5306
rect 22252 4930 22268 5306
rect 22202 4918 22268 4930
rect 22298 5306 22364 5318
rect 22298 4930 22314 5306
rect 22348 4930 22364 5306
rect 22298 4918 22364 4930
rect 22394 5306 22460 5318
rect 22394 4930 22410 5306
rect 22444 4930 22460 5306
rect 22394 4918 22460 4930
rect 22490 5306 22556 5318
rect 22490 4930 22506 5306
rect 22540 4930 22556 5306
rect 22490 4918 22556 4930
rect 22586 5306 22652 5318
rect 22586 4930 22602 5306
rect 22636 4930 22652 5306
rect 22586 4918 22652 4930
rect 22682 5306 22748 5318
rect 22682 4930 22698 5306
rect 22732 4930 22748 5306
rect 22682 4918 22748 4930
rect 22778 5306 22844 5318
rect 22778 4930 22794 5306
rect 22828 4930 22844 5306
rect 22778 4918 22844 4930
rect 22874 5306 22940 5318
rect 22874 4930 22890 5306
rect 22924 4930 22940 5306
rect 22874 4918 22940 4930
rect 22970 5306 23036 5318
rect 22970 4930 22986 5306
rect 23020 4930 23036 5306
rect 22970 4918 23036 4930
rect 23066 5306 23132 5318
rect 23066 4930 23082 5306
rect 23116 4930 23132 5306
rect 23066 4918 23132 4930
rect 23162 5306 23228 5318
rect 23162 4930 23178 5306
rect 23212 4930 23228 5306
rect 23162 4918 23228 4930
rect 23258 5306 23324 5318
rect 23258 4930 23274 5306
rect 23308 4930 23324 5306
rect 23258 4918 23324 4930
rect 23354 5306 23420 5318
rect 23354 4930 23370 5306
rect 23404 4930 23420 5306
rect 23354 4918 23420 4930
rect 23450 5306 23516 5318
rect 23450 4930 23466 5306
rect 23500 4930 23516 5306
rect 23450 4918 23516 4930
rect 23546 5306 23612 5318
rect 23546 4930 23562 5306
rect 23596 4930 23612 5306
rect 23546 4918 23612 4930
rect 23642 5306 23708 5318
rect 23642 4930 23658 5306
rect 23692 4930 23708 5306
rect 23642 4918 23708 4930
rect 23738 5306 23804 5318
rect 23738 4930 23754 5306
rect 23788 4930 23804 5306
rect 23738 4918 23804 4930
rect 23834 5306 23900 5318
rect 23834 4930 23850 5306
rect 23884 4930 23900 5306
rect 23834 4918 23900 4930
rect 23930 5306 23992 5318
rect 23930 4930 23946 5306
rect 23980 4930 23992 5306
rect 23930 4918 23992 4930
rect 214 3716 272 3728
rect 214 3340 226 3716
rect 260 3340 272 3716
rect 214 3328 272 3340
rect 472 3716 530 3728
rect 472 3340 484 3716
rect 518 3340 530 3716
rect 472 3328 530 3340
rect 730 3716 788 3728
rect 730 3340 742 3716
rect 776 3340 788 3716
rect 730 3328 788 3340
rect 988 3716 1046 3728
rect 988 3340 1000 3716
rect 1034 3340 1046 3716
rect 988 3328 1046 3340
rect 1246 3716 1304 3728
rect 1246 3340 1258 3716
rect 1292 3340 1304 3716
rect 1246 3328 1304 3340
rect 1504 3716 1562 3728
rect 1504 3340 1516 3716
rect 1550 3340 1562 3716
rect 1504 3328 1562 3340
rect 214 3098 272 3110
rect 214 2722 226 3098
rect 260 2722 272 3098
rect 214 2710 272 2722
rect 472 3098 530 3110
rect 472 2722 484 3098
rect 518 2722 530 3098
rect 472 2710 530 2722
rect 730 3098 788 3110
rect 730 2722 742 3098
rect 776 2722 788 3098
rect 730 2710 788 2722
rect 988 3098 1046 3110
rect 988 2722 1000 3098
rect 1034 2722 1046 3098
rect 988 2710 1046 2722
rect 1246 3098 1304 3110
rect 1246 2722 1258 3098
rect 1292 2722 1304 3098
rect 1246 2710 1304 2722
rect 1504 3098 1562 3110
rect 1504 2722 1516 3098
rect 1550 2722 1562 3098
rect 1504 2710 1562 2722
rect 214 2480 272 2492
rect 214 2104 226 2480
rect 260 2104 272 2480
rect 214 2092 272 2104
rect 472 2480 530 2492
rect 472 2104 484 2480
rect 518 2104 530 2480
rect 472 2092 530 2104
rect 730 2480 788 2492
rect 730 2104 742 2480
rect 776 2104 788 2480
rect 730 2092 788 2104
rect 988 2480 1046 2492
rect 988 2104 1000 2480
rect 1034 2104 1046 2480
rect 988 2092 1046 2104
rect 1246 2480 1304 2492
rect 1246 2104 1258 2480
rect 1292 2104 1304 2480
rect 1246 2092 1304 2104
rect 1504 2480 1562 2492
rect 1504 2104 1516 2480
rect 1550 2104 1562 2480
rect 1504 2092 1562 2104
rect 214 1862 272 1874
rect 214 1486 226 1862
rect 260 1486 272 1862
rect 214 1474 272 1486
rect 472 1862 530 1874
rect 472 1486 484 1862
rect 518 1486 530 1862
rect 472 1474 530 1486
rect 730 1862 788 1874
rect 730 1486 742 1862
rect 776 1486 788 1862
rect 730 1474 788 1486
rect 988 1862 1046 1874
rect 988 1486 1000 1862
rect 1034 1486 1046 1862
rect 988 1474 1046 1486
rect 1246 1862 1304 1874
rect 1246 1486 1258 1862
rect 1292 1486 1304 1862
rect 1246 1474 1304 1486
rect 1504 1862 1562 1874
rect 1504 1486 1516 1862
rect 1550 1486 1562 1862
rect 1504 1474 1562 1486
rect 214 1244 272 1256
rect 214 868 226 1244
rect 260 868 272 1244
rect 214 856 272 868
rect 472 1244 530 1256
rect 472 868 484 1244
rect 518 868 530 1244
rect 472 856 530 868
rect 730 1244 788 1256
rect 730 868 742 1244
rect 776 868 788 1244
rect 730 856 788 868
rect 988 1244 1046 1256
rect 988 868 1000 1244
rect 1034 868 1046 1244
rect 988 856 1046 868
rect 1246 1244 1304 1256
rect 1246 868 1258 1244
rect 1292 868 1304 1244
rect 1246 856 1304 868
rect 1504 1244 1562 1256
rect 1504 868 1516 1244
rect 1550 868 1562 1244
rect 1504 856 1562 868
rect 214 626 272 638
rect 214 250 226 626
rect 260 250 272 626
rect 214 238 272 250
rect 472 626 530 638
rect 472 250 484 626
rect 518 250 530 626
rect 472 238 530 250
rect 730 626 788 638
rect 730 250 742 626
rect 776 250 788 626
rect 730 238 788 250
rect 988 626 1046 638
rect 988 250 1000 626
rect 1034 250 1046 626
rect 988 238 1046 250
rect 1246 626 1304 638
rect 1246 250 1258 626
rect 1292 250 1304 626
rect 1246 238 1304 250
rect 1504 626 1562 638
rect 1504 250 1516 626
rect 1550 250 1562 626
rect 1504 238 1562 250
rect 2014 3716 2072 3728
rect 2014 3340 2026 3716
rect 2060 3340 2072 3716
rect 2014 3328 2072 3340
rect 2272 3716 2330 3728
rect 2272 3340 2284 3716
rect 2318 3340 2330 3716
rect 2272 3328 2330 3340
rect 2530 3716 2588 3728
rect 2530 3340 2542 3716
rect 2576 3340 2588 3716
rect 2530 3328 2588 3340
rect 2788 3716 2846 3728
rect 2788 3340 2800 3716
rect 2834 3340 2846 3716
rect 2788 3328 2846 3340
rect 3046 3716 3104 3728
rect 3046 3340 3058 3716
rect 3092 3340 3104 3716
rect 3046 3328 3104 3340
rect 3304 3716 3362 3728
rect 3304 3340 3316 3716
rect 3350 3340 3362 3716
rect 3304 3328 3362 3340
rect 2014 3098 2072 3110
rect 2014 2722 2026 3098
rect 2060 2722 2072 3098
rect 2014 2710 2072 2722
rect 2272 3098 2330 3110
rect 2272 2722 2284 3098
rect 2318 2722 2330 3098
rect 2272 2710 2330 2722
rect 2530 3098 2588 3110
rect 2530 2722 2542 3098
rect 2576 2722 2588 3098
rect 2530 2710 2588 2722
rect 2788 3098 2846 3110
rect 2788 2722 2800 3098
rect 2834 2722 2846 3098
rect 2788 2710 2846 2722
rect 3046 3098 3104 3110
rect 3046 2722 3058 3098
rect 3092 2722 3104 3098
rect 3046 2710 3104 2722
rect 3304 3098 3362 3110
rect 3304 2722 3316 3098
rect 3350 2722 3362 3098
rect 3304 2710 3362 2722
rect 2014 2480 2072 2492
rect 2014 2104 2026 2480
rect 2060 2104 2072 2480
rect 2014 2092 2072 2104
rect 2272 2480 2330 2492
rect 2272 2104 2284 2480
rect 2318 2104 2330 2480
rect 2272 2092 2330 2104
rect 2530 2480 2588 2492
rect 2530 2104 2542 2480
rect 2576 2104 2588 2480
rect 2530 2092 2588 2104
rect 2788 2480 2846 2492
rect 2788 2104 2800 2480
rect 2834 2104 2846 2480
rect 2788 2092 2846 2104
rect 3046 2480 3104 2492
rect 3046 2104 3058 2480
rect 3092 2104 3104 2480
rect 3046 2092 3104 2104
rect 3304 2480 3362 2492
rect 3304 2104 3316 2480
rect 3350 2104 3362 2480
rect 3304 2092 3362 2104
rect 2014 1862 2072 1874
rect 2014 1486 2026 1862
rect 2060 1486 2072 1862
rect 2014 1474 2072 1486
rect 2272 1862 2330 1874
rect 2272 1486 2284 1862
rect 2318 1486 2330 1862
rect 2272 1474 2330 1486
rect 2530 1862 2588 1874
rect 2530 1486 2542 1862
rect 2576 1486 2588 1862
rect 2530 1474 2588 1486
rect 2788 1862 2846 1874
rect 2788 1486 2800 1862
rect 2834 1486 2846 1862
rect 2788 1474 2846 1486
rect 3046 1862 3104 1874
rect 3046 1486 3058 1862
rect 3092 1486 3104 1862
rect 3046 1474 3104 1486
rect 3304 1862 3362 1874
rect 3304 1486 3316 1862
rect 3350 1486 3362 1862
rect 3304 1474 3362 1486
rect 2014 1244 2072 1256
rect 2014 868 2026 1244
rect 2060 868 2072 1244
rect 2014 856 2072 868
rect 2272 1244 2330 1256
rect 2272 868 2284 1244
rect 2318 868 2330 1244
rect 2272 856 2330 868
rect 2530 1244 2588 1256
rect 2530 868 2542 1244
rect 2576 868 2588 1244
rect 2530 856 2588 868
rect 2788 1244 2846 1256
rect 2788 868 2800 1244
rect 2834 868 2846 1244
rect 2788 856 2846 868
rect 3046 1244 3104 1256
rect 3046 868 3058 1244
rect 3092 868 3104 1244
rect 3046 856 3104 868
rect 3304 1244 3362 1256
rect 3304 868 3316 1244
rect 3350 868 3362 1244
rect 3304 856 3362 868
rect 2014 626 2072 638
rect 2014 250 2026 626
rect 2060 250 2072 626
rect 2014 238 2072 250
rect 2272 626 2330 638
rect 2272 250 2284 626
rect 2318 250 2330 626
rect 2272 238 2330 250
rect 2530 626 2588 638
rect 2530 250 2542 626
rect 2576 250 2588 626
rect 2530 238 2588 250
rect 2788 626 2846 638
rect 2788 250 2800 626
rect 2834 250 2846 626
rect 2788 238 2846 250
rect 3046 626 3104 638
rect 3046 250 3058 626
rect 3092 250 3104 626
rect 3046 238 3104 250
rect 3304 626 3362 638
rect 3304 250 3316 626
rect 3350 250 3362 626
rect 3304 238 3362 250
rect 3814 3716 3872 3728
rect 3814 3340 3826 3716
rect 3860 3340 3872 3716
rect 3814 3328 3872 3340
rect 4072 3716 4130 3728
rect 4072 3340 4084 3716
rect 4118 3340 4130 3716
rect 4072 3328 4130 3340
rect 4330 3716 4388 3728
rect 4330 3340 4342 3716
rect 4376 3340 4388 3716
rect 4330 3328 4388 3340
rect 4588 3716 4646 3728
rect 4588 3340 4600 3716
rect 4634 3340 4646 3716
rect 4588 3328 4646 3340
rect 4846 3716 4904 3728
rect 4846 3340 4858 3716
rect 4892 3340 4904 3716
rect 4846 3328 4904 3340
rect 5104 3716 5162 3728
rect 5104 3340 5116 3716
rect 5150 3340 5162 3716
rect 5104 3328 5162 3340
rect 3814 3098 3872 3110
rect 3814 2722 3826 3098
rect 3860 2722 3872 3098
rect 3814 2710 3872 2722
rect 4072 3098 4130 3110
rect 4072 2722 4084 3098
rect 4118 2722 4130 3098
rect 4072 2710 4130 2722
rect 4330 3098 4388 3110
rect 4330 2722 4342 3098
rect 4376 2722 4388 3098
rect 4330 2710 4388 2722
rect 4588 3098 4646 3110
rect 4588 2722 4600 3098
rect 4634 2722 4646 3098
rect 4588 2710 4646 2722
rect 4846 3098 4904 3110
rect 4846 2722 4858 3098
rect 4892 2722 4904 3098
rect 4846 2710 4904 2722
rect 5104 3098 5162 3110
rect 5104 2722 5116 3098
rect 5150 2722 5162 3098
rect 5104 2710 5162 2722
rect 3814 2480 3872 2492
rect 3814 2104 3826 2480
rect 3860 2104 3872 2480
rect 3814 2092 3872 2104
rect 4072 2480 4130 2492
rect 4072 2104 4084 2480
rect 4118 2104 4130 2480
rect 4072 2092 4130 2104
rect 4330 2480 4388 2492
rect 4330 2104 4342 2480
rect 4376 2104 4388 2480
rect 4330 2092 4388 2104
rect 4588 2480 4646 2492
rect 4588 2104 4600 2480
rect 4634 2104 4646 2480
rect 4588 2092 4646 2104
rect 4846 2480 4904 2492
rect 4846 2104 4858 2480
rect 4892 2104 4904 2480
rect 4846 2092 4904 2104
rect 5104 2480 5162 2492
rect 5104 2104 5116 2480
rect 5150 2104 5162 2480
rect 5104 2092 5162 2104
rect 3814 1862 3872 1874
rect 3814 1486 3826 1862
rect 3860 1486 3872 1862
rect 3814 1474 3872 1486
rect 4072 1862 4130 1874
rect 4072 1486 4084 1862
rect 4118 1486 4130 1862
rect 4072 1474 4130 1486
rect 4330 1862 4388 1874
rect 4330 1486 4342 1862
rect 4376 1486 4388 1862
rect 4330 1474 4388 1486
rect 4588 1862 4646 1874
rect 4588 1486 4600 1862
rect 4634 1486 4646 1862
rect 4588 1474 4646 1486
rect 4846 1862 4904 1874
rect 4846 1486 4858 1862
rect 4892 1486 4904 1862
rect 4846 1474 4904 1486
rect 5104 1862 5162 1874
rect 5104 1486 5116 1862
rect 5150 1486 5162 1862
rect 5104 1474 5162 1486
rect 3814 1244 3872 1256
rect 3814 868 3826 1244
rect 3860 868 3872 1244
rect 3814 856 3872 868
rect 4072 1244 4130 1256
rect 4072 868 4084 1244
rect 4118 868 4130 1244
rect 4072 856 4130 868
rect 4330 1244 4388 1256
rect 4330 868 4342 1244
rect 4376 868 4388 1244
rect 4330 856 4388 868
rect 4588 1244 4646 1256
rect 4588 868 4600 1244
rect 4634 868 4646 1244
rect 4588 856 4646 868
rect 4846 1244 4904 1256
rect 4846 868 4858 1244
rect 4892 868 4904 1244
rect 4846 856 4904 868
rect 5104 1244 5162 1256
rect 5104 868 5116 1244
rect 5150 868 5162 1244
rect 5104 856 5162 868
rect 3814 626 3872 638
rect 3814 250 3826 626
rect 3860 250 3872 626
rect 3814 238 3872 250
rect 4072 626 4130 638
rect 4072 250 4084 626
rect 4118 250 4130 626
rect 4072 238 4130 250
rect 4330 626 4388 638
rect 4330 250 4342 626
rect 4376 250 4388 626
rect 4330 238 4388 250
rect 4588 626 4646 638
rect 4588 250 4600 626
rect 4634 250 4646 626
rect 4588 238 4646 250
rect 4846 626 4904 638
rect 4846 250 4858 626
rect 4892 250 4904 626
rect 4846 238 4904 250
rect 5104 626 5162 638
rect 5104 250 5116 626
rect 5150 250 5162 626
rect 5104 238 5162 250
rect 5614 3716 5672 3728
rect 5614 3340 5626 3716
rect 5660 3340 5672 3716
rect 5614 3328 5672 3340
rect 5872 3716 5930 3728
rect 5872 3340 5884 3716
rect 5918 3340 5930 3716
rect 5872 3328 5930 3340
rect 6130 3716 6188 3728
rect 6130 3340 6142 3716
rect 6176 3340 6188 3716
rect 6130 3328 6188 3340
rect 6388 3716 6446 3728
rect 6388 3340 6400 3716
rect 6434 3340 6446 3716
rect 6388 3328 6446 3340
rect 6646 3716 6704 3728
rect 6646 3340 6658 3716
rect 6692 3340 6704 3716
rect 6646 3328 6704 3340
rect 6904 3716 6962 3728
rect 6904 3340 6916 3716
rect 6950 3340 6962 3716
rect 6904 3328 6962 3340
rect 5614 3098 5672 3110
rect 5614 2722 5626 3098
rect 5660 2722 5672 3098
rect 5614 2710 5672 2722
rect 5872 3098 5930 3110
rect 5872 2722 5884 3098
rect 5918 2722 5930 3098
rect 5872 2710 5930 2722
rect 6130 3098 6188 3110
rect 6130 2722 6142 3098
rect 6176 2722 6188 3098
rect 6130 2710 6188 2722
rect 6388 3098 6446 3110
rect 6388 2722 6400 3098
rect 6434 2722 6446 3098
rect 6388 2710 6446 2722
rect 6646 3098 6704 3110
rect 6646 2722 6658 3098
rect 6692 2722 6704 3098
rect 6646 2710 6704 2722
rect 6904 3098 6962 3110
rect 6904 2722 6916 3098
rect 6950 2722 6962 3098
rect 6904 2710 6962 2722
rect 5614 2480 5672 2492
rect 5614 2104 5626 2480
rect 5660 2104 5672 2480
rect 5614 2092 5672 2104
rect 5872 2480 5930 2492
rect 5872 2104 5884 2480
rect 5918 2104 5930 2480
rect 5872 2092 5930 2104
rect 6130 2480 6188 2492
rect 6130 2104 6142 2480
rect 6176 2104 6188 2480
rect 6130 2092 6188 2104
rect 6388 2480 6446 2492
rect 6388 2104 6400 2480
rect 6434 2104 6446 2480
rect 6388 2092 6446 2104
rect 6646 2480 6704 2492
rect 6646 2104 6658 2480
rect 6692 2104 6704 2480
rect 6646 2092 6704 2104
rect 6904 2480 6962 2492
rect 6904 2104 6916 2480
rect 6950 2104 6962 2480
rect 6904 2092 6962 2104
rect 5614 1862 5672 1874
rect 5614 1486 5626 1862
rect 5660 1486 5672 1862
rect 5614 1474 5672 1486
rect 5872 1862 5930 1874
rect 5872 1486 5884 1862
rect 5918 1486 5930 1862
rect 5872 1474 5930 1486
rect 6130 1862 6188 1874
rect 6130 1486 6142 1862
rect 6176 1486 6188 1862
rect 6130 1474 6188 1486
rect 6388 1862 6446 1874
rect 6388 1486 6400 1862
rect 6434 1486 6446 1862
rect 6388 1474 6446 1486
rect 6646 1862 6704 1874
rect 6646 1486 6658 1862
rect 6692 1486 6704 1862
rect 6646 1474 6704 1486
rect 6904 1862 6962 1874
rect 6904 1486 6916 1862
rect 6950 1486 6962 1862
rect 6904 1474 6962 1486
rect 5614 1244 5672 1256
rect 5614 868 5626 1244
rect 5660 868 5672 1244
rect 5614 856 5672 868
rect 5872 1244 5930 1256
rect 5872 868 5884 1244
rect 5918 868 5930 1244
rect 5872 856 5930 868
rect 6130 1244 6188 1256
rect 6130 868 6142 1244
rect 6176 868 6188 1244
rect 6130 856 6188 868
rect 6388 1244 6446 1256
rect 6388 868 6400 1244
rect 6434 868 6446 1244
rect 6388 856 6446 868
rect 6646 1244 6704 1256
rect 6646 868 6658 1244
rect 6692 868 6704 1244
rect 6646 856 6704 868
rect 6904 1244 6962 1256
rect 6904 868 6916 1244
rect 6950 868 6962 1244
rect 6904 856 6962 868
rect 5614 626 5672 638
rect 5614 250 5626 626
rect 5660 250 5672 626
rect 5614 238 5672 250
rect 5872 626 5930 638
rect 5872 250 5884 626
rect 5918 250 5930 626
rect 5872 238 5930 250
rect 6130 626 6188 638
rect 6130 250 6142 626
rect 6176 250 6188 626
rect 6130 238 6188 250
rect 6388 626 6446 638
rect 6388 250 6400 626
rect 6434 250 6446 626
rect 6388 238 6446 250
rect 6646 626 6704 638
rect 6646 250 6658 626
rect 6692 250 6704 626
rect 6646 238 6704 250
rect 6904 626 6962 638
rect 6904 250 6916 626
rect 6950 250 6962 626
rect 6904 238 6962 250
rect 14614 3716 14672 3728
rect 14614 3340 14626 3716
rect 14660 3340 14672 3716
rect 14614 3328 14672 3340
rect 14872 3716 14930 3728
rect 14872 3340 14884 3716
rect 14918 3340 14930 3716
rect 14872 3328 14930 3340
rect 15130 3716 15188 3728
rect 15130 3340 15142 3716
rect 15176 3340 15188 3716
rect 15130 3328 15188 3340
rect 15388 3716 15446 3728
rect 15388 3340 15400 3716
rect 15434 3340 15446 3716
rect 15388 3328 15446 3340
rect 15646 3716 15704 3728
rect 15646 3340 15658 3716
rect 15692 3340 15704 3716
rect 15646 3328 15704 3340
rect 15904 3716 15962 3728
rect 15904 3340 15916 3716
rect 15950 3340 15962 3716
rect 15904 3328 15962 3340
rect 14614 3098 14672 3110
rect 14614 2722 14626 3098
rect 14660 2722 14672 3098
rect 14614 2710 14672 2722
rect 14872 3098 14930 3110
rect 14872 2722 14884 3098
rect 14918 2722 14930 3098
rect 14872 2710 14930 2722
rect 15130 3098 15188 3110
rect 15130 2722 15142 3098
rect 15176 2722 15188 3098
rect 15130 2710 15188 2722
rect 15388 3098 15446 3110
rect 15388 2722 15400 3098
rect 15434 2722 15446 3098
rect 15388 2710 15446 2722
rect 15646 3098 15704 3110
rect 15646 2722 15658 3098
rect 15692 2722 15704 3098
rect 15646 2710 15704 2722
rect 15904 3098 15962 3110
rect 15904 2722 15916 3098
rect 15950 2722 15962 3098
rect 15904 2710 15962 2722
rect 14614 2480 14672 2492
rect 14614 2104 14626 2480
rect 14660 2104 14672 2480
rect 14614 2092 14672 2104
rect 14872 2480 14930 2492
rect 14872 2104 14884 2480
rect 14918 2104 14930 2480
rect 14872 2092 14930 2104
rect 15130 2480 15188 2492
rect 15130 2104 15142 2480
rect 15176 2104 15188 2480
rect 15130 2092 15188 2104
rect 15388 2480 15446 2492
rect 15388 2104 15400 2480
rect 15434 2104 15446 2480
rect 15388 2092 15446 2104
rect 15646 2480 15704 2492
rect 15646 2104 15658 2480
rect 15692 2104 15704 2480
rect 15646 2092 15704 2104
rect 15904 2480 15962 2492
rect 15904 2104 15916 2480
rect 15950 2104 15962 2480
rect 15904 2092 15962 2104
rect 14614 1862 14672 1874
rect 14614 1486 14626 1862
rect 14660 1486 14672 1862
rect 14614 1474 14672 1486
rect 14872 1862 14930 1874
rect 14872 1486 14884 1862
rect 14918 1486 14930 1862
rect 14872 1474 14930 1486
rect 15130 1862 15188 1874
rect 15130 1486 15142 1862
rect 15176 1486 15188 1862
rect 15130 1474 15188 1486
rect 15388 1862 15446 1874
rect 15388 1486 15400 1862
rect 15434 1486 15446 1862
rect 15388 1474 15446 1486
rect 15646 1862 15704 1874
rect 15646 1486 15658 1862
rect 15692 1486 15704 1862
rect 15646 1474 15704 1486
rect 15904 1862 15962 1874
rect 15904 1486 15916 1862
rect 15950 1486 15962 1862
rect 15904 1474 15962 1486
rect 14614 1244 14672 1256
rect 14614 868 14626 1244
rect 14660 868 14672 1244
rect 14614 856 14672 868
rect 14872 1244 14930 1256
rect 14872 868 14884 1244
rect 14918 868 14930 1244
rect 14872 856 14930 868
rect 15130 1244 15188 1256
rect 15130 868 15142 1244
rect 15176 868 15188 1244
rect 15130 856 15188 868
rect 15388 1244 15446 1256
rect 15388 868 15400 1244
rect 15434 868 15446 1244
rect 15388 856 15446 868
rect 15646 1244 15704 1256
rect 15646 868 15658 1244
rect 15692 868 15704 1244
rect 15646 856 15704 868
rect 15904 1244 15962 1256
rect 15904 868 15916 1244
rect 15950 868 15962 1244
rect 15904 856 15962 868
rect 14614 626 14672 638
rect 14614 250 14626 626
rect 14660 250 14672 626
rect 14614 238 14672 250
rect 14872 626 14930 638
rect 14872 250 14884 626
rect 14918 250 14930 626
rect 14872 238 14930 250
rect 15130 626 15188 638
rect 15130 250 15142 626
rect 15176 250 15188 626
rect 15130 238 15188 250
rect 15388 626 15446 638
rect 15388 250 15400 626
rect 15434 250 15446 626
rect 15388 238 15446 250
rect 15646 626 15704 638
rect 15646 250 15658 626
rect 15692 250 15704 626
rect 15646 238 15704 250
rect 15904 626 15962 638
rect 15904 250 15916 626
rect 15950 250 15962 626
rect 15904 238 15962 250
rect 16414 3716 16472 3728
rect 16414 3340 16426 3716
rect 16460 3340 16472 3716
rect 16414 3328 16472 3340
rect 16672 3716 16730 3728
rect 16672 3340 16684 3716
rect 16718 3340 16730 3716
rect 16672 3328 16730 3340
rect 16930 3716 16988 3728
rect 16930 3340 16942 3716
rect 16976 3340 16988 3716
rect 16930 3328 16988 3340
rect 17188 3716 17246 3728
rect 17188 3340 17200 3716
rect 17234 3340 17246 3716
rect 17188 3328 17246 3340
rect 17446 3716 17504 3728
rect 17446 3340 17458 3716
rect 17492 3340 17504 3716
rect 17446 3328 17504 3340
rect 17704 3716 17762 3728
rect 17704 3340 17716 3716
rect 17750 3340 17762 3716
rect 17704 3328 17762 3340
rect 16414 3098 16472 3110
rect 16414 2722 16426 3098
rect 16460 2722 16472 3098
rect 16414 2710 16472 2722
rect 16672 3098 16730 3110
rect 16672 2722 16684 3098
rect 16718 2722 16730 3098
rect 16672 2710 16730 2722
rect 16930 3098 16988 3110
rect 16930 2722 16942 3098
rect 16976 2722 16988 3098
rect 16930 2710 16988 2722
rect 17188 3098 17246 3110
rect 17188 2722 17200 3098
rect 17234 2722 17246 3098
rect 17188 2710 17246 2722
rect 17446 3098 17504 3110
rect 17446 2722 17458 3098
rect 17492 2722 17504 3098
rect 17446 2710 17504 2722
rect 17704 3098 17762 3110
rect 17704 2722 17716 3098
rect 17750 2722 17762 3098
rect 17704 2710 17762 2722
rect 16414 2480 16472 2492
rect 16414 2104 16426 2480
rect 16460 2104 16472 2480
rect 16414 2092 16472 2104
rect 16672 2480 16730 2492
rect 16672 2104 16684 2480
rect 16718 2104 16730 2480
rect 16672 2092 16730 2104
rect 16930 2480 16988 2492
rect 16930 2104 16942 2480
rect 16976 2104 16988 2480
rect 16930 2092 16988 2104
rect 17188 2480 17246 2492
rect 17188 2104 17200 2480
rect 17234 2104 17246 2480
rect 17188 2092 17246 2104
rect 17446 2480 17504 2492
rect 17446 2104 17458 2480
rect 17492 2104 17504 2480
rect 17446 2092 17504 2104
rect 17704 2480 17762 2492
rect 17704 2104 17716 2480
rect 17750 2104 17762 2480
rect 17704 2092 17762 2104
rect 16414 1862 16472 1874
rect 16414 1486 16426 1862
rect 16460 1486 16472 1862
rect 16414 1474 16472 1486
rect 16672 1862 16730 1874
rect 16672 1486 16684 1862
rect 16718 1486 16730 1862
rect 16672 1474 16730 1486
rect 16930 1862 16988 1874
rect 16930 1486 16942 1862
rect 16976 1486 16988 1862
rect 16930 1474 16988 1486
rect 17188 1862 17246 1874
rect 17188 1486 17200 1862
rect 17234 1486 17246 1862
rect 17188 1474 17246 1486
rect 17446 1862 17504 1874
rect 17446 1486 17458 1862
rect 17492 1486 17504 1862
rect 17446 1474 17504 1486
rect 17704 1862 17762 1874
rect 17704 1486 17716 1862
rect 17750 1486 17762 1862
rect 17704 1474 17762 1486
rect 16414 1244 16472 1256
rect 16414 868 16426 1244
rect 16460 868 16472 1244
rect 16414 856 16472 868
rect 16672 1244 16730 1256
rect 16672 868 16684 1244
rect 16718 868 16730 1244
rect 16672 856 16730 868
rect 16930 1244 16988 1256
rect 16930 868 16942 1244
rect 16976 868 16988 1244
rect 16930 856 16988 868
rect 17188 1244 17246 1256
rect 17188 868 17200 1244
rect 17234 868 17246 1244
rect 17188 856 17246 868
rect 17446 1244 17504 1256
rect 17446 868 17458 1244
rect 17492 868 17504 1244
rect 17446 856 17504 868
rect 17704 1244 17762 1256
rect 17704 868 17716 1244
rect 17750 868 17762 1244
rect 17704 856 17762 868
rect 16414 626 16472 638
rect 16414 250 16426 626
rect 16460 250 16472 626
rect 16414 238 16472 250
rect 16672 626 16730 638
rect 16672 250 16684 626
rect 16718 250 16730 626
rect 16672 238 16730 250
rect 16930 626 16988 638
rect 16930 250 16942 626
rect 16976 250 16988 626
rect 16930 238 16988 250
rect 17188 626 17246 638
rect 17188 250 17200 626
rect 17234 250 17246 626
rect 17188 238 17246 250
rect 17446 626 17504 638
rect 17446 250 17458 626
rect 17492 250 17504 626
rect 17446 238 17504 250
rect 17704 626 17762 638
rect 17704 250 17716 626
rect 17750 250 17762 626
rect 17704 238 17762 250
rect 18214 3716 18272 3728
rect 18214 3340 18226 3716
rect 18260 3340 18272 3716
rect 18214 3328 18272 3340
rect 18472 3716 18530 3728
rect 18472 3340 18484 3716
rect 18518 3340 18530 3716
rect 18472 3328 18530 3340
rect 18730 3716 18788 3728
rect 18730 3340 18742 3716
rect 18776 3340 18788 3716
rect 18730 3328 18788 3340
rect 18988 3716 19046 3728
rect 18988 3340 19000 3716
rect 19034 3340 19046 3716
rect 18988 3328 19046 3340
rect 19246 3716 19304 3728
rect 19246 3340 19258 3716
rect 19292 3340 19304 3716
rect 19246 3328 19304 3340
rect 19504 3716 19562 3728
rect 19504 3340 19516 3716
rect 19550 3340 19562 3716
rect 19504 3328 19562 3340
rect 18214 3098 18272 3110
rect 18214 2722 18226 3098
rect 18260 2722 18272 3098
rect 18214 2710 18272 2722
rect 18472 3098 18530 3110
rect 18472 2722 18484 3098
rect 18518 2722 18530 3098
rect 18472 2710 18530 2722
rect 18730 3098 18788 3110
rect 18730 2722 18742 3098
rect 18776 2722 18788 3098
rect 18730 2710 18788 2722
rect 18988 3098 19046 3110
rect 18988 2722 19000 3098
rect 19034 2722 19046 3098
rect 18988 2710 19046 2722
rect 19246 3098 19304 3110
rect 19246 2722 19258 3098
rect 19292 2722 19304 3098
rect 19246 2710 19304 2722
rect 19504 3098 19562 3110
rect 19504 2722 19516 3098
rect 19550 2722 19562 3098
rect 19504 2710 19562 2722
rect 18214 2480 18272 2492
rect 18214 2104 18226 2480
rect 18260 2104 18272 2480
rect 18214 2092 18272 2104
rect 18472 2480 18530 2492
rect 18472 2104 18484 2480
rect 18518 2104 18530 2480
rect 18472 2092 18530 2104
rect 18730 2480 18788 2492
rect 18730 2104 18742 2480
rect 18776 2104 18788 2480
rect 18730 2092 18788 2104
rect 18988 2480 19046 2492
rect 18988 2104 19000 2480
rect 19034 2104 19046 2480
rect 18988 2092 19046 2104
rect 19246 2480 19304 2492
rect 19246 2104 19258 2480
rect 19292 2104 19304 2480
rect 19246 2092 19304 2104
rect 19504 2480 19562 2492
rect 19504 2104 19516 2480
rect 19550 2104 19562 2480
rect 19504 2092 19562 2104
rect 18214 1862 18272 1874
rect 18214 1486 18226 1862
rect 18260 1486 18272 1862
rect 18214 1474 18272 1486
rect 18472 1862 18530 1874
rect 18472 1486 18484 1862
rect 18518 1486 18530 1862
rect 18472 1474 18530 1486
rect 18730 1862 18788 1874
rect 18730 1486 18742 1862
rect 18776 1486 18788 1862
rect 18730 1474 18788 1486
rect 18988 1862 19046 1874
rect 18988 1486 19000 1862
rect 19034 1486 19046 1862
rect 18988 1474 19046 1486
rect 19246 1862 19304 1874
rect 19246 1486 19258 1862
rect 19292 1486 19304 1862
rect 19246 1474 19304 1486
rect 19504 1862 19562 1874
rect 19504 1486 19516 1862
rect 19550 1486 19562 1862
rect 19504 1474 19562 1486
rect 18214 1244 18272 1256
rect 18214 868 18226 1244
rect 18260 868 18272 1244
rect 18214 856 18272 868
rect 18472 1244 18530 1256
rect 18472 868 18484 1244
rect 18518 868 18530 1244
rect 18472 856 18530 868
rect 18730 1244 18788 1256
rect 18730 868 18742 1244
rect 18776 868 18788 1244
rect 18730 856 18788 868
rect 18988 1244 19046 1256
rect 18988 868 19000 1244
rect 19034 868 19046 1244
rect 18988 856 19046 868
rect 19246 1244 19304 1256
rect 19246 868 19258 1244
rect 19292 868 19304 1244
rect 19246 856 19304 868
rect 19504 1244 19562 1256
rect 19504 868 19516 1244
rect 19550 868 19562 1244
rect 19504 856 19562 868
rect 18214 626 18272 638
rect 18214 250 18226 626
rect 18260 250 18272 626
rect 18214 238 18272 250
rect 18472 626 18530 638
rect 18472 250 18484 626
rect 18518 250 18530 626
rect 18472 238 18530 250
rect 18730 626 18788 638
rect 18730 250 18742 626
rect 18776 250 18788 626
rect 18730 238 18788 250
rect 18988 626 19046 638
rect 18988 250 19000 626
rect 19034 250 19046 626
rect 18988 238 19046 250
rect 19246 626 19304 638
rect 19246 250 19258 626
rect 19292 250 19304 626
rect 19246 238 19304 250
rect 19504 626 19562 638
rect 19504 250 19516 626
rect 19550 250 19562 626
rect 19504 238 19562 250
rect 20014 3716 20072 3728
rect 20014 3340 20026 3716
rect 20060 3340 20072 3716
rect 20014 3328 20072 3340
rect 20272 3716 20330 3728
rect 20272 3340 20284 3716
rect 20318 3340 20330 3716
rect 20272 3328 20330 3340
rect 20530 3716 20588 3728
rect 20530 3340 20542 3716
rect 20576 3340 20588 3716
rect 20530 3328 20588 3340
rect 20788 3716 20846 3728
rect 20788 3340 20800 3716
rect 20834 3340 20846 3716
rect 20788 3328 20846 3340
rect 21046 3716 21104 3728
rect 21046 3340 21058 3716
rect 21092 3340 21104 3716
rect 21046 3328 21104 3340
rect 21304 3716 21362 3728
rect 21304 3340 21316 3716
rect 21350 3340 21362 3716
rect 21304 3328 21362 3340
rect 20014 3098 20072 3110
rect 20014 2722 20026 3098
rect 20060 2722 20072 3098
rect 20014 2710 20072 2722
rect 20272 3098 20330 3110
rect 20272 2722 20284 3098
rect 20318 2722 20330 3098
rect 20272 2710 20330 2722
rect 20530 3098 20588 3110
rect 20530 2722 20542 3098
rect 20576 2722 20588 3098
rect 20530 2710 20588 2722
rect 20788 3098 20846 3110
rect 20788 2722 20800 3098
rect 20834 2722 20846 3098
rect 20788 2710 20846 2722
rect 21046 3098 21104 3110
rect 21046 2722 21058 3098
rect 21092 2722 21104 3098
rect 21046 2710 21104 2722
rect 21304 3098 21362 3110
rect 21304 2722 21316 3098
rect 21350 2722 21362 3098
rect 21304 2710 21362 2722
rect 20014 2480 20072 2492
rect 20014 2104 20026 2480
rect 20060 2104 20072 2480
rect 20014 2092 20072 2104
rect 20272 2480 20330 2492
rect 20272 2104 20284 2480
rect 20318 2104 20330 2480
rect 20272 2092 20330 2104
rect 20530 2480 20588 2492
rect 20530 2104 20542 2480
rect 20576 2104 20588 2480
rect 20530 2092 20588 2104
rect 20788 2480 20846 2492
rect 20788 2104 20800 2480
rect 20834 2104 20846 2480
rect 20788 2092 20846 2104
rect 21046 2480 21104 2492
rect 21046 2104 21058 2480
rect 21092 2104 21104 2480
rect 21046 2092 21104 2104
rect 21304 2480 21362 2492
rect 21304 2104 21316 2480
rect 21350 2104 21362 2480
rect 21304 2092 21362 2104
rect 20014 1862 20072 1874
rect 20014 1486 20026 1862
rect 20060 1486 20072 1862
rect 20014 1474 20072 1486
rect 20272 1862 20330 1874
rect 20272 1486 20284 1862
rect 20318 1486 20330 1862
rect 20272 1474 20330 1486
rect 20530 1862 20588 1874
rect 20530 1486 20542 1862
rect 20576 1486 20588 1862
rect 20530 1474 20588 1486
rect 20788 1862 20846 1874
rect 20788 1486 20800 1862
rect 20834 1486 20846 1862
rect 20788 1474 20846 1486
rect 21046 1862 21104 1874
rect 21046 1486 21058 1862
rect 21092 1486 21104 1862
rect 21046 1474 21104 1486
rect 21304 1862 21362 1874
rect 21304 1486 21316 1862
rect 21350 1486 21362 1862
rect 21304 1474 21362 1486
rect 20014 1244 20072 1256
rect 20014 868 20026 1244
rect 20060 868 20072 1244
rect 20014 856 20072 868
rect 20272 1244 20330 1256
rect 20272 868 20284 1244
rect 20318 868 20330 1244
rect 20272 856 20330 868
rect 20530 1244 20588 1256
rect 20530 868 20542 1244
rect 20576 868 20588 1244
rect 20530 856 20588 868
rect 20788 1244 20846 1256
rect 20788 868 20800 1244
rect 20834 868 20846 1244
rect 20788 856 20846 868
rect 21046 1244 21104 1256
rect 21046 868 21058 1244
rect 21092 868 21104 1244
rect 21046 856 21104 868
rect 21304 1244 21362 1256
rect 21304 868 21316 1244
rect 21350 868 21362 1244
rect 21304 856 21362 868
rect 20014 626 20072 638
rect 20014 250 20026 626
rect 20060 250 20072 626
rect 20014 238 20072 250
rect 20272 626 20330 638
rect 20272 250 20284 626
rect 20318 250 20330 626
rect 20272 238 20330 250
rect 20530 626 20588 638
rect 20530 250 20542 626
rect 20576 250 20588 626
rect 20530 238 20588 250
rect 20788 626 20846 638
rect 20788 250 20800 626
rect 20834 250 20846 626
rect 20788 238 20846 250
rect 21046 626 21104 638
rect 21046 250 21058 626
rect 21092 250 21104 626
rect 21046 238 21104 250
rect 21304 626 21362 638
rect 21304 250 21316 626
rect 21350 250 21362 626
rect 21304 238 21362 250
<< pdiff >>
rect 6478 27075 6536 27087
rect 6478 26699 6490 27075
rect 6524 26699 6536 27075
rect 6478 26687 6536 26699
rect 6636 27075 6694 27087
rect 6636 26699 6648 27075
rect 6682 26699 6694 27075
rect 6636 26687 6694 26699
rect 6794 27075 6852 27087
rect 6794 26699 6806 27075
rect 6840 26699 6852 27075
rect 6794 26687 6852 26699
rect 6952 27075 7010 27087
rect 6952 26699 6964 27075
rect 6998 26699 7010 27075
rect 6952 26687 7010 26699
rect 7110 27075 7168 27087
rect 7110 26699 7122 27075
rect 7156 26699 7168 27075
rect 7110 26687 7168 26699
rect 7268 27075 7326 27087
rect 7268 26699 7280 27075
rect 7314 26699 7326 27075
rect 7268 26687 7326 26699
rect 7426 27075 7484 27087
rect 7426 26699 7438 27075
rect 7472 26699 7484 27075
rect 7426 26687 7484 26699
rect 7584 27075 7642 27087
rect 7584 26699 7596 27075
rect 7630 26699 7642 27075
rect 7584 26687 7642 26699
rect 7742 27075 7800 27087
rect 7742 26699 7754 27075
rect 7788 26699 7800 27075
rect 7742 26687 7800 26699
rect 7900 27075 7958 27087
rect 7900 26699 7912 27075
rect 7946 26699 7958 27075
rect 7900 26687 7958 26699
rect 8058 27075 8116 27087
rect 8058 26699 8070 27075
rect 8104 26699 8116 27075
rect 8058 26687 8116 26699
rect 6478 26439 6536 26451
rect 6478 26063 6490 26439
rect 6524 26063 6536 26439
rect 6478 26051 6536 26063
rect 6636 26439 6694 26451
rect 6636 26063 6648 26439
rect 6682 26063 6694 26439
rect 6636 26051 6694 26063
rect 6794 26439 6852 26451
rect 6794 26063 6806 26439
rect 6840 26063 6852 26439
rect 6794 26051 6852 26063
rect 6952 26439 7010 26451
rect 6952 26063 6964 26439
rect 6998 26063 7010 26439
rect 6952 26051 7010 26063
rect 7110 26439 7168 26451
rect 7110 26063 7122 26439
rect 7156 26063 7168 26439
rect 7110 26051 7168 26063
rect 7268 26439 7326 26451
rect 7268 26063 7280 26439
rect 7314 26063 7326 26439
rect 7268 26051 7326 26063
rect 7426 26439 7484 26451
rect 7426 26063 7438 26439
rect 7472 26063 7484 26439
rect 7426 26051 7484 26063
rect 7584 26439 7642 26451
rect 7584 26063 7596 26439
rect 7630 26063 7642 26439
rect 7584 26051 7642 26063
rect 7742 26439 7800 26451
rect 7742 26063 7754 26439
rect 7788 26063 7800 26439
rect 7742 26051 7800 26063
rect 7900 26439 7958 26451
rect 7900 26063 7912 26439
rect 7946 26063 7958 26439
rect 7900 26051 7958 26063
rect 8058 26439 8116 26451
rect 8058 26063 8070 26439
rect 8104 26063 8116 26439
rect 8058 26051 8116 26063
rect 6478 25803 6536 25815
rect 6478 25427 6490 25803
rect 6524 25427 6536 25803
rect 6478 25415 6536 25427
rect 6636 25803 6694 25815
rect 6636 25427 6648 25803
rect 6682 25427 6694 25803
rect 6636 25415 6694 25427
rect 6794 25803 6852 25815
rect 6794 25427 6806 25803
rect 6840 25427 6852 25803
rect 6794 25415 6852 25427
rect 6952 25803 7010 25815
rect 6952 25427 6964 25803
rect 6998 25427 7010 25803
rect 6952 25415 7010 25427
rect 7110 25803 7168 25815
rect 7110 25427 7122 25803
rect 7156 25427 7168 25803
rect 7110 25415 7168 25427
rect 7268 25803 7326 25815
rect 7268 25427 7280 25803
rect 7314 25427 7326 25803
rect 7268 25415 7326 25427
rect 7426 25803 7484 25815
rect 7426 25427 7438 25803
rect 7472 25427 7484 25803
rect 7426 25415 7484 25427
rect 7584 25803 7642 25815
rect 7584 25427 7596 25803
rect 7630 25427 7642 25803
rect 7584 25415 7642 25427
rect 7742 25803 7800 25815
rect 7742 25427 7754 25803
rect 7788 25427 7800 25803
rect 7742 25415 7800 25427
rect 7900 25803 7958 25815
rect 7900 25427 7912 25803
rect 7946 25427 7958 25803
rect 7900 25415 7958 25427
rect 8058 25803 8116 25815
rect 8058 25427 8070 25803
rect 8104 25427 8116 25803
rect 8058 25415 8116 25427
rect 8698 27075 8756 27087
rect 8698 26699 8710 27075
rect 8744 26699 8756 27075
rect 8698 26687 8756 26699
rect 8856 27075 8914 27087
rect 8856 26699 8868 27075
rect 8902 26699 8914 27075
rect 8856 26687 8914 26699
rect 9014 27075 9072 27087
rect 9014 26699 9026 27075
rect 9060 26699 9072 27075
rect 9014 26687 9072 26699
rect 9172 27075 9230 27087
rect 9172 26699 9184 27075
rect 9218 26699 9230 27075
rect 9172 26687 9230 26699
rect 9330 27075 9388 27087
rect 9330 26699 9342 27075
rect 9376 26699 9388 27075
rect 9330 26687 9388 26699
rect 9488 27075 9546 27087
rect 9488 26699 9500 27075
rect 9534 26699 9546 27075
rect 9488 26687 9546 26699
rect 9646 27075 9704 27087
rect 9646 26699 9658 27075
rect 9692 26699 9704 27075
rect 9646 26687 9704 26699
rect 9804 27075 9862 27087
rect 9804 26699 9816 27075
rect 9850 26699 9862 27075
rect 9804 26687 9862 26699
rect 9962 27075 10020 27087
rect 9962 26699 9974 27075
rect 10008 26699 10020 27075
rect 9962 26687 10020 26699
rect 10120 27075 10178 27087
rect 10120 26699 10132 27075
rect 10166 26699 10178 27075
rect 10120 26687 10178 26699
rect 10278 27075 10336 27087
rect 10278 26699 10290 27075
rect 10324 26699 10336 27075
rect 10278 26687 10336 26699
rect 8698 26439 8756 26451
rect 8698 26063 8710 26439
rect 8744 26063 8756 26439
rect 8698 26051 8756 26063
rect 8856 26439 8914 26451
rect 8856 26063 8868 26439
rect 8902 26063 8914 26439
rect 8856 26051 8914 26063
rect 9014 26439 9072 26451
rect 9014 26063 9026 26439
rect 9060 26063 9072 26439
rect 9014 26051 9072 26063
rect 9172 26439 9230 26451
rect 9172 26063 9184 26439
rect 9218 26063 9230 26439
rect 9172 26051 9230 26063
rect 9330 26439 9388 26451
rect 9330 26063 9342 26439
rect 9376 26063 9388 26439
rect 9330 26051 9388 26063
rect 9488 26439 9546 26451
rect 9488 26063 9500 26439
rect 9534 26063 9546 26439
rect 9488 26051 9546 26063
rect 9646 26439 9704 26451
rect 9646 26063 9658 26439
rect 9692 26063 9704 26439
rect 9646 26051 9704 26063
rect 9804 26439 9862 26451
rect 9804 26063 9816 26439
rect 9850 26063 9862 26439
rect 9804 26051 9862 26063
rect 9962 26439 10020 26451
rect 9962 26063 9974 26439
rect 10008 26063 10020 26439
rect 9962 26051 10020 26063
rect 10120 26439 10178 26451
rect 10120 26063 10132 26439
rect 10166 26063 10178 26439
rect 10120 26051 10178 26063
rect 10278 26439 10336 26451
rect 10278 26063 10290 26439
rect 10324 26063 10336 26439
rect 10278 26051 10336 26063
rect 8698 25803 8756 25815
rect 8698 25427 8710 25803
rect 8744 25427 8756 25803
rect 8698 25415 8756 25427
rect 8856 25803 8914 25815
rect 8856 25427 8868 25803
rect 8902 25427 8914 25803
rect 8856 25415 8914 25427
rect 9014 25803 9072 25815
rect 9014 25427 9026 25803
rect 9060 25427 9072 25803
rect 9014 25415 9072 25427
rect 9172 25803 9230 25815
rect 9172 25427 9184 25803
rect 9218 25427 9230 25803
rect 9172 25415 9230 25427
rect 9330 25803 9388 25815
rect 9330 25427 9342 25803
rect 9376 25427 9388 25803
rect 9330 25415 9388 25427
rect 9488 25803 9546 25815
rect 9488 25427 9500 25803
rect 9534 25427 9546 25803
rect 9488 25415 9546 25427
rect 9646 25803 9704 25815
rect 9646 25427 9658 25803
rect 9692 25427 9704 25803
rect 9646 25415 9704 25427
rect 9804 25803 9862 25815
rect 9804 25427 9816 25803
rect 9850 25427 9862 25803
rect 9804 25415 9862 25427
rect 9962 25803 10020 25815
rect 9962 25427 9974 25803
rect 10008 25427 10020 25803
rect 9962 25415 10020 25427
rect 10120 25803 10178 25815
rect 10120 25427 10132 25803
rect 10166 25427 10178 25803
rect 10120 25415 10178 25427
rect 10278 25803 10336 25815
rect 10278 25427 10290 25803
rect 10324 25427 10336 25803
rect 10278 25415 10336 25427
rect 10878 27075 10936 27087
rect 10878 26699 10890 27075
rect 10924 26699 10936 27075
rect 10878 26687 10936 26699
rect 11036 27075 11094 27087
rect 11036 26699 11048 27075
rect 11082 26699 11094 27075
rect 11036 26687 11094 26699
rect 11194 27075 11252 27087
rect 11194 26699 11206 27075
rect 11240 26699 11252 27075
rect 11194 26687 11252 26699
rect 11352 27075 11410 27087
rect 11352 26699 11364 27075
rect 11398 26699 11410 27075
rect 11352 26687 11410 26699
rect 11510 27075 11568 27087
rect 11510 26699 11522 27075
rect 11556 26699 11568 27075
rect 11510 26687 11568 26699
rect 11668 27075 11726 27087
rect 11668 26699 11680 27075
rect 11714 26699 11726 27075
rect 11668 26687 11726 26699
rect 11826 27075 11884 27087
rect 11826 26699 11838 27075
rect 11872 26699 11884 27075
rect 11826 26687 11884 26699
rect 11984 27075 12042 27087
rect 11984 26699 11996 27075
rect 12030 26699 12042 27075
rect 11984 26687 12042 26699
rect 12142 27075 12200 27087
rect 12142 26699 12154 27075
rect 12188 26699 12200 27075
rect 12142 26687 12200 26699
rect 12300 27075 12358 27087
rect 12300 26699 12312 27075
rect 12346 26699 12358 27075
rect 12300 26687 12358 26699
rect 12458 27075 12516 27087
rect 12458 26699 12470 27075
rect 12504 26699 12516 27075
rect 12458 26687 12516 26699
rect 10878 26439 10936 26451
rect 10878 26063 10890 26439
rect 10924 26063 10936 26439
rect 10878 26051 10936 26063
rect 11036 26439 11094 26451
rect 11036 26063 11048 26439
rect 11082 26063 11094 26439
rect 11036 26051 11094 26063
rect 11194 26439 11252 26451
rect 11194 26063 11206 26439
rect 11240 26063 11252 26439
rect 11194 26051 11252 26063
rect 11352 26439 11410 26451
rect 11352 26063 11364 26439
rect 11398 26063 11410 26439
rect 11352 26051 11410 26063
rect 11510 26439 11568 26451
rect 11510 26063 11522 26439
rect 11556 26063 11568 26439
rect 11510 26051 11568 26063
rect 11668 26439 11726 26451
rect 11668 26063 11680 26439
rect 11714 26063 11726 26439
rect 11668 26051 11726 26063
rect 11826 26439 11884 26451
rect 11826 26063 11838 26439
rect 11872 26063 11884 26439
rect 11826 26051 11884 26063
rect 11984 26439 12042 26451
rect 11984 26063 11996 26439
rect 12030 26063 12042 26439
rect 11984 26051 12042 26063
rect 12142 26439 12200 26451
rect 12142 26063 12154 26439
rect 12188 26063 12200 26439
rect 12142 26051 12200 26063
rect 12300 26439 12358 26451
rect 12300 26063 12312 26439
rect 12346 26063 12358 26439
rect 12300 26051 12358 26063
rect 12458 26439 12516 26451
rect 12458 26063 12470 26439
rect 12504 26063 12516 26439
rect 12458 26051 12516 26063
rect 10878 25803 10936 25815
rect 10878 25427 10890 25803
rect 10924 25427 10936 25803
rect 10878 25415 10936 25427
rect 11036 25803 11094 25815
rect 11036 25427 11048 25803
rect 11082 25427 11094 25803
rect 11036 25415 11094 25427
rect 11194 25803 11252 25815
rect 11194 25427 11206 25803
rect 11240 25427 11252 25803
rect 11194 25415 11252 25427
rect 11352 25803 11410 25815
rect 11352 25427 11364 25803
rect 11398 25427 11410 25803
rect 11352 25415 11410 25427
rect 11510 25803 11568 25815
rect 11510 25427 11522 25803
rect 11556 25427 11568 25803
rect 11510 25415 11568 25427
rect 11668 25803 11726 25815
rect 11668 25427 11680 25803
rect 11714 25427 11726 25803
rect 11668 25415 11726 25427
rect 11826 25803 11884 25815
rect 11826 25427 11838 25803
rect 11872 25427 11884 25803
rect 11826 25415 11884 25427
rect 11984 25803 12042 25815
rect 11984 25427 11996 25803
rect 12030 25427 12042 25803
rect 11984 25415 12042 25427
rect 12142 25803 12200 25815
rect 12142 25427 12154 25803
rect 12188 25427 12200 25803
rect 12142 25415 12200 25427
rect 12300 25803 12358 25815
rect 12300 25427 12312 25803
rect 12346 25427 12358 25803
rect 12300 25415 12358 25427
rect 12458 25803 12516 25815
rect 12458 25427 12470 25803
rect 12504 25427 12516 25803
rect 12458 25415 12516 25427
rect 13058 27075 13116 27087
rect 13058 26699 13070 27075
rect 13104 26699 13116 27075
rect 13058 26687 13116 26699
rect 13216 27075 13274 27087
rect 13216 26699 13228 27075
rect 13262 26699 13274 27075
rect 13216 26687 13274 26699
rect 13374 27075 13432 27087
rect 13374 26699 13386 27075
rect 13420 26699 13432 27075
rect 13374 26687 13432 26699
rect 13532 27075 13590 27087
rect 13532 26699 13544 27075
rect 13578 26699 13590 27075
rect 13532 26687 13590 26699
rect 13690 27075 13748 27087
rect 13690 26699 13702 27075
rect 13736 26699 13748 27075
rect 13690 26687 13748 26699
rect 13848 27075 13906 27087
rect 13848 26699 13860 27075
rect 13894 26699 13906 27075
rect 13848 26687 13906 26699
rect 14006 27075 14064 27087
rect 14006 26699 14018 27075
rect 14052 26699 14064 27075
rect 14006 26687 14064 26699
rect 14164 27075 14222 27087
rect 14164 26699 14176 27075
rect 14210 26699 14222 27075
rect 14164 26687 14222 26699
rect 14322 27075 14380 27087
rect 14322 26699 14334 27075
rect 14368 26699 14380 27075
rect 14322 26687 14380 26699
rect 14480 27075 14538 27087
rect 14480 26699 14492 27075
rect 14526 26699 14538 27075
rect 14480 26687 14538 26699
rect 14638 27075 14696 27087
rect 14638 26699 14650 27075
rect 14684 26699 14696 27075
rect 14638 26687 14696 26699
rect 13058 26439 13116 26451
rect 13058 26063 13070 26439
rect 13104 26063 13116 26439
rect 13058 26051 13116 26063
rect 13216 26439 13274 26451
rect 13216 26063 13228 26439
rect 13262 26063 13274 26439
rect 13216 26051 13274 26063
rect 13374 26439 13432 26451
rect 13374 26063 13386 26439
rect 13420 26063 13432 26439
rect 13374 26051 13432 26063
rect 13532 26439 13590 26451
rect 13532 26063 13544 26439
rect 13578 26063 13590 26439
rect 13532 26051 13590 26063
rect 13690 26439 13748 26451
rect 13690 26063 13702 26439
rect 13736 26063 13748 26439
rect 13690 26051 13748 26063
rect 13848 26439 13906 26451
rect 13848 26063 13860 26439
rect 13894 26063 13906 26439
rect 13848 26051 13906 26063
rect 14006 26439 14064 26451
rect 14006 26063 14018 26439
rect 14052 26063 14064 26439
rect 14006 26051 14064 26063
rect 14164 26439 14222 26451
rect 14164 26063 14176 26439
rect 14210 26063 14222 26439
rect 14164 26051 14222 26063
rect 14322 26439 14380 26451
rect 14322 26063 14334 26439
rect 14368 26063 14380 26439
rect 14322 26051 14380 26063
rect 14480 26439 14538 26451
rect 14480 26063 14492 26439
rect 14526 26063 14538 26439
rect 14480 26051 14538 26063
rect 14638 26439 14696 26451
rect 14638 26063 14650 26439
rect 14684 26063 14696 26439
rect 14638 26051 14696 26063
rect 13058 25803 13116 25815
rect 13058 25427 13070 25803
rect 13104 25427 13116 25803
rect 13058 25415 13116 25427
rect 13216 25803 13274 25815
rect 13216 25427 13228 25803
rect 13262 25427 13274 25803
rect 13216 25415 13274 25427
rect 13374 25803 13432 25815
rect 13374 25427 13386 25803
rect 13420 25427 13432 25803
rect 13374 25415 13432 25427
rect 13532 25803 13590 25815
rect 13532 25427 13544 25803
rect 13578 25427 13590 25803
rect 13532 25415 13590 25427
rect 13690 25803 13748 25815
rect 13690 25427 13702 25803
rect 13736 25427 13748 25803
rect 13690 25415 13748 25427
rect 13848 25803 13906 25815
rect 13848 25427 13860 25803
rect 13894 25427 13906 25803
rect 13848 25415 13906 25427
rect 14006 25803 14064 25815
rect 14006 25427 14018 25803
rect 14052 25427 14064 25803
rect 14006 25415 14064 25427
rect 14164 25803 14222 25815
rect 14164 25427 14176 25803
rect 14210 25427 14222 25803
rect 14164 25415 14222 25427
rect 14322 25803 14380 25815
rect 14322 25427 14334 25803
rect 14368 25427 14380 25803
rect 14322 25415 14380 25427
rect 14480 25803 14538 25815
rect 14480 25427 14492 25803
rect 14526 25427 14538 25803
rect 14480 25415 14538 25427
rect 14638 25803 14696 25815
rect 14638 25427 14650 25803
rect 14684 25427 14696 25803
rect 14638 25415 14696 25427
rect 15258 27075 15316 27087
rect 15258 26699 15270 27075
rect 15304 26699 15316 27075
rect 15258 26687 15316 26699
rect 15416 27075 15474 27087
rect 15416 26699 15428 27075
rect 15462 26699 15474 27075
rect 15416 26687 15474 26699
rect 15574 27075 15632 27087
rect 15574 26699 15586 27075
rect 15620 26699 15632 27075
rect 15574 26687 15632 26699
rect 15732 27075 15790 27087
rect 15732 26699 15744 27075
rect 15778 26699 15790 27075
rect 15732 26687 15790 26699
rect 15890 27075 15948 27087
rect 15890 26699 15902 27075
rect 15936 26699 15948 27075
rect 15890 26687 15948 26699
rect 16048 27075 16106 27087
rect 16048 26699 16060 27075
rect 16094 26699 16106 27075
rect 16048 26687 16106 26699
rect 16206 27075 16264 27087
rect 16206 26699 16218 27075
rect 16252 26699 16264 27075
rect 16206 26687 16264 26699
rect 16364 27075 16422 27087
rect 16364 26699 16376 27075
rect 16410 26699 16422 27075
rect 16364 26687 16422 26699
rect 16522 27075 16580 27087
rect 16522 26699 16534 27075
rect 16568 26699 16580 27075
rect 16522 26687 16580 26699
rect 16680 27075 16738 27087
rect 16680 26699 16692 27075
rect 16726 26699 16738 27075
rect 16680 26687 16738 26699
rect 16838 27075 16896 27087
rect 16838 26699 16850 27075
rect 16884 26699 16896 27075
rect 16838 26687 16896 26699
rect 15258 26439 15316 26451
rect 15258 26063 15270 26439
rect 15304 26063 15316 26439
rect 15258 26051 15316 26063
rect 15416 26439 15474 26451
rect 15416 26063 15428 26439
rect 15462 26063 15474 26439
rect 15416 26051 15474 26063
rect 15574 26439 15632 26451
rect 15574 26063 15586 26439
rect 15620 26063 15632 26439
rect 15574 26051 15632 26063
rect 15732 26439 15790 26451
rect 15732 26063 15744 26439
rect 15778 26063 15790 26439
rect 15732 26051 15790 26063
rect 15890 26439 15948 26451
rect 15890 26063 15902 26439
rect 15936 26063 15948 26439
rect 15890 26051 15948 26063
rect 16048 26439 16106 26451
rect 16048 26063 16060 26439
rect 16094 26063 16106 26439
rect 16048 26051 16106 26063
rect 16206 26439 16264 26451
rect 16206 26063 16218 26439
rect 16252 26063 16264 26439
rect 16206 26051 16264 26063
rect 16364 26439 16422 26451
rect 16364 26063 16376 26439
rect 16410 26063 16422 26439
rect 16364 26051 16422 26063
rect 16522 26439 16580 26451
rect 16522 26063 16534 26439
rect 16568 26063 16580 26439
rect 16522 26051 16580 26063
rect 16680 26439 16738 26451
rect 16680 26063 16692 26439
rect 16726 26063 16738 26439
rect 16680 26051 16738 26063
rect 16838 26439 16896 26451
rect 16838 26063 16850 26439
rect 16884 26063 16896 26439
rect 16838 26051 16896 26063
rect 15258 25803 15316 25815
rect 15258 25427 15270 25803
rect 15304 25427 15316 25803
rect 15258 25415 15316 25427
rect 15416 25803 15474 25815
rect 15416 25427 15428 25803
rect 15462 25427 15474 25803
rect 15416 25415 15474 25427
rect 15574 25803 15632 25815
rect 15574 25427 15586 25803
rect 15620 25427 15632 25803
rect 15574 25415 15632 25427
rect 15732 25803 15790 25815
rect 15732 25427 15744 25803
rect 15778 25427 15790 25803
rect 15732 25415 15790 25427
rect 15890 25803 15948 25815
rect 15890 25427 15902 25803
rect 15936 25427 15948 25803
rect 15890 25415 15948 25427
rect 16048 25803 16106 25815
rect 16048 25427 16060 25803
rect 16094 25427 16106 25803
rect 16048 25415 16106 25427
rect 16206 25803 16264 25815
rect 16206 25427 16218 25803
rect 16252 25427 16264 25803
rect 16206 25415 16264 25427
rect 16364 25803 16422 25815
rect 16364 25427 16376 25803
rect 16410 25427 16422 25803
rect 16364 25415 16422 25427
rect 16522 25803 16580 25815
rect 16522 25427 16534 25803
rect 16568 25427 16580 25803
rect 16522 25415 16580 25427
rect 16680 25803 16738 25815
rect 16680 25427 16692 25803
rect 16726 25427 16738 25803
rect 16680 25415 16738 25427
rect 16838 25803 16896 25815
rect 16838 25427 16850 25803
rect 16884 25427 16896 25803
rect 16838 25415 16896 25427
rect 6478 24979 6540 24991
rect 6478 24603 6490 24979
rect 6524 24603 6540 24979
rect 6478 24591 6540 24603
rect 6570 24979 6636 24991
rect 6570 24603 6586 24979
rect 6620 24603 6636 24979
rect 6570 24591 6636 24603
rect 6666 24979 6732 24991
rect 6666 24603 6682 24979
rect 6716 24603 6732 24979
rect 6666 24591 6732 24603
rect 6762 24979 6828 24991
rect 6762 24603 6778 24979
rect 6812 24603 6828 24979
rect 6762 24591 6828 24603
rect 6858 24979 6924 24991
rect 6858 24603 6874 24979
rect 6908 24603 6924 24979
rect 6858 24591 6924 24603
rect 6954 24979 7020 24991
rect 6954 24603 6970 24979
rect 7004 24603 7020 24979
rect 6954 24591 7020 24603
rect 7050 24979 7116 24991
rect 7050 24603 7066 24979
rect 7100 24603 7116 24979
rect 7050 24591 7116 24603
rect 7146 24979 7212 24991
rect 7146 24603 7162 24979
rect 7196 24603 7212 24979
rect 7146 24591 7212 24603
rect 7242 24979 7308 24991
rect 7242 24603 7258 24979
rect 7292 24603 7308 24979
rect 7242 24591 7308 24603
rect 7338 24979 7404 24991
rect 7338 24603 7354 24979
rect 7388 24603 7404 24979
rect 7338 24591 7404 24603
rect 7434 24979 7500 24991
rect 7434 24603 7450 24979
rect 7484 24603 7500 24979
rect 7434 24591 7500 24603
rect 7530 24979 7596 24991
rect 7530 24603 7546 24979
rect 7580 24603 7596 24979
rect 7530 24591 7596 24603
rect 7626 24979 7692 24991
rect 7626 24603 7642 24979
rect 7676 24603 7692 24979
rect 7626 24591 7692 24603
rect 7722 24979 7788 24991
rect 7722 24603 7738 24979
rect 7772 24603 7788 24979
rect 7722 24591 7788 24603
rect 7818 24979 7884 24991
rect 7818 24603 7834 24979
rect 7868 24603 7884 24979
rect 7818 24591 7884 24603
rect 7914 24979 7976 24991
rect 7914 24603 7930 24979
rect 7964 24603 7976 24979
rect 7914 24591 7976 24603
rect 6478 24343 6540 24355
rect 6478 23967 6490 24343
rect 6524 23967 6540 24343
rect 6478 23955 6540 23967
rect 6570 24343 6636 24355
rect 6570 23967 6586 24343
rect 6620 23967 6636 24343
rect 6570 23955 6636 23967
rect 6666 24343 6732 24355
rect 6666 23967 6682 24343
rect 6716 23967 6732 24343
rect 6666 23955 6732 23967
rect 6762 24343 6828 24355
rect 6762 23967 6778 24343
rect 6812 23967 6828 24343
rect 6762 23955 6828 23967
rect 6858 24343 6924 24355
rect 6858 23967 6874 24343
rect 6908 23967 6924 24343
rect 6858 23955 6924 23967
rect 6954 24343 7020 24355
rect 6954 23967 6970 24343
rect 7004 23967 7020 24343
rect 6954 23955 7020 23967
rect 7050 24343 7116 24355
rect 7050 23967 7066 24343
rect 7100 23967 7116 24343
rect 7050 23955 7116 23967
rect 7146 24343 7212 24355
rect 7146 23967 7162 24343
rect 7196 23967 7212 24343
rect 7146 23955 7212 23967
rect 7242 24343 7308 24355
rect 7242 23967 7258 24343
rect 7292 23967 7308 24343
rect 7242 23955 7308 23967
rect 7338 24343 7404 24355
rect 7338 23967 7354 24343
rect 7388 23967 7404 24343
rect 7338 23955 7404 23967
rect 7434 24343 7500 24355
rect 7434 23967 7450 24343
rect 7484 23967 7500 24343
rect 7434 23955 7500 23967
rect 7530 24343 7596 24355
rect 7530 23967 7546 24343
rect 7580 23967 7596 24343
rect 7530 23955 7596 23967
rect 7626 24343 7692 24355
rect 7626 23967 7642 24343
rect 7676 23967 7692 24343
rect 7626 23955 7692 23967
rect 7722 24343 7788 24355
rect 7722 23967 7738 24343
rect 7772 23967 7788 24343
rect 7722 23955 7788 23967
rect 7818 24343 7884 24355
rect 7818 23967 7834 24343
rect 7868 23967 7884 24343
rect 7818 23955 7884 23967
rect 7914 24343 7976 24355
rect 7914 23967 7930 24343
rect 7964 23967 7976 24343
rect 7914 23955 7976 23967
rect 8698 24979 8760 24991
rect 8698 24603 8710 24979
rect 8744 24603 8760 24979
rect 8698 24591 8760 24603
rect 8790 24979 8856 24991
rect 8790 24603 8806 24979
rect 8840 24603 8856 24979
rect 8790 24591 8856 24603
rect 8886 24979 8952 24991
rect 8886 24603 8902 24979
rect 8936 24603 8952 24979
rect 8886 24591 8952 24603
rect 8982 24979 9048 24991
rect 8982 24603 8998 24979
rect 9032 24603 9048 24979
rect 8982 24591 9048 24603
rect 9078 24979 9144 24991
rect 9078 24603 9094 24979
rect 9128 24603 9144 24979
rect 9078 24591 9144 24603
rect 9174 24979 9240 24991
rect 9174 24603 9190 24979
rect 9224 24603 9240 24979
rect 9174 24591 9240 24603
rect 9270 24979 9336 24991
rect 9270 24603 9286 24979
rect 9320 24603 9336 24979
rect 9270 24591 9336 24603
rect 9366 24979 9432 24991
rect 9366 24603 9382 24979
rect 9416 24603 9432 24979
rect 9366 24591 9432 24603
rect 9462 24979 9528 24991
rect 9462 24603 9478 24979
rect 9512 24603 9528 24979
rect 9462 24591 9528 24603
rect 9558 24979 9624 24991
rect 9558 24603 9574 24979
rect 9608 24603 9624 24979
rect 9558 24591 9624 24603
rect 9654 24979 9720 24991
rect 9654 24603 9670 24979
rect 9704 24603 9720 24979
rect 9654 24591 9720 24603
rect 9750 24979 9816 24991
rect 9750 24603 9766 24979
rect 9800 24603 9816 24979
rect 9750 24591 9816 24603
rect 9846 24979 9912 24991
rect 9846 24603 9862 24979
rect 9896 24603 9912 24979
rect 9846 24591 9912 24603
rect 9942 24979 10008 24991
rect 9942 24603 9958 24979
rect 9992 24603 10008 24979
rect 9942 24591 10008 24603
rect 10038 24979 10104 24991
rect 10038 24603 10054 24979
rect 10088 24603 10104 24979
rect 10038 24591 10104 24603
rect 10134 24979 10196 24991
rect 10134 24603 10150 24979
rect 10184 24603 10196 24979
rect 10134 24591 10196 24603
rect 8698 24343 8760 24355
rect 8698 23967 8710 24343
rect 8744 23967 8760 24343
rect 8698 23955 8760 23967
rect 8790 24343 8856 24355
rect 8790 23967 8806 24343
rect 8840 23967 8856 24343
rect 8790 23955 8856 23967
rect 8886 24343 8952 24355
rect 8886 23967 8902 24343
rect 8936 23967 8952 24343
rect 8886 23955 8952 23967
rect 8982 24343 9048 24355
rect 8982 23967 8998 24343
rect 9032 23967 9048 24343
rect 8982 23955 9048 23967
rect 9078 24343 9144 24355
rect 9078 23967 9094 24343
rect 9128 23967 9144 24343
rect 9078 23955 9144 23967
rect 9174 24343 9240 24355
rect 9174 23967 9190 24343
rect 9224 23967 9240 24343
rect 9174 23955 9240 23967
rect 9270 24343 9336 24355
rect 9270 23967 9286 24343
rect 9320 23967 9336 24343
rect 9270 23955 9336 23967
rect 9366 24343 9432 24355
rect 9366 23967 9382 24343
rect 9416 23967 9432 24343
rect 9366 23955 9432 23967
rect 9462 24343 9528 24355
rect 9462 23967 9478 24343
rect 9512 23967 9528 24343
rect 9462 23955 9528 23967
rect 9558 24343 9624 24355
rect 9558 23967 9574 24343
rect 9608 23967 9624 24343
rect 9558 23955 9624 23967
rect 9654 24343 9720 24355
rect 9654 23967 9670 24343
rect 9704 23967 9720 24343
rect 9654 23955 9720 23967
rect 9750 24343 9816 24355
rect 9750 23967 9766 24343
rect 9800 23967 9816 24343
rect 9750 23955 9816 23967
rect 9846 24343 9912 24355
rect 9846 23967 9862 24343
rect 9896 23967 9912 24343
rect 9846 23955 9912 23967
rect 9942 24343 10008 24355
rect 9942 23967 9958 24343
rect 9992 23967 10008 24343
rect 9942 23955 10008 23967
rect 10038 24343 10104 24355
rect 10038 23967 10054 24343
rect 10088 23967 10104 24343
rect 10038 23955 10104 23967
rect 10134 24343 10196 24355
rect 10134 23967 10150 24343
rect 10184 23967 10196 24343
rect 10134 23955 10196 23967
rect 10878 24979 10940 24991
rect 10878 24603 10890 24979
rect 10924 24603 10940 24979
rect 10878 24591 10940 24603
rect 10970 24979 11036 24991
rect 10970 24603 10986 24979
rect 11020 24603 11036 24979
rect 10970 24591 11036 24603
rect 11066 24979 11132 24991
rect 11066 24603 11082 24979
rect 11116 24603 11132 24979
rect 11066 24591 11132 24603
rect 11162 24979 11228 24991
rect 11162 24603 11178 24979
rect 11212 24603 11228 24979
rect 11162 24591 11228 24603
rect 11258 24979 11324 24991
rect 11258 24603 11274 24979
rect 11308 24603 11324 24979
rect 11258 24591 11324 24603
rect 11354 24979 11420 24991
rect 11354 24603 11370 24979
rect 11404 24603 11420 24979
rect 11354 24591 11420 24603
rect 11450 24979 11516 24991
rect 11450 24603 11466 24979
rect 11500 24603 11516 24979
rect 11450 24591 11516 24603
rect 11546 24979 11612 24991
rect 11546 24603 11562 24979
rect 11596 24603 11612 24979
rect 11546 24591 11612 24603
rect 11642 24979 11708 24991
rect 11642 24603 11658 24979
rect 11692 24603 11708 24979
rect 11642 24591 11708 24603
rect 11738 24979 11804 24991
rect 11738 24603 11754 24979
rect 11788 24603 11804 24979
rect 11738 24591 11804 24603
rect 11834 24979 11900 24991
rect 11834 24603 11850 24979
rect 11884 24603 11900 24979
rect 11834 24591 11900 24603
rect 11930 24979 11996 24991
rect 11930 24603 11946 24979
rect 11980 24603 11996 24979
rect 11930 24591 11996 24603
rect 12026 24979 12092 24991
rect 12026 24603 12042 24979
rect 12076 24603 12092 24979
rect 12026 24591 12092 24603
rect 12122 24979 12188 24991
rect 12122 24603 12138 24979
rect 12172 24603 12188 24979
rect 12122 24591 12188 24603
rect 12218 24979 12284 24991
rect 12218 24603 12234 24979
rect 12268 24603 12284 24979
rect 12218 24591 12284 24603
rect 12314 24979 12376 24991
rect 12314 24603 12330 24979
rect 12364 24603 12376 24979
rect 12314 24591 12376 24603
rect 10878 24343 10940 24355
rect 10878 23967 10890 24343
rect 10924 23967 10940 24343
rect 10878 23955 10940 23967
rect 10970 24343 11036 24355
rect 10970 23967 10986 24343
rect 11020 23967 11036 24343
rect 10970 23955 11036 23967
rect 11066 24343 11132 24355
rect 11066 23967 11082 24343
rect 11116 23967 11132 24343
rect 11066 23955 11132 23967
rect 11162 24343 11228 24355
rect 11162 23967 11178 24343
rect 11212 23967 11228 24343
rect 11162 23955 11228 23967
rect 11258 24343 11324 24355
rect 11258 23967 11274 24343
rect 11308 23967 11324 24343
rect 11258 23955 11324 23967
rect 11354 24343 11420 24355
rect 11354 23967 11370 24343
rect 11404 23967 11420 24343
rect 11354 23955 11420 23967
rect 11450 24343 11516 24355
rect 11450 23967 11466 24343
rect 11500 23967 11516 24343
rect 11450 23955 11516 23967
rect 11546 24343 11612 24355
rect 11546 23967 11562 24343
rect 11596 23967 11612 24343
rect 11546 23955 11612 23967
rect 11642 24343 11708 24355
rect 11642 23967 11658 24343
rect 11692 23967 11708 24343
rect 11642 23955 11708 23967
rect 11738 24343 11804 24355
rect 11738 23967 11754 24343
rect 11788 23967 11804 24343
rect 11738 23955 11804 23967
rect 11834 24343 11900 24355
rect 11834 23967 11850 24343
rect 11884 23967 11900 24343
rect 11834 23955 11900 23967
rect 11930 24343 11996 24355
rect 11930 23967 11946 24343
rect 11980 23967 11996 24343
rect 11930 23955 11996 23967
rect 12026 24343 12092 24355
rect 12026 23967 12042 24343
rect 12076 23967 12092 24343
rect 12026 23955 12092 23967
rect 12122 24343 12188 24355
rect 12122 23967 12138 24343
rect 12172 23967 12188 24343
rect 12122 23955 12188 23967
rect 12218 24343 12284 24355
rect 12218 23967 12234 24343
rect 12268 23967 12284 24343
rect 12218 23955 12284 23967
rect 12314 24343 12376 24355
rect 12314 23967 12330 24343
rect 12364 23967 12376 24343
rect 12314 23955 12376 23967
rect 13058 24979 13120 24991
rect 13058 24603 13070 24979
rect 13104 24603 13120 24979
rect 13058 24591 13120 24603
rect 13150 24979 13216 24991
rect 13150 24603 13166 24979
rect 13200 24603 13216 24979
rect 13150 24591 13216 24603
rect 13246 24979 13312 24991
rect 13246 24603 13262 24979
rect 13296 24603 13312 24979
rect 13246 24591 13312 24603
rect 13342 24979 13408 24991
rect 13342 24603 13358 24979
rect 13392 24603 13408 24979
rect 13342 24591 13408 24603
rect 13438 24979 13504 24991
rect 13438 24603 13454 24979
rect 13488 24603 13504 24979
rect 13438 24591 13504 24603
rect 13534 24979 13600 24991
rect 13534 24603 13550 24979
rect 13584 24603 13600 24979
rect 13534 24591 13600 24603
rect 13630 24979 13696 24991
rect 13630 24603 13646 24979
rect 13680 24603 13696 24979
rect 13630 24591 13696 24603
rect 13726 24979 13792 24991
rect 13726 24603 13742 24979
rect 13776 24603 13792 24979
rect 13726 24591 13792 24603
rect 13822 24979 13888 24991
rect 13822 24603 13838 24979
rect 13872 24603 13888 24979
rect 13822 24591 13888 24603
rect 13918 24979 13984 24991
rect 13918 24603 13934 24979
rect 13968 24603 13984 24979
rect 13918 24591 13984 24603
rect 14014 24979 14080 24991
rect 14014 24603 14030 24979
rect 14064 24603 14080 24979
rect 14014 24591 14080 24603
rect 14110 24979 14176 24991
rect 14110 24603 14126 24979
rect 14160 24603 14176 24979
rect 14110 24591 14176 24603
rect 14206 24979 14272 24991
rect 14206 24603 14222 24979
rect 14256 24603 14272 24979
rect 14206 24591 14272 24603
rect 14302 24979 14368 24991
rect 14302 24603 14318 24979
rect 14352 24603 14368 24979
rect 14302 24591 14368 24603
rect 14398 24979 14464 24991
rect 14398 24603 14414 24979
rect 14448 24603 14464 24979
rect 14398 24591 14464 24603
rect 14494 24979 14556 24991
rect 14494 24603 14510 24979
rect 14544 24603 14556 24979
rect 14494 24591 14556 24603
rect 13058 24343 13120 24355
rect 13058 23967 13070 24343
rect 13104 23967 13120 24343
rect 13058 23955 13120 23967
rect 13150 24343 13216 24355
rect 13150 23967 13166 24343
rect 13200 23967 13216 24343
rect 13150 23955 13216 23967
rect 13246 24343 13312 24355
rect 13246 23967 13262 24343
rect 13296 23967 13312 24343
rect 13246 23955 13312 23967
rect 13342 24343 13408 24355
rect 13342 23967 13358 24343
rect 13392 23967 13408 24343
rect 13342 23955 13408 23967
rect 13438 24343 13504 24355
rect 13438 23967 13454 24343
rect 13488 23967 13504 24343
rect 13438 23955 13504 23967
rect 13534 24343 13600 24355
rect 13534 23967 13550 24343
rect 13584 23967 13600 24343
rect 13534 23955 13600 23967
rect 13630 24343 13696 24355
rect 13630 23967 13646 24343
rect 13680 23967 13696 24343
rect 13630 23955 13696 23967
rect 13726 24343 13792 24355
rect 13726 23967 13742 24343
rect 13776 23967 13792 24343
rect 13726 23955 13792 23967
rect 13822 24343 13888 24355
rect 13822 23967 13838 24343
rect 13872 23967 13888 24343
rect 13822 23955 13888 23967
rect 13918 24343 13984 24355
rect 13918 23967 13934 24343
rect 13968 23967 13984 24343
rect 13918 23955 13984 23967
rect 14014 24343 14080 24355
rect 14014 23967 14030 24343
rect 14064 23967 14080 24343
rect 14014 23955 14080 23967
rect 14110 24343 14176 24355
rect 14110 23967 14126 24343
rect 14160 23967 14176 24343
rect 14110 23955 14176 23967
rect 14206 24343 14272 24355
rect 14206 23967 14222 24343
rect 14256 23967 14272 24343
rect 14206 23955 14272 23967
rect 14302 24343 14368 24355
rect 14302 23967 14318 24343
rect 14352 23967 14368 24343
rect 14302 23955 14368 23967
rect 14398 24343 14464 24355
rect 14398 23967 14414 24343
rect 14448 23967 14464 24343
rect 14398 23955 14464 23967
rect 14494 24343 14556 24355
rect 14494 23967 14510 24343
rect 14544 23967 14556 24343
rect 14494 23955 14556 23967
rect 15258 24979 15320 24991
rect 15258 24603 15270 24979
rect 15304 24603 15320 24979
rect 15258 24591 15320 24603
rect 15350 24979 15416 24991
rect 15350 24603 15366 24979
rect 15400 24603 15416 24979
rect 15350 24591 15416 24603
rect 15446 24979 15512 24991
rect 15446 24603 15462 24979
rect 15496 24603 15512 24979
rect 15446 24591 15512 24603
rect 15542 24979 15608 24991
rect 15542 24603 15558 24979
rect 15592 24603 15608 24979
rect 15542 24591 15608 24603
rect 15638 24979 15704 24991
rect 15638 24603 15654 24979
rect 15688 24603 15704 24979
rect 15638 24591 15704 24603
rect 15734 24979 15800 24991
rect 15734 24603 15750 24979
rect 15784 24603 15800 24979
rect 15734 24591 15800 24603
rect 15830 24979 15896 24991
rect 15830 24603 15846 24979
rect 15880 24603 15896 24979
rect 15830 24591 15896 24603
rect 15926 24979 15992 24991
rect 15926 24603 15942 24979
rect 15976 24603 15992 24979
rect 15926 24591 15992 24603
rect 16022 24979 16088 24991
rect 16022 24603 16038 24979
rect 16072 24603 16088 24979
rect 16022 24591 16088 24603
rect 16118 24979 16184 24991
rect 16118 24603 16134 24979
rect 16168 24603 16184 24979
rect 16118 24591 16184 24603
rect 16214 24979 16280 24991
rect 16214 24603 16230 24979
rect 16264 24603 16280 24979
rect 16214 24591 16280 24603
rect 16310 24979 16376 24991
rect 16310 24603 16326 24979
rect 16360 24603 16376 24979
rect 16310 24591 16376 24603
rect 16406 24979 16472 24991
rect 16406 24603 16422 24979
rect 16456 24603 16472 24979
rect 16406 24591 16472 24603
rect 16502 24979 16568 24991
rect 16502 24603 16518 24979
rect 16552 24603 16568 24979
rect 16502 24591 16568 24603
rect 16598 24979 16664 24991
rect 16598 24603 16614 24979
rect 16648 24603 16664 24979
rect 16598 24591 16664 24603
rect 16694 24979 16756 24991
rect 16694 24603 16710 24979
rect 16744 24603 16756 24979
rect 16694 24591 16756 24603
rect 15258 24343 15320 24355
rect 15258 23967 15270 24343
rect 15304 23967 15320 24343
rect 15258 23955 15320 23967
rect 15350 24343 15416 24355
rect 15350 23967 15366 24343
rect 15400 23967 15416 24343
rect 15350 23955 15416 23967
rect 15446 24343 15512 24355
rect 15446 23967 15462 24343
rect 15496 23967 15512 24343
rect 15446 23955 15512 23967
rect 15542 24343 15608 24355
rect 15542 23967 15558 24343
rect 15592 23967 15608 24343
rect 15542 23955 15608 23967
rect 15638 24343 15704 24355
rect 15638 23967 15654 24343
rect 15688 23967 15704 24343
rect 15638 23955 15704 23967
rect 15734 24343 15800 24355
rect 15734 23967 15750 24343
rect 15784 23967 15800 24343
rect 15734 23955 15800 23967
rect 15830 24343 15896 24355
rect 15830 23967 15846 24343
rect 15880 23967 15896 24343
rect 15830 23955 15896 23967
rect 15926 24343 15992 24355
rect 15926 23967 15942 24343
rect 15976 23967 15992 24343
rect 15926 23955 15992 23967
rect 16022 24343 16088 24355
rect 16022 23967 16038 24343
rect 16072 23967 16088 24343
rect 16022 23955 16088 23967
rect 16118 24343 16184 24355
rect 16118 23967 16134 24343
rect 16168 23967 16184 24343
rect 16118 23955 16184 23967
rect 16214 24343 16280 24355
rect 16214 23967 16230 24343
rect 16264 23967 16280 24343
rect 16214 23955 16280 23967
rect 16310 24343 16376 24355
rect 16310 23967 16326 24343
rect 16360 23967 16376 24343
rect 16310 23955 16376 23967
rect 16406 24343 16472 24355
rect 16406 23967 16422 24343
rect 16456 23967 16472 24343
rect 16406 23955 16472 23967
rect 16502 24343 16568 24355
rect 16502 23967 16518 24343
rect 16552 23967 16568 24343
rect 16502 23955 16568 23967
rect 16598 24343 16664 24355
rect 16598 23967 16614 24343
rect 16648 23967 16664 24343
rect 16598 23955 16664 23967
rect 16694 24343 16756 24355
rect 16694 23967 16710 24343
rect 16744 23967 16756 24343
rect 16694 23955 16756 23967
rect 19039 25082 19239 25094
rect 19039 25048 19051 25082
rect 19227 25048 19239 25082
rect 19039 25036 19239 25048
rect 19039 23424 19239 23436
rect 19039 23390 19051 23424
rect 19227 23390 19239 23424
rect 19039 23378 19239 23390
rect 18298 23011 18360 23023
rect 18298 22635 18310 23011
rect 18344 22635 18360 23011
rect 18298 22623 18360 22635
rect 18390 23011 18456 23023
rect 18390 22635 18406 23011
rect 18440 22635 18456 23011
rect 18390 22623 18456 22635
rect 18486 23011 18552 23023
rect 18486 22635 18502 23011
rect 18536 22635 18552 23011
rect 18486 22623 18552 22635
rect 18582 23011 18648 23023
rect 18582 22635 18598 23011
rect 18632 22635 18648 23011
rect 18582 22623 18648 22635
rect 18678 23011 18744 23023
rect 18678 22635 18694 23011
rect 18728 22635 18744 23011
rect 18678 22623 18744 22635
rect 18774 23011 18840 23023
rect 18774 22635 18790 23011
rect 18824 22635 18840 23011
rect 18774 22623 18840 22635
rect 18870 23011 18936 23023
rect 18870 22635 18886 23011
rect 18920 22635 18936 23011
rect 18870 22623 18936 22635
rect 18966 23011 19032 23023
rect 18966 22635 18982 23011
rect 19016 22635 19032 23011
rect 18966 22623 19032 22635
rect 19062 23011 19128 23023
rect 19062 22635 19078 23011
rect 19112 22635 19128 23011
rect 19062 22623 19128 22635
rect 19158 23011 19224 23023
rect 19158 22635 19174 23011
rect 19208 22635 19224 23011
rect 19158 22623 19224 22635
rect 19254 23011 19316 23023
rect 19254 22635 19270 23011
rect 19304 22635 19316 23011
rect 19254 22623 19316 22635
rect 5114 10271 5176 10283
rect 5114 9895 5126 10271
rect 5160 9895 5176 10271
rect 5114 9883 5176 9895
rect 5206 10271 5272 10283
rect 5206 9895 5222 10271
rect 5256 9895 5272 10271
rect 5206 9883 5272 9895
rect 5302 10271 5368 10283
rect 5302 9895 5318 10271
rect 5352 9895 5368 10271
rect 5302 9883 5368 9895
rect 5398 10271 5464 10283
rect 5398 9895 5414 10271
rect 5448 9895 5464 10271
rect 5398 9883 5464 9895
rect 5494 10271 5560 10283
rect 5494 9895 5510 10271
rect 5544 9895 5560 10271
rect 5494 9883 5560 9895
rect 5590 10271 5656 10283
rect 5590 9895 5606 10271
rect 5640 9895 5656 10271
rect 5590 9883 5656 9895
rect 5686 10271 5752 10283
rect 5686 9895 5702 10271
rect 5736 9895 5752 10271
rect 5686 9883 5752 9895
rect 5782 10271 5848 10283
rect 5782 9895 5798 10271
rect 5832 9895 5848 10271
rect 5782 9883 5848 9895
rect 5878 10271 5944 10283
rect 5878 9895 5894 10271
rect 5928 9895 5944 10271
rect 5878 9883 5944 9895
rect 5974 10271 6040 10283
rect 5974 9895 5990 10271
rect 6024 9895 6040 10271
rect 5974 9883 6040 9895
rect 6070 10271 6136 10283
rect 6070 9895 6086 10271
rect 6120 9895 6136 10271
rect 6070 9883 6136 9895
rect 6166 10271 6232 10283
rect 6166 9895 6182 10271
rect 6216 9895 6232 10271
rect 6166 9883 6232 9895
rect 6262 10271 6328 10283
rect 6262 9895 6278 10271
rect 6312 9895 6328 10271
rect 6262 9883 6328 9895
rect 6358 10271 6424 10283
rect 6358 9895 6374 10271
rect 6408 9895 6424 10271
rect 6358 9883 6424 9895
rect 6454 10271 6520 10283
rect 6454 9895 6470 10271
rect 6504 9895 6520 10271
rect 6454 9883 6520 9895
rect 6550 10271 6616 10283
rect 6550 9895 6566 10271
rect 6600 9895 6616 10271
rect 6550 9883 6616 9895
rect 6646 10271 6712 10283
rect 6646 9895 6662 10271
rect 6696 9895 6712 10271
rect 6646 9883 6712 9895
rect 6742 10271 6808 10283
rect 6742 9895 6758 10271
rect 6792 9895 6808 10271
rect 6742 9883 6808 9895
rect 6838 10271 6904 10283
rect 6838 9895 6854 10271
rect 6888 9895 6904 10271
rect 6838 9883 6904 9895
rect 6934 10271 7000 10283
rect 6934 9895 6950 10271
rect 6984 9895 7000 10271
rect 6934 9883 7000 9895
rect 7030 10271 7092 10283
rect 7030 9895 7046 10271
rect 7080 9895 7092 10271
rect 7030 9883 7092 9895
rect 5114 9635 5176 9647
rect 5114 9259 5126 9635
rect 5160 9259 5176 9635
rect 5114 9247 5176 9259
rect 5206 9635 5272 9647
rect 5206 9259 5222 9635
rect 5256 9259 5272 9635
rect 5206 9247 5272 9259
rect 5302 9635 5368 9647
rect 5302 9259 5318 9635
rect 5352 9259 5368 9635
rect 5302 9247 5368 9259
rect 5398 9635 5464 9647
rect 5398 9259 5414 9635
rect 5448 9259 5464 9635
rect 5398 9247 5464 9259
rect 5494 9635 5560 9647
rect 5494 9259 5510 9635
rect 5544 9259 5560 9635
rect 5494 9247 5560 9259
rect 5590 9635 5656 9647
rect 5590 9259 5606 9635
rect 5640 9259 5656 9635
rect 5590 9247 5656 9259
rect 5686 9635 5752 9647
rect 5686 9259 5702 9635
rect 5736 9259 5752 9635
rect 5686 9247 5752 9259
rect 5782 9635 5848 9647
rect 5782 9259 5798 9635
rect 5832 9259 5848 9635
rect 5782 9247 5848 9259
rect 5878 9635 5944 9647
rect 5878 9259 5894 9635
rect 5928 9259 5944 9635
rect 5878 9247 5944 9259
rect 5974 9635 6040 9647
rect 5974 9259 5990 9635
rect 6024 9259 6040 9635
rect 5974 9247 6040 9259
rect 6070 9635 6136 9647
rect 6070 9259 6086 9635
rect 6120 9259 6136 9635
rect 6070 9247 6136 9259
rect 6166 9635 6232 9647
rect 6166 9259 6182 9635
rect 6216 9259 6232 9635
rect 6166 9247 6232 9259
rect 6262 9635 6328 9647
rect 6262 9259 6278 9635
rect 6312 9259 6328 9635
rect 6262 9247 6328 9259
rect 6358 9635 6424 9647
rect 6358 9259 6374 9635
rect 6408 9259 6424 9635
rect 6358 9247 6424 9259
rect 6454 9635 6520 9647
rect 6454 9259 6470 9635
rect 6504 9259 6520 9635
rect 6454 9247 6520 9259
rect 6550 9635 6616 9647
rect 6550 9259 6566 9635
rect 6600 9259 6616 9635
rect 6550 9247 6616 9259
rect 6646 9635 6712 9647
rect 6646 9259 6662 9635
rect 6696 9259 6712 9635
rect 6646 9247 6712 9259
rect 6742 9635 6808 9647
rect 6742 9259 6758 9635
rect 6792 9259 6808 9635
rect 6742 9247 6808 9259
rect 6838 9635 6904 9647
rect 6838 9259 6854 9635
rect 6888 9259 6904 9635
rect 6838 9247 6904 9259
rect 6934 9635 7000 9647
rect 6934 9259 6950 9635
rect 6984 9259 7000 9635
rect 6934 9247 7000 9259
rect 7030 9635 7092 9647
rect 7030 9259 7046 9635
rect 7080 9259 7092 9635
rect 7030 9247 7092 9259
rect 19514 10271 19576 10283
rect 19514 9895 19526 10271
rect 19560 9895 19576 10271
rect 19514 9883 19576 9895
rect 19606 10271 19672 10283
rect 19606 9895 19622 10271
rect 19656 9895 19672 10271
rect 19606 9883 19672 9895
rect 19702 10271 19768 10283
rect 19702 9895 19718 10271
rect 19752 9895 19768 10271
rect 19702 9883 19768 9895
rect 19798 10271 19864 10283
rect 19798 9895 19814 10271
rect 19848 9895 19864 10271
rect 19798 9883 19864 9895
rect 19894 10271 19960 10283
rect 19894 9895 19910 10271
rect 19944 9895 19960 10271
rect 19894 9883 19960 9895
rect 19990 10271 20056 10283
rect 19990 9895 20006 10271
rect 20040 9895 20056 10271
rect 19990 9883 20056 9895
rect 20086 10271 20152 10283
rect 20086 9895 20102 10271
rect 20136 9895 20152 10271
rect 20086 9883 20152 9895
rect 20182 10271 20248 10283
rect 20182 9895 20198 10271
rect 20232 9895 20248 10271
rect 20182 9883 20248 9895
rect 20278 10271 20344 10283
rect 20278 9895 20294 10271
rect 20328 9895 20344 10271
rect 20278 9883 20344 9895
rect 20374 10271 20440 10283
rect 20374 9895 20390 10271
rect 20424 9895 20440 10271
rect 20374 9883 20440 9895
rect 20470 10271 20536 10283
rect 20470 9895 20486 10271
rect 20520 9895 20536 10271
rect 20470 9883 20536 9895
rect 20566 10271 20632 10283
rect 20566 9895 20582 10271
rect 20616 9895 20632 10271
rect 20566 9883 20632 9895
rect 20662 10271 20728 10283
rect 20662 9895 20678 10271
rect 20712 9895 20728 10271
rect 20662 9883 20728 9895
rect 20758 10271 20824 10283
rect 20758 9895 20774 10271
rect 20808 9895 20824 10271
rect 20758 9883 20824 9895
rect 20854 10271 20920 10283
rect 20854 9895 20870 10271
rect 20904 9895 20920 10271
rect 20854 9883 20920 9895
rect 20950 10271 21016 10283
rect 20950 9895 20966 10271
rect 21000 9895 21016 10271
rect 20950 9883 21016 9895
rect 21046 10271 21112 10283
rect 21046 9895 21062 10271
rect 21096 9895 21112 10271
rect 21046 9883 21112 9895
rect 21142 10271 21208 10283
rect 21142 9895 21158 10271
rect 21192 9895 21208 10271
rect 21142 9883 21208 9895
rect 21238 10271 21304 10283
rect 21238 9895 21254 10271
rect 21288 9895 21304 10271
rect 21238 9883 21304 9895
rect 21334 10271 21400 10283
rect 21334 9895 21350 10271
rect 21384 9895 21400 10271
rect 21334 9883 21400 9895
rect 21430 10271 21492 10283
rect 21430 9895 21446 10271
rect 21480 9895 21492 10271
rect 21430 9883 21492 9895
rect 19514 9635 19576 9647
rect 19514 9259 19526 9635
rect 19560 9259 19576 9635
rect 19514 9247 19576 9259
rect 19606 9635 19672 9647
rect 19606 9259 19622 9635
rect 19656 9259 19672 9635
rect 19606 9247 19672 9259
rect 19702 9635 19768 9647
rect 19702 9259 19718 9635
rect 19752 9259 19768 9635
rect 19702 9247 19768 9259
rect 19798 9635 19864 9647
rect 19798 9259 19814 9635
rect 19848 9259 19864 9635
rect 19798 9247 19864 9259
rect 19894 9635 19960 9647
rect 19894 9259 19910 9635
rect 19944 9259 19960 9635
rect 19894 9247 19960 9259
rect 19990 9635 20056 9647
rect 19990 9259 20006 9635
rect 20040 9259 20056 9635
rect 19990 9247 20056 9259
rect 20086 9635 20152 9647
rect 20086 9259 20102 9635
rect 20136 9259 20152 9635
rect 20086 9247 20152 9259
rect 20182 9635 20248 9647
rect 20182 9259 20198 9635
rect 20232 9259 20248 9635
rect 20182 9247 20248 9259
rect 20278 9635 20344 9647
rect 20278 9259 20294 9635
rect 20328 9259 20344 9635
rect 20278 9247 20344 9259
rect 20374 9635 20440 9647
rect 20374 9259 20390 9635
rect 20424 9259 20440 9635
rect 20374 9247 20440 9259
rect 20470 9635 20536 9647
rect 20470 9259 20486 9635
rect 20520 9259 20536 9635
rect 20470 9247 20536 9259
rect 20566 9635 20632 9647
rect 20566 9259 20582 9635
rect 20616 9259 20632 9635
rect 20566 9247 20632 9259
rect 20662 9635 20728 9647
rect 20662 9259 20678 9635
rect 20712 9259 20728 9635
rect 20662 9247 20728 9259
rect 20758 9635 20824 9647
rect 20758 9259 20774 9635
rect 20808 9259 20824 9635
rect 20758 9247 20824 9259
rect 20854 9635 20920 9647
rect 20854 9259 20870 9635
rect 20904 9259 20920 9635
rect 20854 9247 20920 9259
rect 20950 9635 21016 9647
rect 20950 9259 20966 9635
rect 21000 9259 21016 9635
rect 20950 9247 21016 9259
rect 21046 9635 21112 9647
rect 21046 9259 21062 9635
rect 21096 9259 21112 9635
rect 21046 9247 21112 9259
rect 21142 9635 21208 9647
rect 21142 9259 21158 9635
rect 21192 9259 21208 9635
rect 21142 9247 21208 9259
rect 21238 9635 21304 9647
rect 21238 9259 21254 9635
rect 21288 9259 21304 9635
rect 21238 9247 21304 9259
rect 21334 9635 21400 9647
rect 21334 9259 21350 9635
rect 21384 9259 21400 9635
rect 21334 9247 21400 9259
rect 21430 9635 21492 9647
rect 21430 9259 21446 9635
rect 21480 9259 21492 9635
rect 21430 9247 21492 9259
<< ndiffc >>
rect 6610 23034 6644 23410
rect 6706 23034 6740 23410
rect 6802 23034 6836 23410
rect 6898 23034 6932 23410
rect 6994 23034 7028 23410
rect 7090 23034 7124 23410
rect 7186 23034 7220 23410
rect 7282 23034 7316 23410
rect 7378 23034 7412 23410
rect 7474 23034 7508 23410
rect 7570 23034 7604 23410
rect 6610 22416 6644 22792
rect 6706 22416 6740 22792
rect 6802 22416 6836 22792
rect 6898 22416 6932 22792
rect 6994 22416 7028 22792
rect 7090 22416 7124 22792
rect 7186 22416 7220 22792
rect 7282 22416 7316 22792
rect 7378 22416 7412 22792
rect 7474 22416 7508 22792
rect 7570 22416 7604 22792
rect 6610 21798 6644 22174
rect 6706 21798 6740 22174
rect 6802 21798 6836 22174
rect 6898 21798 6932 22174
rect 6994 21798 7028 22174
rect 7090 21798 7124 22174
rect 7186 21798 7220 22174
rect 7282 21798 7316 22174
rect 7378 21798 7412 22174
rect 7474 21798 7508 22174
rect 7570 21798 7604 22174
rect 8330 23034 8364 23410
rect 8426 23034 8460 23410
rect 8522 23034 8556 23410
rect 8618 23034 8652 23410
rect 8714 23034 8748 23410
rect 8810 23034 8844 23410
rect 8906 23034 8940 23410
rect 9002 23034 9036 23410
rect 9098 23034 9132 23410
rect 9194 23034 9228 23410
rect 9290 23034 9324 23410
rect 8330 22416 8364 22792
rect 8426 22416 8460 22792
rect 8522 22416 8556 22792
rect 8618 22416 8652 22792
rect 8714 22416 8748 22792
rect 8810 22416 8844 22792
rect 8906 22416 8940 22792
rect 9002 22416 9036 22792
rect 9098 22416 9132 22792
rect 9194 22416 9228 22792
rect 9290 22416 9324 22792
rect 8330 21798 8364 22174
rect 8426 21798 8460 22174
rect 8522 21798 8556 22174
rect 8618 21798 8652 22174
rect 8714 21798 8748 22174
rect 8810 21798 8844 22174
rect 8906 21798 8940 22174
rect 9002 21798 9036 22174
rect 9098 21798 9132 22174
rect 9194 21798 9228 22174
rect 9290 21798 9324 22174
rect 6610 20888 6644 21264
rect 6868 20888 6902 21264
rect 7126 20888 7160 21264
rect 7384 20888 7418 21264
rect 7642 20888 7676 21264
rect 7900 20888 7934 21264
rect 6610 20270 6644 20646
rect 6868 20270 6902 20646
rect 7126 20270 7160 20646
rect 7384 20270 7418 20646
rect 7642 20270 7676 20646
rect 7900 20270 7934 20646
rect 6610 19652 6644 20028
rect 6868 19652 6902 20028
rect 7126 19652 7160 20028
rect 7384 19652 7418 20028
rect 7642 19652 7676 20028
rect 7900 19652 7934 20028
rect 6610 19034 6644 19410
rect 6868 19034 6902 19410
rect 7126 19034 7160 19410
rect 7384 19034 7418 19410
rect 7642 19034 7676 19410
rect 7900 19034 7934 19410
rect 6610 18416 6644 18792
rect 6868 18416 6902 18792
rect 7126 18416 7160 18792
rect 7384 18416 7418 18792
rect 7642 18416 7676 18792
rect 7900 18416 7934 18792
rect 6610 17798 6644 18174
rect 6868 17798 6902 18174
rect 7126 17798 7160 18174
rect 7384 17798 7418 18174
rect 7642 17798 7676 18174
rect 7900 17798 7934 18174
rect 8330 20888 8364 21264
rect 8588 20888 8622 21264
rect 8846 20888 8880 21264
rect 9104 20888 9138 21264
rect 9362 20888 9396 21264
rect 9620 20888 9654 21264
rect 8330 20270 8364 20646
rect 8588 20270 8622 20646
rect 8846 20270 8880 20646
rect 9104 20270 9138 20646
rect 9362 20270 9396 20646
rect 9620 20270 9654 20646
rect 8330 19652 8364 20028
rect 8588 19652 8622 20028
rect 8846 19652 8880 20028
rect 9104 19652 9138 20028
rect 9362 19652 9396 20028
rect 9620 19652 9654 20028
rect 8330 19034 8364 19410
rect 8588 19034 8622 19410
rect 8846 19034 8880 19410
rect 9104 19034 9138 19410
rect 9362 19034 9396 19410
rect 9620 19034 9654 19410
rect 8330 18416 8364 18792
rect 8588 18416 8622 18792
rect 8846 18416 8880 18792
rect 9104 18416 9138 18792
rect 9362 18416 9396 18792
rect 9620 18416 9654 18792
rect 8330 17798 8364 18174
rect 8588 17798 8622 18174
rect 8846 17798 8880 18174
rect 9104 17798 9138 18174
rect 9362 17798 9396 18174
rect 9620 17798 9654 18174
rect 18310 21776 18344 22152
rect 18406 21776 18440 22152
rect 18502 21776 18536 22152
rect 18598 21776 18632 22152
rect 18694 21776 18728 22152
rect 18790 21776 18824 22152
rect 18886 21776 18920 22152
rect 18982 21776 19016 22152
rect 19078 21776 19112 22152
rect 19174 21776 19208 22152
rect 19270 21776 19304 22152
rect 18310 21158 18344 21534
rect 18406 21158 18440 21534
rect 18502 21158 18536 21534
rect 18598 21158 18632 21534
rect 18694 21158 18728 21534
rect 18790 21158 18824 21534
rect 18886 21158 18920 21534
rect 18982 21158 19016 21534
rect 19078 21158 19112 21534
rect 19174 21158 19208 21534
rect 19270 21158 19304 21534
rect 10170 19338 10204 19714
rect 10266 19338 10300 19714
rect 10362 19338 10396 19714
rect 10458 19338 10492 19714
rect 10554 19338 10588 19714
rect 10650 19338 10684 19714
rect 10746 19338 10780 19714
rect 10842 19338 10876 19714
rect 10170 18416 10204 18792
rect 10266 18416 10300 18792
rect 10362 18416 10396 18792
rect 10458 18416 10492 18792
rect 10554 18416 10588 18792
rect 10650 18416 10684 18792
rect 10746 18416 10780 18792
rect 10842 18416 10876 18792
rect 10938 18416 10972 18792
rect 11034 18416 11068 18792
rect 11130 18416 11164 18792
rect 10170 17798 10204 18174
rect 10266 17798 10300 18174
rect 10362 17798 10396 18174
rect 10458 17798 10492 18174
rect 10554 17798 10588 18174
rect 10650 17798 10684 18174
rect 10746 17798 10780 18174
rect 10842 17798 10876 18174
rect 10938 17798 10972 18174
rect 11034 17798 11068 18174
rect 11130 17798 11164 18174
rect 18310 20292 18344 20668
rect 18568 20292 18602 20668
rect 18826 20292 18860 20668
rect 19084 20292 19118 20668
rect 19342 20292 19376 20668
rect 19600 20292 19634 20668
rect 18310 19674 18344 20050
rect 18568 19674 18602 20050
rect 18826 19674 18860 20050
rect 19084 19674 19118 20050
rect 19342 19674 19376 20050
rect 19600 19674 19634 20050
rect 18310 19056 18344 19432
rect 18568 19056 18602 19432
rect 18826 19056 18860 19432
rect 19084 19056 19118 19432
rect 19342 19056 19376 19432
rect 19600 19056 19634 19432
rect 18310 18438 18344 18814
rect 18568 18438 18602 18814
rect 18826 18438 18860 18814
rect 19084 18438 19118 18814
rect 19342 18438 19376 18814
rect 19600 18438 19634 18814
rect -10050 7846 -10016 8222
rect -9954 7846 -9920 8222
rect -9858 7846 -9824 8222
rect -9762 7846 -9728 8222
rect -9666 7846 -9632 8222
rect -9570 7846 -9536 8222
rect -9474 7846 -9440 8222
rect -9378 7846 -9344 8222
rect -9282 7846 -9248 8222
rect -9186 7846 -9152 8222
rect -9090 7846 -9056 8222
rect -10050 7228 -10016 7604
rect -9954 7228 -9920 7604
rect -9858 7228 -9824 7604
rect -9762 7228 -9728 7604
rect -9666 7228 -9632 7604
rect -9570 7228 -9536 7604
rect -9474 7228 -9440 7604
rect -9378 7228 -9344 7604
rect -9282 7228 -9248 7604
rect -9186 7228 -9152 7604
rect -9090 7228 -9056 7604
rect -10050 6610 -10016 6986
rect -9954 6610 -9920 6986
rect -9858 6610 -9824 6986
rect -9762 6610 -9728 6986
rect -9666 6610 -9632 6986
rect -9570 6610 -9536 6986
rect -9474 6610 -9440 6986
rect -9378 6610 -9344 6986
rect -9282 6610 -9248 6986
rect -9186 6610 -9152 6986
rect -9090 6610 -9056 6986
rect -8658 8196 -8482 8230
rect -8658 6538 -8482 6572
rect -10050 5766 -10016 6142
rect -9954 5766 -9920 6142
rect -9858 5766 -9824 6142
rect -9762 5766 -9728 6142
rect -9666 5766 -9632 6142
rect -9570 5766 -9536 6142
rect -9474 5766 -9440 6142
rect -9378 5766 -9344 6142
rect -9282 5766 -9248 6142
rect -9186 5766 -9152 6142
rect -9090 5766 -9056 6142
rect -10050 5148 -10016 5524
rect -9954 5148 -9920 5524
rect -9858 5148 -9824 5524
rect -9762 5148 -9728 5524
rect -9666 5148 -9632 5524
rect -9570 5148 -9536 5524
rect -9474 5148 -9440 5524
rect -9378 5148 -9344 5524
rect -9282 5148 -9248 5524
rect -9186 5148 -9152 5524
rect -9090 5148 -9056 5524
rect -10050 4530 -10016 4906
rect -9954 4530 -9920 4906
rect -9858 4530 -9824 4906
rect -9762 4530 -9728 4906
rect -9666 4530 -9632 4906
rect -9570 4530 -9536 4906
rect -9474 4530 -9440 4906
rect -9378 4530 -9344 4906
rect -9282 4530 -9248 4906
rect -9186 4530 -9152 4906
rect -9090 4530 -9056 4906
rect 1690 8342 1724 8718
rect 1786 8342 1820 8718
rect 1882 8342 1916 8718
rect 1978 8342 2012 8718
rect 2074 8342 2108 8718
rect 2170 8342 2204 8718
rect 2266 8342 2300 8718
rect 2362 8342 2396 8718
rect 2458 8342 2492 8718
rect 2554 8342 2588 8718
rect 2650 8342 2684 8718
rect 2746 8342 2780 8718
rect 2842 8342 2876 8718
rect 2938 8342 2972 8718
rect 3034 8342 3068 8718
rect 3130 8342 3164 8718
rect 3226 8342 3260 8718
rect 3322 8342 3356 8718
rect 3418 8342 3452 8718
rect 3514 8342 3548 8718
rect 3610 8342 3644 8718
rect 1690 7522 1724 7898
rect 1786 7522 1820 7898
rect 1882 7522 1916 7898
rect 1978 7522 2012 7898
rect 2074 7522 2108 7898
rect 2170 7522 2204 7898
rect 2266 7522 2300 7898
rect 2362 7522 2396 7898
rect 2458 7522 2492 7898
rect 2554 7522 2588 7898
rect 2650 7522 2684 7898
rect 2746 7522 2780 7898
rect 2842 7522 2876 7898
rect 2938 7522 2972 7898
rect 3034 7522 3068 7898
rect 3130 7522 3164 7898
rect 3226 7522 3260 7898
rect 3322 7522 3356 7898
rect 3418 7522 3452 7898
rect 3514 7522 3548 7898
rect 3610 7522 3644 7898
rect 1690 6702 1724 7078
rect 1786 6702 1820 7078
rect 1882 6702 1916 7078
rect 1978 6702 2012 7078
rect 2074 6702 2108 7078
rect 2170 6702 2204 7078
rect 2266 6702 2300 7078
rect 2362 6702 2396 7078
rect 2458 6702 2492 7078
rect 2554 6702 2588 7078
rect 2650 6702 2684 7078
rect 2746 6702 2780 7078
rect 2842 6702 2876 7078
rect 2938 6702 2972 7078
rect 3034 6702 3068 7078
rect 3130 6702 3164 7078
rect 3226 6702 3260 7078
rect 3322 6702 3356 7078
rect 3418 6702 3452 7078
rect 3514 6702 3548 7078
rect 3610 6702 3644 7078
rect 5126 8308 5160 8684
rect 5222 8308 5256 8684
rect 5318 8308 5352 8684
rect 5414 8308 5448 8684
rect 5510 8308 5544 8684
rect 5606 8308 5640 8684
rect 5702 8308 5736 8684
rect 5798 8308 5832 8684
rect 5894 8308 5928 8684
rect 5990 8308 6024 8684
rect 6086 8308 6120 8684
rect 6182 8308 6216 8684
rect 6278 8308 6312 8684
rect 6374 8308 6408 8684
rect 6470 8308 6504 8684
rect 6566 8308 6600 8684
rect 6662 8308 6696 8684
rect 6758 8308 6792 8684
rect 6854 8308 6888 8684
rect 6950 8308 6984 8684
rect 7046 8308 7080 8684
rect 5126 7690 5160 8066
rect 5222 7690 5256 8066
rect 5318 7690 5352 8066
rect 5414 7690 5448 8066
rect 5510 7690 5544 8066
rect 5606 7690 5640 8066
rect 5702 7690 5736 8066
rect 5798 7690 5832 8066
rect 5894 7690 5928 8066
rect 5990 7690 6024 8066
rect 6086 7690 6120 8066
rect 6182 7690 6216 8066
rect 6278 7690 6312 8066
rect 6374 7690 6408 8066
rect 6470 7690 6504 8066
rect 6566 7690 6600 8066
rect 6662 7690 6696 8066
rect 6758 7690 6792 8066
rect 6854 7690 6888 8066
rect 6950 7690 6984 8066
rect 7046 7690 7080 8066
rect -10050 3620 -10016 3996
rect -9792 3620 -9758 3996
rect -9534 3620 -9500 3996
rect -9276 3620 -9242 3996
rect -9018 3620 -8984 3996
rect -8760 3620 -8726 3996
rect -10050 3002 -10016 3378
rect -9792 3002 -9758 3378
rect -9534 3002 -9500 3378
rect -9276 3002 -9242 3378
rect -9018 3002 -8984 3378
rect -8760 3002 -8726 3378
rect -10050 2384 -10016 2760
rect -9792 2384 -9758 2760
rect -9534 2384 -9500 2760
rect -9276 2384 -9242 2760
rect -9018 2384 -8984 2760
rect -8760 2384 -8726 2760
rect -10050 1766 -10016 2142
rect -9792 1766 -9758 2142
rect -9534 1766 -9500 2142
rect -9276 1766 -9242 2142
rect -9018 1766 -8984 2142
rect -8760 1766 -8726 2142
rect -10050 1148 -10016 1524
rect -9792 1148 -9758 1524
rect -9534 1148 -9500 1524
rect -9276 1148 -9242 1524
rect -9018 1148 -8984 1524
rect -8760 1148 -8726 1524
rect -10050 530 -10016 906
rect -9792 530 -9758 906
rect -9534 530 -9500 906
rect -9276 530 -9242 906
rect -9018 530 -8984 906
rect -8760 530 -8726 906
rect 226 5486 260 5862
rect 322 5486 356 5862
rect 418 5486 452 5862
rect 514 5486 548 5862
rect 610 5486 644 5862
rect 706 5486 740 5862
rect 802 5486 836 5862
rect 898 5486 932 5862
rect 994 5486 1028 5862
rect 1090 5486 1124 5862
rect 1186 5486 1220 5862
rect 226 4868 260 5244
rect 322 4868 356 5244
rect 418 4868 452 5244
rect 514 4868 548 5244
rect 610 4868 644 5244
rect 706 4868 740 5244
rect 802 4868 836 5244
rect 898 4868 932 5244
rect 994 4868 1028 5244
rect 1090 4868 1124 5244
rect 1186 4868 1220 5244
rect 226 4250 260 4626
rect 322 4250 356 4626
rect 418 4250 452 4626
rect 514 4250 548 4626
rect 610 4250 644 4626
rect 706 4250 740 4626
rect 802 4250 836 4626
rect 898 4250 932 4626
rect 994 4250 1028 4626
rect 1090 4250 1124 4626
rect 1186 4250 1220 4626
rect 2026 5486 2060 5862
rect 2122 5486 2156 5862
rect 2218 5486 2252 5862
rect 2314 5486 2348 5862
rect 2410 5486 2444 5862
rect 2506 5486 2540 5862
rect 2602 5486 2636 5862
rect 2698 5486 2732 5862
rect 2794 5486 2828 5862
rect 2890 5486 2924 5862
rect 2986 5486 3020 5862
rect 2026 4868 2060 5244
rect 2122 4868 2156 5244
rect 2218 4868 2252 5244
rect 2314 4868 2348 5244
rect 2410 4868 2444 5244
rect 2506 4868 2540 5244
rect 2602 4868 2636 5244
rect 2698 4868 2732 5244
rect 2794 4868 2828 5244
rect 2890 4868 2924 5244
rect 2986 4868 3020 5244
rect 2026 4250 2060 4626
rect 2122 4250 2156 4626
rect 2218 4250 2252 4626
rect 2314 4250 2348 4626
rect 2410 4250 2444 4626
rect 2506 4250 2540 4626
rect 2602 4250 2636 4626
rect 2698 4250 2732 4626
rect 2794 4250 2828 4626
rect 2890 4250 2924 4626
rect 2986 4250 3020 4626
rect 3826 5486 3860 5862
rect 3922 5486 3956 5862
rect 4018 5486 4052 5862
rect 4114 5486 4148 5862
rect 4210 5486 4244 5862
rect 4306 5486 4340 5862
rect 4402 5486 4436 5862
rect 4498 5486 4532 5862
rect 4594 5486 4628 5862
rect 4690 5486 4724 5862
rect 4786 5486 4820 5862
rect 3826 4868 3860 5244
rect 3922 4868 3956 5244
rect 4018 4868 4052 5244
rect 4114 4868 4148 5244
rect 4210 4868 4244 5244
rect 4306 4868 4340 5244
rect 4402 4868 4436 5244
rect 4498 4868 4532 5244
rect 4594 4868 4628 5244
rect 4690 4868 4724 5244
rect 4786 4868 4820 5244
rect 3826 4250 3860 4626
rect 3922 4250 3956 4626
rect 4018 4250 4052 4626
rect 4114 4250 4148 4626
rect 4210 4250 4244 4626
rect 4306 4250 4340 4626
rect 4402 4250 4436 4626
rect 4498 4250 4532 4626
rect 4594 4250 4628 4626
rect 4690 4250 4724 4626
rect 4786 4250 4820 4626
rect 5626 5486 5660 5862
rect 5722 5486 5756 5862
rect 5818 5486 5852 5862
rect 5914 5486 5948 5862
rect 6010 5486 6044 5862
rect 6106 5486 6140 5862
rect 6202 5486 6236 5862
rect 6298 5486 6332 5862
rect 6394 5486 6428 5862
rect 6490 5486 6524 5862
rect 6586 5486 6620 5862
rect 5626 4868 5660 5244
rect 5722 4868 5756 5244
rect 5818 4868 5852 5244
rect 5914 4868 5948 5244
rect 6010 4868 6044 5244
rect 6106 4868 6140 5244
rect 6202 4868 6236 5244
rect 6298 4868 6332 5244
rect 6394 4868 6428 5244
rect 6490 4868 6524 5244
rect 6586 4868 6620 5244
rect 5626 4250 5660 4626
rect 5722 4250 5756 4626
rect 5818 4250 5852 4626
rect 5914 4250 5948 4626
rect 6010 4250 6044 4626
rect 6106 4250 6140 4626
rect 6202 4250 6236 4626
rect 6298 4250 6332 4626
rect 6394 4250 6428 4626
rect 6490 4250 6524 4626
rect 6586 4250 6620 4626
rect 7626 9874 7660 10250
rect 7722 9874 7756 10250
rect 7818 9874 7852 10250
rect 7914 9874 7948 10250
rect 8010 9874 8044 10250
rect 8106 9874 8140 10250
rect 8202 9874 8236 10250
rect 8298 9874 8332 10250
rect 8394 9874 8428 10250
rect 8490 9874 8524 10250
rect 8586 9874 8620 10250
rect 8682 9874 8716 10250
rect 8778 9874 8812 10250
rect 8874 9874 8908 10250
rect 8970 9874 9004 10250
rect 9066 9874 9100 10250
rect 9162 9874 9196 10250
rect 9258 9874 9292 10250
rect 9354 9874 9388 10250
rect 9450 9874 9484 10250
rect 9546 9874 9580 10250
rect 7626 9256 7660 9632
rect 7722 9256 7756 9632
rect 7818 9256 7852 9632
rect 7914 9256 7948 9632
rect 8010 9256 8044 9632
rect 8106 9256 8140 9632
rect 8202 9256 8236 9632
rect 8298 9256 8332 9632
rect 8394 9256 8428 9632
rect 8490 9256 8524 9632
rect 8586 9256 8620 9632
rect 8682 9256 8716 9632
rect 8778 9256 8812 9632
rect 8874 9256 8908 9632
rect 8970 9256 9004 9632
rect 9066 9256 9100 9632
rect 9162 9256 9196 9632
rect 9258 9256 9292 9632
rect 9354 9256 9388 9632
rect 9450 9256 9484 9632
rect 9546 9256 9580 9632
rect 7626 8638 7660 9014
rect 7722 8638 7756 9014
rect 7818 8638 7852 9014
rect 7914 8638 7948 9014
rect 8010 8638 8044 9014
rect 8106 8638 8140 9014
rect 8202 8638 8236 9014
rect 8298 8638 8332 9014
rect 8394 8638 8428 9014
rect 8490 8638 8524 9014
rect 8586 8638 8620 9014
rect 8682 8638 8716 9014
rect 8778 8638 8812 9014
rect 8874 8638 8908 9014
rect 8970 8638 9004 9014
rect 9066 8638 9100 9014
rect 9162 8638 9196 9014
rect 9258 8638 9292 9014
rect 9354 8638 9388 9014
rect 9450 8638 9484 9014
rect 9546 8638 9580 9014
rect 7626 8020 7660 8396
rect 7722 8020 7756 8396
rect 7818 8020 7852 8396
rect 7914 8020 7948 8396
rect 8010 8020 8044 8396
rect 8106 8020 8140 8396
rect 8202 8020 8236 8396
rect 8298 8020 8332 8396
rect 8394 8020 8428 8396
rect 8490 8020 8524 8396
rect 8586 8020 8620 8396
rect 8682 8020 8716 8396
rect 8778 8020 8812 8396
rect 8874 8020 8908 8396
rect 8970 8020 9004 8396
rect 9066 8020 9100 8396
rect 9162 8020 9196 8396
rect 9258 8020 9292 8396
rect 9354 8020 9388 8396
rect 9450 8020 9484 8396
rect 9546 8020 9580 8396
rect 7626 7402 7660 7778
rect 7722 7402 7756 7778
rect 7818 7402 7852 7778
rect 7914 7402 7948 7778
rect 8010 7402 8044 7778
rect 8106 7402 8140 7778
rect 8202 7402 8236 7778
rect 8298 7402 8332 7778
rect 8394 7402 8428 7778
rect 8490 7402 8524 7778
rect 8586 7402 8620 7778
rect 8682 7402 8716 7778
rect 8778 7402 8812 7778
rect 8874 7402 8908 7778
rect 8970 7402 9004 7778
rect 9066 7402 9100 7778
rect 9162 7402 9196 7778
rect 9258 7402 9292 7778
rect 9354 7402 9388 7778
rect 9450 7402 9484 7778
rect 9546 7402 9580 7778
rect 7626 6784 7660 7160
rect 7722 6784 7756 7160
rect 7818 6784 7852 7160
rect 7914 6784 7948 7160
rect 8010 6784 8044 7160
rect 8106 6784 8140 7160
rect 8202 6784 8236 7160
rect 8298 6784 8332 7160
rect 8394 6784 8428 7160
rect 8490 6784 8524 7160
rect 8586 6784 8620 7160
rect 8682 6784 8716 7160
rect 8778 6784 8812 7160
rect 8874 6784 8908 7160
rect 8970 6784 9004 7160
rect 9066 6784 9100 7160
rect 9162 6784 9196 7160
rect 9258 6784 9292 7160
rect 9354 6784 9388 7160
rect 9450 6784 9484 7160
rect 9546 6784 9580 7160
rect 7626 6166 7660 6542
rect 7722 6166 7756 6542
rect 7818 6166 7852 6542
rect 7914 6166 7948 6542
rect 8010 6166 8044 6542
rect 8106 6166 8140 6542
rect 8202 6166 8236 6542
rect 8298 6166 8332 6542
rect 8394 6166 8428 6542
rect 8490 6166 8524 6542
rect 8586 6166 8620 6542
rect 8682 6166 8716 6542
rect 8778 6166 8812 6542
rect 8874 6166 8908 6542
rect 8970 6166 9004 6542
rect 9066 6166 9100 6542
rect 9162 6166 9196 6542
rect 9258 6166 9292 6542
rect 9354 6166 9388 6542
rect 9450 6166 9484 6542
rect 9546 6166 9580 6542
rect 7626 5548 7660 5924
rect 7722 5548 7756 5924
rect 7818 5548 7852 5924
rect 7914 5548 7948 5924
rect 8010 5548 8044 5924
rect 8106 5548 8140 5924
rect 8202 5548 8236 5924
rect 8298 5548 8332 5924
rect 8394 5548 8428 5924
rect 8490 5548 8524 5924
rect 8586 5548 8620 5924
rect 8682 5548 8716 5924
rect 8778 5548 8812 5924
rect 8874 5548 8908 5924
rect 8970 5548 9004 5924
rect 9066 5548 9100 5924
rect 9162 5548 9196 5924
rect 9258 5548 9292 5924
rect 9354 5548 9388 5924
rect 9450 5548 9484 5924
rect 9546 5548 9580 5924
rect 7626 4930 7660 5306
rect 7722 4930 7756 5306
rect 7818 4930 7852 5306
rect 7914 4930 7948 5306
rect 8010 4930 8044 5306
rect 8106 4930 8140 5306
rect 8202 4930 8236 5306
rect 8298 4930 8332 5306
rect 8394 4930 8428 5306
rect 8490 4930 8524 5306
rect 8586 4930 8620 5306
rect 8682 4930 8716 5306
rect 8778 4930 8812 5306
rect 8874 4930 8908 5306
rect 8970 4930 9004 5306
rect 9066 4930 9100 5306
rect 9162 4930 9196 5306
rect 9258 4930 9292 5306
rect 9354 4930 9388 5306
rect 9450 4930 9484 5306
rect 9546 4930 9580 5306
rect 16090 8342 16124 8718
rect 16186 8342 16220 8718
rect 16282 8342 16316 8718
rect 16378 8342 16412 8718
rect 16474 8342 16508 8718
rect 16570 8342 16604 8718
rect 16666 8342 16700 8718
rect 16762 8342 16796 8718
rect 16858 8342 16892 8718
rect 16954 8342 16988 8718
rect 17050 8342 17084 8718
rect 17146 8342 17180 8718
rect 17242 8342 17276 8718
rect 17338 8342 17372 8718
rect 17434 8342 17468 8718
rect 17530 8342 17564 8718
rect 17626 8342 17660 8718
rect 17722 8342 17756 8718
rect 17818 8342 17852 8718
rect 17914 8342 17948 8718
rect 18010 8342 18044 8718
rect 16090 7522 16124 7898
rect 16186 7522 16220 7898
rect 16282 7522 16316 7898
rect 16378 7522 16412 7898
rect 16474 7522 16508 7898
rect 16570 7522 16604 7898
rect 16666 7522 16700 7898
rect 16762 7522 16796 7898
rect 16858 7522 16892 7898
rect 16954 7522 16988 7898
rect 17050 7522 17084 7898
rect 17146 7522 17180 7898
rect 17242 7522 17276 7898
rect 17338 7522 17372 7898
rect 17434 7522 17468 7898
rect 17530 7522 17564 7898
rect 17626 7522 17660 7898
rect 17722 7522 17756 7898
rect 17818 7522 17852 7898
rect 17914 7522 17948 7898
rect 18010 7522 18044 7898
rect 16090 6702 16124 7078
rect 16186 6702 16220 7078
rect 16282 6702 16316 7078
rect 16378 6702 16412 7078
rect 16474 6702 16508 7078
rect 16570 6702 16604 7078
rect 16666 6702 16700 7078
rect 16762 6702 16796 7078
rect 16858 6702 16892 7078
rect 16954 6702 16988 7078
rect 17050 6702 17084 7078
rect 17146 6702 17180 7078
rect 17242 6702 17276 7078
rect 17338 6702 17372 7078
rect 17434 6702 17468 7078
rect 17530 6702 17564 7078
rect 17626 6702 17660 7078
rect 17722 6702 17756 7078
rect 17818 6702 17852 7078
rect 17914 6702 17948 7078
rect 18010 6702 18044 7078
rect 19526 8308 19560 8684
rect 19622 8308 19656 8684
rect 19718 8308 19752 8684
rect 19814 8308 19848 8684
rect 19910 8308 19944 8684
rect 20006 8308 20040 8684
rect 20102 8308 20136 8684
rect 20198 8308 20232 8684
rect 20294 8308 20328 8684
rect 20390 8308 20424 8684
rect 20486 8308 20520 8684
rect 20582 8308 20616 8684
rect 20678 8308 20712 8684
rect 20774 8308 20808 8684
rect 20870 8308 20904 8684
rect 20966 8308 21000 8684
rect 21062 8308 21096 8684
rect 21158 8308 21192 8684
rect 21254 8308 21288 8684
rect 21350 8308 21384 8684
rect 21446 8308 21480 8684
rect 19526 7690 19560 8066
rect 19622 7690 19656 8066
rect 19718 7690 19752 8066
rect 19814 7690 19848 8066
rect 19910 7690 19944 8066
rect 20006 7690 20040 8066
rect 20102 7690 20136 8066
rect 20198 7690 20232 8066
rect 20294 7690 20328 8066
rect 20390 7690 20424 8066
rect 20486 7690 20520 8066
rect 20582 7690 20616 8066
rect 20678 7690 20712 8066
rect 20774 7690 20808 8066
rect 20870 7690 20904 8066
rect 20966 7690 21000 8066
rect 21062 7690 21096 8066
rect 21158 7690 21192 8066
rect 21254 7690 21288 8066
rect 21350 7690 21384 8066
rect 21446 7690 21480 8066
rect 14626 5486 14660 5862
rect 14722 5486 14756 5862
rect 14818 5486 14852 5862
rect 14914 5486 14948 5862
rect 15010 5486 15044 5862
rect 15106 5486 15140 5862
rect 15202 5486 15236 5862
rect 15298 5486 15332 5862
rect 15394 5486 15428 5862
rect 15490 5486 15524 5862
rect 15586 5486 15620 5862
rect 14626 4868 14660 5244
rect 14722 4868 14756 5244
rect 14818 4868 14852 5244
rect 14914 4868 14948 5244
rect 15010 4868 15044 5244
rect 15106 4868 15140 5244
rect 15202 4868 15236 5244
rect 15298 4868 15332 5244
rect 15394 4868 15428 5244
rect 15490 4868 15524 5244
rect 15586 4868 15620 5244
rect 14626 4250 14660 4626
rect 14722 4250 14756 4626
rect 14818 4250 14852 4626
rect 14914 4250 14948 4626
rect 15010 4250 15044 4626
rect 15106 4250 15140 4626
rect 15202 4250 15236 4626
rect 15298 4250 15332 4626
rect 15394 4250 15428 4626
rect 15490 4250 15524 4626
rect 15586 4250 15620 4626
rect 16426 5486 16460 5862
rect 16522 5486 16556 5862
rect 16618 5486 16652 5862
rect 16714 5486 16748 5862
rect 16810 5486 16844 5862
rect 16906 5486 16940 5862
rect 17002 5486 17036 5862
rect 17098 5486 17132 5862
rect 17194 5486 17228 5862
rect 17290 5486 17324 5862
rect 17386 5486 17420 5862
rect 16426 4868 16460 5244
rect 16522 4868 16556 5244
rect 16618 4868 16652 5244
rect 16714 4868 16748 5244
rect 16810 4868 16844 5244
rect 16906 4868 16940 5244
rect 17002 4868 17036 5244
rect 17098 4868 17132 5244
rect 17194 4868 17228 5244
rect 17290 4868 17324 5244
rect 17386 4868 17420 5244
rect 16426 4250 16460 4626
rect 16522 4250 16556 4626
rect 16618 4250 16652 4626
rect 16714 4250 16748 4626
rect 16810 4250 16844 4626
rect 16906 4250 16940 4626
rect 17002 4250 17036 4626
rect 17098 4250 17132 4626
rect 17194 4250 17228 4626
rect 17290 4250 17324 4626
rect 17386 4250 17420 4626
rect 18226 5486 18260 5862
rect 18322 5486 18356 5862
rect 18418 5486 18452 5862
rect 18514 5486 18548 5862
rect 18610 5486 18644 5862
rect 18706 5486 18740 5862
rect 18802 5486 18836 5862
rect 18898 5486 18932 5862
rect 18994 5486 19028 5862
rect 19090 5486 19124 5862
rect 19186 5486 19220 5862
rect 18226 4868 18260 5244
rect 18322 4868 18356 5244
rect 18418 4868 18452 5244
rect 18514 4868 18548 5244
rect 18610 4868 18644 5244
rect 18706 4868 18740 5244
rect 18802 4868 18836 5244
rect 18898 4868 18932 5244
rect 18994 4868 19028 5244
rect 19090 4868 19124 5244
rect 19186 4868 19220 5244
rect 18226 4250 18260 4626
rect 18322 4250 18356 4626
rect 18418 4250 18452 4626
rect 18514 4250 18548 4626
rect 18610 4250 18644 4626
rect 18706 4250 18740 4626
rect 18802 4250 18836 4626
rect 18898 4250 18932 4626
rect 18994 4250 19028 4626
rect 19090 4250 19124 4626
rect 19186 4250 19220 4626
rect 20026 5486 20060 5862
rect 20122 5486 20156 5862
rect 20218 5486 20252 5862
rect 20314 5486 20348 5862
rect 20410 5486 20444 5862
rect 20506 5486 20540 5862
rect 20602 5486 20636 5862
rect 20698 5486 20732 5862
rect 20794 5486 20828 5862
rect 20890 5486 20924 5862
rect 20986 5486 21020 5862
rect 20026 4868 20060 5244
rect 20122 4868 20156 5244
rect 20218 4868 20252 5244
rect 20314 4868 20348 5244
rect 20410 4868 20444 5244
rect 20506 4868 20540 5244
rect 20602 4868 20636 5244
rect 20698 4868 20732 5244
rect 20794 4868 20828 5244
rect 20890 4868 20924 5244
rect 20986 4868 21020 5244
rect 20026 4250 20060 4626
rect 20122 4250 20156 4626
rect 20218 4250 20252 4626
rect 20314 4250 20348 4626
rect 20410 4250 20444 4626
rect 20506 4250 20540 4626
rect 20602 4250 20636 4626
rect 20698 4250 20732 4626
rect 20794 4250 20828 4626
rect 20890 4250 20924 4626
rect 20986 4250 21020 4626
rect 22026 9874 22060 10250
rect 22122 9874 22156 10250
rect 22218 9874 22252 10250
rect 22314 9874 22348 10250
rect 22410 9874 22444 10250
rect 22506 9874 22540 10250
rect 22602 9874 22636 10250
rect 22698 9874 22732 10250
rect 22794 9874 22828 10250
rect 22890 9874 22924 10250
rect 22986 9874 23020 10250
rect 23082 9874 23116 10250
rect 23178 9874 23212 10250
rect 23274 9874 23308 10250
rect 23370 9874 23404 10250
rect 23466 9874 23500 10250
rect 23562 9874 23596 10250
rect 23658 9874 23692 10250
rect 23754 9874 23788 10250
rect 23850 9874 23884 10250
rect 23946 9874 23980 10250
rect 22026 9256 22060 9632
rect 22122 9256 22156 9632
rect 22218 9256 22252 9632
rect 22314 9256 22348 9632
rect 22410 9256 22444 9632
rect 22506 9256 22540 9632
rect 22602 9256 22636 9632
rect 22698 9256 22732 9632
rect 22794 9256 22828 9632
rect 22890 9256 22924 9632
rect 22986 9256 23020 9632
rect 23082 9256 23116 9632
rect 23178 9256 23212 9632
rect 23274 9256 23308 9632
rect 23370 9256 23404 9632
rect 23466 9256 23500 9632
rect 23562 9256 23596 9632
rect 23658 9256 23692 9632
rect 23754 9256 23788 9632
rect 23850 9256 23884 9632
rect 23946 9256 23980 9632
rect 22026 8638 22060 9014
rect 22122 8638 22156 9014
rect 22218 8638 22252 9014
rect 22314 8638 22348 9014
rect 22410 8638 22444 9014
rect 22506 8638 22540 9014
rect 22602 8638 22636 9014
rect 22698 8638 22732 9014
rect 22794 8638 22828 9014
rect 22890 8638 22924 9014
rect 22986 8638 23020 9014
rect 23082 8638 23116 9014
rect 23178 8638 23212 9014
rect 23274 8638 23308 9014
rect 23370 8638 23404 9014
rect 23466 8638 23500 9014
rect 23562 8638 23596 9014
rect 23658 8638 23692 9014
rect 23754 8638 23788 9014
rect 23850 8638 23884 9014
rect 23946 8638 23980 9014
rect 22026 8020 22060 8396
rect 22122 8020 22156 8396
rect 22218 8020 22252 8396
rect 22314 8020 22348 8396
rect 22410 8020 22444 8396
rect 22506 8020 22540 8396
rect 22602 8020 22636 8396
rect 22698 8020 22732 8396
rect 22794 8020 22828 8396
rect 22890 8020 22924 8396
rect 22986 8020 23020 8396
rect 23082 8020 23116 8396
rect 23178 8020 23212 8396
rect 23274 8020 23308 8396
rect 23370 8020 23404 8396
rect 23466 8020 23500 8396
rect 23562 8020 23596 8396
rect 23658 8020 23692 8396
rect 23754 8020 23788 8396
rect 23850 8020 23884 8396
rect 23946 8020 23980 8396
rect 22026 7402 22060 7778
rect 22122 7402 22156 7778
rect 22218 7402 22252 7778
rect 22314 7402 22348 7778
rect 22410 7402 22444 7778
rect 22506 7402 22540 7778
rect 22602 7402 22636 7778
rect 22698 7402 22732 7778
rect 22794 7402 22828 7778
rect 22890 7402 22924 7778
rect 22986 7402 23020 7778
rect 23082 7402 23116 7778
rect 23178 7402 23212 7778
rect 23274 7402 23308 7778
rect 23370 7402 23404 7778
rect 23466 7402 23500 7778
rect 23562 7402 23596 7778
rect 23658 7402 23692 7778
rect 23754 7402 23788 7778
rect 23850 7402 23884 7778
rect 23946 7402 23980 7778
rect 22026 6784 22060 7160
rect 22122 6784 22156 7160
rect 22218 6784 22252 7160
rect 22314 6784 22348 7160
rect 22410 6784 22444 7160
rect 22506 6784 22540 7160
rect 22602 6784 22636 7160
rect 22698 6784 22732 7160
rect 22794 6784 22828 7160
rect 22890 6784 22924 7160
rect 22986 6784 23020 7160
rect 23082 6784 23116 7160
rect 23178 6784 23212 7160
rect 23274 6784 23308 7160
rect 23370 6784 23404 7160
rect 23466 6784 23500 7160
rect 23562 6784 23596 7160
rect 23658 6784 23692 7160
rect 23754 6784 23788 7160
rect 23850 6784 23884 7160
rect 23946 6784 23980 7160
rect 22026 6166 22060 6542
rect 22122 6166 22156 6542
rect 22218 6166 22252 6542
rect 22314 6166 22348 6542
rect 22410 6166 22444 6542
rect 22506 6166 22540 6542
rect 22602 6166 22636 6542
rect 22698 6166 22732 6542
rect 22794 6166 22828 6542
rect 22890 6166 22924 6542
rect 22986 6166 23020 6542
rect 23082 6166 23116 6542
rect 23178 6166 23212 6542
rect 23274 6166 23308 6542
rect 23370 6166 23404 6542
rect 23466 6166 23500 6542
rect 23562 6166 23596 6542
rect 23658 6166 23692 6542
rect 23754 6166 23788 6542
rect 23850 6166 23884 6542
rect 23946 6166 23980 6542
rect 22026 5548 22060 5924
rect 22122 5548 22156 5924
rect 22218 5548 22252 5924
rect 22314 5548 22348 5924
rect 22410 5548 22444 5924
rect 22506 5548 22540 5924
rect 22602 5548 22636 5924
rect 22698 5548 22732 5924
rect 22794 5548 22828 5924
rect 22890 5548 22924 5924
rect 22986 5548 23020 5924
rect 23082 5548 23116 5924
rect 23178 5548 23212 5924
rect 23274 5548 23308 5924
rect 23370 5548 23404 5924
rect 23466 5548 23500 5924
rect 23562 5548 23596 5924
rect 23658 5548 23692 5924
rect 23754 5548 23788 5924
rect 23850 5548 23884 5924
rect 23946 5548 23980 5924
rect 22026 4930 22060 5306
rect 22122 4930 22156 5306
rect 22218 4930 22252 5306
rect 22314 4930 22348 5306
rect 22410 4930 22444 5306
rect 22506 4930 22540 5306
rect 22602 4930 22636 5306
rect 22698 4930 22732 5306
rect 22794 4930 22828 5306
rect 22890 4930 22924 5306
rect 22986 4930 23020 5306
rect 23082 4930 23116 5306
rect 23178 4930 23212 5306
rect 23274 4930 23308 5306
rect 23370 4930 23404 5306
rect 23466 4930 23500 5306
rect 23562 4930 23596 5306
rect 23658 4930 23692 5306
rect 23754 4930 23788 5306
rect 23850 4930 23884 5306
rect 23946 4930 23980 5306
rect 226 3340 260 3716
rect 484 3340 518 3716
rect 742 3340 776 3716
rect 1000 3340 1034 3716
rect 1258 3340 1292 3716
rect 1516 3340 1550 3716
rect 226 2722 260 3098
rect 484 2722 518 3098
rect 742 2722 776 3098
rect 1000 2722 1034 3098
rect 1258 2722 1292 3098
rect 1516 2722 1550 3098
rect 226 2104 260 2480
rect 484 2104 518 2480
rect 742 2104 776 2480
rect 1000 2104 1034 2480
rect 1258 2104 1292 2480
rect 1516 2104 1550 2480
rect 226 1486 260 1862
rect 484 1486 518 1862
rect 742 1486 776 1862
rect 1000 1486 1034 1862
rect 1258 1486 1292 1862
rect 1516 1486 1550 1862
rect 226 868 260 1244
rect 484 868 518 1244
rect 742 868 776 1244
rect 1000 868 1034 1244
rect 1258 868 1292 1244
rect 1516 868 1550 1244
rect 226 250 260 626
rect 484 250 518 626
rect 742 250 776 626
rect 1000 250 1034 626
rect 1258 250 1292 626
rect 1516 250 1550 626
rect 2026 3340 2060 3716
rect 2284 3340 2318 3716
rect 2542 3340 2576 3716
rect 2800 3340 2834 3716
rect 3058 3340 3092 3716
rect 3316 3340 3350 3716
rect 2026 2722 2060 3098
rect 2284 2722 2318 3098
rect 2542 2722 2576 3098
rect 2800 2722 2834 3098
rect 3058 2722 3092 3098
rect 3316 2722 3350 3098
rect 2026 2104 2060 2480
rect 2284 2104 2318 2480
rect 2542 2104 2576 2480
rect 2800 2104 2834 2480
rect 3058 2104 3092 2480
rect 3316 2104 3350 2480
rect 2026 1486 2060 1862
rect 2284 1486 2318 1862
rect 2542 1486 2576 1862
rect 2800 1486 2834 1862
rect 3058 1486 3092 1862
rect 3316 1486 3350 1862
rect 2026 868 2060 1244
rect 2284 868 2318 1244
rect 2542 868 2576 1244
rect 2800 868 2834 1244
rect 3058 868 3092 1244
rect 3316 868 3350 1244
rect 2026 250 2060 626
rect 2284 250 2318 626
rect 2542 250 2576 626
rect 2800 250 2834 626
rect 3058 250 3092 626
rect 3316 250 3350 626
rect 3826 3340 3860 3716
rect 4084 3340 4118 3716
rect 4342 3340 4376 3716
rect 4600 3340 4634 3716
rect 4858 3340 4892 3716
rect 5116 3340 5150 3716
rect 3826 2722 3860 3098
rect 4084 2722 4118 3098
rect 4342 2722 4376 3098
rect 4600 2722 4634 3098
rect 4858 2722 4892 3098
rect 5116 2722 5150 3098
rect 3826 2104 3860 2480
rect 4084 2104 4118 2480
rect 4342 2104 4376 2480
rect 4600 2104 4634 2480
rect 4858 2104 4892 2480
rect 5116 2104 5150 2480
rect 3826 1486 3860 1862
rect 4084 1486 4118 1862
rect 4342 1486 4376 1862
rect 4600 1486 4634 1862
rect 4858 1486 4892 1862
rect 5116 1486 5150 1862
rect 3826 868 3860 1244
rect 4084 868 4118 1244
rect 4342 868 4376 1244
rect 4600 868 4634 1244
rect 4858 868 4892 1244
rect 5116 868 5150 1244
rect 3826 250 3860 626
rect 4084 250 4118 626
rect 4342 250 4376 626
rect 4600 250 4634 626
rect 4858 250 4892 626
rect 5116 250 5150 626
rect 5626 3340 5660 3716
rect 5884 3340 5918 3716
rect 6142 3340 6176 3716
rect 6400 3340 6434 3716
rect 6658 3340 6692 3716
rect 6916 3340 6950 3716
rect 5626 2722 5660 3098
rect 5884 2722 5918 3098
rect 6142 2722 6176 3098
rect 6400 2722 6434 3098
rect 6658 2722 6692 3098
rect 6916 2722 6950 3098
rect 5626 2104 5660 2480
rect 5884 2104 5918 2480
rect 6142 2104 6176 2480
rect 6400 2104 6434 2480
rect 6658 2104 6692 2480
rect 6916 2104 6950 2480
rect 5626 1486 5660 1862
rect 5884 1486 5918 1862
rect 6142 1486 6176 1862
rect 6400 1486 6434 1862
rect 6658 1486 6692 1862
rect 6916 1486 6950 1862
rect 5626 868 5660 1244
rect 5884 868 5918 1244
rect 6142 868 6176 1244
rect 6400 868 6434 1244
rect 6658 868 6692 1244
rect 6916 868 6950 1244
rect 5626 250 5660 626
rect 5884 250 5918 626
rect 6142 250 6176 626
rect 6400 250 6434 626
rect 6658 250 6692 626
rect 6916 250 6950 626
rect 14626 3340 14660 3716
rect 14884 3340 14918 3716
rect 15142 3340 15176 3716
rect 15400 3340 15434 3716
rect 15658 3340 15692 3716
rect 15916 3340 15950 3716
rect 14626 2722 14660 3098
rect 14884 2722 14918 3098
rect 15142 2722 15176 3098
rect 15400 2722 15434 3098
rect 15658 2722 15692 3098
rect 15916 2722 15950 3098
rect 14626 2104 14660 2480
rect 14884 2104 14918 2480
rect 15142 2104 15176 2480
rect 15400 2104 15434 2480
rect 15658 2104 15692 2480
rect 15916 2104 15950 2480
rect 14626 1486 14660 1862
rect 14884 1486 14918 1862
rect 15142 1486 15176 1862
rect 15400 1486 15434 1862
rect 15658 1486 15692 1862
rect 15916 1486 15950 1862
rect 14626 868 14660 1244
rect 14884 868 14918 1244
rect 15142 868 15176 1244
rect 15400 868 15434 1244
rect 15658 868 15692 1244
rect 15916 868 15950 1244
rect 14626 250 14660 626
rect 14884 250 14918 626
rect 15142 250 15176 626
rect 15400 250 15434 626
rect 15658 250 15692 626
rect 15916 250 15950 626
rect 16426 3340 16460 3716
rect 16684 3340 16718 3716
rect 16942 3340 16976 3716
rect 17200 3340 17234 3716
rect 17458 3340 17492 3716
rect 17716 3340 17750 3716
rect 16426 2722 16460 3098
rect 16684 2722 16718 3098
rect 16942 2722 16976 3098
rect 17200 2722 17234 3098
rect 17458 2722 17492 3098
rect 17716 2722 17750 3098
rect 16426 2104 16460 2480
rect 16684 2104 16718 2480
rect 16942 2104 16976 2480
rect 17200 2104 17234 2480
rect 17458 2104 17492 2480
rect 17716 2104 17750 2480
rect 16426 1486 16460 1862
rect 16684 1486 16718 1862
rect 16942 1486 16976 1862
rect 17200 1486 17234 1862
rect 17458 1486 17492 1862
rect 17716 1486 17750 1862
rect 16426 868 16460 1244
rect 16684 868 16718 1244
rect 16942 868 16976 1244
rect 17200 868 17234 1244
rect 17458 868 17492 1244
rect 17716 868 17750 1244
rect 16426 250 16460 626
rect 16684 250 16718 626
rect 16942 250 16976 626
rect 17200 250 17234 626
rect 17458 250 17492 626
rect 17716 250 17750 626
rect 18226 3340 18260 3716
rect 18484 3340 18518 3716
rect 18742 3340 18776 3716
rect 19000 3340 19034 3716
rect 19258 3340 19292 3716
rect 19516 3340 19550 3716
rect 18226 2722 18260 3098
rect 18484 2722 18518 3098
rect 18742 2722 18776 3098
rect 19000 2722 19034 3098
rect 19258 2722 19292 3098
rect 19516 2722 19550 3098
rect 18226 2104 18260 2480
rect 18484 2104 18518 2480
rect 18742 2104 18776 2480
rect 19000 2104 19034 2480
rect 19258 2104 19292 2480
rect 19516 2104 19550 2480
rect 18226 1486 18260 1862
rect 18484 1486 18518 1862
rect 18742 1486 18776 1862
rect 19000 1486 19034 1862
rect 19258 1486 19292 1862
rect 19516 1486 19550 1862
rect 18226 868 18260 1244
rect 18484 868 18518 1244
rect 18742 868 18776 1244
rect 19000 868 19034 1244
rect 19258 868 19292 1244
rect 19516 868 19550 1244
rect 18226 250 18260 626
rect 18484 250 18518 626
rect 18742 250 18776 626
rect 19000 250 19034 626
rect 19258 250 19292 626
rect 19516 250 19550 626
rect 20026 3340 20060 3716
rect 20284 3340 20318 3716
rect 20542 3340 20576 3716
rect 20800 3340 20834 3716
rect 21058 3340 21092 3716
rect 21316 3340 21350 3716
rect 20026 2722 20060 3098
rect 20284 2722 20318 3098
rect 20542 2722 20576 3098
rect 20800 2722 20834 3098
rect 21058 2722 21092 3098
rect 21316 2722 21350 3098
rect 20026 2104 20060 2480
rect 20284 2104 20318 2480
rect 20542 2104 20576 2480
rect 20800 2104 20834 2480
rect 21058 2104 21092 2480
rect 21316 2104 21350 2480
rect 20026 1486 20060 1862
rect 20284 1486 20318 1862
rect 20542 1486 20576 1862
rect 20800 1486 20834 1862
rect 21058 1486 21092 1862
rect 21316 1486 21350 1862
rect 20026 868 20060 1244
rect 20284 868 20318 1244
rect 20542 868 20576 1244
rect 20800 868 20834 1244
rect 21058 868 21092 1244
rect 21316 868 21350 1244
rect 20026 250 20060 626
rect 20284 250 20318 626
rect 20542 250 20576 626
rect 20800 250 20834 626
rect 21058 250 21092 626
rect 21316 250 21350 626
<< pdiffc >>
rect 6490 26699 6524 27075
rect 6648 26699 6682 27075
rect 6806 26699 6840 27075
rect 6964 26699 6998 27075
rect 7122 26699 7156 27075
rect 7280 26699 7314 27075
rect 7438 26699 7472 27075
rect 7596 26699 7630 27075
rect 7754 26699 7788 27075
rect 7912 26699 7946 27075
rect 8070 26699 8104 27075
rect 6490 26063 6524 26439
rect 6648 26063 6682 26439
rect 6806 26063 6840 26439
rect 6964 26063 6998 26439
rect 7122 26063 7156 26439
rect 7280 26063 7314 26439
rect 7438 26063 7472 26439
rect 7596 26063 7630 26439
rect 7754 26063 7788 26439
rect 7912 26063 7946 26439
rect 8070 26063 8104 26439
rect 6490 25427 6524 25803
rect 6648 25427 6682 25803
rect 6806 25427 6840 25803
rect 6964 25427 6998 25803
rect 7122 25427 7156 25803
rect 7280 25427 7314 25803
rect 7438 25427 7472 25803
rect 7596 25427 7630 25803
rect 7754 25427 7788 25803
rect 7912 25427 7946 25803
rect 8070 25427 8104 25803
rect 8710 26699 8744 27075
rect 8868 26699 8902 27075
rect 9026 26699 9060 27075
rect 9184 26699 9218 27075
rect 9342 26699 9376 27075
rect 9500 26699 9534 27075
rect 9658 26699 9692 27075
rect 9816 26699 9850 27075
rect 9974 26699 10008 27075
rect 10132 26699 10166 27075
rect 10290 26699 10324 27075
rect 8710 26063 8744 26439
rect 8868 26063 8902 26439
rect 9026 26063 9060 26439
rect 9184 26063 9218 26439
rect 9342 26063 9376 26439
rect 9500 26063 9534 26439
rect 9658 26063 9692 26439
rect 9816 26063 9850 26439
rect 9974 26063 10008 26439
rect 10132 26063 10166 26439
rect 10290 26063 10324 26439
rect 8710 25427 8744 25803
rect 8868 25427 8902 25803
rect 9026 25427 9060 25803
rect 9184 25427 9218 25803
rect 9342 25427 9376 25803
rect 9500 25427 9534 25803
rect 9658 25427 9692 25803
rect 9816 25427 9850 25803
rect 9974 25427 10008 25803
rect 10132 25427 10166 25803
rect 10290 25427 10324 25803
rect 10890 26699 10924 27075
rect 11048 26699 11082 27075
rect 11206 26699 11240 27075
rect 11364 26699 11398 27075
rect 11522 26699 11556 27075
rect 11680 26699 11714 27075
rect 11838 26699 11872 27075
rect 11996 26699 12030 27075
rect 12154 26699 12188 27075
rect 12312 26699 12346 27075
rect 12470 26699 12504 27075
rect 10890 26063 10924 26439
rect 11048 26063 11082 26439
rect 11206 26063 11240 26439
rect 11364 26063 11398 26439
rect 11522 26063 11556 26439
rect 11680 26063 11714 26439
rect 11838 26063 11872 26439
rect 11996 26063 12030 26439
rect 12154 26063 12188 26439
rect 12312 26063 12346 26439
rect 12470 26063 12504 26439
rect 10890 25427 10924 25803
rect 11048 25427 11082 25803
rect 11206 25427 11240 25803
rect 11364 25427 11398 25803
rect 11522 25427 11556 25803
rect 11680 25427 11714 25803
rect 11838 25427 11872 25803
rect 11996 25427 12030 25803
rect 12154 25427 12188 25803
rect 12312 25427 12346 25803
rect 12470 25427 12504 25803
rect 13070 26699 13104 27075
rect 13228 26699 13262 27075
rect 13386 26699 13420 27075
rect 13544 26699 13578 27075
rect 13702 26699 13736 27075
rect 13860 26699 13894 27075
rect 14018 26699 14052 27075
rect 14176 26699 14210 27075
rect 14334 26699 14368 27075
rect 14492 26699 14526 27075
rect 14650 26699 14684 27075
rect 13070 26063 13104 26439
rect 13228 26063 13262 26439
rect 13386 26063 13420 26439
rect 13544 26063 13578 26439
rect 13702 26063 13736 26439
rect 13860 26063 13894 26439
rect 14018 26063 14052 26439
rect 14176 26063 14210 26439
rect 14334 26063 14368 26439
rect 14492 26063 14526 26439
rect 14650 26063 14684 26439
rect 13070 25427 13104 25803
rect 13228 25427 13262 25803
rect 13386 25427 13420 25803
rect 13544 25427 13578 25803
rect 13702 25427 13736 25803
rect 13860 25427 13894 25803
rect 14018 25427 14052 25803
rect 14176 25427 14210 25803
rect 14334 25427 14368 25803
rect 14492 25427 14526 25803
rect 14650 25427 14684 25803
rect 15270 26699 15304 27075
rect 15428 26699 15462 27075
rect 15586 26699 15620 27075
rect 15744 26699 15778 27075
rect 15902 26699 15936 27075
rect 16060 26699 16094 27075
rect 16218 26699 16252 27075
rect 16376 26699 16410 27075
rect 16534 26699 16568 27075
rect 16692 26699 16726 27075
rect 16850 26699 16884 27075
rect 15270 26063 15304 26439
rect 15428 26063 15462 26439
rect 15586 26063 15620 26439
rect 15744 26063 15778 26439
rect 15902 26063 15936 26439
rect 16060 26063 16094 26439
rect 16218 26063 16252 26439
rect 16376 26063 16410 26439
rect 16534 26063 16568 26439
rect 16692 26063 16726 26439
rect 16850 26063 16884 26439
rect 15270 25427 15304 25803
rect 15428 25427 15462 25803
rect 15586 25427 15620 25803
rect 15744 25427 15778 25803
rect 15902 25427 15936 25803
rect 16060 25427 16094 25803
rect 16218 25427 16252 25803
rect 16376 25427 16410 25803
rect 16534 25427 16568 25803
rect 16692 25427 16726 25803
rect 16850 25427 16884 25803
rect 6490 24603 6524 24979
rect 6586 24603 6620 24979
rect 6682 24603 6716 24979
rect 6778 24603 6812 24979
rect 6874 24603 6908 24979
rect 6970 24603 7004 24979
rect 7066 24603 7100 24979
rect 7162 24603 7196 24979
rect 7258 24603 7292 24979
rect 7354 24603 7388 24979
rect 7450 24603 7484 24979
rect 7546 24603 7580 24979
rect 7642 24603 7676 24979
rect 7738 24603 7772 24979
rect 7834 24603 7868 24979
rect 7930 24603 7964 24979
rect 6490 23967 6524 24343
rect 6586 23967 6620 24343
rect 6682 23967 6716 24343
rect 6778 23967 6812 24343
rect 6874 23967 6908 24343
rect 6970 23967 7004 24343
rect 7066 23967 7100 24343
rect 7162 23967 7196 24343
rect 7258 23967 7292 24343
rect 7354 23967 7388 24343
rect 7450 23967 7484 24343
rect 7546 23967 7580 24343
rect 7642 23967 7676 24343
rect 7738 23967 7772 24343
rect 7834 23967 7868 24343
rect 7930 23967 7964 24343
rect 8710 24603 8744 24979
rect 8806 24603 8840 24979
rect 8902 24603 8936 24979
rect 8998 24603 9032 24979
rect 9094 24603 9128 24979
rect 9190 24603 9224 24979
rect 9286 24603 9320 24979
rect 9382 24603 9416 24979
rect 9478 24603 9512 24979
rect 9574 24603 9608 24979
rect 9670 24603 9704 24979
rect 9766 24603 9800 24979
rect 9862 24603 9896 24979
rect 9958 24603 9992 24979
rect 10054 24603 10088 24979
rect 10150 24603 10184 24979
rect 8710 23967 8744 24343
rect 8806 23967 8840 24343
rect 8902 23967 8936 24343
rect 8998 23967 9032 24343
rect 9094 23967 9128 24343
rect 9190 23967 9224 24343
rect 9286 23967 9320 24343
rect 9382 23967 9416 24343
rect 9478 23967 9512 24343
rect 9574 23967 9608 24343
rect 9670 23967 9704 24343
rect 9766 23967 9800 24343
rect 9862 23967 9896 24343
rect 9958 23967 9992 24343
rect 10054 23967 10088 24343
rect 10150 23967 10184 24343
rect 10890 24603 10924 24979
rect 10986 24603 11020 24979
rect 11082 24603 11116 24979
rect 11178 24603 11212 24979
rect 11274 24603 11308 24979
rect 11370 24603 11404 24979
rect 11466 24603 11500 24979
rect 11562 24603 11596 24979
rect 11658 24603 11692 24979
rect 11754 24603 11788 24979
rect 11850 24603 11884 24979
rect 11946 24603 11980 24979
rect 12042 24603 12076 24979
rect 12138 24603 12172 24979
rect 12234 24603 12268 24979
rect 12330 24603 12364 24979
rect 10890 23967 10924 24343
rect 10986 23967 11020 24343
rect 11082 23967 11116 24343
rect 11178 23967 11212 24343
rect 11274 23967 11308 24343
rect 11370 23967 11404 24343
rect 11466 23967 11500 24343
rect 11562 23967 11596 24343
rect 11658 23967 11692 24343
rect 11754 23967 11788 24343
rect 11850 23967 11884 24343
rect 11946 23967 11980 24343
rect 12042 23967 12076 24343
rect 12138 23967 12172 24343
rect 12234 23967 12268 24343
rect 12330 23967 12364 24343
rect 13070 24603 13104 24979
rect 13166 24603 13200 24979
rect 13262 24603 13296 24979
rect 13358 24603 13392 24979
rect 13454 24603 13488 24979
rect 13550 24603 13584 24979
rect 13646 24603 13680 24979
rect 13742 24603 13776 24979
rect 13838 24603 13872 24979
rect 13934 24603 13968 24979
rect 14030 24603 14064 24979
rect 14126 24603 14160 24979
rect 14222 24603 14256 24979
rect 14318 24603 14352 24979
rect 14414 24603 14448 24979
rect 14510 24603 14544 24979
rect 13070 23967 13104 24343
rect 13166 23967 13200 24343
rect 13262 23967 13296 24343
rect 13358 23967 13392 24343
rect 13454 23967 13488 24343
rect 13550 23967 13584 24343
rect 13646 23967 13680 24343
rect 13742 23967 13776 24343
rect 13838 23967 13872 24343
rect 13934 23967 13968 24343
rect 14030 23967 14064 24343
rect 14126 23967 14160 24343
rect 14222 23967 14256 24343
rect 14318 23967 14352 24343
rect 14414 23967 14448 24343
rect 14510 23967 14544 24343
rect 15270 24603 15304 24979
rect 15366 24603 15400 24979
rect 15462 24603 15496 24979
rect 15558 24603 15592 24979
rect 15654 24603 15688 24979
rect 15750 24603 15784 24979
rect 15846 24603 15880 24979
rect 15942 24603 15976 24979
rect 16038 24603 16072 24979
rect 16134 24603 16168 24979
rect 16230 24603 16264 24979
rect 16326 24603 16360 24979
rect 16422 24603 16456 24979
rect 16518 24603 16552 24979
rect 16614 24603 16648 24979
rect 16710 24603 16744 24979
rect 15270 23967 15304 24343
rect 15366 23967 15400 24343
rect 15462 23967 15496 24343
rect 15558 23967 15592 24343
rect 15654 23967 15688 24343
rect 15750 23967 15784 24343
rect 15846 23967 15880 24343
rect 15942 23967 15976 24343
rect 16038 23967 16072 24343
rect 16134 23967 16168 24343
rect 16230 23967 16264 24343
rect 16326 23967 16360 24343
rect 16422 23967 16456 24343
rect 16518 23967 16552 24343
rect 16614 23967 16648 24343
rect 16710 23967 16744 24343
rect 19051 25048 19227 25082
rect 19051 23390 19227 23424
rect 18310 22635 18344 23011
rect 18406 22635 18440 23011
rect 18502 22635 18536 23011
rect 18598 22635 18632 23011
rect 18694 22635 18728 23011
rect 18790 22635 18824 23011
rect 18886 22635 18920 23011
rect 18982 22635 19016 23011
rect 19078 22635 19112 23011
rect 19174 22635 19208 23011
rect 19270 22635 19304 23011
rect 5126 9895 5160 10271
rect 5222 9895 5256 10271
rect 5318 9895 5352 10271
rect 5414 9895 5448 10271
rect 5510 9895 5544 10271
rect 5606 9895 5640 10271
rect 5702 9895 5736 10271
rect 5798 9895 5832 10271
rect 5894 9895 5928 10271
rect 5990 9895 6024 10271
rect 6086 9895 6120 10271
rect 6182 9895 6216 10271
rect 6278 9895 6312 10271
rect 6374 9895 6408 10271
rect 6470 9895 6504 10271
rect 6566 9895 6600 10271
rect 6662 9895 6696 10271
rect 6758 9895 6792 10271
rect 6854 9895 6888 10271
rect 6950 9895 6984 10271
rect 7046 9895 7080 10271
rect 5126 9259 5160 9635
rect 5222 9259 5256 9635
rect 5318 9259 5352 9635
rect 5414 9259 5448 9635
rect 5510 9259 5544 9635
rect 5606 9259 5640 9635
rect 5702 9259 5736 9635
rect 5798 9259 5832 9635
rect 5894 9259 5928 9635
rect 5990 9259 6024 9635
rect 6086 9259 6120 9635
rect 6182 9259 6216 9635
rect 6278 9259 6312 9635
rect 6374 9259 6408 9635
rect 6470 9259 6504 9635
rect 6566 9259 6600 9635
rect 6662 9259 6696 9635
rect 6758 9259 6792 9635
rect 6854 9259 6888 9635
rect 6950 9259 6984 9635
rect 7046 9259 7080 9635
rect 19526 9895 19560 10271
rect 19622 9895 19656 10271
rect 19718 9895 19752 10271
rect 19814 9895 19848 10271
rect 19910 9895 19944 10271
rect 20006 9895 20040 10271
rect 20102 9895 20136 10271
rect 20198 9895 20232 10271
rect 20294 9895 20328 10271
rect 20390 9895 20424 10271
rect 20486 9895 20520 10271
rect 20582 9895 20616 10271
rect 20678 9895 20712 10271
rect 20774 9895 20808 10271
rect 20870 9895 20904 10271
rect 20966 9895 21000 10271
rect 21062 9895 21096 10271
rect 21158 9895 21192 10271
rect 21254 9895 21288 10271
rect 21350 9895 21384 10271
rect 21446 9895 21480 10271
rect 19526 9259 19560 9635
rect 19622 9259 19656 9635
rect 19718 9259 19752 9635
rect 19814 9259 19848 9635
rect 19910 9259 19944 9635
rect 20006 9259 20040 9635
rect 20102 9259 20136 9635
rect 20198 9259 20232 9635
rect 20294 9259 20328 9635
rect 20390 9259 20424 9635
rect 20486 9259 20520 9635
rect 20582 9259 20616 9635
rect 20678 9259 20712 9635
rect 20774 9259 20808 9635
rect 20870 9259 20904 9635
rect 20966 9259 21000 9635
rect 21062 9259 21096 9635
rect 21158 9259 21192 9635
rect 21254 9259 21288 9635
rect 21350 9259 21384 9635
rect 21446 9259 21480 9635
<< psubdiff >>
rect 18196 25182 18292 25216
rect 18642 25182 18738 25216
rect 18196 25120 18230 25182
rect 6496 23562 6592 23596
rect 7622 23562 7718 23596
rect 6496 23500 6530 23562
rect 7684 23500 7718 23562
rect 6496 21646 6530 21708
rect 7684 21646 7718 21708
rect 6496 21612 6592 21646
rect 7622 21612 7718 21646
rect 8216 23562 8312 23596
rect 9342 23562 9438 23596
rect 8216 23500 8250 23562
rect 9404 23500 9438 23562
rect 8216 21646 8250 21708
rect 18704 25120 18738 25182
rect 18196 23326 18230 23388
rect 18704 23326 18738 23388
rect 18196 23292 18292 23326
rect 18642 23292 18738 23326
rect 9404 21646 9438 21708
rect 8216 21612 8312 21646
rect 9342 21612 9438 21646
rect 18196 22304 18292 22338
rect 19322 22304 19418 22338
rect 18196 22242 18230 22304
rect 6496 21416 6592 21450
rect 7952 21416 8048 21450
rect 6496 21354 6530 21416
rect 8014 21354 8048 21416
rect 6496 17646 6530 17708
rect 8014 17646 8048 17708
rect 6496 17612 6592 17646
rect 7952 17612 8048 17646
rect 8216 21416 8312 21450
rect 9672 21416 9768 21450
rect 8216 21354 8250 21416
rect 9734 21354 9768 21416
rect 8216 17646 8250 17708
rect 19384 22242 19418 22304
rect 18196 21006 18230 21068
rect 19384 21006 19418 21068
rect 18196 20972 18292 21006
rect 19322 20972 19418 21006
rect 18196 20820 18292 20854
rect 19652 20820 19748 20854
rect 18196 20758 18230 20820
rect 10056 19866 10152 19900
rect 10894 19866 10990 19900
rect 10056 19804 10090 19866
rect 10956 19804 10990 19866
rect 10056 19186 10090 19248
rect 10956 19186 10990 19248
rect 10056 19152 10152 19186
rect 10894 19152 10990 19186
rect 9734 17646 9768 17708
rect 8216 17612 8312 17646
rect 9672 17612 9768 17646
rect 10056 18944 10152 18978
rect 11182 18944 11278 18978
rect 10056 18882 10090 18944
rect 11244 18882 11278 18944
rect 10056 17646 10090 17708
rect 19714 20758 19748 20820
rect 18196 18286 18230 18348
rect 19714 18286 19748 18348
rect 18196 18252 18292 18286
rect 19652 18252 19748 18286
rect 11244 17646 11278 17708
rect 10056 17612 10152 17646
rect 11182 17612 11278 17646
rect 2472 11214 2568 11248
rect 4808 11214 4904 11248
rect 2472 11152 2506 11214
rect 4870 11152 4904 11214
rect 2472 9358 2506 9420
rect 16872 11214 16968 11248
rect 19208 11214 19304 11248
rect 16872 11152 16906 11214
rect 4870 9358 4904 9420
rect 2472 9324 2568 9358
rect 4808 9324 4904 9358
rect -10164 8374 -10068 8408
rect -9038 8374 -8942 8408
rect -10164 8312 -10130 8374
rect -8976 8312 -8942 8374
rect -10164 6458 -10130 6520
rect -8976 6458 -8942 6520
rect -10164 6424 -10068 6458
rect -9038 6424 -8942 6458
rect -8844 8310 -8748 8344
rect -8392 8310 -8296 8344
rect -8844 8248 -8810 8310
rect -8330 8248 -8296 8310
rect -8844 6458 -8810 6520
rect -8330 6458 -8296 6520
rect -8844 6424 -8748 6458
rect -8392 6424 -8296 6458
rect -10164 6294 -10068 6328
rect -9038 6294 -8942 6328
rect -10164 6232 -10130 6294
rect -8976 6232 -8942 6294
rect -10164 4378 -10130 4440
rect 1576 8870 1672 8904
rect 3662 8870 3758 8904
rect 1576 8808 1610 8870
rect 3724 8808 3758 8870
rect 1576 8190 1610 8252
rect 3724 8190 3758 8252
rect 1576 8156 1672 8190
rect 3662 8156 3758 8190
rect 1576 8050 1672 8084
rect 3662 8050 3758 8084
rect 1576 7988 1610 8050
rect 3724 7988 3758 8050
rect 1576 7370 1610 7432
rect 3724 7370 3758 7432
rect 1576 7336 1672 7370
rect 3662 7336 3758 7370
rect 1576 7230 1672 7264
rect 3662 7230 3758 7264
rect 1576 7168 1610 7230
rect 3724 7168 3758 7230
rect 1576 6550 1610 6612
rect 3724 6550 3758 6612
rect 1576 6516 1672 6550
rect 3662 6516 3758 6550
rect 7512 10402 7608 10436
rect 9598 10402 9694 10436
rect 7512 10340 7546 10402
rect 5012 8836 5108 8870
rect 7098 8836 7194 8870
rect 5012 8774 5046 8836
rect 7160 8774 7194 8836
rect 5012 7538 5046 7600
rect 7160 7538 7194 7600
rect 5012 7504 5108 7538
rect 7098 7504 7194 7538
rect -8976 4378 -8942 4440
rect -10164 4344 -10068 4378
rect -9038 4344 -8942 4378
rect 112 6014 208 6048
rect 1238 6014 1334 6048
rect 112 5952 146 6014
rect -10164 4148 -10068 4182
rect -8708 4148 -8612 4182
rect -10164 4086 -10130 4148
rect -8646 4086 -8612 4148
rect -10164 378 -10130 440
rect 1300 5952 1334 6014
rect 112 4098 146 4160
rect 1300 4098 1334 4160
rect 112 4064 208 4098
rect 1238 4064 1334 4098
rect 1912 6014 2008 6048
rect 3038 6014 3134 6048
rect 1912 5952 1946 6014
rect 3100 5952 3134 6014
rect 1912 4098 1946 4160
rect 3100 4098 3134 4160
rect 1912 4064 2008 4098
rect 3038 4064 3134 4098
rect 3712 6014 3808 6048
rect 4838 6014 4934 6048
rect 3712 5952 3746 6014
rect 4900 5952 4934 6014
rect 3712 4098 3746 4160
rect 4900 4098 4934 4160
rect 3712 4064 3808 4098
rect 4838 4064 4934 4098
rect 5512 6014 5608 6048
rect 6638 6014 6734 6048
rect 5512 5952 5546 6014
rect 6700 5952 6734 6014
rect 5512 4098 5546 4160
rect 9660 10340 9694 10402
rect 7512 4778 7546 4840
rect 19270 11152 19304 11214
rect 16872 9358 16906 9420
rect 19270 9358 19304 9420
rect 16872 9324 16968 9358
rect 19208 9324 19304 9358
rect 15976 8870 16072 8904
rect 18062 8870 18158 8904
rect 15976 8808 16010 8870
rect 18124 8808 18158 8870
rect 15976 8190 16010 8252
rect 18124 8190 18158 8252
rect 15976 8156 16072 8190
rect 18062 8156 18158 8190
rect 15976 8050 16072 8084
rect 18062 8050 18158 8084
rect 15976 7988 16010 8050
rect 18124 7988 18158 8050
rect 15976 7370 16010 7432
rect 18124 7370 18158 7432
rect 15976 7336 16072 7370
rect 18062 7336 18158 7370
rect 15976 7230 16072 7264
rect 18062 7230 18158 7264
rect 15976 7168 16010 7230
rect 18124 7168 18158 7230
rect 15976 6550 16010 6612
rect 18124 6550 18158 6612
rect 15976 6516 16072 6550
rect 18062 6516 18158 6550
rect 21912 10402 22008 10436
rect 23998 10402 24094 10436
rect 21912 10340 21946 10402
rect 19412 8836 19508 8870
rect 21498 8836 21594 8870
rect 19412 8774 19446 8836
rect 21560 8774 21594 8836
rect 19412 7538 19446 7600
rect 21560 7538 21594 7600
rect 19412 7504 19508 7538
rect 21498 7504 21594 7538
rect 9660 4778 9694 4840
rect 7512 4744 7608 4778
rect 9598 4744 9694 4778
rect 14512 6014 14608 6048
rect 15638 6014 15734 6048
rect 14512 5952 14546 6014
rect 6700 4098 6734 4160
rect 5512 4064 5608 4098
rect 6638 4064 6734 4098
rect 15700 5952 15734 6014
rect 14512 4098 14546 4160
rect 15700 4098 15734 4160
rect 14512 4064 14608 4098
rect 15638 4064 15734 4098
rect 16312 6014 16408 6048
rect 17438 6014 17534 6048
rect 16312 5952 16346 6014
rect 17500 5952 17534 6014
rect 16312 4098 16346 4160
rect 17500 4098 17534 4160
rect 16312 4064 16408 4098
rect 17438 4064 17534 4098
rect 18112 6014 18208 6048
rect 19238 6014 19334 6048
rect 18112 5952 18146 6014
rect 19300 5952 19334 6014
rect 18112 4098 18146 4160
rect 19300 4098 19334 4160
rect 18112 4064 18208 4098
rect 19238 4064 19334 4098
rect 19912 6014 20008 6048
rect 21038 6014 21134 6048
rect 19912 5952 19946 6014
rect 21100 5952 21134 6014
rect 19912 4098 19946 4160
rect 24060 10340 24094 10402
rect 21912 4778 21946 4840
rect 24060 4778 24094 4840
rect 21912 4744 22008 4778
rect 23998 4744 24094 4778
rect 21100 4098 21134 4160
rect 19912 4064 20008 4098
rect 21038 4064 21134 4098
rect 112 3868 208 3902
rect 1568 3868 1664 3902
rect 112 3806 146 3868
rect -8500 958 -8290 982
rect -8500 684 -8290 708
rect -8646 378 -8612 440
rect -10164 344 -10068 378
rect -8708 344 -8612 378
rect 1630 3806 1664 3868
rect 112 98 146 160
rect 1630 98 1664 160
rect 112 64 208 98
rect 1568 64 1664 98
rect 1912 3868 2008 3902
rect 3368 3868 3464 3902
rect 1912 3806 1946 3868
rect 3430 3806 3464 3868
rect 1912 98 1946 160
rect 3430 98 3464 160
rect 1912 64 2008 98
rect 3368 64 3464 98
rect 3712 3868 3808 3902
rect 5168 3868 5264 3902
rect 3712 3806 3746 3868
rect 5230 3806 5264 3868
rect 3712 98 3746 160
rect 5230 98 5264 160
rect 3712 64 3808 98
rect 5168 64 5264 98
rect 5512 3868 5608 3902
rect 6968 3868 7064 3902
rect 5512 3806 5546 3868
rect 7030 3806 7064 3868
rect 5512 98 5546 160
rect 7030 98 7064 160
rect 5512 64 5608 98
rect 6968 64 7064 98
rect 14512 3868 14608 3902
rect 15968 3868 16064 3902
rect 14512 3806 14546 3868
rect 16030 3806 16064 3868
rect 14512 98 14546 160
rect 16030 98 16064 160
rect 14512 64 14608 98
rect 15968 64 16064 98
rect 16312 3868 16408 3902
rect 17768 3868 17864 3902
rect 16312 3806 16346 3868
rect 17830 3806 17864 3868
rect 16312 98 16346 160
rect 17830 98 17864 160
rect 16312 64 16408 98
rect 17768 64 17864 98
rect 18112 3868 18208 3902
rect 19568 3868 19664 3902
rect 18112 3806 18146 3868
rect 19630 3806 19664 3868
rect 18112 98 18146 160
rect 19630 98 19664 160
rect 18112 64 18208 98
rect 19568 64 19664 98
rect 19912 3868 20008 3902
rect 21368 3868 21464 3902
rect 19912 3806 19946 3868
rect 21430 3806 21464 3868
rect 19912 98 19946 160
rect 21430 98 21464 160
rect 19912 64 20008 98
rect 21368 64 21464 98
rect -2792 -1188 -2768 -382
rect -1960 -1188 -1936 -382
rect 11608 -1188 11632 -382
rect 12440 -1188 12464 -382
<< nsubdiff >>
rect 6376 27236 6472 27270
rect 8122 27236 8218 27270
rect 6376 27174 6410 27236
rect 8184 27174 8218 27236
rect 6376 25266 6410 25328
rect 8184 25266 8218 25328
rect 6376 25232 6472 25266
rect 8122 25232 8218 25266
rect 8596 27236 8692 27270
rect 10342 27236 10438 27270
rect 8596 27174 8630 27236
rect 10404 27174 10438 27236
rect 8596 25266 8630 25328
rect 10404 25266 10438 25328
rect 8596 25232 8692 25266
rect 10342 25232 10438 25266
rect 10776 27236 10872 27270
rect 12522 27236 12618 27270
rect 10776 27174 10810 27236
rect 12584 27174 12618 27236
rect 10776 25266 10810 25328
rect 12584 25266 12618 25328
rect 10776 25232 10872 25266
rect 12522 25232 12618 25266
rect 12956 27236 13052 27270
rect 14702 27236 14798 27270
rect 12956 27174 12990 27236
rect 14764 27174 14798 27236
rect 12956 25266 12990 25328
rect 14764 25266 14798 25328
rect 12956 25232 13052 25266
rect 14702 25232 14798 25266
rect 15156 27236 15252 27270
rect 16902 27236 16998 27270
rect 15156 27174 15190 27236
rect 16964 27174 16998 27236
rect 15156 25266 15190 25328
rect 16964 25266 16998 25328
rect 15156 25232 15252 25266
rect 16902 25232 16998 25266
rect 6376 25140 6472 25174
rect 7982 25140 8078 25174
rect 6376 25078 6410 25140
rect 8044 25078 8078 25140
rect 6376 23806 6410 23868
rect 8044 23806 8078 23868
rect 6376 23772 6472 23806
rect 7982 23772 8078 23806
rect 8596 25140 8692 25174
rect 10202 25140 10298 25174
rect 8596 25078 8630 25140
rect 10264 25078 10298 25140
rect 8596 23806 8630 23868
rect 10264 23806 10298 23868
rect 8596 23772 8692 23806
rect 10202 23772 10298 23806
rect 10776 25140 10872 25174
rect 12382 25140 12478 25174
rect 10776 25078 10810 25140
rect 12444 25078 12478 25140
rect 10776 23806 10810 23868
rect 12444 23806 12478 23868
rect 10776 23772 10872 23806
rect 12382 23772 12478 23806
rect 12956 25140 13052 25174
rect 14562 25140 14658 25174
rect 12956 25078 12990 25140
rect 14624 25078 14658 25140
rect 12956 23806 12990 23868
rect 14624 23806 14658 23868
rect 12956 23772 13052 23806
rect 14562 23772 14658 23806
rect 15156 25140 15252 25174
rect 16762 25140 16858 25174
rect 15156 25078 15190 25140
rect 16824 25078 16858 25140
rect 15156 23806 15190 23868
rect 16824 23806 16858 23868
rect 15156 23772 15252 23806
rect 16762 23772 16858 23806
rect 18856 25162 18952 25196
rect 19326 25162 19422 25196
rect 18856 25100 18890 25162
rect 19388 25100 19422 25162
rect 18856 23310 18890 23372
rect 19388 23310 19422 23372
rect 18856 23276 18952 23310
rect 19326 23276 19422 23310
rect 18196 23172 18292 23206
rect 19322 23172 19418 23206
rect 18196 23110 18230 23172
rect 19384 23110 19418 23172
rect 18196 22474 18230 22536
rect 19384 22474 19418 22536
rect 18196 22440 18292 22474
rect 19322 22440 19418 22474
rect 5012 10432 5108 10466
rect 7098 10432 7194 10466
rect 5012 10370 5046 10432
rect 1277 9183 4063 9203
rect 1277 9149 1357 9183
rect 3983 9149 4063 9183
rect 1277 9129 4063 9149
rect 1277 9123 1351 9129
rect 1277 6297 1297 9123
rect 1331 6297 1351 9123
rect 3989 9123 4063 9129
rect 1277 6291 1351 6297
rect 3989 6297 4009 9123
rect 4043 6297 4063 9123
rect 7160 10370 7194 10432
rect 5012 9098 5046 9160
rect 7160 9098 7194 9160
rect 5012 9064 5108 9098
rect 7098 9064 7194 9098
rect 3989 6291 4063 6297
rect 1277 6271 4063 6291
rect 1277 6237 1357 6271
rect 3983 6237 4063 6271
rect 1277 6217 4063 6237
rect 19412 10432 19508 10466
rect 21498 10432 21594 10466
rect 19412 10370 19446 10432
rect 15677 9183 18463 9203
rect 15677 9149 15757 9183
rect 18383 9149 18463 9183
rect 15677 9129 18463 9149
rect 15677 9123 15751 9129
rect 15677 6297 15697 9123
rect 15731 6297 15751 9123
rect 18389 9123 18463 9129
rect 15677 6291 15751 6297
rect 18389 6297 18409 9123
rect 18443 6297 18463 9123
rect 21560 10370 21594 10432
rect 19412 9098 19446 9160
rect 21560 9098 21594 9160
rect 19412 9064 19508 9098
rect 21498 9064 21594 9098
rect 18389 6291 18463 6297
rect 15677 6271 18463 6291
rect 15677 6237 15757 6271
rect 18383 6237 18463 6271
rect 15677 6217 18463 6237
<< psubdiffcont >>
rect 18292 25182 18642 25216
rect 6592 23562 7622 23596
rect 6496 21708 6530 23500
rect 7684 21708 7718 23500
rect 6592 21612 7622 21646
rect 8312 23562 9342 23596
rect 8216 21708 8250 23500
rect 9404 21708 9438 23500
rect 18196 23388 18230 25120
rect 18704 23388 18738 25120
rect 18292 23292 18642 23326
rect 8312 21612 9342 21646
rect 18292 22304 19322 22338
rect 6592 21416 7952 21450
rect 6496 17708 6530 21354
rect 8014 17708 8048 21354
rect 6592 17612 7952 17646
rect 8312 21416 9672 21450
rect 8216 17708 8250 21354
rect 9734 17708 9768 21354
rect 18196 21068 18230 22242
rect 19384 21068 19418 22242
rect 18292 20972 19322 21006
rect 18292 20820 19652 20854
rect 10152 19866 10894 19900
rect 10056 19248 10090 19804
rect 10956 19248 10990 19804
rect 10152 19152 10894 19186
rect 8312 17612 9672 17646
rect 10152 18944 11182 18978
rect 10056 17708 10090 18882
rect 11244 17708 11278 18882
rect 18196 18348 18230 20758
rect 19714 18348 19748 20758
rect 18292 18252 19652 18286
rect 10152 17612 11182 17646
rect 2568 11214 4808 11248
rect 2472 9420 2506 11152
rect 4870 9420 4904 11152
rect 16968 11214 19208 11248
rect 2568 9324 4808 9358
rect -10068 8374 -9038 8408
rect -10164 6520 -10130 8312
rect -8976 6520 -8942 8312
rect -10068 6424 -9038 6458
rect -8748 8310 -8392 8344
rect -8844 6520 -8810 8248
rect -8330 6520 -8296 8248
rect -8748 6424 -8392 6458
rect -10068 6294 -9038 6328
rect -10164 4440 -10130 6232
rect -8976 4440 -8942 6232
rect 1672 8870 3662 8904
rect 1576 8252 1610 8808
rect 3724 8252 3758 8808
rect 1672 8156 3662 8190
rect 1672 8050 3662 8084
rect 1576 7432 1610 7988
rect 3724 7432 3758 7988
rect 1672 7336 3662 7370
rect 1672 7230 3662 7264
rect 1576 6612 1610 7168
rect 3724 6612 3758 7168
rect 1672 6516 3662 6550
rect 7608 10402 9598 10436
rect 5108 8836 7098 8870
rect 5012 7600 5046 8774
rect 7160 7600 7194 8774
rect 5108 7504 7098 7538
rect -10068 4344 -9038 4378
rect 208 6014 1238 6048
rect -10068 4148 -8708 4182
rect -10164 440 -10130 4086
rect -8646 440 -8612 4086
rect 112 4160 146 5952
rect 1300 4160 1334 5952
rect 208 4064 1238 4098
rect 2008 6014 3038 6048
rect 1912 4160 1946 5952
rect 3100 4160 3134 5952
rect 2008 4064 3038 4098
rect 3808 6014 4838 6048
rect 3712 4160 3746 5952
rect 4900 4160 4934 5952
rect 3808 4064 4838 4098
rect 5608 6014 6638 6048
rect 5512 4160 5546 5952
rect 6700 4160 6734 5952
rect 7512 4840 7546 10340
rect 9660 4840 9694 10340
rect 16872 9420 16906 11152
rect 19270 9420 19304 11152
rect 16968 9324 19208 9358
rect 16072 8870 18062 8904
rect 15976 8252 16010 8808
rect 18124 8252 18158 8808
rect 16072 8156 18062 8190
rect 16072 8050 18062 8084
rect 15976 7432 16010 7988
rect 18124 7432 18158 7988
rect 16072 7336 18062 7370
rect 16072 7230 18062 7264
rect 15976 6612 16010 7168
rect 18124 6612 18158 7168
rect 16072 6516 18062 6550
rect 22008 10402 23998 10436
rect 19508 8836 21498 8870
rect 19412 7600 19446 8774
rect 21560 7600 21594 8774
rect 19508 7504 21498 7538
rect 7608 4744 9598 4778
rect 14608 6014 15638 6048
rect 5608 4064 6638 4098
rect 14512 4160 14546 5952
rect 15700 4160 15734 5952
rect 14608 4064 15638 4098
rect 16408 6014 17438 6048
rect 16312 4160 16346 5952
rect 17500 4160 17534 5952
rect 16408 4064 17438 4098
rect 18208 6014 19238 6048
rect 18112 4160 18146 5952
rect 19300 4160 19334 5952
rect 18208 4064 19238 4098
rect 20008 6014 21038 6048
rect 19912 4160 19946 5952
rect 21100 4160 21134 5952
rect 21912 4840 21946 10340
rect 24060 4840 24094 10340
rect 22008 4744 23998 4778
rect 20008 4064 21038 4098
rect 208 3868 1568 3902
rect -8500 708 -8290 958
rect -10068 344 -8708 378
rect 112 160 146 3806
rect 1630 160 1664 3806
rect 208 64 1568 98
rect 2008 3868 3368 3902
rect 1912 160 1946 3806
rect 3430 160 3464 3806
rect 2008 64 3368 98
rect 3808 3868 5168 3902
rect 3712 160 3746 3806
rect 5230 160 5264 3806
rect 3808 64 5168 98
rect 5608 3868 6968 3902
rect 5512 160 5546 3806
rect 7030 160 7064 3806
rect 5608 64 6968 98
rect 14608 3868 15968 3902
rect 14512 160 14546 3806
rect 16030 160 16064 3806
rect 14608 64 15968 98
rect 16408 3868 17768 3902
rect 16312 160 16346 3806
rect 17830 160 17864 3806
rect 16408 64 17768 98
rect 18208 3868 19568 3902
rect 18112 160 18146 3806
rect 19630 160 19664 3806
rect 18208 64 19568 98
rect 20008 3868 21368 3902
rect 19912 160 19946 3806
rect 21430 160 21464 3806
rect 20008 64 21368 98
rect -2768 -1188 -1960 -382
rect 11632 -1188 12440 -382
<< nsubdiffcont >>
rect 6472 27236 8122 27270
rect 6376 25328 6410 27174
rect 8184 25328 8218 27174
rect 6472 25232 8122 25266
rect 8692 27236 10342 27270
rect 8596 25328 8630 27174
rect 10404 25328 10438 27174
rect 8692 25232 10342 25266
rect 10872 27236 12522 27270
rect 10776 25328 10810 27174
rect 12584 25328 12618 27174
rect 10872 25232 12522 25266
rect 13052 27236 14702 27270
rect 12956 25328 12990 27174
rect 14764 25328 14798 27174
rect 13052 25232 14702 25266
rect 15252 27236 16902 27270
rect 15156 25328 15190 27174
rect 16964 25328 16998 27174
rect 15252 25232 16902 25266
rect 6472 25140 7982 25174
rect 6376 23868 6410 25078
rect 8044 23868 8078 25078
rect 6472 23772 7982 23806
rect 8692 25140 10202 25174
rect 8596 23868 8630 25078
rect 10264 23868 10298 25078
rect 8692 23772 10202 23806
rect 10872 25140 12382 25174
rect 10776 23868 10810 25078
rect 12444 23868 12478 25078
rect 10872 23772 12382 23806
rect 13052 25140 14562 25174
rect 12956 23868 12990 25078
rect 14624 23868 14658 25078
rect 13052 23772 14562 23806
rect 15252 25140 16762 25174
rect 15156 23868 15190 25078
rect 16824 23868 16858 25078
rect 15252 23772 16762 23806
rect 18952 25162 19326 25196
rect 18856 23372 18890 25100
rect 19388 23372 19422 25100
rect 18952 23276 19326 23310
rect 18292 23172 19322 23206
rect 18196 22536 18230 23110
rect 19384 22536 19418 23110
rect 18292 22440 19322 22474
rect 5108 10432 7098 10466
rect 1357 9149 3983 9183
rect 1297 6297 1331 9123
rect 4009 6297 4043 9123
rect 5012 9160 5046 10370
rect 7160 9160 7194 10370
rect 5108 9064 7098 9098
rect 1357 6237 3983 6271
rect 19508 10432 21498 10466
rect 15757 9149 18383 9183
rect 15697 6297 15731 9123
rect 18409 6297 18443 9123
rect 19412 9160 19446 10370
rect 21560 9160 21594 10370
rect 19508 9064 21498 9098
rect 15757 6237 18383 6271
<< poly >>
rect 6536 27168 6636 27184
rect 6536 27134 6552 27168
rect 6620 27134 6636 27168
rect 6536 27087 6636 27134
rect 6694 27168 6794 27184
rect 6694 27134 6710 27168
rect 6778 27134 6794 27168
rect 6694 27087 6794 27134
rect 6852 27168 6952 27184
rect 6852 27134 6868 27168
rect 6936 27134 6952 27168
rect 6852 27087 6952 27134
rect 7010 27168 7110 27184
rect 7010 27134 7026 27168
rect 7094 27134 7110 27168
rect 7010 27087 7110 27134
rect 7168 27168 7268 27184
rect 7168 27134 7184 27168
rect 7252 27134 7268 27168
rect 7168 27087 7268 27134
rect 7326 27168 7426 27184
rect 7326 27134 7342 27168
rect 7410 27134 7426 27168
rect 7326 27087 7426 27134
rect 7484 27168 7584 27184
rect 7484 27134 7500 27168
rect 7568 27134 7584 27168
rect 7484 27087 7584 27134
rect 7642 27168 7742 27184
rect 7642 27134 7658 27168
rect 7726 27134 7742 27168
rect 7642 27087 7742 27134
rect 7800 27168 7900 27184
rect 7800 27134 7816 27168
rect 7884 27134 7900 27168
rect 7800 27087 7900 27134
rect 7958 27168 8058 27184
rect 7958 27134 7974 27168
rect 8042 27134 8058 27168
rect 7958 27087 8058 27134
rect 6536 26640 6636 26687
rect 6536 26606 6552 26640
rect 6620 26606 6636 26640
rect 6536 26590 6636 26606
rect 6694 26640 6794 26687
rect 6694 26606 6710 26640
rect 6778 26606 6794 26640
rect 6694 26590 6794 26606
rect 6852 26640 6952 26687
rect 6852 26606 6868 26640
rect 6936 26606 6952 26640
rect 6852 26590 6952 26606
rect 7010 26640 7110 26687
rect 7010 26606 7026 26640
rect 7094 26606 7110 26640
rect 7010 26590 7110 26606
rect 7168 26640 7268 26687
rect 7168 26606 7184 26640
rect 7252 26606 7268 26640
rect 7168 26590 7268 26606
rect 7326 26640 7426 26687
rect 7326 26606 7342 26640
rect 7410 26606 7426 26640
rect 7326 26590 7426 26606
rect 7484 26640 7584 26687
rect 7484 26606 7500 26640
rect 7568 26606 7584 26640
rect 7484 26590 7584 26606
rect 7642 26640 7742 26687
rect 7642 26606 7658 26640
rect 7726 26606 7742 26640
rect 7642 26590 7742 26606
rect 7800 26640 7900 26687
rect 7800 26606 7816 26640
rect 7884 26606 7900 26640
rect 7800 26590 7900 26606
rect 7958 26640 8058 26687
rect 7958 26606 7974 26640
rect 8042 26606 8058 26640
rect 7958 26590 8058 26606
rect 6536 26532 6636 26548
rect 6536 26498 6552 26532
rect 6620 26498 6636 26532
rect 6536 26451 6636 26498
rect 6694 26532 6794 26548
rect 6694 26498 6710 26532
rect 6778 26498 6794 26532
rect 6694 26451 6794 26498
rect 6852 26532 6952 26548
rect 6852 26498 6868 26532
rect 6936 26498 6952 26532
rect 6852 26451 6952 26498
rect 7010 26532 7110 26548
rect 7010 26498 7026 26532
rect 7094 26498 7110 26532
rect 7010 26451 7110 26498
rect 7168 26532 7268 26548
rect 7168 26498 7184 26532
rect 7252 26498 7268 26532
rect 7168 26451 7268 26498
rect 7326 26532 7426 26548
rect 7326 26498 7342 26532
rect 7410 26498 7426 26532
rect 7326 26451 7426 26498
rect 7484 26532 7584 26548
rect 7484 26498 7500 26532
rect 7568 26498 7584 26532
rect 7484 26451 7584 26498
rect 7642 26532 7742 26548
rect 7642 26498 7658 26532
rect 7726 26498 7742 26532
rect 7642 26451 7742 26498
rect 7800 26532 7900 26548
rect 7800 26498 7816 26532
rect 7884 26498 7900 26532
rect 7800 26451 7900 26498
rect 7958 26532 8058 26548
rect 7958 26498 7974 26532
rect 8042 26498 8058 26532
rect 7958 26451 8058 26498
rect 6536 26004 6636 26051
rect 6536 25970 6552 26004
rect 6620 25970 6636 26004
rect 6536 25954 6636 25970
rect 6694 26004 6794 26051
rect 6694 25970 6710 26004
rect 6778 25970 6794 26004
rect 6694 25954 6794 25970
rect 6852 26004 6952 26051
rect 6852 25970 6868 26004
rect 6936 25970 6952 26004
rect 6852 25954 6952 25970
rect 7010 26004 7110 26051
rect 7010 25970 7026 26004
rect 7094 25970 7110 26004
rect 7010 25954 7110 25970
rect 7168 26004 7268 26051
rect 7168 25970 7184 26004
rect 7252 25970 7268 26004
rect 7168 25954 7268 25970
rect 7326 26004 7426 26051
rect 7326 25970 7342 26004
rect 7410 25970 7426 26004
rect 7326 25954 7426 25970
rect 7484 26004 7584 26051
rect 7484 25970 7500 26004
rect 7568 25970 7584 26004
rect 7484 25954 7584 25970
rect 7642 26004 7742 26051
rect 7642 25970 7658 26004
rect 7726 25970 7742 26004
rect 7642 25954 7742 25970
rect 7800 26004 7900 26051
rect 7800 25970 7816 26004
rect 7884 25970 7900 26004
rect 7800 25954 7900 25970
rect 7958 26004 8058 26051
rect 7958 25970 7974 26004
rect 8042 25970 8058 26004
rect 7958 25954 8058 25970
rect 6536 25896 6636 25912
rect 6536 25862 6552 25896
rect 6620 25862 6636 25896
rect 6536 25815 6636 25862
rect 6694 25896 6794 25912
rect 6694 25862 6710 25896
rect 6778 25862 6794 25896
rect 6694 25815 6794 25862
rect 6852 25896 6952 25912
rect 6852 25862 6868 25896
rect 6936 25862 6952 25896
rect 6852 25815 6952 25862
rect 7010 25896 7110 25912
rect 7010 25862 7026 25896
rect 7094 25862 7110 25896
rect 7010 25815 7110 25862
rect 7168 25896 7268 25912
rect 7168 25862 7184 25896
rect 7252 25862 7268 25896
rect 7168 25815 7268 25862
rect 7326 25896 7426 25912
rect 7326 25862 7342 25896
rect 7410 25862 7426 25896
rect 7326 25815 7426 25862
rect 7484 25896 7584 25912
rect 7484 25862 7500 25896
rect 7568 25862 7584 25896
rect 7484 25815 7584 25862
rect 7642 25896 7742 25912
rect 7642 25862 7658 25896
rect 7726 25862 7742 25896
rect 7642 25815 7742 25862
rect 7800 25896 7900 25912
rect 7800 25862 7816 25896
rect 7884 25862 7900 25896
rect 7800 25815 7900 25862
rect 7958 25896 8058 25912
rect 7958 25862 7974 25896
rect 8042 25862 8058 25896
rect 7958 25815 8058 25862
rect 6536 25368 6636 25415
rect 6536 25334 6552 25368
rect 6620 25334 6636 25368
rect 6536 25318 6636 25334
rect 6694 25368 6794 25415
rect 6694 25334 6710 25368
rect 6778 25334 6794 25368
rect 6694 25318 6794 25334
rect 6852 25368 6952 25415
rect 6852 25334 6868 25368
rect 6936 25334 6952 25368
rect 6852 25318 6952 25334
rect 7010 25368 7110 25415
rect 7010 25334 7026 25368
rect 7094 25334 7110 25368
rect 7010 25318 7110 25334
rect 7168 25368 7268 25415
rect 7168 25334 7184 25368
rect 7252 25334 7268 25368
rect 7168 25318 7268 25334
rect 7326 25368 7426 25415
rect 7326 25334 7342 25368
rect 7410 25334 7426 25368
rect 7326 25318 7426 25334
rect 7484 25368 7584 25415
rect 7484 25334 7500 25368
rect 7568 25334 7584 25368
rect 7484 25318 7584 25334
rect 7642 25368 7742 25415
rect 7642 25334 7658 25368
rect 7726 25334 7742 25368
rect 7642 25318 7742 25334
rect 7800 25368 7900 25415
rect 7800 25334 7816 25368
rect 7884 25334 7900 25368
rect 7800 25318 7900 25334
rect 7958 25368 8058 25415
rect 7958 25334 7974 25368
rect 8042 25334 8058 25368
rect 7958 25318 8058 25334
rect 8756 27168 8856 27184
rect 8756 27134 8772 27168
rect 8840 27134 8856 27168
rect 8756 27087 8856 27134
rect 8914 27168 9014 27184
rect 8914 27134 8930 27168
rect 8998 27134 9014 27168
rect 8914 27087 9014 27134
rect 9072 27168 9172 27184
rect 9072 27134 9088 27168
rect 9156 27134 9172 27168
rect 9072 27087 9172 27134
rect 9230 27168 9330 27184
rect 9230 27134 9246 27168
rect 9314 27134 9330 27168
rect 9230 27087 9330 27134
rect 9388 27168 9488 27184
rect 9388 27134 9404 27168
rect 9472 27134 9488 27168
rect 9388 27087 9488 27134
rect 9546 27168 9646 27184
rect 9546 27134 9562 27168
rect 9630 27134 9646 27168
rect 9546 27087 9646 27134
rect 9704 27168 9804 27184
rect 9704 27134 9720 27168
rect 9788 27134 9804 27168
rect 9704 27087 9804 27134
rect 9862 27168 9962 27184
rect 9862 27134 9878 27168
rect 9946 27134 9962 27168
rect 9862 27087 9962 27134
rect 10020 27168 10120 27184
rect 10020 27134 10036 27168
rect 10104 27134 10120 27168
rect 10020 27087 10120 27134
rect 10178 27168 10278 27184
rect 10178 27134 10194 27168
rect 10262 27134 10278 27168
rect 10178 27087 10278 27134
rect 8756 26640 8856 26687
rect 8756 26606 8772 26640
rect 8840 26606 8856 26640
rect 8756 26590 8856 26606
rect 8914 26640 9014 26687
rect 8914 26606 8930 26640
rect 8998 26606 9014 26640
rect 8914 26590 9014 26606
rect 9072 26640 9172 26687
rect 9072 26606 9088 26640
rect 9156 26606 9172 26640
rect 9072 26590 9172 26606
rect 9230 26640 9330 26687
rect 9230 26606 9246 26640
rect 9314 26606 9330 26640
rect 9230 26590 9330 26606
rect 9388 26640 9488 26687
rect 9388 26606 9404 26640
rect 9472 26606 9488 26640
rect 9388 26590 9488 26606
rect 9546 26640 9646 26687
rect 9546 26606 9562 26640
rect 9630 26606 9646 26640
rect 9546 26590 9646 26606
rect 9704 26640 9804 26687
rect 9704 26606 9720 26640
rect 9788 26606 9804 26640
rect 9704 26590 9804 26606
rect 9862 26640 9962 26687
rect 9862 26606 9878 26640
rect 9946 26606 9962 26640
rect 9862 26590 9962 26606
rect 10020 26640 10120 26687
rect 10020 26606 10036 26640
rect 10104 26606 10120 26640
rect 10020 26590 10120 26606
rect 10178 26640 10278 26687
rect 10178 26606 10194 26640
rect 10262 26606 10278 26640
rect 10178 26590 10278 26606
rect 8756 26532 8856 26548
rect 8756 26498 8772 26532
rect 8840 26498 8856 26532
rect 8756 26451 8856 26498
rect 8914 26532 9014 26548
rect 8914 26498 8930 26532
rect 8998 26498 9014 26532
rect 8914 26451 9014 26498
rect 9072 26532 9172 26548
rect 9072 26498 9088 26532
rect 9156 26498 9172 26532
rect 9072 26451 9172 26498
rect 9230 26532 9330 26548
rect 9230 26498 9246 26532
rect 9314 26498 9330 26532
rect 9230 26451 9330 26498
rect 9388 26532 9488 26548
rect 9388 26498 9404 26532
rect 9472 26498 9488 26532
rect 9388 26451 9488 26498
rect 9546 26532 9646 26548
rect 9546 26498 9562 26532
rect 9630 26498 9646 26532
rect 9546 26451 9646 26498
rect 9704 26532 9804 26548
rect 9704 26498 9720 26532
rect 9788 26498 9804 26532
rect 9704 26451 9804 26498
rect 9862 26532 9962 26548
rect 9862 26498 9878 26532
rect 9946 26498 9962 26532
rect 9862 26451 9962 26498
rect 10020 26532 10120 26548
rect 10020 26498 10036 26532
rect 10104 26498 10120 26532
rect 10020 26451 10120 26498
rect 10178 26532 10278 26548
rect 10178 26498 10194 26532
rect 10262 26498 10278 26532
rect 10178 26451 10278 26498
rect 8756 26004 8856 26051
rect 8756 25970 8772 26004
rect 8840 25970 8856 26004
rect 8756 25954 8856 25970
rect 8914 26004 9014 26051
rect 8914 25970 8930 26004
rect 8998 25970 9014 26004
rect 8914 25954 9014 25970
rect 9072 26004 9172 26051
rect 9072 25970 9088 26004
rect 9156 25970 9172 26004
rect 9072 25954 9172 25970
rect 9230 26004 9330 26051
rect 9230 25970 9246 26004
rect 9314 25970 9330 26004
rect 9230 25954 9330 25970
rect 9388 26004 9488 26051
rect 9388 25970 9404 26004
rect 9472 25970 9488 26004
rect 9388 25954 9488 25970
rect 9546 26004 9646 26051
rect 9546 25970 9562 26004
rect 9630 25970 9646 26004
rect 9546 25954 9646 25970
rect 9704 26004 9804 26051
rect 9704 25970 9720 26004
rect 9788 25970 9804 26004
rect 9704 25954 9804 25970
rect 9862 26004 9962 26051
rect 9862 25970 9878 26004
rect 9946 25970 9962 26004
rect 9862 25954 9962 25970
rect 10020 26004 10120 26051
rect 10020 25970 10036 26004
rect 10104 25970 10120 26004
rect 10020 25954 10120 25970
rect 10178 26004 10278 26051
rect 10178 25970 10194 26004
rect 10262 25970 10278 26004
rect 10178 25954 10278 25970
rect 8756 25896 8856 25912
rect 8756 25862 8772 25896
rect 8840 25862 8856 25896
rect 8756 25815 8856 25862
rect 8914 25896 9014 25912
rect 8914 25862 8930 25896
rect 8998 25862 9014 25896
rect 8914 25815 9014 25862
rect 9072 25896 9172 25912
rect 9072 25862 9088 25896
rect 9156 25862 9172 25896
rect 9072 25815 9172 25862
rect 9230 25896 9330 25912
rect 9230 25862 9246 25896
rect 9314 25862 9330 25896
rect 9230 25815 9330 25862
rect 9388 25896 9488 25912
rect 9388 25862 9404 25896
rect 9472 25862 9488 25896
rect 9388 25815 9488 25862
rect 9546 25896 9646 25912
rect 9546 25862 9562 25896
rect 9630 25862 9646 25896
rect 9546 25815 9646 25862
rect 9704 25896 9804 25912
rect 9704 25862 9720 25896
rect 9788 25862 9804 25896
rect 9704 25815 9804 25862
rect 9862 25896 9962 25912
rect 9862 25862 9878 25896
rect 9946 25862 9962 25896
rect 9862 25815 9962 25862
rect 10020 25896 10120 25912
rect 10020 25862 10036 25896
rect 10104 25862 10120 25896
rect 10020 25815 10120 25862
rect 10178 25896 10278 25912
rect 10178 25862 10194 25896
rect 10262 25862 10278 25896
rect 10178 25815 10278 25862
rect 8756 25368 8856 25415
rect 8756 25334 8772 25368
rect 8840 25334 8856 25368
rect 8756 25318 8856 25334
rect 8914 25368 9014 25415
rect 8914 25334 8930 25368
rect 8998 25334 9014 25368
rect 8914 25318 9014 25334
rect 9072 25368 9172 25415
rect 9072 25334 9088 25368
rect 9156 25334 9172 25368
rect 9072 25318 9172 25334
rect 9230 25368 9330 25415
rect 9230 25334 9246 25368
rect 9314 25334 9330 25368
rect 9230 25318 9330 25334
rect 9388 25368 9488 25415
rect 9388 25334 9404 25368
rect 9472 25334 9488 25368
rect 9388 25318 9488 25334
rect 9546 25368 9646 25415
rect 9546 25334 9562 25368
rect 9630 25334 9646 25368
rect 9546 25318 9646 25334
rect 9704 25368 9804 25415
rect 9704 25334 9720 25368
rect 9788 25334 9804 25368
rect 9704 25318 9804 25334
rect 9862 25368 9962 25415
rect 9862 25334 9878 25368
rect 9946 25334 9962 25368
rect 9862 25318 9962 25334
rect 10020 25368 10120 25415
rect 10020 25334 10036 25368
rect 10104 25334 10120 25368
rect 10020 25318 10120 25334
rect 10178 25368 10278 25415
rect 10178 25334 10194 25368
rect 10262 25334 10278 25368
rect 10178 25318 10278 25334
rect 10936 27168 11036 27184
rect 10936 27134 10952 27168
rect 11020 27134 11036 27168
rect 10936 27087 11036 27134
rect 11094 27168 11194 27184
rect 11094 27134 11110 27168
rect 11178 27134 11194 27168
rect 11094 27087 11194 27134
rect 11252 27168 11352 27184
rect 11252 27134 11268 27168
rect 11336 27134 11352 27168
rect 11252 27087 11352 27134
rect 11410 27168 11510 27184
rect 11410 27134 11426 27168
rect 11494 27134 11510 27168
rect 11410 27087 11510 27134
rect 11568 27168 11668 27184
rect 11568 27134 11584 27168
rect 11652 27134 11668 27168
rect 11568 27087 11668 27134
rect 11726 27168 11826 27184
rect 11726 27134 11742 27168
rect 11810 27134 11826 27168
rect 11726 27087 11826 27134
rect 11884 27168 11984 27184
rect 11884 27134 11900 27168
rect 11968 27134 11984 27168
rect 11884 27087 11984 27134
rect 12042 27168 12142 27184
rect 12042 27134 12058 27168
rect 12126 27134 12142 27168
rect 12042 27087 12142 27134
rect 12200 27168 12300 27184
rect 12200 27134 12216 27168
rect 12284 27134 12300 27168
rect 12200 27087 12300 27134
rect 12358 27168 12458 27184
rect 12358 27134 12374 27168
rect 12442 27134 12458 27168
rect 12358 27087 12458 27134
rect 10936 26640 11036 26687
rect 10936 26606 10952 26640
rect 11020 26606 11036 26640
rect 10936 26590 11036 26606
rect 11094 26640 11194 26687
rect 11094 26606 11110 26640
rect 11178 26606 11194 26640
rect 11094 26590 11194 26606
rect 11252 26640 11352 26687
rect 11252 26606 11268 26640
rect 11336 26606 11352 26640
rect 11252 26590 11352 26606
rect 11410 26640 11510 26687
rect 11410 26606 11426 26640
rect 11494 26606 11510 26640
rect 11410 26590 11510 26606
rect 11568 26640 11668 26687
rect 11568 26606 11584 26640
rect 11652 26606 11668 26640
rect 11568 26590 11668 26606
rect 11726 26640 11826 26687
rect 11726 26606 11742 26640
rect 11810 26606 11826 26640
rect 11726 26590 11826 26606
rect 11884 26640 11984 26687
rect 11884 26606 11900 26640
rect 11968 26606 11984 26640
rect 11884 26590 11984 26606
rect 12042 26640 12142 26687
rect 12042 26606 12058 26640
rect 12126 26606 12142 26640
rect 12042 26590 12142 26606
rect 12200 26640 12300 26687
rect 12200 26606 12216 26640
rect 12284 26606 12300 26640
rect 12200 26590 12300 26606
rect 12358 26640 12458 26687
rect 12358 26606 12374 26640
rect 12442 26606 12458 26640
rect 12358 26590 12458 26606
rect 10936 26532 11036 26548
rect 10936 26498 10952 26532
rect 11020 26498 11036 26532
rect 10936 26451 11036 26498
rect 11094 26532 11194 26548
rect 11094 26498 11110 26532
rect 11178 26498 11194 26532
rect 11094 26451 11194 26498
rect 11252 26532 11352 26548
rect 11252 26498 11268 26532
rect 11336 26498 11352 26532
rect 11252 26451 11352 26498
rect 11410 26532 11510 26548
rect 11410 26498 11426 26532
rect 11494 26498 11510 26532
rect 11410 26451 11510 26498
rect 11568 26532 11668 26548
rect 11568 26498 11584 26532
rect 11652 26498 11668 26532
rect 11568 26451 11668 26498
rect 11726 26532 11826 26548
rect 11726 26498 11742 26532
rect 11810 26498 11826 26532
rect 11726 26451 11826 26498
rect 11884 26532 11984 26548
rect 11884 26498 11900 26532
rect 11968 26498 11984 26532
rect 11884 26451 11984 26498
rect 12042 26532 12142 26548
rect 12042 26498 12058 26532
rect 12126 26498 12142 26532
rect 12042 26451 12142 26498
rect 12200 26532 12300 26548
rect 12200 26498 12216 26532
rect 12284 26498 12300 26532
rect 12200 26451 12300 26498
rect 12358 26532 12458 26548
rect 12358 26498 12374 26532
rect 12442 26498 12458 26532
rect 12358 26451 12458 26498
rect 10936 26004 11036 26051
rect 10936 25970 10952 26004
rect 11020 25970 11036 26004
rect 10936 25954 11036 25970
rect 11094 26004 11194 26051
rect 11094 25970 11110 26004
rect 11178 25970 11194 26004
rect 11094 25954 11194 25970
rect 11252 26004 11352 26051
rect 11252 25970 11268 26004
rect 11336 25970 11352 26004
rect 11252 25954 11352 25970
rect 11410 26004 11510 26051
rect 11410 25970 11426 26004
rect 11494 25970 11510 26004
rect 11410 25954 11510 25970
rect 11568 26004 11668 26051
rect 11568 25970 11584 26004
rect 11652 25970 11668 26004
rect 11568 25954 11668 25970
rect 11726 26004 11826 26051
rect 11726 25970 11742 26004
rect 11810 25970 11826 26004
rect 11726 25954 11826 25970
rect 11884 26004 11984 26051
rect 11884 25970 11900 26004
rect 11968 25970 11984 26004
rect 11884 25954 11984 25970
rect 12042 26004 12142 26051
rect 12042 25970 12058 26004
rect 12126 25970 12142 26004
rect 12042 25954 12142 25970
rect 12200 26004 12300 26051
rect 12200 25970 12216 26004
rect 12284 25970 12300 26004
rect 12200 25954 12300 25970
rect 12358 26004 12458 26051
rect 12358 25970 12374 26004
rect 12442 25970 12458 26004
rect 12358 25954 12458 25970
rect 10936 25896 11036 25912
rect 10936 25862 10952 25896
rect 11020 25862 11036 25896
rect 10936 25815 11036 25862
rect 11094 25896 11194 25912
rect 11094 25862 11110 25896
rect 11178 25862 11194 25896
rect 11094 25815 11194 25862
rect 11252 25896 11352 25912
rect 11252 25862 11268 25896
rect 11336 25862 11352 25896
rect 11252 25815 11352 25862
rect 11410 25896 11510 25912
rect 11410 25862 11426 25896
rect 11494 25862 11510 25896
rect 11410 25815 11510 25862
rect 11568 25896 11668 25912
rect 11568 25862 11584 25896
rect 11652 25862 11668 25896
rect 11568 25815 11668 25862
rect 11726 25896 11826 25912
rect 11726 25862 11742 25896
rect 11810 25862 11826 25896
rect 11726 25815 11826 25862
rect 11884 25896 11984 25912
rect 11884 25862 11900 25896
rect 11968 25862 11984 25896
rect 11884 25815 11984 25862
rect 12042 25896 12142 25912
rect 12042 25862 12058 25896
rect 12126 25862 12142 25896
rect 12042 25815 12142 25862
rect 12200 25896 12300 25912
rect 12200 25862 12216 25896
rect 12284 25862 12300 25896
rect 12200 25815 12300 25862
rect 12358 25896 12458 25912
rect 12358 25862 12374 25896
rect 12442 25862 12458 25896
rect 12358 25815 12458 25862
rect 10936 25368 11036 25415
rect 10936 25334 10952 25368
rect 11020 25334 11036 25368
rect 10936 25318 11036 25334
rect 11094 25368 11194 25415
rect 11094 25334 11110 25368
rect 11178 25334 11194 25368
rect 11094 25318 11194 25334
rect 11252 25368 11352 25415
rect 11252 25334 11268 25368
rect 11336 25334 11352 25368
rect 11252 25318 11352 25334
rect 11410 25368 11510 25415
rect 11410 25334 11426 25368
rect 11494 25334 11510 25368
rect 11410 25318 11510 25334
rect 11568 25368 11668 25415
rect 11568 25334 11584 25368
rect 11652 25334 11668 25368
rect 11568 25318 11668 25334
rect 11726 25368 11826 25415
rect 11726 25334 11742 25368
rect 11810 25334 11826 25368
rect 11726 25318 11826 25334
rect 11884 25368 11984 25415
rect 11884 25334 11900 25368
rect 11968 25334 11984 25368
rect 11884 25318 11984 25334
rect 12042 25368 12142 25415
rect 12042 25334 12058 25368
rect 12126 25334 12142 25368
rect 12042 25318 12142 25334
rect 12200 25368 12300 25415
rect 12200 25334 12216 25368
rect 12284 25334 12300 25368
rect 12200 25318 12300 25334
rect 12358 25368 12458 25415
rect 12358 25334 12374 25368
rect 12442 25334 12458 25368
rect 12358 25318 12458 25334
rect 13116 27168 13216 27184
rect 13116 27134 13132 27168
rect 13200 27134 13216 27168
rect 13116 27087 13216 27134
rect 13274 27168 13374 27184
rect 13274 27134 13290 27168
rect 13358 27134 13374 27168
rect 13274 27087 13374 27134
rect 13432 27168 13532 27184
rect 13432 27134 13448 27168
rect 13516 27134 13532 27168
rect 13432 27087 13532 27134
rect 13590 27168 13690 27184
rect 13590 27134 13606 27168
rect 13674 27134 13690 27168
rect 13590 27087 13690 27134
rect 13748 27168 13848 27184
rect 13748 27134 13764 27168
rect 13832 27134 13848 27168
rect 13748 27087 13848 27134
rect 13906 27168 14006 27184
rect 13906 27134 13922 27168
rect 13990 27134 14006 27168
rect 13906 27087 14006 27134
rect 14064 27168 14164 27184
rect 14064 27134 14080 27168
rect 14148 27134 14164 27168
rect 14064 27087 14164 27134
rect 14222 27168 14322 27184
rect 14222 27134 14238 27168
rect 14306 27134 14322 27168
rect 14222 27087 14322 27134
rect 14380 27168 14480 27184
rect 14380 27134 14396 27168
rect 14464 27134 14480 27168
rect 14380 27087 14480 27134
rect 14538 27168 14638 27184
rect 14538 27134 14554 27168
rect 14622 27134 14638 27168
rect 14538 27087 14638 27134
rect 13116 26640 13216 26687
rect 13116 26606 13132 26640
rect 13200 26606 13216 26640
rect 13116 26590 13216 26606
rect 13274 26640 13374 26687
rect 13274 26606 13290 26640
rect 13358 26606 13374 26640
rect 13274 26590 13374 26606
rect 13432 26640 13532 26687
rect 13432 26606 13448 26640
rect 13516 26606 13532 26640
rect 13432 26590 13532 26606
rect 13590 26640 13690 26687
rect 13590 26606 13606 26640
rect 13674 26606 13690 26640
rect 13590 26590 13690 26606
rect 13748 26640 13848 26687
rect 13748 26606 13764 26640
rect 13832 26606 13848 26640
rect 13748 26590 13848 26606
rect 13906 26640 14006 26687
rect 13906 26606 13922 26640
rect 13990 26606 14006 26640
rect 13906 26590 14006 26606
rect 14064 26640 14164 26687
rect 14064 26606 14080 26640
rect 14148 26606 14164 26640
rect 14064 26590 14164 26606
rect 14222 26640 14322 26687
rect 14222 26606 14238 26640
rect 14306 26606 14322 26640
rect 14222 26590 14322 26606
rect 14380 26640 14480 26687
rect 14380 26606 14396 26640
rect 14464 26606 14480 26640
rect 14380 26590 14480 26606
rect 14538 26640 14638 26687
rect 14538 26606 14554 26640
rect 14622 26606 14638 26640
rect 14538 26590 14638 26606
rect 13116 26532 13216 26548
rect 13116 26498 13132 26532
rect 13200 26498 13216 26532
rect 13116 26451 13216 26498
rect 13274 26532 13374 26548
rect 13274 26498 13290 26532
rect 13358 26498 13374 26532
rect 13274 26451 13374 26498
rect 13432 26532 13532 26548
rect 13432 26498 13448 26532
rect 13516 26498 13532 26532
rect 13432 26451 13532 26498
rect 13590 26532 13690 26548
rect 13590 26498 13606 26532
rect 13674 26498 13690 26532
rect 13590 26451 13690 26498
rect 13748 26532 13848 26548
rect 13748 26498 13764 26532
rect 13832 26498 13848 26532
rect 13748 26451 13848 26498
rect 13906 26532 14006 26548
rect 13906 26498 13922 26532
rect 13990 26498 14006 26532
rect 13906 26451 14006 26498
rect 14064 26532 14164 26548
rect 14064 26498 14080 26532
rect 14148 26498 14164 26532
rect 14064 26451 14164 26498
rect 14222 26532 14322 26548
rect 14222 26498 14238 26532
rect 14306 26498 14322 26532
rect 14222 26451 14322 26498
rect 14380 26532 14480 26548
rect 14380 26498 14396 26532
rect 14464 26498 14480 26532
rect 14380 26451 14480 26498
rect 14538 26532 14638 26548
rect 14538 26498 14554 26532
rect 14622 26498 14638 26532
rect 14538 26451 14638 26498
rect 13116 26004 13216 26051
rect 13116 25970 13132 26004
rect 13200 25970 13216 26004
rect 13116 25954 13216 25970
rect 13274 26004 13374 26051
rect 13274 25970 13290 26004
rect 13358 25970 13374 26004
rect 13274 25954 13374 25970
rect 13432 26004 13532 26051
rect 13432 25970 13448 26004
rect 13516 25970 13532 26004
rect 13432 25954 13532 25970
rect 13590 26004 13690 26051
rect 13590 25970 13606 26004
rect 13674 25970 13690 26004
rect 13590 25954 13690 25970
rect 13748 26004 13848 26051
rect 13748 25970 13764 26004
rect 13832 25970 13848 26004
rect 13748 25954 13848 25970
rect 13906 26004 14006 26051
rect 13906 25970 13922 26004
rect 13990 25970 14006 26004
rect 13906 25954 14006 25970
rect 14064 26004 14164 26051
rect 14064 25970 14080 26004
rect 14148 25970 14164 26004
rect 14064 25954 14164 25970
rect 14222 26004 14322 26051
rect 14222 25970 14238 26004
rect 14306 25970 14322 26004
rect 14222 25954 14322 25970
rect 14380 26004 14480 26051
rect 14380 25970 14396 26004
rect 14464 25970 14480 26004
rect 14380 25954 14480 25970
rect 14538 26004 14638 26051
rect 14538 25970 14554 26004
rect 14622 25970 14638 26004
rect 14538 25954 14638 25970
rect 13116 25896 13216 25912
rect 13116 25862 13132 25896
rect 13200 25862 13216 25896
rect 13116 25815 13216 25862
rect 13274 25896 13374 25912
rect 13274 25862 13290 25896
rect 13358 25862 13374 25896
rect 13274 25815 13374 25862
rect 13432 25896 13532 25912
rect 13432 25862 13448 25896
rect 13516 25862 13532 25896
rect 13432 25815 13532 25862
rect 13590 25896 13690 25912
rect 13590 25862 13606 25896
rect 13674 25862 13690 25896
rect 13590 25815 13690 25862
rect 13748 25896 13848 25912
rect 13748 25862 13764 25896
rect 13832 25862 13848 25896
rect 13748 25815 13848 25862
rect 13906 25896 14006 25912
rect 13906 25862 13922 25896
rect 13990 25862 14006 25896
rect 13906 25815 14006 25862
rect 14064 25896 14164 25912
rect 14064 25862 14080 25896
rect 14148 25862 14164 25896
rect 14064 25815 14164 25862
rect 14222 25896 14322 25912
rect 14222 25862 14238 25896
rect 14306 25862 14322 25896
rect 14222 25815 14322 25862
rect 14380 25896 14480 25912
rect 14380 25862 14396 25896
rect 14464 25862 14480 25896
rect 14380 25815 14480 25862
rect 14538 25896 14638 25912
rect 14538 25862 14554 25896
rect 14622 25862 14638 25896
rect 14538 25815 14638 25862
rect 13116 25368 13216 25415
rect 13116 25334 13132 25368
rect 13200 25334 13216 25368
rect 13116 25318 13216 25334
rect 13274 25368 13374 25415
rect 13274 25334 13290 25368
rect 13358 25334 13374 25368
rect 13274 25318 13374 25334
rect 13432 25368 13532 25415
rect 13432 25334 13448 25368
rect 13516 25334 13532 25368
rect 13432 25318 13532 25334
rect 13590 25368 13690 25415
rect 13590 25334 13606 25368
rect 13674 25334 13690 25368
rect 13590 25318 13690 25334
rect 13748 25368 13848 25415
rect 13748 25334 13764 25368
rect 13832 25334 13848 25368
rect 13748 25318 13848 25334
rect 13906 25368 14006 25415
rect 13906 25334 13922 25368
rect 13990 25334 14006 25368
rect 13906 25318 14006 25334
rect 14064 25368 14164 25415
rect 14064 25334 14080 25368
rect 14148 25334 14164 25368
rect 14064 25318 14164 25334
rect 14222 25368 14322 25415
rect 14222 25334 14238 25368
rect 14306 25334 14322 25368
rect 14222 25318 14322 25334
rect 14380 25368 14480 25415
rect 14380 25334 14396 25368
rect 14464 25334 14480 25368
rect 14380 25318 14480 25334
rect 14538 25368 14638 25415
rect 14538 25334 14554 25368
rect 14622 25334 14638 25368
rect 14538 25318 14638 25334
rect 15316 27168 15416 27184
rect 15316 27134 15332 27168
rect 15400 27134 15416 27168
rect 15316 27087 15416 27134
rect 15474 27168 15574 27184
rect 15474 27134 15490 27168
rect 15558 27134 15574 27168
rect 15474 27087 15574 27134
rect 15632 27168 15732 27184
rect 15632 27134 15648 27168
rect 15716 27134 15732 27168
rect 15632 27087 15732 27134
rect 15790 27168 15890 27184
rect 15790 27134 15806 27168
rect 15874 27134 15890 27168
rect 15790 27087 15890 27134
rect 15948 27168 16048 27184
rect 15948 27134 15964 27168
rect 16032 27134 16048 27168
rect 15948 27087 16048 27134
rect 16106 27168 16206 27184
rect 16106 27134 16122 27168
rect 16190 27134 16206 27168
rect 16106 27087 16206 27134
rect 16264 27168 16364 27184
rect 16264 27134 16280 27168
rect 16348 27134 16364 27168
rect 16264 27087 16364 27134
rect 16422 27168 16522 27184
rect 16422 27134 16438 27168
rect 16506 27134 16522 27168
rect 16422 27087 16522 27134
rect 16580 27168 16680 27184
rect 16580 27134 16596 27168
rect 16664 27134 16680 27168
rect 16580 27087 16680 27134
rect 16738 27168 16838 27184
rect 16738 27134 16754 27168
rect 16822 27134 16838 27168
rect 16738 27087 16838 27134
rect 15316 26640 15416 26687
rect 15316 26606 15332 26640
rect 15400 26606 15416 26640
rect 15316 26590 15416 26606
rect 15474 26640 15574 26687
rect 15474 26606 15490 26640
rect 15558 26606 15574 26640
rect 15474 26590 15574 26606
rect 15632 26640 15732 26687
rect 15632 26606 15648 26640
rect 15716 26606 15732 26640
rect 15632 26590 15732 26606
rect 15790 26640 15890 26687
rect 15790 26606 15806 26640
rect 15874 26606 15890 26640
rect 15790 26590 15890 26606
rect 15948 26640 16048 26687
rect 15948 26606 15964 26640
rect 16032 26606 16048 26640
rect 15948 26590 16048 26606
rect 16106 26640 16206 26687
rect 16106 26606 16122 26640
rect 16190 26606 16206 26640
rect 16106 26590 16206 26606
rect 16264 26640 16364 26687
rect 16264 26606 16280 26640
rect 16348 26606 16364 26640
rect 16264 26590 16364 26606
rect 16422 26640 16522 26687
rect 16422 26606 16438 26640
rect 16506 26606 16522 26640
rect 16422 26590 16522 26606
rect 16580 26640 16680 26687
rect 16580 26606 16596 26640
rect 16664 26606 16680 26640
rect 16580 26590 16680 26606
rect 16738 26640 16838 26687
rect 16738 26606 16754 26640
rect 16822 26606 16838 26640
rect 16738 26590 16838 26606
rect 15316 26532 15416 26548
rect 15316 26498 15332 26532
rect 15400 26498 15416 26532
rect 15316 26451 15416 26498
rect 15474 26532 15574 26548
rect 15474 26498 15490 26532
rect 15558 26498 15574 26532
rect 15474 26451 15574 26498
rect 15632 26532 15732 26548
rect 15632 26498 15648 26532
rect 15716 26498 15732 26532
rect 15632 26451 15732 26498
rect 15790 26532 15890 26548
rect 15790 26498 15806 26532
rect 15874 26498 15890 26532
rect 15790 26451 15890 26498
rect 15948 26532 16048 26548
rect 15948 26498 15964 26532
rect 16032 26498 16048 26532
rect 15948 26451 16048 26498
rect 16106 26532 16206 26548
rect 16106 26498 16122 26532
rect 16190 26498 16206 26532
rect 16106 26451 16206 26498
rect 16264 26532 16364 26548
rect 16264 26498 16280 26532
rect 16348 26498 16364 26532
rect 16264 26451 16364 26498
rect 16422 26532 16522 26548
rect 16422 26498 16438 26532
rect 16506 26498 16522 26532
rect 16422 26451 16522 26498
rect 16580 26532 16680 26548
rect 16580 26498 16596 26532
rect 16664 26498 16680 26532
rect 16580 26451 16680 26498
rect 16738 26532 16838 26548
rect 16738 26498 16754 26532
rect 16822 26498 16838 26532
rect 16738 26451 16838 26498
rect 15316 26004 15416 26051
rect 15316 25970 15332 26004
rect 15400 25970 15416 26004
rect 15316 25954 15416 25970
rect 15474 26004 15574 26051
rect 15474 25970 15490 26004
rect 15558 25970 15574 26004
rect 15474 25954 15574 25970
rect 15632 26004 15732 26051
rect 15632 25970 15648 26004
rect 15716 25970 15732 26004
rect 15632 25954 15732 25970
rect 15790 26004 15890 26051
rect 15790 25970 15806 26004
rect 15874 25970 15890 26004
rect 15790 25954 15890 25970
rect 15948 26004 16048 26051
rect 15948 25970 15964 26004
rect 16032 25970 16048 26004
rect 15948 25954 16048 25970
rect 16106 26004 16206 26051
rect 16106 25970 16122 26004
rect 16190 25970 16206 26004
rect 16106 25954 16206 25970
rect 16264 26004 16364 26051
rect 16264 25970 16280 26004
rect 16348 25970 16364 26004
rect 16264 25954 16364 25970
rect 16422 26004 16522 26051
rect 16422 25970 16438 26004
rect 16506 25970 16522 26004
rect 16422 25954 16522 25970
rect 16580 26004 16680 26051
rect 16580 25970 16596 26004
rect 16664 25970 16680 26004
rect 16580 25954 16680 25970
rect 16738 26004 16838 26051
rect 16738 25970 16754 26004
rect 16822 25970 16838 26004
rect 16738 25954 16838 25970
rect 15316 25896 15416 25912
rect 15316 25862 15332 25896
rect 15400 25862 15416 25896
rect 15316 25815 15416 25862
rect 15474 25896 15574 25912
rect 15474 25862 15490 25896
rect 15558 25862 15574 25896
rect 15474 25815 15574 25862
rect 15632 25896 15732 25912
rect 15632 25862 15648 25896
rect 15716 25862 15732 25896
rect 15632 25815 15732 25862
rect 15790 25896 15890 25912
rect 15790 25862 15806 25896
rect 15874 25862 15890 25896
rect 15790 25815 15890 25862
rect 15948 25896 16048 25912
rect 15948 25862 15964 25896
rect 16032 25862 16048 25896
rect 15948 25815 16048 25862
rect 16106 25896 16206 25912
rect 16106 25862 16122 25896
rect 16190 25862 16206 25896
rect 16106 25815 16206 25862
rect 16264 25896 16364 25912
rect 16264 25862 16280 25896
rect 16348 25862 16364 25896
rect 16264 25815 16364 25862
rect 16422 25896 16522 25912
rect 16422 25862 16438 25896
rect 16506 25862 16522 25896
rect 16422 25815 16522 25862
rect 16580 25896 16680 25912
rect 16580 25862 16596 25896
rect 16664 25862 16680 25896
rect 16580 25815 16680 25862
rect 16738 25896 16838 25912
rect 16738 25862 16754 25896
rect 16822 25862 16838 25896
rect 16738 25815 16838 25862
rect 15316 25368 15416 25415
rect 15316 25334 15332 25368
rect 15400 25334 15416 25368
rect 15316 25318 15416 25334
rect 15474 25368 15574 25415
rect 15474 25334 15490 25368
rect 15558 25334 15574 25368
rect 15474 25318 15574 25334
rect 15632 25368 15732 25415
rect 15632 25334 15648 25368
rect 15716 25334 15732 25368
rect 15632 25318 15732 25334
rect 15790 25368 15890 25415
rect 15790 25334 15806 25368
rect 15874 25334 15890 25368
rect 15790 25318 15890 25334
rect 15948 25368 16048 25415
rect 15948 25334 15964 25368
rect 16032 25334 16048 25368
rect 15948 25318 16048 25334
rect 16106 25368 16206 25415
rect 16106 25334 16122 25368
rect 16190 25334 16206 25368
rect 16106 25318 16206 25334
rect 16264 25368 16364 25415
rect 16264 25334 16280 25368
rect 16348 25334 16364 25368
rect 16264 25318 16364 25334
rect 16422 25368 16522 25415
rect 16422 25334 16438 25368
rect 16506 25334 16522 25368
rect 16422 25318 16522 25334
rect 16580 25368 16680 25415
rect 16580 25334 16596 25368
rect 16664 25334 16680 25368
rect 16580 25318 16680 25334
rect 16738 25368 16838 25415
rect 16738 25334 16754 25368
rect 16822 25334 16838 25368
rect 16738 25318 16838 25334
rect 6522 25072 6588 25088
rect 6522 25038 6538 25072
rect 6572 25038 6588 25072
rect 6522 25022 6588 25038
rect 6714 25072 6780 25088
rect 6714 25038 6730 25072
rect 6764 25038 6780 25072
rect 6714 25022 6780 25038
rect 6906 25072 6972 25088
rect 6906 25038 6922 25072
rect 6956 25038 6972 25072
rect 6906 25022 6972 25038
rect 7098 25072 7164 25088
rect 7098 25038 7114 25072
rect 7148 25038 7164 25072
rect 7098 25022 7164 25038
rect 7290 25072 7356 25088
rect 7290 25038 7306 25072
rect 7340 25038 7356 25072
rect 7290 25022 7356 25038
rect 7482 25072 7548 25088
rect 7482 25038 7498 25072
rect 7532 25038 7548 25072
rect 7482 25022 7548 25038
rect 7674 25072 7740 25088
rect 7674 25038 7690 25072
rect 7724 25038 7740 25072
rect 7674 25022 7740 25038
rect 7866 25072 7932 25088
rect 7866 25038 7882 25072
rect 7916 25038 7932 25072
rect 7866 25022 7932 25038
rect 6540 24991 6570 25022
rect 6636 24991 6666 25017
rect 6732 24991 6762 25022
rect 6828 24991 6858 25017
rect 6924 24991 6954 25022
rect 7020 24991 7050 25017
rect 7116 24991 7146 25022
rect 7212 24991 7242 25017
rect 7308 24991 7338 25022
rect 7404 24991 7434 25017
rect 7500 24991 7530 25022
rect 7596 24991 7626 25017
rect 7692 24991 7722 25022
rect 7788 24991 7818 25017
rect 7884 24991 7914 25022
rect 6540 24565 6570 24591
rect 6636 24560 6666 24591
rect 6732 24565 6762 24591
rect 6828 24560 6858 24591
rect 6924 24565 6954 24591
rect 7020 24560 7050 24591
rect 7116 24565 7146 24591
rect 7212 24560 7242 24591
rect 7308 24565 7338 24591
rect 7404 24560 7434 24591
rect 7500 24565 7530 24591
rect 7596 24560 7626 24591
rect 7692 24565 7722 24591
rect 7788 24560 7818 24591
rect 7884 24565 7914 24591
rect 6618 24544 6684 24560
rect 6618 24510 6634 24544
rect 6668 24510 6684 24544
rect 6618 24494 6684 24510
rect 6810 24544 6876 24560
rect 6810 24510 6826 24544
rect 6860 24510 6876 24544
rect 6810 24494 6876 24510
rect 7002 24544 7068 24560
rect 7002 24510 7018 24544
rect 7052 24510 7068 24544
rect 7002 24494 7068 24510
rect 7194 24544 7260 24560
rect 7194 24510 7210 24544
rect 7244 24510 7260 24544
rect 7194 24494 7260 24510
rect 7386 24544 7452 24560
rect 7386 24510 7402 24544
rect 7436 24510 7452 24544
rect 7386 24494 7452 24510
rect 7578 24544 7644 24560
rect 7578 24510 7594 24544
rect 7628 24510 7644 24544
rect 7578 24494 7644 24510
rect 7770 24544 7836 24560
rect 7770 24510 7786 24544
rect 7820 24510 7836 24544
rect 7770 24494 7836 24510
rect 6618 24436 6684 24452
rect 6618 24402 6634 24436
rect 6668 24402 6684 24436
rect 6618 24386 6684 24402
rect 6810 24436 6876 24452
rect 6810 24402 6826 24436
rect 6860 24402 6876 24436
rect 6810 24386 6876 24402
rect 7002 24436 7068 24452
rect 7002 24402 7018 24436
rect 7052 24402 7068 24436
rect 7002 24386 7068 24402
rect 7194 24436 7260 24452
rect 7194 24402 7210 24436
rect 7244 24402 7260 24436
rect 7194 24386 7260 24402
rect 7386 24436 7452 24452
rect 7386 24402 7402 24436
rect 7436 24402 7452 24436
rect 7386 24386 7452 24402
rect 7578 24436 7644 24452
rect 7578 24402 7594 24436
rect 7628 24402 7644 24436
rect 7578 24386 7644 24402
rect 7770 24436 7836 24452
rect 7770 24402 7786 24436
rect 7820 24402 7836 24436
rect 7770 24386 7836 24402
rect 6540 24355 6570 24381
rect 6636 24355 6666 24386
rect 6732 24355 6762 24381
rect 6828 24355 6858 24386
rect 6924 24355 6954 24381
rect 7020 24355 7050 24386
rect 7116 24355 7146 24381
rect 7212 24355 7242 24386
rect 7308 24355 7338 24381
rect 7404 24355 7434 24386
rect 7500 24355 7530 24381
rect 7596 24355 7626 24386
rect 7692 24355 7722 24381
rect 7788 24355 7818 24386
rect 7884 24355 7914 24381
rect 6540 23924 6570 23955
rect 6636 23929 6666 23955
rect 6732 23924 6762 23955
rect 6828 23929 6858 23955
rect 6924 23924 6954 23955
rect 7020 23929 7050 23955
rect 7116 23924 7146 23955
rect 7212 23929 7242 23955
rect 7308 23924 7338 23955
rect 7404 23929 7434 23955
rect 7500 23924 7530 23955
rect 7596 23929 7626 23955
rect 7692 23924 7722 23955
rect 7788 23929 7818 23955
rect 7884 23924 7914 23955
rect 6522 23908 6588 23924
rect 6522 23874 6538 23908
rect 6572 23874 6588 23908
rect 6522 23858 6588 23874
rect 6714 23908 6780 23924
rect 6714 23874 6730 23908
rect 6764 23874 6780 23908
rect 6714 23858 6780 23874
rect 6906 23908 6972 23924
rect 6906 23874 6922 23908
rect 6956 23874 6972 23908
rect 6906 23858 6972 23874
rect 7098 23908 7164 23924
rect 7098 23874 7114 23908
rect 7148 23874 7164 23908
rect 7098 23858 7164 23874
rect 7290 23908 7356 23924
rect 7290 23874 7306 23908
rect 7340 23874 7356 23908
rect 7290 23858 7356 23874
rect 7482 23908 7548 23924
rect 7482 23874 7498 23908
rect 7532 23874 7548 23908
rect 7482 23858 7548 23874
rect 7674 23908 7740 23924
rect 7674 23874 7690 23908
rect 7724 23874 7740 23908
rect 7674 23858 7740 23874
rect 7866 23908 7932 23924
rect 7866 23874 7882 23908
rect 7916 23874 7932 23908
rect 7866 23858 7932 23874
rect 8742 25072 8808 25088
rect 8742 25038 8758 25072
rect 8792 25038 8808 25072
rect 8742 25022 8808 25038
rect 8934 25072 9000 25088
rect 8934 25038 8950 25072
rect 8984 25038 9000 25072
rect 8934 25022 9000 25038
rect 9126 25072 9192 25088
rect 9126 25038 9142 25072
rect 9176 25038 9192 25072
rect 9126 25022 9192 25038
rect 9318 25072 9384 25088
rect 9318 25038 9334 25072
rect 9368 25038 9384 25072
rect 9318 25022 9384 25038
rect 9510 25072 9576 25088
rect 9510 25038 9526 25072
rect 9560 25038 9576 25072
rect 9510 25022 9576 25038
rect 9702 25072 9768 25088
rect 9702 25038 9718 25072
rect 9752 25038 9768 25072
rect 9702 25022 9768 25038
rect 9894 25072 9960 25088
rect 9894 25038 9910 25072
rect 9944 25038 9960 25072
rect 9894 25022 9960 25038
rect 10086 25072 10152 25088
rect 10086 25038 10102 25072
rect 10136 25038 10152 25072
rect 10086 25022 10152 25038
rect 8760 24991 8790 25022
rect 8856 24991 8886 25017
rect 8952 24991 8982 25022
rect 9048 24991 9078 25017
rect 9144 24991 9174 25022
rect 9240 24991 9270 25017
rect 9336 24991 9366 25022
rect 9432 24991 9462 25017
rect 9528 24991 9558 25022
rect 9624 24991 9654 25017
rect 9720 24991 9750 25022
rect 9816 24991 9846 25017
rect 9912 24991 9942 25022
rect 10008 24991 10038 25017
rect 10104 24991 10134 25022
rect 8760 24565 8790 24591
rect 8856 24560 8886 24591
rect 8952 24565 8982 24591
rect 9048 24560 9078 24591
rect 9144 24565 9174 24591
rect 9240 24560 9270 24591
rect 9336 24565 9366 24591
rect 9432 24560 9462 24591
rect 9528 24565 9558 24591
rect 9624 24560 9654 24591
rect 9720 24565 9750 24591
rect 9816 24560 9846 24591
rect 9912 24565 9942 24591
rect 10008 24560 10038 24591
rect 10104 24565 10134 24591
rect 8838 24544 8904 24560
rect 8838 24510 8854 24544
rect 8888 24510 8904 24544
rect 8838 24494 8904 24510
rect 9030 24544 9096 24560
rect 9030 24510 9046 24544
rect 9080 24510 9096 24544
rect 9030 24494 9096 24510
rect 9222 24544 9288 24560
rect 9222 24510 9238 24544
rect 9272 24510 9288 24544
rect 9222 24494 9288 24510
rect 9414 24544 9480 24560
rect 9414 24510 9430 24544
rect 9464 24510 9480 24544
rect 9414 24494 9480 24510
rect 9606 24544 9672 24560
rect 9606 24510 9622 24544
rect 9656 24510 9672 24544
rect 9606 24494 9672 24510
rect 9798 24544 9864 24560
rect 9798 24510 9814 24544
rect 9848 24510 9864 24544
rect 9798 24494 9864 24510
rect 9990 24544 10056 24560
rect 9990 24510 10006 24544
rect 10040 24510 10056 24544
rect 9990 24494 10056 24510
rect 8838 24436 8904 24452
rect 8838 24402 8854 24436
rect 8888 24402 8904 24436
rect 8838 24386 8904 24402
rect 9030 24436 9096 24452
rect 9030 24402 9046 24436
rect 9080 24402 9096 24436
rect 9030 24386 9096 24402
rect 9222 24436 9288 24452
rect 9222 24402 9238 24436
rect 9272 24402 9288 24436
rect 9222 24386 9288 24402
rect 9414 24436 9480 24452
rect 9414 24402 9430 24436
rect 9464 24402 9480 24436
rect 9414 24386 9480 24402
rect 9606 24436 9672 24452
rect 9606 24402 9622 24436
rect 9656 24402 9672 24436
rect 9606 24386 9672 24402
rect 9798 24436 9864 24452
rect 9798 24402 9814 24436
rect 9848 24402 9864 24436
rect 9798 24386 9864 24402
rect 9990 24436 10056 24452
rect 9990 24402 10006 24436
rect 10040 24402 10056 24436
rect 9990 24386 10056 24402
rect 8760 24355 8790 24381
rect 8856 24355 8886 24386
rect 8952 24355 8982 24381
rect 9048 24355 9078 24386
rect 9144 24355 9174 24381
rect 9240 24355 9270 24386
rect 9336 24355 9366 24381
rect 9432 24355 9462 24386
rect 9528 24355 9558 24381
rect 9624 24355 9654 24386
rect 9720 24355 9750 24381
rect 9816 24355 9846 24386
rect 9912 24355 9942 24381
rect 10008 24355 10038 24386
rect 10104 24355 10134 24381
rect 8760 23924 8790 23955
rect 8856 23929 8886 23955
rect 8952 23924 8982 23955
rect 9048 23929 9078 23955
rect 9144 23924 9174 23955
rect 9240 23929 9270 23955
rect 9336 23924 9366 23955
rect 9432 23929 9462 23955
rect 9528 23924 9558 23955
rect 9624 23929 9654 23955
rect 9720 23924 9750 23955
rect 9816 23929 9846 23955
rect 9912 23924 9942 23955
rect 10008 23929 10038 23955
rect 10104 23924 10134 23955
rect 8742 23908 8808 23924
rect 8742 23874 8758 23908
rect 8792 23874 8808 23908
rect 8742 23858 8808 23874
rect 8934 23908 9000 23924
rect 8934 23874 8950 23908
rect 8984 23874 9000 23908
rect 8934 23858 9000 23874
rect 9126 23908 9192 23924
rect 9126 23874 9142 23908
rect 9176 23874 9192 23908
rect 9126 23858 9192 23874
rect 9318 23908 9384 23924
rect 9318 23874 9334 23908
rect 9368 23874 9384 23908
rect 9318 23858 9384 23874
rect 9510 23908 9576 23924
rect 9510 23874 9526 23908
rect 9560 23874 9576 23908
rect 9510 23858 9576 23874
rect 9702 23908 9768 23924
rect 9702 23874 9718 23908
rect 9752 23874 9768 23908
rect 9702 23858 9768 23874
rect 9894 23908 9960 23924
rect 9894 23874 9910 23908
rect 9944 23874 9960 23908
rect 9894 23858 9960 23874
rect 10086 23908 10152 23924
rect 10086 23874 10102 23908
rect 10136 23874 10152 23908
rect 10086 23858 10152 23874
rect 10922 25072 10988 25088
rect 10922 25038 10938 25072
rect 10972 25038 10988 25072
rect 10922 25022 10988 25038
rect 11114 25072 11180 25088
rect 11114 25038 11130 25072
rect 11164 25038 11180 25072
rect 11114 25022 11180 25038
rect 11306 25072 11372 25088
rect 11306 25038 11322 25072
rect 11356 25038 11372 25072
rect 11306 25022 11372 25038
rect 11498 25072 11564 25088
rect 11498 25038 11514 25072
rect 11548 25038 11564 25072
rect 11498 25022 11564 25038
rect 11690 25072 11756 25088
rect 11690 25038 11706 25072
rect 11740 25038 11756 25072
rect 11690 25022 11756 25038
rect 11882 25072 11948 25088
rect 11882 25038 11898 25072
rect 11932 25038 11948 25072
rect 11882 25022 11948 25038
rect 12074 25072 12140 25088
rect 12074 25038 12090 25072
rect 12124 25038 12140 25072
rect 12074 25022 12140 25038
rect 12266 25072 12332 25088
rect 12266 25038 12282 25072
rect 12316 25038 12332 25072
rect 12266 25022 12332 25038
rect 10940 24991 10970 25022
rect 11036 24991 11066 25017
rect 11132 24991 11162 25022
rect 11228 24991 11258 25017
rect 11324 24991 11354 25022
rect 11420 24991 11450 25017
rect 11516 24991 11546 25022
rect 11612 24991 11642 25017
rect 11708 24991 11738 25022
rect 11804 24991 11834 25017
rect 11900 24991 11930 25022
rect 11996 24991 12026 25017
rect 12092 24991 12122 25022
rect 12188 24991 12218 25017
rect 12284 24991 12314 25022
rect 10940 24565 10970 24591
rect 11036 24560 11066 24591
rect 11132 24565 11162 24591
rect 11228 24560 11258 24591
rect 11324 24565 11354 24591
rect 11420 24560 11450 24591
rect 11516 24565 11546 24591
rect 11612 24560 11642 24591
rect 11708 24565 11738 24591
rect 11804 24560 11834 24591
rect 11900 24565 11930 24591
rect 11996 24560 12026 24591
rect 12092 24565 12122 24591
rect 12188 24560 12218 24591
rect 12284 24565 12314 24591
rect 11018 24544 11084 24560
rect 11018 24510 11034 24544
rect 11068 24510 11084 24544
rect 11018 24494 11084 24510
rect 11210 24544 11276 24560
rect 11210 24510 11226 24544
rect 11260 24510 11276 24544
rect 11210 24494 11276 24510
rect 11402 24544 11468 24560
rect 11402 24510 11418 24544
rect 11452 24510 11468 24544
rect 11402 24494 11468 24510
rect 11594 24544 11660 24560
rect 11594 24510 11610 24544
rect 11644 24510 11660 24544
rect 11594 24494 11660 24510
rect 11786 24544 11852 24560
rect 11786 24510 11802 24544
rect 11836 24510 11852 24544
rect 11786 24494 11852 24510
rect 11978 24544 12044 24560
rect 11978 24510 11994 24544
rect 12028 24510 12044 24544
rect 11978 24494 12044 24510
rect 12170 24544 12236 24560
rect 12170 24510 12186 24544
rect 12220 24510 12236 24544
rect 12170 24494 12236 24510
rect 11018 24436 11084 24452
rect 11018 24402 11034 24436
rect 11068 24402 11084 24436
rect 11018 24386 11084 24402
rect 11210 24436 11276 24452
rect 11210 24402 11226 24436
rect 11260 24402 11276 24436
rect 11210 24386 11276 24402
rect 11402 24436 11468 24452
rect 11402 24402 11418 24436
rect 11452 24402 11468 24436
rect 11402 24386 11468 24402
rect 11594 24436 11660 24452
rect 11594 24402 11610 24436
rect 11644 24402 11660 24436
rect 11594 24386 11660 24402
rect 11786 24436 11852 24452
rect 11786 24402 11802 24436
rect 11836 24402 11852 24436
rect 11786 24386 11852 24402
rect 11978 24436 12044 24452
rect 11978 24402 11994 24436
rect 12028 24402 12044 24436
rect 11978 24386 12044 24402
rect 12170 24436 12236 24452
rect 12170 24402 12186 24436
rect 12220 24402 12236 24436
rect 12170 24386 12236 24402
rect 10940 24355 10970 24381
rect 11036 24355 11066 24386
rect 11132 24355 11162 24381
rect 11228 24355 11258 24386
rect 11324 24355 11354 24381
rect 11420 24355 11450 24386
rect 11516 24355 11546 24381
rect 11612 24355 11642 24386
rect 11708 24355 11738 24381
rect 11804 24355 11834 24386
rect 11900 24355 11930 24381
rect 11996 24355 12026 24386
rect 12092 24355 12122 24381
rect 12188 24355 12218 24386
rect 12284 24355 12314 24381
rect 10940 23924 10970 23955
rect 11036 23929 11066 23955
rect 11132 23924 11162 23955
rect 11228 23929 11258 23955
rect 11324 23924 11354 23955
rect 11420 23929 11450 23955
rect 11516 23924 11546 23955
rect 11612 23929 11642 23955
rect 11708 23924 11738 23955
rect 11804 23929 11834 23955
rect 11900 23924 11930 23955
rect 11996 23929 12026 23955
rect 12092 23924 12122 23955
rect 12188 23929 12218 23955
rect 12284 23924 12314 23955
rect 10922 23908 10988 23924
rect 10922 23874 10938 23908
rect 10972 23874 10988 23908
rect 10922 23858 10988 23874
rect 11114 23908 11180 23924
rect 11114 23874 11130 23908
rect 11164 23874 11180 23908
rect 11114 23858 11180 23874
rect 11306 23908 11372 23924
rect 11306 23874 11322 23908
rect 11356 23874 11372 23908
rect 11306 23858 11372 23874
rect 11498 23908 11564 23924
rect 11498 23874 11514 23908
rect 11548 23874 11564 23908
rect 11498 23858 11564 23874
rect 11690 23908 11756 23924
rect 11690 23874 11706 23908
rect 11740 23874 11756 23908
rect 11690 23858 11756 23874
rect 11882 23908 11948 23924
rect 11882 23874 11898 23908
rect 11932 23874 11948 23908
rect 11882 23858 11948 23874
rect 12074 23908 12140 23924
rect 12074 23874 12090 23908
rect 12124 23874 12140 23908
rect 12074 23858 12140 23874
rect 12266 23908 12332 23924
rect 12266 23874 12282 23908
rect 12316 23874 12332 23908
rect 12266 23858 12332 23874
rect 13102 25072 13168 25088
rect 13102 25038 13118 25072
rect 13152 25038 13168 25072
rect 13102 25022 13168 25038
rect 13294 25072 13360 25088
rect 13294 25038 13310 25072
rect 13344 25038 13360 25072
rect 13294 25022 13360 25038
rect 13486 25072 13552 25088
rect 13486 25038 13502 25072
rect 13536 25038 13552 25072
rect 13486 25022 13552 25038
rect 13678 25072 13744 25088
rect 13678 25038 13694 25072
rect 13728 25038 13744 25072
rect 13678 25022 13744 25038
rect 13870 25072 13936 25088
rect 13870 25038 13886 25072
rect 13920 25038 13936 25072
rect 13870 25022 13936 25038
rect 14062 25072 14128 25088
rect 14062 25038 14078 25072
rect 14112 25038 14128 25072
rect 14062 25022 14128 25038
rect 14254 25072 14320 25088
rect 14254 25038 14270 25072
rect 14304 25038 14320 25072
rect 14254 25022 14320 25038
rect 14446 25072 14512 25088
rect 14446 25038 14462 25072
rect 14496 25038 14512 25072
rect 14446 25022 14512 25038
rect 13120 24991 13150 25022
rect 13216 24991 13246 25017
rect 13312 24991 13342 25022
rect 13408 24991 13438 25017
rect 13504 24991 13534 25022
rect 13600 24991 13630 25017
rect 13696 24991 13726 25022
rect 13792 24991 13822 25017
rect 13888 24991 13918 25022
rect 13984 24991 14014 25017
rect 14080 24991 14110 25022
rect 14176 24991 14206 25017
rect 14272 24991 14302 25022
rect 14368 24991 14398 25017
rect 14464 24991 14494 25022
rect 13120 24565 13150 24591
rect 13216 24560 13246 24591
rect 13312 24565 13342 24591
rect 13408 24560 13438 24591
rect 13504 24565 13534 24591
rect 13600 24560 13630 24591
rect 13696 24565 13726 24591
rect 13792 24560 13822 24591
rect 13888 24565 13918 24591
rect 13984 24560 14014 24591
rect 14080 24565 14110 24591
rect 14176 24560 14206 24591
rect 14272 24565 14302 24591
rect 14368 24560 14398 24591
rect 14464 24565 14494 24591
rect 13198 24544 13264 24560
rect 13198 24510 13214 24544
rect 13248 24510 13264 24544
rect 13198 24494 13264 24510
rect 13390 24544 13456 24560
rect 13390 24510 13406 24544
rect 13440 24510 13456 24544
rect 13390 24494 13456 24510
rect 13582 24544 13648 24560
rect 13582 24510 13598 24544
rect 13632 24510 13648 24544
rect 13582 24494 13648 24510
rect 13774 24544 13840 24560
rect 13774 24510 13790 24544
rect 13824 24510 13840 24544
rect 13774 24494 13840 24510
rect 13966 24544 14032 24560
rect 13966 24510 13982 24544
rect 14016 24510 14032 24544
rect 13966 24494 14032 24510
rect 14158 24544 14224 24560
rect 14158 24510 14174 24544
rect 14208 24510 14224 24544
rect 14158 24494 14224 24510
rect 14350 24544 14416 24560
rect 14350 24510 14366 24544
rect 14400 24510 14416 24544
rect 14350 24494 14416 24510
rect 13198 24436 13264 24452
rect 13198 24402 13214 24436
rect 13248 24402 13264 24436
rect 13198 24386 13264 24402
rect 13390 24436 13456 24452
rect 13390 24402 13406 24436
rect 13440 24402 13456 24436
rect 13390 24386 13456 24402
rect 13582 24436 13648 24452
rect 13582 24402 13598 24436
rect 13632 24402 13648 24436
rect 13582 24386 13648 24402
rect 13774 24436 13840 24452
rect 13774 24402 13790 24436
rect 13824 24402 13840 24436
rect 13774 24386 13840 24402
rect 13966 24436 14032 24452
rect 13966 24402 13982 24436
rect 14016 24402 14032 24436
rect 13966 24386 14032 24402
rect 14158 24436 14224 24452
rect 14158 24402 14174 24436
rect 14208 24402 14224 24436
rect 14158 24386 14224 24402
rect 14350 24436 14416 24452
rect 14350 24402 14366 24436
rect 14400 24402 14416 24436
rect 14350 24386 14416 24402
rect 13120 24355 13150 24381
rect 13216 24355 13246 24386
rect 13312 24355 13342 24381
rect 13408 24355 13438 24386
rect 13504 24355 13534 24381
rect 13600 24355 13630 24386
rect 13696 24355 13726 24381
rect 13792 24355 13822 24386
rect 13888 24355 13918 24381
rect 13984 24355 14014 24386
rect 14080 24355 14110 24381
rect 14176 24355 14206 24386
rect 14272 24355 14302 24381
rect 14368 24355 14398 24386
rect 14464 24355 14494 24381
rect 13120 23924 13150 23955
rect 13216 23929 13246 23955
rect 13312 23924 13342 23955
rect 13408 23929 13438 23955
rect 13504 23924 13534 23955
rect 13600 23929 13630 23955
rect 13696 23924 13726 23955
rect 13792 23929 13822 23955
rect 13888 23924 13918 23955
rect 13984 23929 14014 23955
rect 14080 23924 14110 23955
rect 14176 23929 14206 23955
rect 14272 23924 14302 23955
rect 14368 23929 14398 23955
rect 14464 23924 14494 23955
rect 13102 23908 13168 23924
rect 13102 23874 13118 23908
rect 13152 23874 13168 23908
rect 13102 23858 13168 23874
rect 13294 23908 13360 23924
rect 13294 23874 13310 23908
rect 13344 23874 13360 23908
rect 13294 23858 13360 23874
rect 13486 23908 13552 23924
rect 13486 23874 13502 23908
rect 13536 23874 13552 23908
rect 13486 23858 13552 23874
rect 13678 23908 13744 23924
rect 13678 23874 13694 23908
rect 13728 23874 13744 23908
rect 13678 23858 13744 23874
rect 13870 23908 13936 23924
rect 13870 23874 13886 23908
rect 13920 23874 13936 23908
rect 13870 23858 13936 23874
rect 14062 23908 14128 23924
rect 14062 23874 14078 23908
rect 14112 23874 14128 23908
rect 14062 23858 14128 23874
rect 14254 23908 14320 23924
rect 14254 23874 14270 23908
rect 14304 23874 14320 23908
rect 14254 23858 14320 23874
rect 14446 23908 14512 23924
rect 14446 23874 14462 23908
rect 14496 23874 14512 23908
rect 14446 23858 14512 23874
rect 15302 25072 15368 25088
rect 15302 25038 15318 25072
rect 15352 25038 15368 25072
rect 15302 25022 15368 25038
rect 15494 25072 15560 25088
rect 15494 25038 15510 25072
rect 15544 25038 15560 25072
rect 15494 25022 15560 25038
rect 15686 25072 15752 25088
rect 15686 25038 15702 25072
rect 15736 25038 15752 25072
rect 15686 25022 15752 25038
rect 15878 25072 15944 25088
rect 15878 25038 15894 25072
rect 15928 25038 15944 25072
rect 15878 25022 15944 25038
rect 16070 25072 16136 25088
rect 16070 25038 16086 25072
rect 16120 25038 16136 25072
rect 16070 25022 16136 25038
rect 16262 25072 16328 25088
rect 16262 25038 16278 25072
rect 16312 25038 16328 25072
rect 16262 25022 16328 25038
rect 16454 25072 16520 25088
rect 16454 25038 16470 25072
rect 16504 25038 16520 25072
rect 16454 25022 16520 25038
rect 16646 25072 16712 25088
rect 16646 25038 16662 25072
rect 16696 25038 16712 25072
rect 16646 25022 16712 25038
rect 15320 24991 15350 25022
rect 15416 24991 15446 25017
rect 15512 24991 15542 25022
rect 15608 24991 15638 25017
rect 15704 24991 15734 25022
rect 15800 24991 15830 25017
rect 15896 24991 15926 25022
rect 15992 24991 16022 25017
rect 16088 24991 16118 25022
rect 16184 24991 16214 25017
rect 16280 24991 16310 25022
rect 16376 24991 16406 25017
rect 16472 24991 16502 25022
rect 16568 24991 16598 25017
rect 16664 24991 16694 25022
rect 15320 24565 15350 24591
rect 15416 24560 15446 24591
rect 15512 24565 15542 24591
rect 15608 24560 15638 24591
rect 15704 24565 15734 24591
rect 15800 24560 15830 24591
rect 15896 24565 15926 24591
rect 15992 24560 16022 24591
rect 16088 24565 16118 24591
rect 16184 24560 16214 24591
rect 16280 24565 16310 24591
rect 16376 24560 16406 24591
rect 16472 24565 16502 24591
rect 16568 24560 16598 24591
rect 16664 24565 16694 24591
rect 15398 24544 15464 24560
rect 15398 24510 15414 24544
rect 15448 24510 15464 24544
rect 15398 24494 15464 24510
rect 15590 24544 15656 24560
rect 15590 24510 15606 24544
rect 15640 24510 15656 24544
rect 15590 24494 15656 24510
rect 15782 24544 15848 24560
rect 15782 24510 15798 24544
rect 15832 24510 15848 24544
rect 15782 24494 15848 24510
rect 15974 24544 16040 24560
rect 15974 24510 15990 24544
rect 16024 24510 16040 24544
rect 15974 24494 16040 24510
rect 16166 24544 16232 24560
rect 16166 24510 16182 24544
rect 16216 24510 16232 24544
rect 16166 24494 16232 24510
rect 16358 24544 16424 24560
rect 16358 24510 16374 24544
rect 16408 24510 16424 24544
rect 16358 24494 16424 24510
rect 16550 24544 16616 24560
rect 16550 24510 16566 24544
rect 16600 24510 16616 24544
rect 16550 24494 16616 24510
rect 15398 24436 15464 24452
rect 15398 24402 15414 24436
rect 15448 24402 15464 24436
rect 15398 24386 15464 24402
rect 15590 24436 15656 24452
rect 15590 24402 15606 24436
rect 15640 24402 15656 24436
rect 15590 24386 15656 24402
rect 15782 24436 15848 24452
rect 15782 24402 15798 24436
rect 15832 24402 15848 24436
rect 15782 24386 15848 24402
rect 15974 24436 16040 24452
rect 15974 24402 15990 24436
rect 16024 24402 16040 24436
rect 15974 24386 16040 24402
rect 16166 24436 16232 24452
rect 16166 24402 16182 24436
rect 16216 24402 16232 24436
rect 16166 24386 16232 24402
rect 16358 24436 16424 24452
rect 16358 24402 16374 24436
rect 16408 24402 16424 24436
rect 16358 24386 16424 24402
rect 16550 24436 16616 24452
rect 16550 24402 16566 24436
rect 16600 24402 16616 24436
rect 16550 24386 16616 24402
rect 15320 24355 15350 24381
rect 15416 24355 15446 24386
rect 15512 24355 15542 24381
rect 15608 24355 15638 24386
rect 15704 24355 15734 24381
rect 15800 24355 15830 24386
rect 15896 24355 15926 24381
rect 15992 24355 16022 24386
rect 16088 24355 16118 24381
rect 16184 24355 16214 24386
rect 16280 24355 16310 24381
rect 16376 24355 16406 24386
rect 16472 24355 16502 24381
rect 16568 24355 16598 24386
rect 16664 24355 16694 24381
rect 15320 23924 15350 23955
rect 15416 23929 15446 23955
rect 15512 23924 15542 23955
rect 15608 23929 15638 23955
rect 15704 23924 15734 23955
rect 15800 23929 15830 23955
rect 15896 23924 15926 23955
rect 15992 23929 16022 23955
rect 16088 23924 16118 23955
rect 16184 23929 16214 23955
rect 16280 23924 16310 23955
rect 16376 23929 16406 23955
rect 16472 23924 16502 23955
rect 16568 23929 16598 23955
rect 16664 23924 16694 23955
rect 15302 23908 15368 23924
rect 15302 23874 15318 23908
rect 15352 23874 15368 23908
rect 15302 23858 15368 23874
rect 15494 23908 15560 23924
rect 15494 23874 15510 23908
rect 15544 23874 15560 23908
rect 15494 23858 15560 23874
rect 15686 23908 15752 23924
rect 15686 23874 15702 23908
rect 15736 23874 15752 23908
rect 15686 23858 15752 23874
rect 15878 23908 15944 23924
rect 15878 23874 15894 23908
rect 15928 23874 15944 23908
rect 15878 23858 15944 23874
rect 16070 23908 16136 23924
rect 16070 23874 16086 23908
rect 16120 23874 16136 23908
rect 16070 23858 16136 23874
rect 16262 23908 16328 23924
rect 16262 23874 16278 23908
rect 16312 23874 16328 23908
rect 16262 23858 16328 23874
rect 16454 23908 16520 23924
rect 16454 23874 16470 23908
rect 16504 23874 16520 23908
rect 16454 23858 16520 23874
rect 16646 23908 16712 23924
rect 16646 23874 16662 23908
rect 16696 23874 16712 23908
rect 16646 23858 16712 23874
rect 6738 23494 6804 23510
rect 6738 23460 6754 23494
rect 6788 23460 6804 23494
rect 6660 23422 6690 23448
rect 6738 23444 6804 23460
rect 6930 23494 6996 23510
rect 6930 23460 6946 23494
rect 6980 23460 6996 23494
rect 6756 23422 6786 23444
rect 6852 23422 6882 23448
rect 6930 23444 6996 23460
rect 7122 23494 7188 23510
rect 7122 23460 7138 23494
rect 7172 23460 7188 23494
rect 6948 23422 6978 23444
rect 7044 23422 7074 23448
rect 7122 23444 7188 23460
rect 7314 23494 7380 23510
rect 7314 23460 7330 23494
rect 7364 23460 7380 23494
rect 7140 23422 7170 23444
rect 7236 23422 7266 23448
rect 7314 23444 7380 23460
rect 7506 23494 7572 23510
rect 7506 23460 7522 23494
rect 7556 23460 7572 23494
rect 7332 23422 7362 23444
rect 7428 23422 7458 23448
rect 7506 23444 7572 23460
rect 7524 23422 7554 23444
rect 6660 23000 6690 23022
rect 6642 22984 6708 23000
rect 6756 22996 6786 23022
rect 6852 23000 6882 23022
rect 6642 22950 6658 22984
rect 6692 22950 6708 22984
rect 6642 22934 6708 22950
rect 6834 22984 6900 23000
rect 6948 22996 6978 23022
rect 7044 23000 7074 23022
rect 6834 22950 6850 22984
rect 6884 22950 6900 22984
rect 6834 22934 6900 22950
rect 7026 22984 7092 23000
rect 7140 22996 7170 23022
rect 7236 23000 7266 23022
rect 7026 22950 7042 22984
rect 7076 22950 7092 22984
rect 7026 22934 7092 22950
rect 7218 22984 7284 23000
rect 7332 22996 7362 23022
rect 7428 23000 7458 23022
rect 7218 22950 7234 22984
rect 7268 22950 7284 22984
rect 7218 22934 7284 22950
rect 7410 22984 7476 23000
rect 7524 22996 7554 23022
rect 7410 22950 7426 22984
rect 7460 22950 7476 22984
rect 7410 22934 7476 22950
rect 6642 22876 6708 22892
rect 6642 22842 6658 22876
rect 6692 22842 6708 22876
rect 6642 22826 6708 22842
rect 6834 22876 6900 22892
rect 6834 22842 6850 22876
rect 6884 22842 6900 22876
rect 6660 22804 6690 22826
rect 6756 22804 6786 22830
rect 6834 22826 6900 22842
rect 7026 22876 7092 22892
rect 7026 22842 7042 22876
rect 7076 22842 7092 22876
rect 6852 22804 6882 22826
rect 6948 22804 6978 22830
rect 7026 22826 7092 22842
rect 7218 22876 7284 22892
rect 7218 22842 7234 22876
rect 7268 22842 7284 22876
rect 7044 22804 7074 22826
rect 7140 22804 7170 22830
rect 7218 22826 7284 22842
rect 7410 22876 7476 22892
rect 7410 22842 7426 22876
rect 7460 22842 7476 22876
rect 7236 22804 7266 22826
rect 7332 22804 7362 22830
rect 7410 22826 7476 22842
rect 7428 22804 7458 22826
rect 7524 22804 7554 22830
rect 6660 22378 6690 22404
rect 6756 22382 6786 22404
rect 6738 22366 6804 22382
rect 6852 22378 6882 22404
rect 6948 22382 6978 22404
rect 6738 22332 6754 22366
rect 6788 22332 6804 22366
rect 6738 22316 6804 22332
rect 6930 22366 6996 22382
rect 7044 22378 7074 22404
rect 7140 22382 7170 22404
rect 6930 22332 6946 22366
rect 6980 22332 6996 22366
rect 6930 22316 6996 22332
rect 7122 22366 7188 22382
rect 7236 22378 7266 22404
rect 7332 22382 7362 22404
rect 7122 22332 7138 22366
rect 7172 22332 7188 22366
rect 7122 22316 7188 22332
rect 7314 22366 7380 22382
rect 7428 22378 7458 22404
rect 7524 22382 7554 22404
rect 7314 22332 7330 22366
rect 7364 22332 7380 22366
rect 7314 22316 7380 22332
rect 7506 22366 7572 22382
rect 7506 22332 7522 22366
rect 7556 22332 7572 22366
rect 7506 22316 7572 22332
rect 6738 22258 6804 22274
rect 6738 22224 6754 22258
rect 6788 22224 6804 22258
rect 6660 22186 6690 22212
rect 6738 22208 6804 22224
rect 6930 22258 6996 22274
rect 6930 22224 6946 22258
rect 6980 22224 6996 22258
rect 6756 22186 6786 22208
rect 6852 22186 6882 22212
rect 6930 22208 6996 22224
rect 7122 22258 7188 22274
rect 7122 22224 7138 22258
rect 7172 22224 7188 22258
rect 6948 22186 6978 22208
rect 7044 22186 7074 22212
rect 7122 22208 7188 22224
rect 7314 22258 7380 22274
rect 7314 22224 7330 22258
rect 7364 22224 7380 22258
rect 7140 22186 7170 22208
rect 7236 22186 7266 22212
rect 7314 22208 7380 22224
rect 7506 22258 7572 22274
rect 7506 22224 7522 22258
rect 7556 22224 7572 22258
rect 7332 22186 7362 22208
rect 7428 22186 7458 22212
rect 7506 22208 7572 22224
rect 7524 22186 7554 22208
rect 6660 21764 6690 21786
rect 6642 21748 6708 21764
rect 6756 21760 6786 21786
rect 6852 21764 6882 21786
rect 6642 21714 6658 21748
rect 6692 21714 6708 21748
rect 6642 21698 6708 21714
rect 6834 21748 6900 21764
rect 6948 21760 6978 21786
rect 7044 21764 7074 21786
rect 6834 21714 6850 21748
rect 6884 21714 6900 21748
rect 6834 21698 6900 21714
rect 7026 21748 7092 21764
rect 7140 21760 7170 21786
rect 7236 21764 7266 21786
rect 7026 21714 7042 21748
rect 7076 21714 7092 21748
rect 7026 21698 7092 21714
rect 7218 21748 7284 21764
rect 7332 21760 7362 21786
rect 7428 21764 7458 21786
rect 7218 21714 7234 21748
rect 7268 21714 7284 21748
rect 7218 21698 7284 21714
rect 7410 21748 7476 21764
rect 7524 21760 7554 21786
rect 7410 21714 7426 21748
rect 7460 21714 7476 21748
rect 7410 21698 7476 21714
rect 8458 23494 8524 23510
rect 8458 23460 8474 23494
rect 8508 23460 8524 23494
rect 8380 23422 8410 23448
rect 8458 23444 8524 23460
rect 8650 23494 8716 23510
rect 8650 23460 8666 23494
rect 8700 23460 8716 23494
rect 8476 23422 8506 23444
rect 8572 23422 8602 23448
rect 8650 23444 8716 23460
rect 8842 23494 8908 23510
rect 8842 23460 8858 23494
rect 8892 23460 8908 23494
rect 8668 23422 8698 23444
rect 8764 23422 8794 23448
rect 8842 23444 8908 23460
rect 9034 23494 9100 23510
rect 9034 23460 9050 23494
rect 9084 23460 9100 23494
rect 8860 23422 8890 23444
rect 8956 23422 8986 23448
rect 9034 23444 9100 23460
rect 9226 23494 9292 23510
rect 9226 23460 9242 23494
rect 9276 23460 9292 23494
rect 9052 23422 9082 23444
rect 9148 23422 9178 23448
rect 9226 23444 9292 23460
rect 9244 23422 9274 23444
rect 8380 23000 8410 23022
rect 8362 22984 8428 23000
rect 8476 22996 8506 23022
rect 8572 23000 8602 23022
rect 8362 22950 8378 22984
rect 8412 22950 8428 22984
rect 8362 22934 8428 22950
rect 8554 22984 8620 23000
rect 8668 22996 8698 23022
rect 8764 23000 8794 23022
rect 8554 22950 8570 22984
rect 8604 22950 8620 22984
rect 8554 22934 8620 22950
rect 8746 22984 8812 23000
rect 8860 22996 8890 23022
rect 8956 23000 8986 23022
rect 8746 22950 8762 22984
rect 8796 22950 8812 22984
rect 8746 22934 8812 22950
rect 8938 22984 9004 23000
rect 9052 22996 9082 23022
rect 9148 23000 9178 23022
rect 8938 22950 8954 22984
rect 8988 22950 9004 22984
rect 8938 22934 9004 22950
rect 9130 22984 9196 23000
rect 9244 22996 9274 23022
rect 9130 22950 9146 22984
rect 9180 22950 9196 22984
rect 9130 22934 9196 22950
rect 8362 22876 8428 22892
rect 8362 22842 8378 22876
rect 8412 22842 8428 22876
rect 8362 22826 8428 22842
rect 8554 22876 8620 22892
rect 8554 22842 8570 22876
rect 8604 22842 8620 22876
rect 8380 22804 8410 22826
rect 8476 22804 8506 22830
rect 8554 22826 8620 22842
rect 8746 22876 8812 22892
rect 8746 22842 8762 22876
rect 8796 22842 8812 22876
rect 8572 22804 8602 22826
rect 8668 22804 8698 22830
rect 8746 22826 8812 22842
rect 8938 22876 9004 22892
rect 8938 22842 8954 22876
rect 8988 22842 9004 22876
rect 8764 22804 8794 22826
rect 8860 22804 8890 22830
rect 8938 22826 9004 22842
rect 9130 22876 9196 22892
rect 9130 22842 9146 22876
rect 9180 22842 9196 22876
rect 8956 22804 8986 22826
rect 9052 22804 9082 22830
rect 9130 22826 9196 22842
rect 9148 22804 9178 22826
rect 9244 22804 9274 22830
rect 8380 22378 8410 22404
rect 8476 22382 8506 22404
rect 8458 22366 8524 22382
rect 8572 22378 8602 22404
rect 8668 22382 8698 22404
rect 8458 22332 8474 22366
rect 8508 22332 8524 22366
rect 8458 22316 8524 22332
rect 8650 22366 8716 22382
rect 8764 22378 8794 22404
rect 8860 22382 8890 22404
rect 8650 22332 8666 22366
rect 8700 22332 8716 22366
rect 8650 22316 8716 22332
rect 8842 22366 8908 22382
rect 8956 22378 8986 22404
rect 9052 22382 9082 22404
rect 8842 22332 8858 22366
rect 8892 22332 8908 22366
rect 8842 22316 8908 22332
rect 9034 22366 9100 22382
rect 9148 22378 9178 22404
rect 9244 22382 9274 22404
rect 9034 22332 9050 22366
rect 9084 22332 9100 22366
rect 9034 22316 9100 22332
rect 9226 22366 9292 22382
rect 9226 22332 9242 22366
rect 9276 22332 9292 22366
rect 9226 22316 9292 22332
rect 8458 22258 8524 22274
rect 8458 22224 8474 22258
rect 8508 22224 8524 22258
rect 8380 22186 8410 22212
rect 8458 22208 8524 22224
rect 8650 22258 8716 22274
rect 8650 22224 8666 22258
rect 8700 22224 8716 22258
rect 8476 22186 8506 22208
rect 8572 22186 8602 22212
rect 8650 22208 8716 22224
rect 8842 22258 8908 22274
rect 8842 22224 8858 22258
rect 8892 22224 8908 22258
rect 8668 22186 8698 22208
rect 8764 22186 8794 22212
rect 8842 22208 8908 22224
rect 9034 22258 9100 22274
rect 9034 22224 9050 22258
rect 9084 22224 9100 22258
rect 8860 22186 8890 22208
rect 8956 22186 8986 22212
rect 9034 22208 9100 22224
rect 9226 22258 9292 22274
rect 9226 22224 9242 22258
rect 9276 22224 9292 22258
rect 9052 22186 9082 22208
rect 9148 22186 9178 22212
rect 9226 22208 9292 22224
rect 9244 22186 9274 22208
rect 8380 21764 8410 21786
rect 8362 21748 8428 21764
rect 8476 21760 8506 21786
rect 8572 21764 8602 21786
rect 8362 21714 8378 21748
rect 8412 21714 8428 21748
rect 8362 21698 8428 21714
rect 8554 21748 8620 21764
rect 8668 21760 8698 21786
rect 8764 21764 8794 21786
rect 8554 21714 8570 21748
rect 8604 21714 8620 21748
rect 8554 21698 8620 21714
rect 8746 21748 8812 21764
rect 8860 21760 8890 21786
rect 8956 21764 8986 21786
rect 8746 21714 8762 21748
rect 8796 21714 8812 21748
rect 8746 21698 8812 21714
rect 8938 21748 9004 21764
rect 9052 21760 9082 21786
rect 9148 21764 9178 21786
rect 8938 21714 8954 21748
rect 8988 21714 9004 21748
rect 8938 21698 9004 21714
rect 9130 21748 9196 21764
rect 9244 21760 9274 21786
rect 9130 21714 9146 21748
rect 9180 21714 9196 21748
rect 9130 21698 9196 21714
rect 18942 25020 19039 25036
rect 18942 23452 18958 25020
rect 18992 23452 19039 25020
rect 18942 23436 19039 23452
rect 19239 25020 19336 25036
rect 19239 23452 19286 25020
rect 19320 23452 19336 25020
rect 19239 23436 19336 23452
rect 18438 23104 18504 23120
rect 18438 23070 18454 23104
rect 18488 23070 18504 23104
rect 18438 23054 18504 23070
rect 18630 23104 18696 23120
rect 18630 23070 18646 23104
rect 18680 23070 18696 23104
rect 18630 23054 18696 23070
rect 18822 23104 18888 23120
rect 18822 23070 18838 23104
rect 18872 23070 18888 23104
rect 18822 23054 18888 23070
rect 19014 23104 19080 23120
rect 19014 23070 19030 23104
rect 19064 23070 19080 23104
rect 19014 23054 19080 23070
rect 19206 23104 19272 23120
rect 19206 23070 19222 23104
rect 19256 23070 19272 23104
rect 19206 23054 19272 23070
rect 18360 23023 18390 23049
rect 18456 23023 18486 23054
rect 18552 23023 18582 23049
rect 18648 23023 18678 23054
rect 18744 23023 18774 23049
rect 18840 23023 18870 23054
rect 18936 23023 18966 23049
rect 19032 23023 19062 23054
rect 19128 23023 19158 23049
rect 19224 23023 19254 23054
rect 18360 22592 18390 22623
rect 18456 22597 18486 22623
rect 18552 22592 18582 22623
rect 18648 22597 18678 22623
rect 18744 22592 18774 22623
rect 18840 22597 18870 22623
rect 18936 22592 18966 22623
rect 19032 22597 19062 22623
rect 19128 22592 19158 22623
rect 19224 22597 19254 22623
rect 18342 22576 18408 22592
rect 18342 22542 18358 22576
rect 18392 22542 18408 22576
rect 18342 22526 18408 22542
rect 18534 22576 18600 22592
rect 18534 22542 18550 22576
rect 18584 22542 18600 22576
rect 18534 22526 18600 22542
rect 18726 22576 18792 22592
rect 18726 22542 18742 22576
rect 18776 22542 18792 22576
rect 18726 22526 18792 22542
rect 18918 22576 18984 22592
rect 18918 22542 18934 22576
rect 18968 22542 18984 22576
rect 18918 22526 18984 22542
rect 19110 22576 19176 22592
rect 19110 22542 19126 22576
rect 19160 22542 19176 22576
rect 19110 22526 19176 22542
rect 6656 21348 6856 21364
rect 6656 21314 6672 21348
rect 6840 21314 6856 21348
rect 6656 21276 6856 21314
rect 6914 21348 7114 21364
rect 6914 21314 6930 21348
rect 7098 21314 7114 21348
rect 6914 21276 7114 21314
rect 7172 21348 7372 21364
rect 7172 21314 7188 21348
rect 7356 21314 7372 21348
rect 7172 21276 7372 21314
rect 7430 21348 7630 21364
rect 7430 21314 7446 21348
rect 7614 21314 7630 21348
rect 7430 21276 7630 21314
rect 7688 21348 7888 21364
rect 7688 21314 7704 21348
rect 7872 21314 7888 21348
rect 7688 21276 7888 21314
rect 6656 20838 6856 20876
rect 6656 20804 6672 20838
rect 6840 20804 6856 20838
rect 6656 20788 6856 20804
rect 6914 20838 7114 20876
rect 6914 20804 6930 20838
rect 7098 20804 7114 20838
rect 6914 20788 7114 20804
rect 7172 20838 7372 20876
rect 7172 20804 7188 20838
rect 7356 20804 7372 20838
rect 7172 20788 7372 20804
rect 7430 20838 7630 20876
rect 7430 20804 7446 20838
rect 7614 20804 7630 20838
rect 7430 20788 7630 20804
rect 7688 20838 7888 20876
rect 7688 20804 7704 20838
rect 7872 20804 7888 20838
rect 7688 20788 7888 20804
rect 6656 20730 6856 20746
rect 6656 20696 6672 20730
rect 6840 20696 6856 20730
rect 6656 20658 6856 20696
rect 6914 20730 7114 20746
rect 6914 20696 6930 20730
rect 7098 20696 7114 20730
rect 6914 20658 7114 20696
rect 7172 20730 7372 20746
rect 7172 20696 7188 20730
rect 7356 20696 7372 20730
rect 7172 20658 7372 20696
rect 7430 20730 7630 20746
rect 7430 20696 7446 20730
rect 7614 20696 7630 20730
rect 7430 20658 7630 20696
rect 7688 20730 7888 20746
rect 7688 20696 7704 20730
rect 7872 20696 7888 20730
rect 7688 20658 7888 20696
rect 6656 20220 6856 20258
rect 6656 20186 6672 20220
rect 6840 20186 6856 20220
rect 6656 20170 6856 20186
rect 6914 20220 7114 20258
rect 6914 20186 6930 20220
rect 7098 20186 7114 20220
rect 6914 20170 7114 20186
rect 7172 20220 7372 20258
rect 7172 20186 7188 20220
rect 7356 20186 7372 20220
rect 7172 20170 7372 20186
rect 7430 20220 7630 20258
rect 7430 20186 7446 20220
rect 7614 20186 7630 20220
rect 7430 20170 7630 20186
rect 7688 20220 7888 20258
rect 7688 20186 7704 20220
rect 7872 20186 7888 20220
rect 7688 20170 7888 20186
rect 6656 20112 6856 20128
rect 6656 20078 6672 20112
rect 6840 20078 6856 20112
rect 6656 20040 6856 20078
rect 6914 20112 7114 20128
rect 6914 20078 6930 20112
rect 7098 20078 7114 20112
rect 6914 20040 7114 20078
rect 7172 20112 7372 20128
rect 7172 20078 7188 20112
rect 7356 20078 7372 20112
rect 7172 20040 7372 20078
rect 7430 20112 7630 20128
rect 7430 20078 7446 20112
rect 7614 20078 7630 20112
rect 7430 20040 7630 20078
rect 7688 20112 7888 20128
rect 7688 20078 7704 20112
rect 7872 20078 7888 20112
rect 7688 20040 7888 20078
rect 6656 19602 6856 19640
rect 6656 19568 6672 19602
rect 6840 19568 6856 19602
rect 6656 19552 6856 19568
rect 6914 19602 7114 19640
rect 6914 19568 6930 19602
rect 7098 19568 7114 19602
rect 6914 19552 7114 19568
rect 7172 19602 7372 19640
rect 7172 19568 7188 19602
rect 7356 19568 7372 19602
rect 7172 19552 7372 19568
rect 7430 19602 7630 19640
rect 7430 19568 7446 19602
rect 7614 19568 7630 19602
rect 7430 19552 7630 19568
rect 7688 19602 7888 19640
rect 7688 19568 7704 19602
rect 7872 19568 7888 19602
rect 7688 19552 7888 19568
rect 6656 19494 6856 19510
rect 6656 19460 6672 19494
rect 6840 19460 6856 19494
rect 6656 19422 6856 19460
rect 6914 19494 7114 19510
rect 6914 19460 6930 19494
rect 7098 19460 7114 19494
rect 6914 19422 7114 19460
rect 7172 19494 7372 19510
rect 7172 19460 7188 19494
rect 7356 19460 7372 19494
rect 7172 19422 7372 19460
rect 7430 19494 7630 19510
rect 7430 19460 7446 19494
rect 7614 19460 7630 19494
rect 7430 19422 7630 19460
rect 7688 19494 7888 19510
rect 7688 19460 7704 19494
rect 7872 19460 7888 19494
rect 7688 19422 7888 19460
rect 6656 18984 6856 19022
rect 6656 18950 6672 18984
rect 6840 18950 6856 18984
rect 6656 18934 6856 18950
rect 6914 18984 7114 19022
rect 6914 18950 6930 18984
rect 7098 18950 7114 18984
rect 6914 18934 7114 18950
rect 7172 18984 7372 19022
rect 7172 18950 7188 18984
rect 7356 18950 7372 18984
rect 7172 18934 7372 18950
rect 7430 18984 7630 19022
rect 7430 18950 7446 18984
rect 7614 18950 7630 18984
rect 7430 18934 7630 18950
rect 7688 18984 7888 19022
rect 7688 18950 7704 18984
rect 7872 18950 7888 18984
rect 7688 18934 7888 18950
rect 6656 18876 6856 18892
rect 6656 18842 6672 18876
rect 6840 18842 6856 18876
rect 6656 18804 6856 18842
rect 6914 18876 7114 18892
rect 6914 18842 6930 18876
rect 7098 18842 7114 18876
rect 6914 18804 7114 18842
rect 7172 18876 7372 18892
rect 7172 18842 7188 18876
rect 7356 18842 7372 18876
rect 7172 18804 7372 18842
rect 7430 18876 7630 18892
rect 7430 18842 7446 18876
rect 7614 18842 7630 18876
rect 7430 18804 7630 18842
rect 7688 18876 7888 18892
rect 7688 18842 7704 18876
rect 7872 18842 7888 18876
rect 7688 18804 7888 18842
rect 6656 18366 6856 18404
rect 6656 18332 6672 18366
rect 6840 18332 6856 18366
rect 6656 18316 6856 18332
rect 6914 18366 7114 18404
rect 6914 18332 6930 18366
rect 7098 18332 7114 18366
rect 6914 18316 7114 18332
rect 7172 18366 7372 18404
rect 7172 18332 7188 18366
rect 7356 18332 7372 18366
rect 7172 18316 7372 18332
rect 7430 18366 7630 18404
rect 7430 18332 7446 18366
rect 7614 18332 7630 18366
rect 7430 18316 7630 18332
rect 7688 18366 7888 18404
rect 7688 18332 7704 18366
rect 7872 18332 7888 18366
rect 7688 18316 7888 18332
rect 6656 18258 6856 18274
rect 6656 18224 6672 18258
rect 6840 18224 6856 18258
rect 6656 18186 6856 18224
rect 6914 18258 7114 18274
rect 6914 18224 6930 18258
rect 7098 18224 7114 18258
rect 6914 18186 7114 18224
rect 7172 18258 7372 18274
rect 7172 18224 7188 18258
rect 7356 18224 7372 18258
rect 7172 18186 7372 18224
rect 7430 18258 7630 18274
rect 7430 18224 7446 18258
rect 7614 18224 7630 18258
rect 7430 18186 7630 18224
rect 7688 18258 7888 18274
rect 7688 18224 7704 18258
rect 7872 18224 7888 18258
rect 7688 18186 7888 18224
rect 6656 17748 6856 17786
rect 6656 17714 6672 17748
rect 6840 17714 6856 17748
rect 6656 17698 6856 17714
rect 6914 17748 7114 17786
rect 6914 17714 6930 17748
rect 7098 17714 7114 17748
rect 6914 17698 7114 17714
rect 7172 17748 7372 17786
rect 7172 17714 7188 17748
rect 7356 17714 7372 17748
rect 7172 17698 7372 17714
rect 7430 17748 7630 17786
rect 7430 17714 7446 17748
rect 7614 17714 7630 17748
rect 7430 17698 7630 17714
rect 7688 17748 7888 17786
rect 7688 17714 7704 17748
rect 7872 17714 7888 17748
rect 7688 17698 7888 17714
rect 8376 21348 8576 21364
rect 8376 21314 8392 21348
rect 8560 21314 8576 21348
rect 8376 21276 8576 21314
rect 8634 21348 8834 21364
rect 8634 21314 8650 21348
rect 8818 21314 8834 21348
rect 8634 21276 8834 21314
rect 8892 21348 9092 21364
rect 8892 21314 8908 21348
rect 9076 21314 9092 21348
rect 8892 21276 9092 21314
rect 9150 21348 9350 21364
rect 9150 21314 9166 21348
rect 9334 21314 9350 21348
rect 9150 21276 9350 21314
rect 9408 21348 9608 21364
rect 9408 21314 9424 21348
rect 9592 21314 9608 21348
rect 9408 21276 9608 21314
rect 8376 20838 8576 20876
rect 8376 20804 8392 20838
rect 8560 20804 8576 20838
rect 8376 20788 8576 20804
rect 8634 20838 8834 20876
rect 8634 20804 8650 20838
rect 8818 20804 8834 20838
rect 8634 20788 8834 20804
rect 8892 20838 9092 20876
rect 8892 20804 8908 20838
rect 9076 20804 9092 20838
rect 8892 20788 9092 20804
rect 9150 20838 9350 20876
rect 9150 20804 9166 20838
rect 9334 20804 9350 20838
rect 9150 20788 9350 20804
rect 9408 20838 9608 20876
rect 9408 20804 9424 20838
rect 9592 20804 9608 20838
rect 9408 20788 9608 20804
rect 8376 20730 8576 20746
rect 8376 20696 8392 20730
rect 8560 20696 8576 20730
rect 8376 20658 8576 20696
rect 8634 20730 8834 20746
rect 8634 20696 8650 20730
rect 8818 20696 8834 20730
rect 8634 20658 8834 20696
rect 8892 20730 9092 20746
rect 8892 20696 8908 20730
rect 9076 20696 9092 20730
rect 8892 20658 9092 20696
rect 9150 20730 9350 20746
rect 9150 20696 9166 20730
rect 9334 20696 9350 20730
rect 9150 20658 9350 20696
rect 9408 20730 9608 20746
rect 9408 20696 9424 20730
rect 9592 20696 9608 20730
rect 9408 20658 9608 20696
rect 8376 20220 8576 20258
rect 8376 20186 8392 20220
rect 8560 20186 8576 20220
rect 8376 20170 8576 20186
rect 8634 20220 8834 20258
rect 8634 20186 8650 20220
rect 8818 20186 8834 20220
rect 8634 20170 8834 20186
rect 8892 20220 9092 20258
rect 8892 20186 8908 20220
rect 9076 20186 9092 20220
rect 8892 20170 9092 20186
rect 9150 20220 9350 20258
rect 9150 20186 9166 20220
rect 9334 20186 9350 20220
rect 9150 20170 9350 20186
rect 9408 20220 9608 20258
rect 9408 20186 9424 20220
rect 9592 20186 9608 20220
rect 9408 20170 9608 20186
rect 8376 20112 8576 20128
rect 8376 20078 8392 20112
rect 8560 20078 8576 20112
rect 8376 20040 8576 20078
rect 8634 20112 8834 20128
rect 8634 20078 8650 20112
rect 8818 20078 8834 20112
rect 8634 20040 8834 20078
rect 8892 20112 9092 20128
rect 8892 20078 8908 20112
rect 9076 20078 9092 20112
rect 8892 20040 9092 20078
rect 9150 20112 9350 20128
rect 9150 20078 9166 20112
rect 9334 20078 9350 20112
rect 9150 20040 9350 20078
rect 9408 20112 9608 20128
rect 9408 20078 9424 20112
rect 9592 20078 9608 20112
rect 9408 20040 9608 20078
rect 8376 19602 8576 19640
rect 8376 19568 8392 19602
rect 8560 19568 8576 19602
rect 8376 19552 8576 19568
rect 8634 19602 8834 19640
rect 8634 19568 8650 19602
rect 8818 19568 8834 19602
rect 8634 19552 8834 19568
rect 8892 19602 9092 19640
rect 8892 19568 8908 19602
rect 9076 19568 9092 19602
rect 8892 19552 9092 19568
rect 9150 19602 9350 19640
rect 9150 19568 9166 19602
rect 9334 19568 9350 19602
rect 9150 19552 9350 19568
rect 9408 19602 9608 19640
rect 9408 19568 9424 19602
rect 9592 19568 9608 19602
rect 9408 19552 9608 19568
rect 8376 19494 8576 19510
rect 8376 19460 8392 19494
rect 8560 19460 8576 19494
rect 8376 19422 8576 19460
rect 8634 19494 8834 19510
rect 8634 19460 8650 19494
rect 8818 19460 8834 19494
rect 8634 19422 8834 19460
rect 8892 19494 9092 19510
rect 8892 19460 8908 19494
rect 9076 19460 9092 19494
rect 8892 19422 9092 19460
rect 9150 19494 9350 19510
rect 9150 19460 9166 19494
rect 9334 19460 9350 19494
rect 9150 19422 9350 19460
rect 9408 19494 9608 19510
rect 9408 19460 9424 19494
rect 9592 19460 9608 19494
rect 9408 19422 9608 19460
rect 8376 18984 8576 19022
rect 8376 18950 8392 18984
rect 8560 18950 8576 18984
rect 8376 18934 8576 18950
rect 8634 18984 8834 19022
rect 8634 18950 8650 18984
rect 8818 18950 8834 18984
rect 8634 18934 8834 18950
rect 8892 18984 9092 19022
rect 8892 18950 8908 18984
rect 9076 18950 9092 18984
rect 8892 18934 9092 18950
rect 9150 18984 9350 19022
rect 9150 18950 9166 18984
rect 9334 18950 9350 18984
rect 9150 18934 9350 18950
rect 9408 18984 9608 19022
rect 9408 18950 9424 18984
rect 9592 18950 9608 18984
rect 9408 18934 9608 18950
rect 8376 18876 8576 18892
rect 8376 18842 8392 18876
rect 8560 18842 8576 18876
rect 8376 18804 8576 18842
rect 8634 18876 8834 18892
rect 8634 18842 8650 18876
rect 8818 18842 8834 18876
rect 8634 18804 8834 18842
rect 8892 18876 9092 18892
rect 8892 18842 8908 18876
rect 9076 18842 9092 18876
rect 8892 18804 9092 18842
rect 9150 18876 9350 18892
rect 9150 18842 9166 18876
rect 9334 18842 9350 18876
rect 9150 18804 9350 18842
rect 9408 18876 9608 18892
rect 9408 18842 9424 18876
rect 9592 18842 9608 18876
rect 9408 18804 9608 18842
rect 8376 18366 8576 18404
rect 8376 18332 8392 18366
rect 8560 18332 8576 18366
rect 8376 18316 8576 18332
rect 8634 18366 8834 18404
rect 8634 18332 8650 18366
rect 8818 18332 8834 18366
rect 8634 18316 8834 18332
rect 8892 18366 9092 18404
rect 8892 18332 8908 18366
rect 9076 18332 9092 18366
rect 8892 18316 9092 18332
rect 9150 18366 9350 18404
rect 9150 18332 9166 18366
rect 9334 18332 9350 18366
rect 9150 18316 9350 18332
rect 9408 18366 9608 18404
rect 9408 18332 9424 18366
rect 9592 18332 9608 18366
rect 9408 18316 9608 18332
rect 8376 18258 8576 18274
rect 8376 18224 8392 18258
rect 8560 18224 8576 18258
rect 8376 18186 8576 18224
rect 8634 18258 8834 18274
rect 8634 18224 8650 18258
rect 8818 18224 8834 18258
rect 8634 18186 8834 18224
rect 8892 18258 9092 18274
rect 8892 18224 8908 18258
rect 9076 18224 9092 18258
rect 8892 18186 9092 18224
rect 9150 18258 9350 18274
rect 9150 18224 9166 18258
rect 9334 18224 9350 18258
rect 9150 18186 9350 18224
rect 9408 18258 9608 18274
rect 9408 18224 9424 18258
rect 9592 18224 9608 18258
rect 9408 18186 9608 18224
rect 8376 17748 8576 17786
rect 8376 17714 8392 17748
rect 8560 17714 8576 17748
rect 8376 17698 8576 17714
rect 8634 17748 8834 17786
rect 8634 17714 8650 17748
rect 8818 17714 8834 17748
rect 8634 17698 8834 17714
rect 8892 17748 9092 17786
rect 8892 17714 8908 17748
rect 9076 17714 9092 17748
rect 8892 17698 9092 17714
rect 9150 17748 9350 17786
rect 9150 17714 9166 17748
rect 9334 17714 9350 17748
rect 9150 17698 9350 17714
rect 9408 17748 9608 17786
rect 9408 17714 9424 17748
rect 9592 17714 9608 17748
rect 9408 17698 9608 17714
rect 18438 22236 18504 22252
rect 18438 22202 18454 22236
rect 18488 22202 18504 22236
rect 18360 22164 18390 22190
rect 18438 22186 18504 22202
rect 18630 22236 18696 22252
rect 18630 22202 18646 22236
rect 18680 22202 18696 22236
rect 18456 22164 18486 22186
rect 18552 22164 18582 22190
rect 18630 22186 18696 22202
rect 18822 22236 18888 22252
rect 18822 22202 18838 22236
rect 18872 22202 18888 22236
rect 18648 22164 18678 22186
rect 18744 22164 18774 22190
rect 18822 22186 18888 22202
rect 19014 22236 19080 22252
rect 19014 22202 19030 22236
rect 19064 22202 19080 22236
rect 18840 22164 18870 22186
rect 18936 22164 18966 22190
rect 19014 22186 19080 22202
rect 19206 22236 19272 22252
rect 19206 22202 19222 22236
rect 19256 22202 19272 22236
rect 19032 22164 19062 22186
rect 19128 22164 19158 22190
rect 19206 22186 19272 22202
rect 19224 22164 19254 22186
rect 18360 21742 18390 21764
rect 18342 21726 18408 21742
rect 18456 21738 18486 21764
rect 18552 21742 18582 21764
rect 18342 21692 18358 21726
rect 18392 21692 18408 21726
rect 18342 21676 18408 21692
rect 18534 21726 18600 21742
rect 18648 21738 18678 21764
rect 18744 21742 18774 21764
rect 18534 21692 18550 21726
rect 18584 21692 18600 21726
rect 18534 21676 18600 21692
rect 18726 21726 18792 21742
rect 18840 21738 18870 21764
rect 18936 21742 18966 21764
rect 18726 21692 18742 21726
rect 18776 21692 18792 21726
rect 18726 21676 18792 21692
rect 18918 21726 18984 21742
rect 19032 21738 19062 21764
rect 19128 21742 19158 21764
rect 18918 21692 18934 21726
rect 18968 21692 18984 21726
rect 18918 21676 18984 21692
rect 19110 21726 19176 21742
rect 19224 21738 19254 21764
rect 19110 21692 19126 21726
rect 19160 21692 19176 21726
rect 19110 21676 19176 21692
rect 18342 21618 18408 21634
rect 18342 21584 18358 21618
rect 18392 21584 18408 21618
rect 18342 21568 18408 21584
rect 18534 21618 18600 21634
rect 18534 21584 18550 21618
rect 18584 21584 18600 21618
rect 18360 21546 18390 21568
rect 18456 21546 18486 21572
rect 18534 21568 18600 21584
rect 18726 21618 18792 21634
rect 18726 21584 18742 21618
rect 18776 21584 18792 21618
rect 18552 21546 18582 21568
rect 18648 21546 18678 21572
rect 18726 21568 18792 21584
rect 18918 21618 18984 21634
rect 18918 21584 18934 21618
rect 18968 21584 18984 21618
rect 18744 21546 18774 21568
rect 18840 21546 18870 21572
rect 18918 21568 18984 21584
rect 19110 21618 19176 21634
rect 19110 21584 19126 21618
rect 19160 21584 19176 21618
rect 18936 21546 18966 21568
rect 19032 21546 19062 21572
rect 19110 21568 19176 21584
rect 19128 21546 19158 21568
rect 19224 21546 19254 21572
rect 18360 21120 18390 21146
rect 18456 21124 18486 21146
rect 18438 21108 18504 21124
rect 18552 21120 18582 21146
rect 18648 21124 18678 21146
rect 18438 21074 18454 21108
rect 18488 21074 18504 21108
rect 18438 21058 18504 21074
rect 18630 21108 18696 21124
rect 18744 21120 18774 21146
rect 18840 21124 18870 21146
rect 18630 21074 18646 21108
rect 18680 21074 18696 21108
rect 18630 21058 18696 21074
rect 18822 21108 18888 21124
rect 18936 21120 18966 21146
rect 19032 21124 19062 21146
rect 18822 21074 18838 21108
rect 18872 21074 18888 21108
rect 18822 21058 18888 21074
rect 19014 21108 19080 21124
rect 19128 21120 19158 21146
rect 19224 21124 19254 21146
rect 19014 21074 19030 21108
rect 19064 21074 19080 21108
rect 19014 21058 19080 21074
rect 19206 21108 19272 21124
rect 19206 21074 19222 21108
rect 19256 21074 19272 21108
rect 19206 21058 19272 21074
rect 10298 19798 10364 19814
rect 10298 19764 10314 19798
rect 10348 19764 10364 19798
rect 10220 19726 10250 19752
rect 10298 19748 10364 19764
rect 10490 19798 10556 19814
rect 10490 19764 10506 19798
rect 10540 19764 10556 19798
rect 10316 19726 10346 19748
rect 10412 19726 10442 19752
rect 10490 19748 10556 19764
rect 10682 19798 10748 19814
rect 10682 19764 10698 19798
rect 10732 19764 10748 19798
rect 10508 19726 10538 19748
rect 10604 19726 10634 19752
rect 10682 19748 10748 19764
rect 10700 19726 10730 19748
rect 10796 19726 10826 19752
rect 10220 19304 10250 19326
rect 10202 19288 10268 19304
rect 10316 19300 10346 19326
rect 10412 19304 10442 19326
rect 10202 19254 10218 19288
rect 10252 19254 10268 19288
rect 10202 19238 10268 19254
rect 10394 19288 10460 19304
rect 10508 19300 10538 19326
rect 10604 19304 10634 19326
rect 10394 19254 10410 19288
rect 10444 19254 10460 19288
rect 10394 19238 10460 19254
rect 10586 19288 10652 19304
rect 10700 19300 10730 19326
rect 10796 19304 10826 19326
rect 10586 19254 10602 19288
rect 10636 19254 10652 19288
rect 10586 19238 10652 19254
rect 10778 19288 10844 19304
rect 10778 19254 10794 19288
rect 10828 19254 10844 19288
rect 10778 19238 10844 19254
rect 10202 18876 10268 18892
rect 10202 18842 10218 18876
rect 10252 18842 10268 18876
rect 10202 18826 10268 18842
rect 10394 18876 10460 18892
rect 10394 18842 10410 18876
rect 10444 18842 10460 18876
rect 10220 18804 10250 18826
rect 10316 18804 10346 18830
rect 10394 18826 10460 18842
rect 10586 18876 10652 18892
rect 10586 18842 10602 18876
rect 10636 18842 10652 18876
rect 10412 18804 10442 18826
rect 10508 18804 10538 18830
rect 10586 18826 10652 18842
rect 10778 18876 10844 18892
rect 10778 18842 10794 18876
rect 10828 18842 10844 18876
rect 10604 18804 10634 18826
rect 10700 18804 10730 18830
rect 10778 18826 10844 18842
rect 10970 18876 11036 18892
rect 10970 18842 10986 18876
rect 11020 18842 11036 18876
rect 10796 18804 10826 18826
rect 10892 18804 10922 18830
rect 10970 18826 11036 18842
rect 10988 18804 11018 18826
rect 11084 18804 11114 18830
rect 10220 18378 10250 18404
rect 10316 18382 10346 18404
rect 10298 18366 10364 18382
rect 10412 18378 10442 18404
rect 10508 18382 10538 18404
rect 10298 18332 10314 18366
rect 10348 18332 10364 18366
rect 10298 18316 10364 18332
rect 10490 18366 10556 18382
rect 10604 18378 10634 18404
rect 10700 18382 10730 18404
rect 10490 18332 10506 18366
rect 10540 18332 10556 18366
rect 10490 18316 10556 18332
rect 10682 18366 10748 18382
rect 10796 18378 10826 18404
rect 10892 18382 10922 18404
rect 10682 18332 10698 18366
rect 10732 18332 10748 18366
rect 10682 18316 10748 18332
rect 10874 18366 10940 18382
rect 10988 18378 11018 18404
rect 11084 18382 11114 18404
rect 10874 18332 10890 18366
rect 10924 18332 10940 18366
rect 10874 18316 10940 18332
rect 11066 18366 11132 18382
rect 11066 18332 11082 18366
rect 11116 18332 11132 18366
rect 11066 18316 11132 18332
rect 10298 18258 10364 18274
rect 10298 18224 10314 18258
rect 10348 18224 10364 18258
rect 10220 18186 10250 18212
rect 10298 18208 10364 18224
rect 10490 18258 10556 18274
rect 10490 18224 10506 18258
rect 10540 18224 10556 18258
rect 10316 18186 10346 18208
rect 10412 18186 10442 18212
rect 10490 18208 10556 18224
rect 10682 18258 10748 18274
rect 10682 18224 10698 18258
rect 10732 18224 10748 18258
rect 10508 18186 10538 18208
rect 10604 18186 10634 18212
rect 10682 18208 10748 18224
rect 10874 18258 10940 18274
rect 10874 18224 10890 18258
rect 10924 18224 10940 18258
rect 10700 18186 10730 18208
rect 10796 18186 10826 18212
rect 10874 18208 10940 18224
rect 11066 18258 11132 18274
rect 11066 18224 11082 18258
rect 11116 18224 11132 18258
rect 10892 18186 10922 18208
rect 10988 18186 11018 18212
rect 11066 18208 11132 18224
rect 11084 18186 11114 18208
rect 10220 17764 10250 17786
rect 10202 17748 10268 17764
rect 10316 17760 10346 17786
rect 10412 17764 10442 17786
rect 10202 17714 10218 17748
rect 10252 17714 10268 17748
rect 10202 17698 10268 17714
rect 10394 17748 10460 17764
rect 10508 17760 10538 17786
rect 10604 17764 10634 17786
rect 10394 17714 10410 17748
rect 10444 17714 10460 17748
rect 10394 17698 10460 17714
rect 10586 17748 10652 17764
rect 10700 17760 10730 17786
rect 10796 17764 10826 17786
rect 10586 17714 10602 17748
rect 10636 17714 10652 17748
rect 10586 17698 10652 17714
rect 10778 17748 10844 17764
rect 10892 17760 10922 17786
rect 10988 17764 11018 17786
rect 10778 17714 10794 17748
rect 10828 17714 10844 17748
rect 10778 17698 10844 17714
rect 10970 17748 11036 17764
rect 11084 17760 11114 17786
rect 10970 17714 10986 17748
rect 11020 17714 11036 17748
rect 10970 17698 11036 17714
rect 18356 20752 18556 20768
rect 18356 20718 18372 20752
rect 18540 20718 18556 20752
rect 18356 20680 18556 20718
rect 18614 20752 18814 20768
rect 18614 20718 18630 20752
rect 18798 20718 18814 20752
rect 18614 20680 18814 20718
rect 18872 20752 19072 20768
rect 18872 20718 18888 20752
rect 19056 20718 19072 20752
rect 18872 20680 19072 20718
rect 19130 20752 19330 20768
rect 19130 20718 19146 20752
rect 19314 20718 19330 20752
rect 19130 20680 19330 20718
rect 19388 20752 19588 20768
rect 19388 20718 19404 20752
rect 19572 20718 19588 20752
rect 19388 20680 19588 20718
rect 18356 20242 18556 20280
rect 18356 20208 18372 20242
rect 18540 20208 18556 20242
rect 18356 20192 18556 20208
rect 18614 20242 18814 20280
rect 18614 20208 18630 20242
rect 18798 20208 18814 20242
rect 18614 20192 18814 20208
rect 18872 20242 19072 20280
rect 18872 20208 18888 20242
rect 19056 20208 19072 20242
rect 18872 20192 19072 20208
rect 19130 20242 19330 20280
rect 19130 20208 19146 20242
rect 19314 20208 19330 20242
rect 19130 20192 19330 20208
rect 19388 20242 19588 20280
rect 19388 20208 19404 20242
rect 19572 20208 19588 20242
rect 19388 20192 19588 20208
rect 18356 20134 18556 20150
rect 18356 20100 18372 20134
rect 18540 20100 18556 20134
rect 18356 20062 18556 20100
rect 18614 20134 18814 20150
rect 18614 20100 18630 20134
rect 18798 20100 18814 20134
rect 18614 20062 18814 20100
rect 18872 20134 19072 20150
rect 18872 20100 18888 20134
rect 19056 20100 19072 20134
rect 18872 20062 19072 20100
rect 19130 20134 19330 20150
rect 19130 20100 19146 20134
rect 19314 20100 19330 20134
rect 19130 20062 19330 20100
rect 19388 20134 19588 20150
rect 19388 20100 19404 20134
rect 19572 20100 19588 20134
rect 19388 20062 19588 20100
rect 18356 19624 18556 19662
rect 18356 19590 18372 19624
rect 18540 19590 18556 19624
rect 18356 19574 18556 19590
rect 18614 19624 18814 19662
rect 18614 19590 18630 19624
rect 18798 19590 18814 19624
rect 18614 19574 18814 19590
rect 18872 19624 19072 19662
rect 18872 19590 18888 19624
rect 19056 19590 19072 19624
rect 18872 19574 19072 19590
rect 19130 19624 19330 19662
rect 19130 19590 19146 19624
rect 19314 19590 19330 19624
rect 19130 19574 19330 19590
rect 19388 19624 19588 19662
rect 19388 19590 19404 19624
rect 19572 19590 19588 19624
rect 19388 19574 19588 19590
rect 18356 19516 18556 19532
rect 18356 19482 18372 19516
rect 18540 19482 18556 19516
rect 18356 19444 18556 19482
rect 18614 19516 18814 19532
rect 18614 19482 18630 19516
rect 18798 19482 18814 19516
rect 18614 19444 18814 19482
rect 18872 19516 19072 19532
rect 18872 19482 18888 19516
rect 19056 19482 19072 19516
rect 18872 19444 19072 19482
rect 19130 19516 19330 19532
rect 19130 19482 19146 19516
rect 19314 19482 19330 19516
rect 19130 19444 19330 19482
rect 19388 19516 19588 19532
rect 19388 19482 19404 19516
rect 19572 19482 19588 19516
rect 19388 19444 19588 19482
rect 18356 19006 18556 19044
rect 18356 18972 18372 19006
rect 18540 18972 18556 19006
rect 18356 18956 18556 18972
rect 18614 19006 18814 19044
rect 18614 18972 18630 19006
rect 18798 18972 18814 19006
rect 18614 18956 18814 18972
rect 18872 19006 19072 19044
rect 18872 18972 18888 19006
rect 19056 18972 19072 19006
rect 18872 18956 19072 18972
rect 19130 19006 19330 19044
rect 19130 18972 19146 19006
rect 19314 18972 19330 19006
rect 19130 18956 19330 18972
rect 19388 19006 19588 19044
rect 19388 18972 19404 19006
rect 19572 18972 19588 19006
rect 19388 18956 19588 18972
rect 18356 18898 18556 18914
rect 18356 18864 18372 18898
rect 18540 18864 18556 18898
rect 18356 18826 18556 18864
rect 18614 18898 18814 18914
rect 18614 18864 18630 18898
rect 18798 18864 18814 18898
rect 18614 18826 18814 18864
rect 18872 18898 19072 18914
rect 18872 18864 18888 18898
rect 19056 18864 19072 18898
rect 18872 18826 19072 18864
rect 19130 18898 19330 18914
rect 19130 18864 19146 18898
rect 19314 18864 19330 18898
rect 19130 18826 19330 18864
rect 19388 18898 19588 18914
rect 19388 18864 19404 18898
rect 19572 18864 19588 18898
rect 19388 18826 19588 18864
rect 18356 18388 18556 18426
rect 18356 18354 18372 18388
rect 18540 18354 18556 18388
rect 18356 18338 18556 18354
rect 18614 18388 18814 18426
rect 18614 18354 18630 18388
rect 18798 18354 18814 18388
rect 18614 18338 18814 18354
rect 18872 18388 19072 18426
rect 18872 18354 18888 18388
rect 19056 18354 19072 18388
rect 18872 18338 19072 18354
rect 19130 18388 19330 18426
rect 19130 18354 19146 18388
rect 19314 18354 19330 18388
rect 19130 18338 19330 18354
rect 19388 18388 19588 18426
rect 19388 18354 19404 18388
rect 19572 18354 19588 18388
rect 19388 18338 19588 18354
rect -9922 8306 -9856 8322
rect -9922 8272 -9906 8306
rect -9872 8272 -9856 8306
rect -10000 8234 -9970 8260
rect -9922 8256 -9856 8272
rect -9730 8306 -9664 8322
rect -9730 8272 -9714 8306
rect -9680 8272 -9664 8306
rect -9904 8234 -9874 8256
rect -9808 8234 -9778 8260
rect -9730 8256 -9664 8272
rect -9538 8306 -9472 8322
rect -9538 8272 -9522 8306
rect -9488 8272 -9472 8306
rect -9712 8234 -9682 8256
rect -9616 8234 -9586 8260
rect -9538 8256 -9472 8272
rect -9346 8306 -9280 8322
rect -9346 8272 -9330 8306
rect -9296 8272 -9280 8306
rect -9520 8234 -9490 8256
rect -9424 8234 -9394 8260
rect -9346 8256 -9280 8272
rect -9154 8306 -9088 8322
rect -9154 8272 -9138 8306
rect -9104 8272 -9088 8306
rect -9328 8234 -9298 8256
rect -9232 8234 -9202 8260
rect -9154 8256 -9088 8272
rect -9136 8234 -9106 8256
rect -10000 7812 -9970 7834
rect -10018 7796 -9952 7812
rect -9904 7808 -9874 7834
rect -9808 7812 -9778 7834
rect -10018 7762 -10002 7796
rect -9968 7762 -9952 7796
rect -10018 7746 -9952 7762
rect -9826 7796 -9760 7812
rect -9712 7808 -9682 7834
rect -9616 7812 -9586 7834
rect -9826 7762 -9810 7796
rect -9776 7762 -9760 7796
rect -9826 7746 -9760 7762
rect -9634 7796 -9568 7812
rect -9520 7808 -9490 7834
rect -9424 7812 -9394 7834
rect -9634 7762 -9618 7796
rect -9584 7762 -9568 7796
rect -9634 7746 -9568 7762
rect -9442 7796 -9376 7812
rect -9328 7808 -9298 7834
rect -9232 7812 -9202 7834
rect -9442 7762 -9426 7796
rect -9392 7762 -9376 7796
rect -9442 7746 -9376 7762
rect -9250 7796 -9184 7812
rect -9136 7808 -9106 7834
rect -9250 7762 -9234 7796
rect -9200 7762 -9184 7796
rect -9250 7746 -9184 7762
rect -10018 7688 -9952 7704
rect -10018 7654 -10002 7688
rect -9968 7654 -9952 7688
rect -10018 7638 -9952 7654
rect -9826 7688 -9760 7704
rect -9826 7654 -9810 7688
rect -9776 7654 -9760 7688
rect -10000 7616 -9970 7638
rect -9904 7616 -9874 7642
rect -9826 7638 -9760 7654
rect -9634 7688 -9568 7704
rect -9634 7654 -9618 7688
rect -9584 7654 -9568 7688
rect -9808 7616 -9778 7638
rect -9712 7616 -9682 7642
rect -9634 7638 -9568 7654
rect -9442 7688 -9376 7704
rect -9442 7654 -9426 7688
rect -9392 7654 -9376 7688
rect -9616 7616 -9586 7638
rect -9520 7616 -9490 7642
rect -9442 7638 -9376 7654
rect -9250 7688 -9184 7704
rect -9250 7654 -9234 7688
rect -9200 7654 -9184 7688
rect -9424 7616 -9394 7638
rect -9328 7616 -9298 7642
rect -9250 7638 -9184 7654
rect -9232 7616 -9202 7638
rect -9136 7616 -9106 7642
rect -10000 7190 -9970 7216
rect -9904 7194 -9874 7216
rect -9922 7178 -9856 7194
rect -9808 7190 -9778 7216
rect -9712 7194 -9682 7216
rect -9922 7144 -9906 7178
rect -9872 7144 -9856 7178
rect -9922 7128 -9856 7144
rect -9730 7178 -9664 7194
rect -9616 7190 -9586 7216
rect -9520 7194 -9490 7216
rect -9730 7144 -9714 7178
rect -9680 7144 -9664 7178
rect -9730 7128 -9664 7144
rect -9538 7178 -9472 7194
rect -9424 7190 -9394 7216
rect -9328 7194 -9298 7216
rect -9538 7144 -9522 7178
rect -9488 7144 -9472 7178
rect -9538 7128 -9472 7144
rect -9346 7178 -9280 7194
rect -9232 7190 -9202 7216
rect -9136 7194 -9106 7216
rect -9346 7144 -9330 7178
rect -9296 7144 -9280 7178
rect -9346 7128 -9280 7144
rect -9154 7178 -9088 7194
rect -9154 7144 -9138 7178
rect -9104 7144 -9088 7178
rect -9154 7128 -9088 7144
rect -9922 7070 -9856 7086
rect -9922 7036 -9906 7070
rect -9872 7036 -9856 7070
rect -10000 6998 -9970 7024
rect -9922 7020 -9856 7036
rect -9730 7070 -9664 7086
rect -9730 7036 -9714 7070
rect -9680 7036 -9664 7070
rect -9904 6998 -9874 7020
rect -9808 6998 -9778 7024
rect -9730 7020 -9664 7036
rect -9538 7070 -9472 7086
rect -9538 7036 -9522 7070
rect -9488 7036 -9472 7070
rect -9712 6998 -9682 7020
rect -9616 6998 -9586 7024
rect -9538 7020 -9472 7036
rect -9346 7070 -9280 7086
rect -9346 7036 -9330 7070
rect -9296 7036 -9280 7070
rect -9520 6998 -9490 7020
rect -9424 6998 -9394 7024
rect -9346 7020 -9280 7036
rect -9154 7070 -9088 7086
rect -9154 7036 -9138 7070
rect -9104 7036 -9088 7070
rect -9328 6998 -9298 7020
rect -9232 6998 -9202 7024
rect -9154 7020 -9088 7036
rect -9136 6998 -9106 7020
rect -10000 6576 -9970 6598
rect -10018 6560 -9952 6576
rect -9904 6572 -9874 6598
rect -9808 6576 -9778 6598
rect -10018 6526 -10002 6560
rect -9968 6526 -9952 6560
rect -10018 6510 -9952 6526
rect -9826 6560 -9760 6576
rect -9712 6572 -9682 6598
rect -9616 6576 -9586 6598
rect -9826 6526 -9810 6560
rect -9776 6526 -9760 6560
rect -9826 6510 -9760 6526
rect -9634 6560 -9568 6576
rect -9520 6572 -9490 6598
rect -9424 6576 -9394 6598
rect -9634 6526 -9618 6560
rect -9584 6526 -9568 6560
rect -9634 6510 -9568 6526
rect -9442 6560 -9376 6576
rect -9328 6572 -9298 6598
rect -9232 6576 -9202 6598
rect -9442 6526 -9426 6560
rect -9392 6526 -9376 6560
rect -9442 6510 -9376 6526
rect -9250 6560 -9184 6576
rect -9136 6572 -9106 6598
rect -9250 6526 -9234 6560
rect -9200 6526 -9184 6560
rect -9250 6510 -9184 6526
rect -8758 8168 -8670 8184
rect -8758 6600 -8742 8168
rect -8708 6600 -8670 8168
rect -8758 6584 -8670 6600
rect -8470 8168 -8382 8184
rect -8470 6600 -8432 8168
rect -8398 6600 -8382 8168
rect -8470 6584 -8382 6600
rect -9922 6226 -9856 6242
rect -9922 6192 -9906 6226
rect -9872 6192 -9856 6226
rect -10000 6154 -9970 6180
rect -9922 6176 -9856 6192
rect -9730 6226 -9664 6242
rect -9730 6192 -9714 6226
rect -9680 6192 -9664 6226
rect -9904 6154 -9874 6176
rect -9808 6154 -9778 6180
rect -9730 6176 -9664 6192
rect -9538 6226 -9472 6242
rect -9538 6192 -9522 6226
rect -9488 6192 -9472 6226
rect -9712 6154 -9682 6176
rect -9616 6154 -9586 6180
rect -9538 6176 -9472 6192
rect -9346 6226 -9280 6242
rect -9346 6192 -9330 6226
rect -9296 6192 -9280 6226
rect -9520 6154 -9490 6176
rect -9424 6154 -9394 6180
rect -9346 6176 -9280 6192
rect -9154 6226 -9088 6242
rect -9154 6192 -9138 6226
rect -9104 6192 -9088 6226
rect -9328 6154 -9298 6176
rect -9232 6154 -9202 6180
rect -9154 6176 -9088 6192
rect -9136 6154 -9106 6176
rect -10000 5732 -9970 5754
rect -10018 5716 -9952 5732
rect -9904 5728 -9874 5754
rect -9808 5732 -9778 5754
rect -10018 5682 -10002 5716
rect -9968 5682 -9952 5716
rect -10018 5666 -9952 5682
rect -9826 5716 -9760 5732
rect -9712 5728 -9682 5754
rect -9616 5732 -9586 5754
rect -9826 5682 -9810 5716
rect -9776 5682 -9760 5716
rect -9826 5666 -9760 5682
rect -9634 5716 -9568 5732
rect -9520 5728 -9490 5754
rect -9424 5732 -9394 5754
rect -9634 5682 -9618 5716
rect -9584 5682 -9568 5716
rect -9634 5666 -9568 5682
rect -9442 5716 -9376 5732
rect -9328 5728 -9298 5754
rect -9232 5732 -9202 5754
rect -9442 5682 -9426 5716
rect -9392 5682 -9376 5716
rect -9442 5666 -9376 5682
rect -9250 5716 -9184 5732
rect -9136 5728 -9106 5754
rect -9250 5682 -9234 5716
rect -9200 5682 -9184 5716
rect -9250 5666 -9184 5682
rect -10018 5608 -9952 5624
rect -10018 5574 -10002 5608
rect -9968 5574 -9952 5608
rect -10018 5558 -9952 5574
rect -9826 5608 -9760 5624
rect -9826 5574 -9810 5608
rect -9776 5574 -9760 5608
rect -10000 5536 -9970 5558
rect -9904 5536 -9874 5562
rect -9826 5558 -9760 5574
rect -9634 5608 -9568 5624
rect -9634 5574 -9618 5608
rect -9584 5574 -9568 5608
rect -9808 5536 -9778 5558
rect -9712 5536 -9682 5562
rect -9634 5558 -9568 5574
rect -9442 5608 -9376 5624
rect -9442 5574 -9426 5608
rect -9392 5574 -9376 5608
rect -9616 5536 -9586 5558
rect -9520 5536 -9490 5562
rect -9442 5558 -9376 5574
rect -9250 5608 -9184 5624
rect -9250 5574 -9234 5608
rect -9200 5574 -9184 5608
rect -9424 5536 -9394 5558
rect -9328 5536 -9298 5562
rect -9250 5558 -9184 5574
rect -9232 5536 -9202 5558
rect -9136 5536 -9106 5562
rect -10000 5110 -9970 5136
rect -9904 5114 -9874 5136
rect -9922 5098 -9856 5114
rect -9808 5110 -9778 5136
rect -9712 5114 -9682 5136
rect -9922 5064 -9906 5098
rect -9872 5064 -9856 5098
rect -9922 5048 -9856 5064
rect -9730 5098 -9664 5114
rect -9616 5110 -9586 5136
rect -9520 5114 -9490 5136
rect -9730 5064 -9714 5098
rect -9680 5064 -9664 5098
rect -9730 5048 -9664 5064
rect -9538 5098 -9472 5114
rect -9424 5110 -9394 5136
rect -9328 5114 -9298 5136
rect -9538 5064 -9522 5098
rect -9488 5064 -9472 5098
rect -9538 5048 -9472 5064
rect -9346 5098 -9280 5114
rect -9232 5110 -9202 5136
rect -9136 5114 -9106 5136
rect -9346 5064 -9330 5098
rect -9296 5064 -9280 5098
rect -9346 5048 -9280 5064
rect -9154 5098 -9088 5114
rect -9154 5064 -9138 5098
rect -9104 5064 -9088 5098
rect -9154 5048 -9088 5064
rect -9922 4990 -9856 5006
rect -9922 4956 -9906 4990
rect -9872 4956 -9856 4990
rect -10000 4918 -9970 4944
rect -9922 4940 -9856 4956
rect -9730 4990 -9664 5006
rect -9730 4956 -9714 4990
rect -9680 4956 -9664 4990
rect -9904 4918 -9874 4940
rect -9808 4918 -9778 4944
rect -9730 4940 -9664 4956
rect -9538 4990 -9472 5006
rect -9538 4956 -9522 4990
rect -9488 4956 -9472 4990
rect -9712 4918 -9682 4940
rect -9616 4918 -9586 4944
rect -9538 4940 -9472 4956
rect -9346 4990 -9280 5006
rect -9346 4956 -9330 4990
rect -9296 4956 -9280 4990
rect -9520 4918 -9490 4940
rect -9424 4918 -9394 4944
rect -9346 4940 -9280 4956
rect -9154 4990 -9088 5006
rect -9154 4956 -9138 4990
rect -9104 4956 -9088 4990
rect -9328 4918 -9298 4940
rect -9232 4918 -9202 4944
rect -9154 4940 -9088 4956
rect -9136 4918 -9106 4940
rect -10000 4496 -9970 4518
rect -10018 4480 -9952 4496
rect -9904 4492 -9874 4518
rect -9808 4496 -9778 4518
rect -10018 4446 -10002 4480
rect -9968 4446 -9952 4480
rect -10018 4430 -9952 4446
rect -9826 4480 -9760 4496
rect -9712 4492 -9682 4518
rect -9616 4496 -9586 4518
rect -9826 4446 -9810 4480
rect -9776 4446 -9760 4480
rect -9826 4430 -9760 4446
rect -9634 4480 -9568 4496
rect -9520 4492 -9490 4518
rect -9424 4496 -9394 4518
rect -9634 4446 -9618 4480
rect -9584 4446 -9568 4480
rect -9634 4430 -9568 4446
rect -9442 4480 -9376 4496
rect -9328 4492 -9298 4518
rect -9232 4496 -9202 4518
rect -9442 4446 -9426 4480
rect -9392 4446 -9376 4480
rect -9442 4430 -9376 4446
rect -9250 4480 -9184 4496
rect -9136 4492 -9106 4518
rect -9250 4446 -9234 4480
rect -9200 4446 -9184 4480
rect -9250 4430 -9184 4446
rect 1818 8802 1884 8818
rect 1818 8768 1834 8802
rect 1868 8768 1884 8802
rect 1740 8730 1770 8756
rect 1818 8752 1884 8768
rect 2010 8802 2076 8818
rect 2010 8768 2026 8802
rect 2060 8768 2076 8802
rect 1836 8730 1866 8752
rect 1932 8730 1962 8756
rect 2010 8752 2076 8768
rect 2202 8802 2268 8818
rect 2202 8768 2218 8802
rect 2252 8768 2268 8802
rect 2028 8730 2058 8752
rect 2124 8730 2154 8756
rect 2202 8752 2268 8768
rect 2394 8802 2460 8818
rect 2394 8768 2410 8802
rect 2444 8768 2460 8802
rect 2220 8730 2250 8752
rect 2316 8730 2346 8756
rect 2394 8752 2460 8768
rect 2586 8802 2652 8818
rect 2586 8768 2602 8802
rect 2636 8768 2652 8802
rect 2412 8730 2442 8752
rect 2508 8730 2538 8756
rect 2586 8752 2652 8768
rect 2778 8802 2844 8818
rect 2778 8768 2794 8802
rect 2828 8768 2844 8802
rect 2604 8730 2634 8752
rect 2700 8730 2730 8756
rect 2778 8752 2844 8768
rect 2970 8802 3036 8818
rect 2970 8768 2986 8802
rect 3020 8768 3036 8802
rect 2796 8730 2826 8752
rect 2892 8730 2922 8756
rect 2970 8752 3036 8768
rect 3162 8802 3228 8818
rect 3162 8768 3178 8802
rect 3212 8768 3228 8802
rect 2988 8730 3018 8752
rect 3084 8730 3114 8756
rect 3162 8752 3228 8768
rect 3354 8802 3420 8818
rect 3354 8768 3370 8802
rect 3404 8768 3420 8802
rect 3180 8730 3210 8752
rect 3276 8730 3306 8756
rect 3354 8752 3420 8768
rect 3546 8802 3612 8818
rect 3546 8768 3562 8802
rect 3596 8768 3612 8802
rect 3372 8730 3402 8752
rect 3468 8730 3498 8756
rect 3546 8752 3612 8768
rect 3564 8730 3594 8752
rect 1740 8308 1770 8330
rect 1722 8292 1788 8308
rect 1836 8304 1866 8330
rect 1932 8308 1962 8330
rect 1722 8258 1738 8292
rect 1772 8258 1788 8292
rect 1722 8242 1788 8258
rect 1914 8292 1980 8308
rect 2028 8304 2058 8330
rect 2124 8308 2154 8330
rect 1914 8258 1930 8292
rect 1964 8258 1980 8292
rect 1914 8242 1980 8258
rect 2106 8292 2172 8308
rect 2220 8304 2250 8330
rect 2316 8308 2346 8330
rect 2106 8258 2122 8292
rect 2156 8258 2172 8292
rect 2106 8242 2172 8258
rect 2298 8292 2364 8308
rect 2412 8304 2442 8330
rect 2508 8308 2538 8330
rect 2298 8258 2314 8292
rect 2348 8258 2364 8292
rect 2298 8242 2364 8258
rect 2490 8292 2556 8308
rect 2604 8304 2634 8330
rect 2700 8308 2730 8330
rect 2490 8258 2506 8292
rect 2540 8258 2556 8292
rect 2490 8242 2556 8258
rect 2682 8292 2748 8308
rect 2796 8304 2826 8330
rect 2892 8308 2922 8330
rect 2682 8258 2698 8292
rect 2732 8258 2748 8292
rect 2682 8242 2748 8258
rect 2874 8292 2940 8308
rect 2988 8304 3018 8330
rect 3084 8308 3114 8330
rect 2874 8258 2890 8292
rect 2924 8258 2940 8292
rect 2874 8242 2940 8258
rect 3066 8292 3132 8308
rect 3180 8304 3210 8330
rect 3276 8308 3306 8330
rect 3066 8258 3082 8292
rect 3116 8258 3132 8292
rect 3066 8242 3132 8258
rect 3258 8292 3324 8308
rect 3372 8304 3402 8330
rect 3468 8308 3498 8330
rect 3258 8258 3274 8292
rect 3308 8258 3324 8292
rect 3258 8242 3324 8258
rect 3450 8292 3516 8308
rect 3564 8304 3594 8330
rect 3450 8258 3466 8292
rect 3500 8258 3516 8292
rect 3450 8242 3516 8258
rect 1818 7982 1884 7998
rect 1818 7948 1834 7982
rect 1868 7948 1884 7982
rect 1740 7910 1770 7936
rect 1818 7932 1884 7948
rect 2010 7982 2076 7998
rect 2010 7948 2026 7982
rect 2060 7948 2076 7982
rect 1836 7910 1866 7932
rect 1932 7910 1962 7936
rect 2010 7932 2076 7948
rect 2202 7982 2268 7998
rect 2202 7948 2218 7982
rect 2252 7948 2268 7982
rect 2028 7910 2058 7932
rect 2124 7910 2154 7936
rect 2202 7932 2268 7948
rect 2394 7982 2460 7998
rect 2394 7948 2410 7982
rect 2444 7948 2460 7982
rect 2220 7910 2250 7932
rect 2316 7910 2346 7936
rect 2394 7932 2460 7948
rect 2586 7982 2652 7998
rect 2586 7948 2602 7982
rect 2636 7948 2652 7982
rect 2412 7910 2442 7932
rect 2508 7910 2538 7936
rect 2586 7932 2652 7948
rect 2778 7982 2844 7998
rect 2778 7948 2794 7982
rect 2828 7948 2844 7982
rect 2604 7910 2634 7932
rect 2700 7910 2730 7936
rect 2778 7932 2844 7948
rect 2970 7982 3036 7998
rect 2970 7948 2986 7982
rect 3020 7948 3036 7982
rect 2796 7910 2826 7932
rect 2892 7910 2922 7936
rect 2970 7932 3036 7948
rect 3162 7982 3228 7998
rect 3162 7948 3178 7982
rect 3212 7948 3228 7982
rect 2988 7910 3018 7932
rect 3084 7910 3114 7936
rect 3162 7932 3228 7948
rect 3354 7982 3420 7998
rect 3354 7948 3370 7982
rect 3404 7948 3420 7982
rect 3180 7910 3210 7932
rect 3276 7910 3306 7936
rect 3354 7932 3420 7948
rect 3546 7982 3612 7998
rect 3546 7948 3562 7982
rect 3596 7948 3612 7982
rect 3372 7910 3402 7932
rect 3468 7910 3498 7936
rect 3546 7932 3612 7948
rect 3564 7910 3594 7932
rect 1740 7488 1770 7510
rect 1722 7472 1788 7488
rect 1836 7484 1866 7510
rect 1932 7488 1962 7510
rect 1722 7438 1738 7472
rect 1772 7438 1788 7472
rect 1722 7422 1788 7438
rect 1914 7472 1980 7488
rect 2028 7484 2058 7510
rect 2124 7488 2154 7510
rect 1914 7438 1930 7472
rect 1964 7438 1980 7472
rect 1914 7422 1980 7438
rect 2106 7472 2172 7488
rect 2220 7484 2250 7510
rect 2316 7488 2346 7510
rect 2106 7438 2122 7472
rect 2156 7438 2172 7472
rect 2106 7422 2172 7438
rect 2298 7472 2364 7488
rect 2412 7484 2442 7510
rect 2508 7488 2538 7510
rect 2298 7438 2314 7472
rect 2348 7438 2364 7472
rect 2298 7422 2364 7438
rect 2490 7472 2556 7488
rect 2604 7484 2634 7510
rect 2700 7488 2730 7510
rect 2490 7438 2506 7472
rect 2540 7438 2556 7472
rect 2490 7422 2556 7438
rect 2682 7472 2748 7488
rect 2796 7484 2826 7510
rect 2892 7488 2922 7510
rect 2682 7438 2698 7472
rect 2732 7438 2748 7472
rect 2682 7422 2748 7438
rect 2874 7472 2940 7488
rect 2988 7484 3018 7510
rect 3084 7488 3114 7510
rect 2874 7438 2890 7472
rect 2924 7438 2940 7472
rect 2874 7422 2940 7438
rect 3066 7472 3132 7488
rect 3180 7484 3210 7510
rect 3276 7488 3306 7510
rect 3066 7438 3082 7472
rect 3116 7438 3132 7472
rect 3066 7422 3132 7438
rect 3258 7472 3324 7488
rect 3372 7484 3402 7510
rect 3468 7488 3498 7510
rect 3258 7438 3274 7472
rect 3308 7438 3324 7472
rect 3258 7422 3324 7438
rect 3450 7472 3516 7488
rect 3564 7484 3594 7510
rect 3450 7438 3466 7472
rect 3500 7438 3516 7472
rect 3450 7422 3516 7438
rect 1818 7162 1884 7178
rect 1818 7128 1834 7162
rect 1868 7128 1884 7162
rect 1740 7090 1770 7116
rect 1818 7112 1884 7128
rect 2010 7162 2076 7178
rect 2010 7128 2026 7162
rect 2060 7128 2076 7162
rect 1836 7090 1866 7112
rect 1932 7090 1962 7116
rect 2010 7112 2076 7128
rect 2202 7162 2268 7178
rect 2202 7128 2218 7162
rect 2252 7128 2268 7162
rect 2028 7090 2058 7112
rect 2124 7090 2154 7116
rect 2202 7112 2268 7128
rect 2394 7162 2460 7178
rect 2394 7128 2410 7162
rect 2444 7128 2460 7162
rect 2220 7090 2250 7112
rect 2316 7090 2346 7116
rect 2394 7112 2460 7128
rect 2586 7162 2652 7178
rect 2586 7128 2602 7162
rect 2636 7128 2652 7162
rect 2412 7090 2442 7112
rect 2508 7090 2538 7116
rect 2586 7112 2652 7128
rect 2778 7162 2844 7178
rect 2778 7128 2794 7162
rect 2828 7128 2844 7162
rect 2604 7090 2634 7112
rect 2700 7090 2730 7116
rect 2778 7112 2844 7128
rect 2970 7162 3036 7178
rect 2970 7128 2986 7162
rect 3020 7128 3036 7162
rect 2796 7090 2826 7112
rect 2892 7090 2922 7116
rect 2970 7112 3036 7128
rect 3162 7162 3228 7178
rect 3162 7128 3178 7162
rect 3212 7128 3228 7162
rect 2988 7090 3018 7112
rect 3084 7090 3114 7116
rect 3162 7112 3228 7128
rect 3354 7162 3420 7178
rect 3354 7128 3370 7162
rect 3404 7128 3420 7162
rect 3180 7090 3210 7112
rect 3276 7090 3306 7116
rect 3354 7112 3420 7128
rect 3546 7162 3612 7178
rect 3546 7128 3562 7162
rect 3596 7128 3612 7162
rect 3372 7090 3402 7112
rect 3468 7090 3498 7116
rect 3546 7112 3612 7128
rect 3564 7090 3594 7112
rect 1740 6668 1770 6690
rect 1722 6652 1788 6668
rect 1836 6664 1866 6690
rect 1932 6668 1962 6690
rect 1722 6618 1738 6652
rect 1772 6618 1788 6652
rect 1722 6602 1788 6618
rect 1914 6652 1980 6668
rect 2028 6664 2058 6690
rect 2124 6668 2154 6690
rect 1914 6618 1930 6652
rect 1964 6618 1980 6652
rect 1914 6602 1980 6618
rect 2106 6652 2172 6668
rect 2220 6664 2250 6690
rect 2316 6668 2346 6690
rect 2106 6618 2122 6652
rect 2156 6618 2172 6652
rect 2106 6602 2172 6618
rect 2298 6652 2364 6668
rect 2412 6664 2442 6690
rect 2508 6668 2538 6690
rect 2298 6618 2314 6652
rect 2348 6618 2364 6652
rect 2298 6602 2364 6618
rect 2490 6652 2556 6668
rect 2604 6664 2634 6690
rect 2700 6668 2730 6690
rect 2490 6618 2506 6652
rect 2540 6618 2556 6652
rect 2490 6602 2556 6618
rect 2682 6652 2748 6668
rect 2796 6664 2826 6690
rect 2892 6668 2922 6690
rect 2682 6618 2698 6652
rect 2732 6618 2748 6652
rect 2682 6602 2748 6618
rect 2874 6652 2940 6668
rect 2988 6664 3018 6690
rect 3084 6668 3114 6690
rect 2874 6618 2890 6652
rect 2924 6618 2940 6652
rect 2874 6602 2940 6618
rect 3066 6652 3132 6668
rect 3180 6664 3210 6690
rect 3276 6668 3306 6690
rect 3066 6618 3082 6652
rect 3116 6618 3132 6652
rect 3066 6602 3132 6618
rect 3258 6652 3324 6668
rect 3372 6664 3402 6690
rect 3468 6668 3498 6690
rect 3258 6618 3274 6652
rect 3308 6618 3324 6652
rect 3258 6602 3324 6618
rect 3450 6652 3516 6668
rect 3564 6664 3594 6690
rect 3450 6618 3466 6652
rect 3500 6618 3516 6652
rect 3450 6602 3516 6618
rect 5158 10364 5224 10380
rect 5158 10330 5174 10364
rect 5208 10330 5224 10364
rect 5158 10314 5224 10330
rect 5350 10364 5416 10380
rect 5350 10330 5366 10364
rect 5400 10330 5416 10364
rect 5350 10314 5416 10330
rect 5542 10364 5608 10380
rect 5542 10330 5558 10364
rect 5592 10330 5608 10364
rect 5542 10314 5608 10330
rect 5734 10364 5800 10380
rect 5734 10330 5750 10364
rect 5784 10330 5800 10364
rect 5734 10314 5800 10330
rect 5926 10364 5992 10380
rect 5926 10330 5942 10364
rect 5976 10330 5992 10364
rect 5926 10314 5992 10330
rect 6118 10364 6184 10380
rect 6118 10330 6134 10364
rect 6168 10330 6184 10364
rect 6118 10314 6184 10330
rect 6310 10364 6376 10380
rect 6310 10330 6326 10364
rect 6360 10330 6376 10364
rect 6310 10314 6376 10330
rect 6502 10364 6568 10380
rect 6502 10330 6518 10364
rect 6552 10330 6568 10364
rect 6502 10314 6568 10330
rect 6694 10364 6760 10380
rect 6694 10330 6710 10364
rect 6744 10330 6760 10364
rect 6694 10314 6760 10330
rect 6886 10364 6952 10380
rect 6886 10330 6902 10364
rect 6936 10330 6952 10364
rect 6886 10314 6952 10330
rect 5176 10283 5206 10314
rect 5272 10283 5302 10309
rect 5368 10283 5398 10314
rect 5464 10283 5494 10309
rect 5560 10283 5590 10314
rect 5656 10283 5686 10309
rect 5752 10283 5782 10314
rect 5848 10283 5878 10309
rect 5944 10283 5974 10314
rect 6040 10283 6070 10309
rect 6136 10283 6166 10314
rect 6232 10283 6262 10309
rect 6328 10283 6358 10314
rect 6424 10283 6454 10309
rect 6520 10283 6550 10314
rect 6616 10283 6646 10309
rect 6712 10283 6742 10314
rect 6808 10283 6838 10309
rect 6904 10283 6934 10314
rect 7000 10283 7030 10309
rect 5176 9857 5206 9883
rect 5272 9852 5302 9883
rect 5368 9857 5398 9883
rect 5464 9852 5494 9883
rect 5560 9857 5590 9883
rect 5656 9852 5686 9883
rect 5752 9857 5782 9883
rect 5848 9852 5878 9883
rect 5944 9857 5974 9883
rect 6040 9852 6070 9883
rect 6136 9857 6166 9883
rect 6232 9852 6262 9883
rect 6328 9857 6358 9883
rect 6424 9852 6454 9883
rect 6520 9857 6550 9883
rect 6616 9852 6646 9883
rect 6712 9857 6742 9883
rect 6808 9852 6838 9883
rect 6904 9857 6934 9883
rect 7000 9852 7030 9883
rect 5254 9836 5320 9852
rect 5254 9802 5270 9836
rect 5304 9802 5320 9836
rect 5254 9786 5320 9802
rect 5446 9836 5512 9852
rect 5446 9802 5462 9836
rect 5496 9802 5512 9836
rect 5446 9786 5512 9802
rect 5638 9836 5704 9852
rect 5638 9802 5654 9836
rect 5688 9802 5704 9836
rect 5638 9786 5704 9802
rect 5830 9836 5896 9852
rect 5830 9802 5846 9836
rect 5880 9802 5896 9836
rect 5830 9786 5896 9802
rect 6022 9836 6088 9852
rect 6022 9802 6038 9836
rect 6072 9802 6088 9836
rect 6022 9786 6088 9802
rect 6214 9836 6280 9852
rect 6214 9802 6230 9836
rect 6264 9802 6280 9836
rect 6214 9786 6280 9802
rect 6406 9836 6472 9852
rect 6406 9802 6422 9836
rect 6456 9802 6472 9836
rect 6406 9786 6472 9802
rect 6598 9836 6664 9852
rect 6598 9802 6614 9836
rect 6648 9802 6664 9836
rect 6598 9786 6664 9802
rect 6790 9836 6856 9852
rect 6790 9802 6806 9836
rect 6840 9802 6856 9836
rect 6790 9786 6856 9802
rect 6982 9836 7048 9852
rect 6982 9802 6998 9836
rect 7032 9802 7048 9836
rect 6982 9786 7048 9802
rect 5254 9728 5320 9744
rect 5254 9694 5270 9728
rect 5304 9694 5320 9728
rect 5254 9678 5320 9694
rect 5446 9728 5512 9744
rect 5446 9694 5462 9728
rect 5496 9694 5512 9728
rect 5446 9678 5512 9694
rect 5638 9728 5704 9744
rect 5638 9694 5654 9728
rect 5688 9694 5704 9728
rect 5638 9678 5704 9694
rect 5830 9728 5896 9744
rect 5830 9694 5846 9728
rect 5880 9694 5896 9728
rect 5830 9678 5896 9694
rect 6022 9728 6088 9744
rect 6022 9694 6038 9728
rect 6072 9694 6088 9728
rect 6022 9678 6088 9694
rect 6214 9728 6280 9744
rect 6214 9694 6230 9728
rect 6264 9694 6280 9728
rect 6214 9678 6280 9694
rect 6406 9728 6472 9744
rect 6406 9694 6422 9728
rect 6456 9694 6472 9728
rect 6406 9678 6472 9694
rect 6598 9728 6664 9744
rect 6598 9694 6614 9728
rect 6648 9694 6664 9728
rect 6598 9678 6664 9694
rect 6790 9728 6856 9744
rect 6790 9694 6806 9728
rect 6840 9694 6856 9728
rect 6790 9678 6856 9694
rect 6982 9728 7048 9744
rect 6982 9694 6998 9728
rect 7032 9694 7048 9728
rect 6982 9678 7048 9694
rect 5176 9647 5206 9673
rect 5272 9647 5302 9678
rect 5368 9647 5398 9673
rect 5464 9647 5494 9678
rect 5560 9647 5590 9673
rect 5656 9647 5686 9678
rect 5752 9647 5782 9673
rect 5848 9647 5878 9678
rect 5944 9647 5974 9673
rect 6040 9647 6070 9678
rect 6136 9647 6166 9673
rect 6232 9647 6262 9678
rect 6328 9647 6358 9673
rect 6424 9647 6454 9678
rect 6520 9647 6550 9673
rect 6616 9647 6646 9678
rect 6712 9647 6742 9673
rect 6808 9647 6838 9678
rect 6904 9647 6934 9673
rect 7000 9647 7030 9678
rect 5176 9216 5206 9247
rect 5272 9221 5302 9247
rect 5368 9216 5398 9247
rect 5464 9221 5494 9247
rect 5560 9216 5590 9247
rect 5656 9221 5686 9247
rect 5752 9216 5782 9247
rect 5848 9221 5878 9247
rect 5944 9216 5974 9247
rect 6040 9221 6070 9247
rect 6136 9216 6166 9247
rect 6232 9221 6262 9247
rect 6328 9216 6358 9247
rect 6424 9221 6454 9247
rect 6520 9216 6550 9247
rect 6616 9221 6646 9247
rect 6712 9216 6742 9247
rect 6808 9221 6838 9247
rect 6904 9216 6934 9247
rect 7000 9221 7030 9247
rect 5158 9200 5224 9216
rect 5158 9166 5174 9200
rect 5208 9166 5224 9200
rect 5158 9150 5224 9166
rect 5350 9200 5416 9216
rect 5350 9166 5366 9200
rect 5400 9166 5416 9200
rect 5350 9150 5416 9166
rect 5542 9200 5608 9216
rect 5542 9166 5558 9200
rect 5592 9166 5608 9200
rect 5542 9150 5608 9166
rect 5734 9200 5800 9216
rect 5734 9166 5750 9200
rect 5784 9166 5800 9200
rect 5734 9150 5800 9166
rect 5926 9200 5992 9216
rect 5926 9166 5942 9200
rect 5976 9166 5992 9200
rect 5926 9150 5992 9166
rect 6118 9200 6184 9216
rect 6118 9166 6134 9200
rect 6168 9166 6184 9200
rect 6118 9150 6184 9166
rect 6310 9200 6376 9216
rect 6310 9166 6326 9200
rect 6360 9166 6376 9200
rect 6310 9150 6376 9166
rect 6502 9200 6568 9216
rect 6502 9166 6518 9200
rect 6552 9166 6568 9200
rect 6502 9150 6568 9166
rect 6694 9200 6760 9216
rect 6694 9166 6710 9200
rect 6744 9166 6760 9200
rect 6694 9150 6760 9166
rect 6886 9200 6952 9216
rect 6886 9166 6902 9200
rect 6936 9166 6952 9200
rect 6886 9150 6952 9166
rect 5158 8768 5224 8784
rect 5158 8734 5174 8768
rect 5208 8734 5224 8768
rect 5158 8718 5224 8734
rect 5350 8768 5416 8784
rect 5350 8734 5366 8768
rect 5400 8734 5416 8768
rect 5176 8696 5206 8718
rect 5272 8696 5302 8722
rect 5350 8718 5416 8734
rect 5542 8768 5608 8784
rect 5542 8734 5558 8768
rect 5592 8734 5608 8768
rect 5368 8696 5398 8718
rect 5464 8696 5494 8722
rect 5542 8718 5608 8734
rect 5734 8768 5800 8784
rect 5734 8734 5750 8768
rect 5784 8734 5800 8768
rect 5560 8696 5590 8718
rect 5656 8696 5686 8722
rect 5734 8718 5800 8734
rect 5926 8768 5992 8784
rect 5926 8734 5942 8768
rect 5976 8734 5992 8768
rect 5752 8696 5782 8718
rect 5848 8696 5878 8722
rect 5926 8718 5992 8734
rect 6118 8768 6184 8784
rect 6118 8734 6134 8768
rect 6168 8734 6184 8768
rect 5944 8696 5974 8718
rect 6040 8696 6070 8722
rect 6118 8718 6184 8734
rect 6310 8768 6376 8784
rect 6310 8734 6326 8768
rect 6360 8734 6376 8768
rect 6136 8696 6166 8718
rect 6232 8696 6262 8722
rect 6310 8718 6376 8734
rect 6502 8768 6568 8784
rect 6502 8734 6518 8768
rect 6552 8734 6568 8768
rect 6328 8696 6358 8718
rect 6424 8696 6454 8722
rect 6502 8718 6568 8734
rect 6694 8768 6760 8784
rect 6694 8734 6710 8768
rect 6744 8734 6760 8768
rect 6520 8696 6550 8718
rect 6616 8696 6646 8722
rect 6694 8718 6760 8734
rect 6886 8768 6952 8784
rect 6886 8734 6902 8768
rect 6936 8734 6952 8768
rect 6712 8696 6742 8718
rect 6808 8696 6838 8722
rect 6886 8718 6952 8734
rect 6904 8696 6934 8718
rect 7000 8696 7030 8722
rect 5176 8270 5206 8296
rect 5272 8274 5302 8296
rect 5254 8258 5320 8274
rect 5368 8270 5398 8296
rect 5464 8274 5494 8296
rect 5254 8224 5270 8258
rect 5304 8224 5320 8258
rect 5254 8208 5320 8224
rect 5446 8258 5512 8274
rect 5560 8270 5590 8296
rect 5656 8274 5686 8296
rect 5446 8224 5462 8258
rect 5496 8224 5512 8258
rect 5446 8208 5512 8224
rect 5638 8258 5704 8274
rect 5752 8270 5782 8296
rect 5848 8274 5878 8296
rect 5638 8224 5654 8258
rect 5688 8224 5704 8258
rect 5638 8208 5704 8224
rect 5830 8258 5896 8274
rect 5944 8270 5974 8296
rect 6040 8274 6070 8296
rect 5830 8224 5846 8258
rect 5880 8224 5896 8258
rect 5830 8208 5896 8224
rect 6022 8258 6088 8274
rect 6136 8270 6166 8296
rect 6232 8274 6262 8296
rect 6022 8224 6038 8258
rect 6072 8224 6088 8258
rect 6022 8208 6088 8224
rect 6214 8258 6280 8274
rect 6328 8270 6358 8296
rect 6424 8274 6454 8296
rect 6214 8224 6230 8258
rect 6264 8224 6280 8258
rect 6214 8208 6280 8224
rect 6406 8258 6472 8274
rect 6520 8270 6550 8296
rect 6616 8274 6646 8296
rect 6406 8224 6422 8258
rect 6456 8224 6472 8258
rect 6406 8208 6472 8224
rect 6598 8258 6664 8274
rect 6712 8270 6742 8296
rect 6808 8274 6838 8296
rect 6598 8224 6614 8258
rect 6648 8224 6664 8258
rect 6598 8208 6664 8224
rect 6790 8258 6856 8274
rect 6904 8270 6934 8296
rect 7000 8274 7030 8296
rect 6790 8224 6806 8258
rect 6840 8224 6856 8258
rect 6790 8208 6856 8224
rect 6982 8258 7048 8274
rect 6982 8224 6998 8258
rect 7032 8224 7048 8258
rect 6982 8208 7048 8224
rect 5254 8150 5320 8166
rect 5254 8116 5270 8150
rect 5304 8116 5320 8150
rect 5176 8078 5206 8104
rect 5254 8100 5320 8116
rect 5446 8150 5512 8166
rect 5446 8116 5462 8150
rect 5496 8116 5512 8150
rect 5272 8078 5302 8100
rect 5368 8078 5398 8104
rect 5446 8100 5512 8116
rect 5638 8150 5704 8166
rect 5638 8116 5654 8150
rect 5688 8116 5704 8150
rect 5464 8078 5494 8100
rect 5560 8078 5590 8104
rect 5638 8100 5704 8116
rect 5830 8150 5896 8166
rect 5830 8116 5846 8150
rect 5880 8116 5896 8150
rect 5656 8078 5686 8100
rect 5752 8078 5782 8104
rect 5830 8100 5896 8116
rect 6022 8150 6088 8166
rect 6022 8116 6038 8150
rect 6072 8116 6088 8150
rect 5848 8078 5878 8100
rect 5944 8078 5974 8104
rect 6022 8100 6088 8116
rect 6214 8150 6280 8166
rect 6214 8116 6230 8150
rect 6264 8116 6280 8150
rect 6040 8078 6070 8100
rect 6136 8078 6166 8104
rect 6214 8100 6280 8116
rect 6406 8150 6472 8166
rect 6406 8116 6422 8150
rect 6456 8116 6472 8150
rect 6232 8078 6262 8100
rect 6328 8078 6358 8104
rect 6406 8100 6472 8116
rect 6598 8150 6664 8166
rect 6598 8116 6614 8150
rect 6648 8116 6664 8150
rect 6424 8078 6454 8100
rect 6520 8078 6550 8104
rect 6598 8100 6664 8116
rect 6790 8150 6856 8166
rect 6790 8116 6806 8150
rect 6840 8116 6856 8150
rect 6616 8078 6646 8100
rect 6712 8078 6742 8104
rect 6790 8100 6856 8116
rect 6982 8150 7048 8166
rect 6982 8116 6998 8150
rect 7032 8116 7048 8150
rect 6808 8078 6838 8100
rect 6904 8078 6934 8104
rect 6982 8100 7048 8116
rect 7000 8078 7030 8100
rect 5176 7656 5206 7678
rect 5158 7640 5224 7656
rect 5272 7652 5302 7678
rect 5368 7656 5398 7678
rect 5158 7606 5174 7640
rect 5208 7606 5224 7640
rect 5158 7590 5224 7606
rect 5350 7640 5416 7656
rect 5464 7652 5494 7678
rect 5560 7656 5590 7678
rect 5350 7606 5366 7640
rect 5400 7606 5416 7640
rect 5350 7590 5416 7606
rect 5542 7640 5608 7656
rect 5656 7652 5686 7678
rect 5752 7656 5782 7678
rect 5542 7606 5558 7640
rect 5592 7606 5608 7640
rect 5542 7590 5608 7606
rect 5734 7640 5800 7656
rect 5848 7652 5878 7678
rect 5944 7656 5974 7678
rect 5734 7606 5750 7640
rect 5784 7606 5800 7640
rect 5734 7590 5800 7606
rect 5926 7640 5992 7656
rect 6040 7652 6070 7678
rect 6136 7656 6166 7678
rect 5926 7606 5942 7640
rect 5976 7606 5992 7640
rect 5926 7590 5992 7606
rect 6118 7640 6184 7656
rect 6232 7652 6262 7678
rect 6328 7656 6358 7678
rect 6118 7606 6134 7640
rect 6168 7606 6184 7640
rect 6118 7590 6184 7606
rect 6310 7640 6376 7656
rect 6424 7652 6454 7678
rect 6520 7656 6550 7678
rect 6310 7606 6326 7640
rect 6360 7606 6376 7640
rect 6310 7590 6376 7606
rect 6502 7640 6568 7656
rect 6616 7652 6646 7678
rect 6712 7656 6742 7678
rect 6502 7606 6518 7640
rect 6552 7606 6568 7640
rect 6502 7590 6568 7606
rect 6694 7640 6760 7656
rect 6808 7652 6838 7678
rect 6904 7656 6934 7678
rect 6694 7606 6710 7640
rect 6744 7606 6760 7640
rect 6694 7590 6760 7606
rect 6886 7640 6952 7656
rect 7000 7652 7030 7678
rect 6886 7606 6902 7640
rect 6936 7606 6952 7640
rect 6886 7590 6952 7606
rect -10004 4080 -9804 4096
rect -10004 4046 -9988 4080
rect -9820 4046 -9804 4080
rect -10004 4008 -9804 4046
rect -9746 4080 -9546 4096
rect -9746 4046 -9730 4080
rect -9562 4046 -9546 4080
rect -9746 4008 -9546 4046
rect -9488 4080 -9288 4096
rect -9488 4046 -9472 4080
rect -9304 4046 -9288 4080
rect -9488 4008 -9288 4046
rect -9230 4080 -9030 4096
rect -9230 4046 -9214 4080
rect -9046 4046 -9030 4080
rect -9230 4008 -9030 4046
rect -8972 4080 -8772 4096
rect -8972 4046 -8956 4080
rect -8788 4046 -8772 4080
rect -8972 4008 -8772 4046
rect -10004 3570 -9804 3608
rect -10004 3536 -9988 3570
rect -9820 3536 -9804 3570
rect -10004 3520 -9804 3536
rect -9746 3570 -9546 3608
rect -9746 3536 -9730 3570
rect -9562 3536 -9546 3570
rect -9746 3520 -9546 3536
rect -9488 3570 -9288 3608
rect -9488 3536 -9472 3570
rect -9304 3536 -9288 3570
rect -9488 3520 -9288 3536
rect -9230 3570 -9030 3608
rect -9230 3536 -9214 3570
rect -9046 3536 -9030 3570
rect -9230 3520 -9030 3536
rect -8972 3570 -8772 3608
rect -8972 3536 -8956 3570
rect -8788 3536 -8772 3570
rect -8972 3520 -8772 3536
rect -10004 3462 -9804 3478
rect -10004 3428 -9988 3462
rect -9820 3428 -9804 3462
rect -10004 3390 -9804 3428
rect -9746 3462 -9546 3478
rect -9746 3428 -9730 3462
rect -9562 3428 -9546 3462
rect -9746 3390 -9546 3428
rect -9488 3462 -9288 3478
rect -9488 3428 -9472 3462
rect -9304 3428 -9288 3462
rect -9488 3390 -9288 3428
rect -9230 3462 -9030 3478
rect -9230 3428 -9214 3462
rect -9046 3428 -9030 3462
rect -9230 3390 -9030 3428
rect -8972 3462 -8772 3478
rect -8972 3428 -8956 3462
rect -8788 3428 -8772 3462
rect -8972 3390 -8772 3428
rect -10004 2952 -9804 2990
rect -10004 2918 -9988 2952
rect -9820 2918 -9804 2952
rect -10004 2902 -9804 2918
rect -9746 2952 -9546 2990
rect -9746 2918 -9730 2952
rect -9562 2918 -9546 2952
rect -9746 2902 -9546 2918
rect -9488 2952 -9288 2990
rect -9488 2918 -9472 2952
rect -9304 2918 -9288 2952
rect -9488 2902 -9288 2918
rect -9230 2952 -9030 2990
rect -9230 2918 -9214 2952
rect -9046 2918 -9030 2952
rect -9230 2902 -9030 2918
rect -8972 2952 -8772 2990
rect -8972 2918 -8956 2952
rect -8788 2918 -8772 2952
rect -8972 2902 -8772 2918
rect -10004 2844 -9804 2860
rect -10004 2810 -9988 2844
rect -9820 2810 -9804 2844
rect -10004 2772 -9804 2810
rect -9746 2844 -9546 2860
rect -9746 2810 -9730 2844
rect -9562 2810 -9546 2844
rect -9746 2772 -9546 2810
rect -9488 2844 -9288 2860
rect -9488 2810 -9472 2844
rect -9304 2810 -9288 2844
rect -9488 2772 -9288 2810
rect -9230 2844 -9030 2860
rect -9230 2810 -9214 2844
rect -9046 2810 -9030 2844
rect -9230 2772 -9030 2810
rect -8972 2844 -8772 2860
rect -8972 2810 -8956 2844
rect -8788 2810 -8772 2844
rect -8972 2772 -8772 2810
rect -10004 2334 -9804 2372
rect -10004 2300 -9988 2334
rect -9820 2300 -9804 2334
rect -10004 2284 -9804 2300
rect -9746 2334 -9546 2372
rect -9746 2300 -9730 2334
rect -9562 2300 -9546 2334
rect -9746 2284 -9546 2300
rect -9488 2334 -9288 2372
rect -9488 2300 -9472 2334
rect -9304 2300 -9288 2334
rect -9488 2284 -9288 2300
rect -9230 2334 -9030 2372
rect -9230 2300 -9214 2334
rect -9046 2300 -9030 2334
rect -9230 2284 -9030 2300
rect -8972 2334 -8772 2372
rect -8972 2300 -8956 2334
rect -8788 2300 -8772 2334
rect -8972 2284 -8772 2300
rect -10004 2226 -9804 2242
rect -10004 2192 -9988 2226
rect -9820 2192 -9804 2226
rect -10004 2154 -9804 2192
rect -9746 2226 -9546 2242
rect -9746 2192 -9730 2226
rect -9562 2192 -9546 2226
rect -9746 2154 -9546 2192
rect -9488 2226 -9288 2242
rect -9488 2192 -9472 2226
rect -9304 2192 -9288 2226
rect -9488 2154 -9288 2192
rect -9230 2226 -9030 2242
rect -9230 2192 -9214 2226
rect -9046 2192 -9030 2226
rect -9230 2154 -9030 2192
rect -8972 2226 -8772 2242
rect -8972 2192 -8956 2226
rect -8788 2192 -8772 2226
rect -8972 2154 -8772 2192
rect -10004 1716 -9804 1754
rect -10004 1682 -9988 1716
rect -9820 1682 -9804 1716
rect -10004 1666 -9804 1682
rect -9746 1716 -9546 1754
rect -9746 1682 -9730 1716
rect -9562 1682 -9546 1716
rect -9746 1666 -9546 1682
rect -9488 1716 -9288 1754
rect -9488 1682 -9472 1716
rect -9304 1682 -9288 1716
rect -9488 1666 -9288 1682
rect -9230 1716 -9030 1754
rect -9230 1682 -9214 1716
rect -9046 1682 -9030 1716
rect -9230 1666 -9030 1682
rect -8972 1716 -8772 1754
rect -8972 1682 -8956 1716
rect -8788 1682 -8772 1716
rect -8972 1666 -8772 1682
rect -10004 1608 -9804 1624
rect -10004 1574 -9988 1608
rect -9820 1574 -9804 1608
rect -10004 1536 -9804 1574
rect -9746 1608 -9546 1624
rect -9746 1574 -9730 1608
rect -9562 1574 -9546 1608
rect -9746 1536 -9546 1574
rect -9488 1608 -9288 1624
rect -9488 1574 -9472 1608
rect -9304 1574 -9288 1608
rect -9488 1536 -9288 1574
rect -9230 1608 -9030 1624
rect -9230 1574 -9214 1608
rect -9046 1574 -9030 1608
rect -9230 1536 -9030 1574
rect -8972 1608 -8772 1624
rect -8972 1574 -8956 1608
rect -8788 1574 -8772 1608
rect -8972 1536 -8772 1574
rect -10004 1098 -9804 1136
rect -10004 1064 -9988 1098
rect -9820 1064 -9804 1098
rect -10004 1048 -9804 1064
rect -9746 1098 -9546 1136
rect -9746 1064 -9730 1098
rect -9562 1064 -9546 1098
rect -9746 1048 -9546 1064
rect -9488 1098 -9288 1136
rect -9488 1064 -9472 1098
rect -9304 1064 -9288 1098
rect -9488 1048 -9288 1064
rect -9230 1098 -9030 1136
rect -9230 1064 -9214 1098
rect -9046 1064 -9030 1098
rect -9230 1048 -9030 1064
rect -8972 1098 -8772 1136
rect -8972 1064 -8956 1098
rect -8788 1064 -8772 1098
rect -8972 1048 -8772 1064
rect -10004 990 -9804 1006
rect -10004 956 -9988 990
rect -9820 956 -9804 990
rect -10004 918 -9804 956
rect -9746 990 -9546 1006
rect -9746 956 -9730 990
rect -9562 956 -9546 990
rect -9746 918 -9546 956
rect -9488 990 -9288 1006
rect -9488 956 -9472 990
rect -9304 956 -9288 990
rect -9488 918 -9288 956
rect -9230 990 -9030 1006
rect -9230 956 -9214 990
rect -9046 956 -9030 990
rect -9230 918 -9030 956
rect -8972 990 -8772 1006
rect -8972 956 -8956 990
rect -8788 956 -8772 990
rect -8972 918 -8772 956
rect -10004 480 -9804 518
rect -10004 446 -9988 480
rect -9820 446 -9804 480
rect -10004 430 -9804 446
rect -9746 480 -9546 518
rect -9746 446 -9730 480
rect -9562 446 -9546 480
rect -9746 430 -9546 446
rect -9488 480 -9288 518
rect -9488 446 -9472 480
rect -9304 446 -9288 480
rect -9488 430 -9288 446
rect -9230 480 -9030 518
rect -9230 446 -9214 480
rect -9046 446 -9030 480
rect -9230 430 -9030 446
rect -8972 480 -8772 518
rect -8972 446 -8956 480
rect -8788 446 -8772 480
rect -8972 430 -8772 446
rect 354 5946 420 5962
rect 354 5912 370 5946
rect 404 5912 420 5946
rect 276 5874 306 5900
rect 354 5896 420 5912
rect 546 5946 612 5962
rect 546 5912 562 5946
rect 596 5912 612 5946
rect 372 5874 402 5896
rect 468 5874 498 5900
rect 546 5896 612 5912
rect 738 5946 804 5962
rect 738 5912 754 5946
rect 788 5912 804 5946
rect 564 5874 594 5896
rect 660 5874 690 5900
rect 738 5896 804 5912
rect 930 5946 996 5962
rect 930 5912 946 5946
rect 980 5912 996 5946
rect 756 5874 786 5896
rect 852 5874 882 5900
rect 930 5896 996 5912
rect 1122 5946 1188 5962
rect 1122 5912 1138 5946
rect 1172 5912 1188 5946
rect 948 5874 978 5896
rect 1044 5874 1074 5900
rect 1122 5896 1188 5912
rect 1140 5874 1170 5896
rect 276 5452 306 5474
rect 258 5436 324 5452
rect 372 5448 402 5474
rect 468 5452 498 5474
rect 258 5402 274 5436
rect 308 5402 324 5436
rect 258 5386 324 5402
rect 450 5436 516 5452
rect 564 5448 594 5474
rect 660 5452 690 5474
rect 450 5402 466 5436
rect 500 5402 516 5436
rect 450 5386 516 5402
rect 642 5436 708 5452
rect 756 5448 786 5474
rect 852 5452 882 5474
rect 642 5402 658 5436
rect 692 5402 708 5436
rect 642 5386 708 5402
rect 834 5436 900 5452
rect 948 5448 978 5474
rect 1044 5452 1074 5474
rect 834 5402 850 5436
rect 884 5402 900 5436
rect 834 5386 900 5402
rect 1026 5436 1092 5452
rect 1140 5448 1170 5474
rect 1026 5402 1042 5436
rect 1076 5402 1092 5436
rect 1026 5386 1092 5402
rect 258 5328 324 5344
rect 258 5294 274 5328
rect 308 5294 324 5328
rect 258 5278 324 5294
rect 450 5328 516 5344
rect 450 5294 466 5328
rect 500 5294 516 5328
rect 276 5256 306 5278
rect 372 5256 402 5282
rect 450 5278 516 5294
rect 642 5328 708 5344
rect 642 5294 658 5328
rect 692 5294 708 5328
rect 468 5256 498 5278
rect 564 5256 594 5282
rect 642 5278 708 5294
rect 834 5328 900 5344
rect 834 5294 850 5328
rect 884 5294 900 5328
rect 660 5256 690 5278
rect 756 5256 786 5282
rect 834 5278 900 5294
rect 1026 5328 1092 5344
rect 1026 5294 1042 5328
rect 1076 5294 1092 5328
rect 852 5256 882 5278
rect 948 5256 978 5282
rect 1026 5278 1092 5294
rect 1044 5256 1074 5278
rect 1140 5256 1170 5282
rect 276 4830 306 4856
rect 372 4834 402 4856
rect 354 4818 420 4834
rect 468 4830 498 4856
rect 564 4834 594 4856
rect 354 4784 370 4818
rect 404 4784 420 4818
rect 354 4768 420 4784
rect 546 4818 612 4834
rect 660 4830 690 4856
rect 756 4834 786 4856
rect 546 4784 562 4818
rect 596 4784 612 4818
rect 546 4768 612 4784
rect 738 4818 804 4834
rect 852 4830 882 4856
rect 948 4834 978 4856
rect 738 4784 754 4818
rect 788 4784 804 4818
rect 738 4768 804 4784
rect 930 4818 996 4834
rect 1044 4830 1074 4856
rect 1140 4834 1170 4856
rect 930 4784 946 4818
rect 980 4784 996 4818
rect 930 4768 996 4784
rect 1122 4818 1188 4834
rect 1122 4784 1138 4818
rect 1172 4784 1188 4818
rect 1122 4768 1188 4784
rect 354 4710 420 4726
rect 354 4676 370 4710
rect 404 4676 420 4710
rect 276 4638 306 4664
rect 354 4660 420 4676
rect 546 4710 612 4726
rect 546 4676 562 4710
rect 596 4676 612 4710
rect 372 4638 402 4660
rect 468 4638 498 4664
rect 546 4660 612 4676
rect 738 4710 804 4726
rect 738 4676 754 4710
rect 788 4676 804 4710
rect 564 4638 594 4660
rect 660 4638 690 4664
rect 738 4660 804 4676
rect 930 4710 996 4726
rect 930 4676 946 4710
rect 980 4676 996 4710
rect 756 4638 786 4660
rect 852 4638 882 4664
rect 930 4660 996 4676
rect 1122 4710 1188 4726
rect 1122 4676 1138 4710
rect 1172 4676 1188 4710
rect 948 4638 978 4660
rect 1044 4638 1074 4664
rect 1122 4660 1188 4676
rect 1140 4638 1170 4660
rect 276 4216 306 4238
rect 258 4200 324 4216
rect 372 4212 402 4238
rect 468 4216 498 4238
rect 258 4166 274 4200
rect 308 4166 324 4200
rect 258 4150 324 4166
rect 450 4200 516 4216
rect 564 4212 594 4238
rect 660 4216 690 4238
rect 450 4166 466 4200
rect 500 4166 516 4200
rect 450 4150 516 4166
rect 642 4200 708 4216
rect 756 4212 786 4238
rect 852 4216 882 4238
rect 642 4166 658 4200
rect 692 4166 708 4200
rect 642 4150 708 4166
rect 834 4200 900 4216
rect 948 4212 978 4238
rect 1044 4216 1074 4238
rect 834 4166 850 4200
rect 884 4166 900 4200
rect 834 4150 900 4166
rect 1026 4200 1092 4216
rect 1140 4212 1170 4238
rect 1026 4166 1042 4200
rect 1076 4166 1092 4200
rect 1026 4150 1092 4166
rect 2154 5946 2220 5962
rect 2154 5912 2170 5946
rect 2204 5912 2220 5946
rect 2076 5874 2106 5900
rect 2154 5896 2220 5912
rect 2346 5946 2412 5962
rect 2346 5912 2362 5946
rect 2396 5912 2412 5946
rect 2172 5874 2202 5896
rect 2268 5874 2298 5900
rect 2346 5896 2412 5912
rect 2538 5946 2604 5962
rect 2538 5912 2554 5946
rect 2588 5912 2604 5946
rect 2364 5874 2394 5896
rect 2460 5874 2490 5900
rect 2538 5896 2604 5912
rect 2730 5946 2796 5962
rect 2730 5912 2746 5946
rect 2780 5912 2796 5946
rect 2556 5874 2586 5896
rect 2652 5874 2682 5900
rect 2730 5896 2796 5912
rect 2922 5946 2988 5962
rect 2922 5912 2938 5946
rect 2972 5912 2988 5946
rect 2748 5874 2778 5896
rect 2844 5874 2874 5900
rect 2922 5896 2988 5912
rect 2940 5874 2970 5896
rect 2076 5452 2106 5474
rect 2058 5436 2124 5452
rect 2172 5448 2202 5474
rect 2268 5452 2298 5474
rect 2058 5402 2074 5436
rect 2108 5402 2124 5436
rect 2058 5386 2124 5402
rect 2250 5436 2316 5452
rect 2364 5448 2394 5474
rect 2460 5452 2490 5474
rect 2250 5402 2266 5436
rect 2300 5402 2316 5436
rect 2250 5386 2316 5402
rect 2442 5436 2508 5452
rect 2556 5448 2586 5474
rect 2652 5452 2682 5474
rect 2442 5402 2458 5436
rect 2492 5402 2508 5436
rect 2442 5386 2508 5402
rect 2634 5436 2700 5452
rect 2748 5448 2778 5474
rect 2844 5452 2874 5474
rect 2634 5402 2650 5436
rect 2684 5402 2700 5436
rect 2634 5386 2700 5402
rect 2826 5436 2892 5452
rect 2940 5448 2970 5474
rect 2826 5402 2842 5436
rect 2876 5402 2892 5436
rect 2826 5386 2892 5402
rect 2058 5328 2124 5344
rect 2058 5294 2074 5328
rect 2108 5294 2124 5328
rect 2058 5278 2124 5294
rect 2250 5328 2316 5344
rect 2250 5294 2266 5328
rect 2300 5294 2316 5328
rect 2076 5256 2106 5278
rect 2172 5256 2202 5282
rect 2250 5278 2316 5294
rect 2442 5328 2508 5344
rect 2442 5294 2458 5328
rect 2492 5294 2508 5328
rect 2268 5256 2298 5278
rect 2364 5256 2394 5282
rect 2442 5278 2508 5294
rect 2634 5328 2700 5344
rect 2634 5294 2650 5328
rect 2684 5294 2700 5328
rect 2460 5256 2490 5278
rect 2556 5256 2586 5282
rect 2634 5278 2700 5294
rect 2826 5328 2892 5344
rect 2826 5294 2842 5328
rect 2876 5294 2892 5328
rect 2652 5256 2682 5278
rect 2748 5256 2778 5282
rect 2826 5278 2892 5294
rect 2844 5256 2874 5278
rect 2940 5256 2970 5282
rect 2076 4830 2106 4856
rect 2172 4834 2202 4856
rect 2154 4818 2220 4834
rect 2268 4830 2298 4856
rect 2364 4834 2394 4856
rect 2154 4784 2170 4818
rect 2204 4784 2220 4818
rect 2154 4768 2220 4784
rect 2346 4818 2412 4834
rect 2460 4830 2490 4856
rect 2556 4834 2586 4856
rect 2346 4784 2362 4818
rect 2396 4784 2412 4818
rect 2346 4768 2412 4784
rect 2538 4818 2604 4834
rect 2652 4830 2682 4856
rect 2748 4834 2778 4856
rect 2538 4784 2554 4818
rect 2588 4784 2604 4818
rect 2538 4768 2604 4784
rect 2730 4818 2796 4834
rect 2844 4830 2874 4856
rect 2940 4834 2970 4856
rect 2730 4784 2746 4818
rect 2780 4784 2796 4818
rect 2730 4768 2796 4784
rect 2922 4818 2988 4834
rect 2922 4784 2938 4818
rect 2972 4784 2988 4818
rect 2922 4768 2988 4784
rect 2154 4710 2220 4726
rect 2154 4676 2170 4710
rect 2204 4676 2220 4710
rect 2076 4638 2106 4664
rect 2154 4660 2220 4676
rect 2346 4710 2412 4726
rect 2346 4676 2362 4710
rect 2396 4676 2412 4710
rect 2172 4638 2202 4660
rect 2268 4638 2298 4664
rect 2346 4660 2412 4676
rect 2538 4710 2604 4726
rect 2538 4676 2554 4710
rect 2588 4676 2604 4710
rect 2364 4638 2394 4660
rect 2460 4638 2490 4664
rect 2538 4660 2604 4676
rect 2730 4710 2796 4726
rect 2730 4676 2746 4710
rect 2780 4676 2796 4710
rect 2556 4638 2586 4660
rect 2652 4638 2682 4664
rect 2730 4660 2796 4676
rect 2922 4710 2988 4726
rect 2922 4676 2938 4710
rect 2972 4676 2988 4710
rect 2748 4638 2778 4660
rect 2844 4638 2874 4664
rect 2922 4660 2988 4676
rect 2940 4638 2970 4660
rect 2076 4216 2106 4238
rect 2058 4200 2124 4216
rect 2172 4212 2202 4238
rect 2268 4216 2298 4238
rect 2058 4166 2074 4200
rect 2108 4166 2124 4200
rect 2058 4150 2124 4166
rect 2250 4200 2316 4216
rect 2364 4212 2394 4238
rect 2460 4216 2490 4238
rect 2250 4166 2266 4200
rect 2300 4166 2316 4200
rect 2250 4150 2316 4166
rect 2442 4200 2508 4216
rect 2556 4212 2586 4238
rect 2652 4216 2682 4238
rect 2442 4166 2458 4200
rect 2492 4166 2508 4200
rect 2442 4150 2508 4166
rect 2634 4200 2700 4216
rect 2748 4212 2778 4238
rect 2844 4216 2874 4238
rect 2634 4166 2650 4200
rect 2684 4166 2700 4200
rect 2634 4150 2700 4166
rect 2826 4200 2892 4216
rect 2940 4212 2970 4238
rect 2826 4166 2842 4200
rect 2876 4166 2892 4200
rect 2826 4150 2892 4166
rect 3954 5946 4020 5962
rect 3954 5912 3970 5946
rect 4004 5912 4020 5946
rect 3876 5874 3906 5900
rect 3954 5896 4020 5912
rect 4146 5946 4212 5962
rect 4146 5912 4162 5946
rect 4196 5912 4212 5946
rect 3972 5874 4002 5896
rect 4068 5874 4098 5900
rect 4146 5896 4212 5912
rect 4338 5946 4404 5962
rect 4338 5912 4354 5946
rect 4388 5912 4404 5946
rect 4164 5874 4194 5896
rect 4260 5874 4290 5900
rect 4338 5896 4404 5912
rect 4530 5946 4596 5962
rect 4530 5912 4546 5946
rect 4580 5912 4596 5946
rect 4356 5874 4386 5896
rect 4452 5874 4482 5900
rect 4530 5896 4596 5912
rect 4722 5946 4788 5962
rect 4722 5912 4738 5946
rect 4772 5912 4788 5946
rect 4548 5874 4578 5896
rect 4644 5874 4674 5900
rect 4722 5896 4788 5912
rect 4740 5874 4770 5896
rect 3876 5452 3906 5474
rect 3858 5436 3924 5452
rect 3972 5448 4002 5474
rect 4068 5452 4098 5474
rect 3858 5402 3874 5436
rect 3908 5402 3924 5436
rect 3858 5386 3924 5402
rect 4050 5436 4116 5452
rect 4164 5448 4194 5474
rect 4260 5452 4290 5474
rect 4050 5402 4066 5436
rect 4100 5402 4116 5436
rect 4050 5386 4116 5402
rect 4242 5436 4308 5452
rect 4356 5448 4386 5474
rect 4452 5452 4482 5474
rect 4242 5402 4258 5436
rect 4292 5402 4308 5436
rect 4242 5386 4308 5402
rect 4434 5436 4500 5452
rect 4548 5448 4578 5474
rect 4644 5452 4674 5474
rect 4434 5402 4450 5436
rect 4484 5402 4500 5436
rect 4434 5386 4500 5402
rect 4626 5436 4692 5452
rect 4740 5448 4770 5474
rect 4626 5402 4642 5436
rect 4676 5402 4692 5436
rect 4626 5386 4692 5402
rect 3858 5328 3924 5344
rect 3858 5294 3874 5328
rect 3908 5294 3924 5328
rect 3858 5278 3924 5294
rect 4050 5328 4116 5344
rect 4050 5294 4066 5328
rect 4100 5294 4116 5328
rect 3876 5256 3906 5278
rect 3972 5256 4002 5282
rect 4050 5278 4116 5294
rect 4242 5328 4308 5344
rect 4242 5294 4258 5328
rect 4292 5294 4308 5328
rect 4068 5256 4098 5278
rect 4164 5256 4194 5282
rect 4242 5278 4308 5294
rect 4434 5328 4500 5344
rect 4434 5294 4450 5328
rect 4484 5294 4500 5328
rect 4260 5256 4290 5278
rect 4356 5256 4386 5282
rect 4434 5278 4500 5294
rect 4626 5328 4692 5344
rect 4626 5294 4642 5328
rect 4676 5294 4692 5328
rect 4452 5256 4482 5278
rect 4548 5256 4578 5282
rect 4626 5278 4692 5294
rect 4644 5256 4674 5278
rect 4740 5256 4770 5282
rect 3876 4830 3906 4856
rect 3972 4834 4002 4856
rect 3954 4818 4020 4834
rect 4068 4830 4098 4856
rect 4164 4834 4194 4856
rect 3954 4784 3970 4818
rect 4004 4784 4020 4818
rect 3954 4768 4020 4784
rect 4146 4818 4212 4834
rect 4260 4830 4290 4856
rect 4356 4834 4386 4856
rect 4146 4784 4162 4818
rect 4196 4784 4212 4818
rect 4146 4768 4212 4784
rect 4338 4818 4404 4834
rect 4452 4830 4482 4856
rect 4548 4834 4578 4856
rect 4338 4784 4354 4818
rect 4388 4784 4404 4818
rect 4338 4768 4404 4784
rect 4530 4818 4596 4834
rect 4644 4830 4674 4856
rect 4740 4834 4770 4856
rect 4530 4784 4546 4818
rect 4580 4784 4596 4818
rect 4530 4768 4596 4784
rect 4722 4818 4788 4834
rect 4722 4784 4738 4818
rect 4772 4784 4788 4818
rect 4722 4768 4788 4784
rect 3954 4710 4020 4726
rect 3954 4676 3970 4710
rect 4004 4676 4020 4710
rect 3876 4638 3906 4664
rect 3954 4660 4020 4676
rect 4146 4710 4212 4726
rect 4146 4676 4162 4710
rect 4196 4676 4212 4710
rect 3972 4638 4002 4660
rect 4068 4638 4098 4664
rect 4146 4660 4212 4676
rect 4338 4710 4404 4726
rect 4338 4676 4354 4710
rect 4388 4676 4404 4710
rect 4164 4638 4194 4660
rect 4260 4638 4290 4664
rect 4338 4660 4404 4676
rect 4530 4710 4596 4726
rect 4530 4676 4546 4710
rect 4580 4676 4596 4710
rect 4356 4638 4386 4660
rect 4452 4638 4482 4664
rect 4530 4660 4596 4676
rect 4722 4710 4788 4726
rect 4722 4676 4738 4710
rect 4772 4676 4788 4710
rect 4548 4638 4578 4660
rect 4644 4638 4674 4664
rect 4722 4660 4788 4676
rect 4740 4638 4770 4660
rect 3876 4216 3906 4238
rect 3858 4200 3924 4216
rect 3972 4212 4002 4238
rect 4068 4216 4098 4238
rect 3858 4166 3874 4200
rect 3908 4166 3924 4200
rect 3858 4150 3924 4166
rect 4050 4200 4116 4216
rect 4164 4212 4194 4238
rect 4260 4216 4290 4238
rect 4050 4166 4066 4200
rect 4100 4166 4116 4200
rect 4050 4150 4116 4166
rect 4242 4200 4308 4216
rect 4356 4212 4386 4238
rect 4452 4216 4482 4238
rect 4242 4166 4258 4200
rect 4292 4166 4308 4200
rect 4242 4150 4308 4166
rect 4434 4200 4500 4216
rect 4548 4212 4578 4238
rect 4644 4216 4674 4238
rect 4434 4166 4450 4200
rect 4484 4166 4500 4200
rect 4434 4150 4500 4166
rect 4626 4200 4692 4216
rect 4740 4212 4770 4238
rect 4626 4166 4642 4200
rect 4676 4166 4692 4200
rect 4626 4150 4692 4166
rect 5754 5946 5820 5962
rect 5754 5912 5770 5946
rect 5804 5912 5820 5946
rect 5676 5874 5706 5900
rect 5754 5896 5820 5912
rect 5946 5946 6012 5962
rect 5946 5912 5962 5946
rect 5996 5912 6012 5946
rect 5772 5874 5802 5896
rect 5868 5874 5898 5900
rect 5946 5896 6012 5912
rect 6138 5946 6204 5962
rect 6138 5912 6154 5946
rect 6188 5912 6204 5946
rect 5964 5874 5994 5896
rect 6060 5874 6090 5900
rect 6138 5896 6204 5912
rect 6330 5946 6396 5962
rect 6330 5912 6346 5946
rect 6380 5912 6396 5946
rect 6156 5874 6186 5896
rect 6252 5874 6282 5900
rect 6330 5896 6396 5912
rect 6522 5946 6588 5962
rect 6522 5912 6538 5946
rect 6572 5912 6588 5946
rect 6348 5874 6378 5896
rect 6444 5874 6474 5900
rect 6522 5896 6588 5912
rect 6540 5874 6570 5896
rect 5676 5452 5706 5474
rect 5658 5436 5724 5452
rect 5772 5448 5802 5474
rect 5868 5452 5898 5474
rect 5658 5402 5674 5436
rect 5708 5402 5724 5436
rect 5658 5386 5724 5402
rect 5850 5436 5916 5452
rect 5964 5448 5994 5474
rect 6060 5452 6090 5474
rect 5850 5402 5866 5436
rect 5900 5402 5916 5436
rect 5850 5386 5916 5402
rect 6042 5436 6108 5452
rect 6156 5448 6186 5474
rect 6252 5452 6282 5474
rect 6042 5402 6058 5436
rect 6092 5402 6108 5436
rect 6042 5386 6108 5402
rect 6234 5436 6300 5452
rect 6348 5448 6378 5474
rect 6444 5452 6474 5474
rect 6234 5402 6250 5436
rect 6284 5402 6300 5436
rect 6234 5386 6300 5402
rect 6426 5436 6492 5452
rect 6540 5448 6570 5474
rect 6426 5402 6442 5436
rect 6476 5402 6492 5436
rect 6426 5386 6492 5402
rect 5658 5328 5724 5344
rect 5658 5294 5674 5328
rect 5708 5294 5724 5328
rect 5658 5278 5724 5294
rect 5850 5328 5916 5344
rect 5850 5294 5866 5328
rect 5900 5294 5916 5328
rect 5676 5256 5706 5278
rect 5772 5256 5802 5282
rect 5850 5278 5916 5294
rect 6042 5328 6108 5344
rect 6042 5294 6058 5328
rect 6092 5294 6108 5328
rect 5868 5256 5898 5278
rect 5964 5256 5994 5282
rect 6042 5278 6108 5294
rect 6234 5328 6300 5344
rect 6234 5294 6250 5328
rect 6284 5294 6300 5328
rect 6060 5256 6090 5278
rect 6156 5256 6186 5282
rect 6234 5278 6300 5294
rect 6426 5328 6492 5344
rect 6426 5294 6442 5328
rect 6476 5294 6492 5328
rect 6252 5256 6282 5278
rect 6348 5256 6378 5282
rect 6426 5278 6492 5294
rect 6444 5256 6474 5278
rect 6540 5256 6570 5282
rect 5676 4830 5706 4856
rect 5772 4834 5802 4856
rect 5754 4818 5820 4834
rect 5868 4830 5898 4856
rect 5964 4834 5994 4856
rect 5754 4784 5770 4818
rect 5804 4784 5820 4818
rect 5754 4768 5820 4784
rect 5946 4818 6012 4834
rect 6060 4830 6090 4856
rect 6156 4834 6186 4856
rect 5946 4784 5962 4818
rect 5996 4784 6012 4818
rect 5946 4768 6012 4784
rect 6138 4818 6204 4834
rect 6252 4830 6282 4856
rect 6348 4834 6378 4856
rect 6138 4784 6154 4818
rect 6188 4784 6204 4818
rect 6138 4768 6204 4784
rect 6330 4818 6396 4834
rect 6444 4830 6474 4856
rect 6540 4834 6570 4856
rect 6330 4784 6346 4818
rect 6380 4784 6396 4818
rect 6330 4768 6396 4784
rect 6522 4818 6588 4834
rect 6522 4784 6538 4818
rect 6572 4784 6588 4818
rect 6522 4768 6588 4784
rect 5754 4710 5820 4726
rect 5754 4676 5770 4710
rect 5804 4676 5820 4710
rect 5676 4638 5706 4664
rect 5754 4660 5820 4676
rect 5946 4710 6012 4726
rect 5946 4676 5962 4710
rect 5996 4676 6012 4710
rect 5772 4638 5802 4660
rect 5868 4638 5898 4664
rect 5946 4660 6012 4676
rect 6138 4710 6204 4726
rect 6138 4676 6154 4710
rect 6188 4676 6204 4710
rect 5964 4638 5994 4660
rect 6060 4638 6090 4664
rect 6138 4660 6204 4676
rect 6330 4710 6396 4726
rect 6330 4676 6346 4710
rect 6380 4676 6396 4710
rect 6156 4638 6186 4660
rect 6252 4638 6282 4664
rect 6330 4660 6396 4676
rect 6522 4710 6588 4726
rect 6522 4676 6538 4710
rect 6572 4676 6588 4710
rect 6348 4638 6378 4660
rect 6444 4638 6474 4664
rect 6522 4660 6588 4676
rect 6540 4638 6570 4660
rect 5676 4216 5706 4238
rect 5658 4200 5724 4216
rect 5772 4212 5802 4238
rect 5868 4216 5898 4238
rect 5658 4166 5674 4200
rect 5708 4166 5724 4200
rect 5658 4150 5724 4166
rect 5850 4200 5916 4216
rect 5964 4212 5994 4238
rect 6060 4216 6090 4238
rect 5850 4166 5866 4200
rect 5900 4166 5916 4200
rect 5850 4150 5916 4166
rect 6042 4200 6108 4216
rect 6156 4212 6186 4238
rect 6252 4216 6282 4238
rect 6042 4166 6058 4200
rect 6092 4166 6108 4200
rect 6042 4150 6108 4166
rect 6234 4200 6300 4216
rect 6348 4212 6378 4238
rect 6444 4216 6474 4238
rect 6234 4166 6250 4200
rect 6284 4166 6300 4200
rect 6234 4150 6300 4166
rect 6426 4200 6492 4216
rect 6540 4212 6570 4238
rect 6426 4166 6442 4200
rect 6476 4166 6492 4200
rect 6426 4150 6492 4166
rect 7754 10334 7820 10350
rect 7754 10300 7770 10334
rect 7804 10300 7820 10334
rect 7676 10262 7706 10288
rect 7754 10284 7820 10300
rect 7946 10334 8012 10350
rect 7946 10300 7962 10334
rect 7996 10300 8012 10334
rect 7772 10262 7802 10284
rect 7868 10262 7898 10288
rect 7946 10284 8012 10300
rect 8138 10334 8204 10350
rect 8138 10300 8154 10334
rect 8188 10300 8204 10334
rect 7964 10262 7994 10284
rect 8060 10262 8090 10288
rect 8138 10284 8204 10300
rect 8330 10334 8396 10350
rect 8330 10300 8346 10334
rect 8380 10300 8396 10334
rect 8156 10262 8186 10284
rect 8252 10262 8282 10288
rect 8330 10284 8396 10300
rect 8522 10334 8588 10350
rect 8522 10300 8538 10334
rect 8572 10300 8588 10334
rect 8348 10262 8378 10284
rect 8444 10262 8474 10288
rect 8522 10284 8588 10300
rect 8714 10334 8780 10350
rect 8714 10300 8730 10334
rect 8764 10300 8780 10334
rect 8540 10262 8570 10284
rect 8636 10262 8666 10288
rect 8714 10284 8780 10300
rect 8906 10334 8972 10350
rect 8906 10300 8922 10334
rect 8956 10300 8972 10334
rect 8732 10262 8762 10284
rect 8828 10262 8858 10288
rect 8906 10284 8972 10300
rect 9098 10334 9164 10350
rect 9098 10300 9114 10334
rect 9148 10300 9164 10334
rect 8924 10262 8954 10284
rect 9020 10262 9050 10288
rect 9098 10284 9164 10300
rect 9290 10334 9356 10350
rect 9290 10300 9306 10334
rect 9340 10300 9356 10334
rect 9116 10262 9146 10284
rect 9212 10262 9242 10288
rect 9290 10284 9356 10300
rect 9482 10334 9548 10350
rect 9482 10300 9498 10334
rect 9532 10300 9548 10334
rect 9308 10262 9338 10284
rect 9404 10262 9434 10288
rect 9482 10284 9548 10300
rect 9500 10262 9530 10284
rect 7676 9840 7706 9862
rect 7658 9824 7724 9840
rect 7772 9836 7802 9862
rect 7868 9840 7898 9862
rect 7658 9790 7674 9824
rect 7708 9790 7724 9824
rect 7658 9774 7724 9790
rect 7850 9824 7916 9840
rect 7964 9836 7994 9862
rect 8060 9840 8090 9862
rect 7850 9790 7866 9824
rect 7900 9790 7916 9824
rect 7850 9774 7916 9790
rect 8042 9824 8108 9840
rect 8156 9836 8186 9862
rect 8252 9840 8282 9862
rect 8042 9790 8058 9824
rect 8092 9790 8108 9824
rect 8042 9774 8108 9790
rect 8234 9824 8300 9840
rect 8348 9836 8378 9862
rect 8444 9840 8474 9862
rect 8234 9790 8250 9824
rect 8284 9790 8300 9824
rect 8234 9774 8300 9790
rect 8426 9824 8492 9840
rect 8540 9836 8570 9862
rect 8636 9840 8666 9862
rect 8426 9790 8442 9824
rect 8476 9790 8492 9824
rect 8426 9774 8492 9790
rect 8618 9824 8684 9840
rect 8732 9836 8762 9862
rect 8828 9840 8858 9862
rect 8618 9790 8634 9824
rect 8668 9790 8684 9824
rect 8618 9774 8684 9790
rect 8810 9824 8876 9840
rect 8924 9836 8954 9862
rect 9020 9840 9050 9862
rect 8810 9790 8826 9824
rect 8860 9790 8876 9824
rect 8810 9774 8876 9790
rect 9002 9824 9068 9840
rect 9116 9836 9146 9862
rect 9212 9840 9242 9862
rect 9002 9790 9018 9824
rect 9052 9790 9068 9824
rect 9002 9774 9068 9790
rect 9194 9824 9260 9840
rect 9308 9836 9338 9862
rect 9404 9840 9434 9862
rect 9194 9790 9210 9824
rect 9244 9790 9260 9824
rect 9194 9774 9260 9790
rect 9386 9824 9452 9840
rect 9500 9836 9530 9862
rect 9386 9790 9402 9824
rect 9436 9790 9452 9824
rect 9386 9774 9452 9790
rect 7658 9716 7724 9732
rect 7658 9682 7674 9716
rect 7708 9682 7724 9716
rect 7658 9666 7724 9682
rect 7850 9716 7916 9732
rect 7850 9682 7866 9716
rect 7900 9682 7916 9716
rect 7676 9644 7706 9666
rect 7772 9644 7802 9670
rect 7850 9666 7916 9682
rect 8042 9716 8108 9732
rect 8042 9682 8058 9716
rect 8092 9682 8108 9716
rect 7868 9644 7898 9666
rect 7964 9644 7994 9670
rect 8042 9666 8108 9682
rect 8234 9716 8300 9732
rect 8234 9682 8250 9716
rect 8284 9682 8300 9716
rect 8060 9644 8090 9666
rect 8156 9644 8186 9670
rect 8234 9666 8300 9682
rect 8426 9716 8492 9732
rect 8426 9682 8442 9716
rect 8476 9682 8492 9716
rect 8252 9644 8282 9666
rect 8348 9644 8378 9670
rect 8426 9666 8492 9682
rect 8618 9716 8684 9732
rect 8618 9682 8634 9716
rect 8668 9682 8684 9716
rect 8444 9644 8474 9666
rect 8540 9644 8570 9670
rect 8618 9666 8684 9682
rect 8810 9716 8876 9732
rect 8810 9682 8826 9716
rect 8860 9682 8876 9716
rect 8636 9644 8666 9666
rect 8732 9644 8762 9670
rect 8810 9666 8876 9682
rect 9002 9716 9068 9732
rect 9002 9682 9018 9716
rect 9052 9682 9068 9716
rect 8828 9644 8858 9666
rect 8924 9644 8954 9670
rect 9002 9666 9068 9682
rect 9194 9716 9260 9732
rect 9194 9682 9210 9716
rect 9244 9682 9260 9716
rect 9020 9644 9050 9666
rect 9116 9644 9146 9670
rect 9194 9666 9260 9682
rect 9386 9716 9452 9732
rect 9386 9682 9402 9716
rect 9436 9682 9452 9716
rect 9212 9644 9242 9666
rect 9308 9644 9338 9670
rect 9386 9666 9452 9682
rect 9404 9644 9434 9666
rect 9500 9644 9530 9670
rect 7676 9218 7706 9244
rect 7772 9222 7802 9244
rect 7754 9206 7820 9222
rect 7868 9218 7898 9244
rect 7964 9222 7994 9244
rect 7754 9172 7770 9206
rect 7804 9172 7820 9206
rect 7754 9156 7820 9172
rect 7946 9206 8012 9222
rect 8060 9218 8090 9244
rect 8156 9222 8186 9244
rect 7946 9172 7962 9206
rect 7996 9172 8012 9206
rect 7946 9156 8012 9172
rect 8138 9206 8204 9222
rect 8252 9218 8282 9244
rect 8348 9222 8378 9244
rect 8138 9172 8154 9206
rect 8188 9172 8204 9206
rect 8138 9156 8204 9172
rect 8330 9206 8396 9222
rect 8444 9218 8474 9244
rect 8540 9222 8570 9244
rect 8330 9172 8346 9206
rect 8380 9172 8396 9206
rect 8330 9156 8396 9172
rect 8522 9206 8588 9222
rect 8636 9218 8666 9244
rect 8732 9222 8762 9244
rect 8522 9172 8538 9206
rect 8572 9172 8588 9206
rect 8522 9156 8588 9172
rect 8714 9206 8780 9222
rect 8828 9218 8858 9244
rect 8924 9222 8954 9244
rect 8714 9172 8730 9206
rect 8764 9172 8780 9206
rect 8714 9156 8780 9172
rect 8906 9206 8972 9222
rect 9020 9218 9050 9244
rect 9116 9222 9146 9244
rect 8906 9172 8922 9206
rect 8956 9172 8972 9206
rect 8906 9156 8972 9172
rect 9098 9206 9164 9222
rect 9212 9218 9242 9244
rect 9308 9222 9338 9244
rect 9098 9172 9114 9206
rect 9148 9172 9164 9206
rect 9098 9156 9164 9172
rect 9290 9206 9356 9222
rect 9404 9218 9434 9244
rect 9500 9222 9530 9244
rect 9290 9172 9306 9206
rect 9340 9172 9356 9206
rect 9290 9156 9356 9172
rect 9482 9206 9548 9222
rect 9482 9172 9498 9206
rect 9532 9172 9548 9206
rect 9482 9156 9548 9172
rect 7754 9098 7820 9114
rect 7754 9064 7770 9098
rect 7804 9064 7820 9098
rect 7676 9026 7706 9052
rect 7754 9048 7820 9064
rect 7946 9098 8012 9114
rect 7946 9064 7962 9098
rect 7996 9064 8012 9098
rect 7772 9026 7802 9048
rect 7868 9026 7898 9052
rect 7946 9048 8012 9064
rect 8138 9098 8204 9114
rect 8138 9064 8154 9098
rect 8188 9064 8204 9098
rect 7964 9026 7994 9048
rect 8060 9026 8090 9052
rect 8138 9048 8204 9064
rect 8330 9098 8396 9114
rect 8330 9064 8346 9098
rect 8380 9064 8396 9098
rect 8156 9026 8186 9048
rect 8252 9026 8282 9052
rect 8330 9048 8396 9064
rect 8522 9098 8588 9114
rect 8522 9064 8538 9098
rect 8572 9064 8588 9098
rect 8348 9026 8378 9048
rect 8444 9026 8474 9052
rect 8522 9048 8588 9064
rect 8714 9098 8780 9114
rect 8714 9064 8730 9098
rect 8764 9064 8780 9098
rect 8540 9026 8570 9048
rect 8636 9026 8666 9052
rect 8714 9048 8780 9064
rect 8906 9098 8972 9114
rect 8906 9064 8922 9098
rect 8956 9064 8972 9098
rect 8732 9026 8762 9048
rect 8828 9026 8858 9052
rect 8906 9048 8972 9064
rect 9098 9098 9164 9114
rect 9098 9064 9114 9098
rect 9148 9064 9164 9098
rect 8924 9026 8954 9048
rect 9020 9026 9050 9052
rect 9098 9048 9164 9064
rect 9290 9098 9356 9114
rect 9290 9064 9306 9098
rect 9340 9064 9356 9098
rect 9116 9026 9146 9048
rect 9212 9026 9242 9052
rect 9290 9048 9356 9064
rect 9482 9098 9548 9114
rect 9482 9064 9498 9098
rect 9532 9064 9548 9098
rect 9308 9026 9338 9048
rect 9404 9026 9434 9052
rect 9482 9048 9548 9064
rect 9500 9026 9530 9048
rect 7676 8604 7706 8626
rect 7658 8588 7724 8604
rect 7772 8600 7802 8626
rect 7868 8604 7898 8626
rect 7658 8554 7674 8588
rect 7708 8554 7724 8588
rect 7658 8538 7724 8554
rect 7850 8588 7916 8604
rect 7964 8600 7994 8626
rect 8060 8604 8090 8626
rect 7850 8554 7866 8588
rect 7900 8554 7916 8588
rect 7850 8538 7916 8554
rect 8042 8588 8108 8604
rect 8156 8600 8186 8626
rect 8252 8604 8282 8626
rect 8042 8554 8058 8588
rect 8092 8554 8108 8588
rect 8042 8538 8108 8554
rect 8234 8588 8300 8604
rect 8348 8600 8378 8626
rect 8444 8604 8474 8626
rect 8234 8554 8250 8588
rect 8284 8554 8300 8588
rect 8234 8538 8300 8554
rect 8426 8588 8492 8604
rect 8540 8600 8570 8626
rect 8636 8604 8666 8626
rect 8426 8554 8442 8588
rect 8476 8554 8492 8588
rect 8426 8538 8492 8554
rect 8618 8588 8684 8604
rect 8732 8600 8762 8626
rect 8828 8604 8858 8626
rect 8618 8554 8634 8588
rect 8668 8554 8684 8588
rect 8618 8538 8684 8554
rect 8810 8588 8876 8604
rect 8924 8600 8954 8626
rect 9020 8604 9050 8626
rect 8810 8554 8826 8588
rect 8860 8554 8876 8588
rect 8810 8538 8876 8554
rect 9002 8588 9068 8604
rect 9116 8600 9146 8626
rect 9212 8604 9242 8626
rect 9002 8554 9018 8588
rect 9052 8554 9068 8588
rect 9002 8538 9068 8554
rect 9194 8588 9260 8604
rect 9308 8600 9338 8626
rect 9404 8604 9434 8626
rect 9194 8554 9210 8588
rect 9244 8554 9260 8588
rect 9194 8538 9260 8554
rect 9386 8588 9452 8604
rect 9500 8600 9530 8626
rect 9386 8554 9402 8588
rect 9436 8554 9452 8588
rect 9386 8538 9452 8554
rect 7658 8480 7724 8496
rect 7658 8446 7674 8480
rect 7708 8446 7724 8480
rect 7658 8430 7724 8446
rect 7850 8480 7916 8496
rect 7850 8446 7866 8480
rect 7900 8446 7916 8480
rect 7676 8408 7706 8430
rect 7772 8408 7802 8434
rect 7850 8430 7916 8446
rect 8042 8480 8108 8496
rect 8042 8446 8058 8480
rect 8092 8446 8108 8480
rect 7868 8408 7898 8430
rect 7964 8408 7994 8434
rect 8042 8430 8108 8446
rect 8234 8480 8300 8496
rect 8234 8446 8250 8480
rect 8284 8446 8300 8480
rect 8060 8408 8090 8430
rect 8156 8408 8186 8434
rect 8234 8430 8300 8446
rect 8426 8480 8492 8496
rect 8426 8446 8442 8480
rect 8476 8446 8492 8480
rect 8252 8408 8282 8430
rect 8348 8408 8378 8434
rect 8426 8430 8492 8446
rect 8618 8480 8684 8496
rect 8618 8446 8634 8480
rect 8668 8446 8684 8480
rect 8444 8408 8474 8430
rect 8540 8408 8570 8434
rect 8618 8430 8684 8446
rect 8810 8480 8876 8496
rect 8810 8446 8826 8480
rect 8860 8446 8876 8480
rect 8636 8408 8666 8430
rect 8732 8408 8762 8434
rect 8810 8430 8876 8446
rect 9002 8480 9068 8496
rect 9002 8446 9018 8480
rect 9052 8446 9068 8480
rect 8828 8408 8858 8430
rect 8924 8408 8954 8434
rect 9002 8430 9068 8446
rect 9194 8480 9260 8496
rect 9194 8446 9210 8480
rect 9244 8446 9260 8480
rect 9020 8408 9050 8430
rect 9116 8408 9146 8434
rect 9194 8430 9260 8446
rect 9386 8480 9452 8496
rect 9386 8446 9402 8480
rect 9436 8446 9452 8480
rect 9212 8408 9242 8430
rect 9308 8408 9338 8434
rect 9386 8430 9452 8446
rect 9404 8408 9434 8430
rect 9500 8408 9530 8434
rect 7676 7982 7706 8008
rect 7772 7986 7802 8008
rect 7754 7970 7820 7986
rect 7868 7982 7898 8008
rect 7964 7986 7994 8008
rect 7754 7936 7770 7970
rect 7804 7936 7820 7970
rect 7754 7920 7820 7936
rect 7946 7970 8012 7986
rect 8060 7982 8090 8008
rect 8156 7986 8186 8008
rect 7946 7936 7962 7970
rect 7996 7936 8012 7970
rect 7946 7920 8012 7936
rect 8138 7970 8204 7986
rect 8252 7982 8282 8008
rect 8348 7986 8378 8008
rect 8138 7936 8154 7970
rect 8188 7936 8204 7970
rect 8138 7920 8204 7936
rect 8330 7970 8396 7986
rect 8444 7982 8474 8008
rect 8540 7986 8570 8008
rect 8330 7936 8346 7970
rect 8380 7936 8396 7970
rect 8330 7920 8396 7936
rect 8522 7970 8588 7986
rect 8636 7982 8666 8008
rect 8732 7986 8762 8008
rect 8522 7936 8538 7970
rect 8572 7936 8588 7970
rect 8522 7920 8588 7936
rect 8714 7970 8780 7986
rect 8828 7982 8858 8008
rect 8924 7986 8954 8008
rect 8714 7936 8730 7970
rect 8764 7936 8780 7970
rect 8714 7920 8780 7936
rect 8906 7970 8972 7986
rect 9020 7982 9050 8008
rect 9116 7986 9146 8008
rect 8906 7936 8922 7970
rect 8956 7936 8972 7970
rect 8906 7920 8972 7936
rect 9098 7970 9164 7986
rect 9212 7982 9242 8008
rect 9308 7986 9338 8008
rect 9098 7936 9114 7970
rect 9148 7936 9164 7970
rect 9098 7920 9164 7936
rect 9290 7970 9356 7986
rect 9404 7982 9434 8008
rect 9500 7986 9530 8008
rect 9290 7936 9306 7970
rect 9340 7936 9356 7970
rect 9290 7920 9356 7936
rect 9482 7970 9548 7986
rect 9482 7936 9498 7970
rect 9532 7936 9548 7970
rect 9482 7920 9548 7936
rect 7754 7862 7820 7878
rect 7754 7828 7770 7862
rect 7804 7828 7820 7862
rect 7676 7790 7706 7816
rect 7754 7812 7820 7828
rect 7946 7862 8012 7878
rect 7946 7828 7962 7862
rect 7996 7828 8012 7862
rect 7772 7790 7802 7812
rect 7868 7790 7898 7816
rect 7946 7812 8012 7828
rect 8138 7862 8204 7878
rect 8138 7828 8154 7862
rect 8188 7828 8204 7862
rect 7964 7790 7994 7812
rect 8060 7790 8090 7816
rect 8138 7812 8204 7828
rect 8330 7862 8396 7878
rect 8330 7828 8346 7862
rect 8380 7828 8396 7862
rect 8156 7790 8186 7812
rect 8252 7790 8282 7816
rect 8330 7812 8396 7828
rect 8522 7862 8588 7878
rect 8522 7828 8538 7862
rect 8572 7828 8588 7862
rect 8348 7790 8378 7812
rect 8444 7790 8474 7816
rect 8522 7812 8588 7828
rect 8714 7862 8780 7878
rect 8714 7828 8730 7862
rect 8764 7828 8780 7862
rect 8540 7790 8570 7812
rect 8636 7790 8666 7816
rect 8714 7812 8780 7828
rect 8906 7862 8972 7878
rect 8906 7828 8922 7862
rect 8956 7828 8972 7862
rect 8732 7790 8762 7812
rect 8828 7790 8858 7816
rect 8906 7812 8972 7828
rect 9098 7862 9164 7878
rect 9098 7828 9114 7862
rect 9148 7828 9164 7862
rect 8924 7790 8954 7812
rect 9020 7790 9050 7816
rect 9098 7812 9164 7828
rect 9290 7862 9356 7878
rect 9290 7828 9306 7862
rect 9340 7828 9356 7862
rect 9116 7790 9146 7812
rect 9212 7790 9242 7816
rect 9290 7812 9356 7828
rect 9482 7862 9548 7878
rect 9482 7828 9498 7862
rect 9532 7828 9548 7862
rect 9308 7790 9338 7812
rect 9404 7790 9434 7816
rect 9482 7812 9548 7828
rect 9500 7790 9530 7812
rect 7676 7368 7706 7390
rect 7658 7352 7724 7368
rect 7772 7364 7802 7390
rect 7868 7368 7898 7390
rect 7658 7318 7674 7352
rect 7708 7318 7724 7352
rect 7658 7302 7724 7318
rect 7850 7352 7916 7368
rect 7964 7364 7994 7390
rect 8060 7368 8090 7390
rect 7850 7318 7866 7352
rect 7900 7318 7916 7352
rect 7850 7302 7916 7318
rect 8042 7352 8108 7368
rect 8156 7364 8186 7390
rect 8252 7368 8282 7390
rect 8042 7318 8058 7352
rect 8092 7318 8108 7352
rect 8042 7302 8108 7318
rect 8234 7352 8300 7368
rect 8348 7364 8378 7390
rect 8444 7368 8474 7390
rect 8234 7318 8250 7352
rect 8284 7318 8300 7352
rect 8234 7302 8300 7318
rect 8426 7352 8492 7368
rect 8540 7364 8570 7390
rect 8636 7368 8666 7390
rect 8426 7318 8442 7352
rect 8476 7318 8492 7352
rect 8426 7302 8492 7318
rect 8618 7352 8684 7368
rect 8732 7364 8762 7390
rect 8828 7368 8858 7390
rect 8618 7318 8634 7352
rect 8668 7318 8684 7352
rect 8618 7302 8684 7318
rect 8810 7352 8876 7368
rect 8924 7364 8954 7390
rect 9020 7368 9050 7390
rect 8810 7318 8826 7352
rect 8860 7318 8876 7352
rect 8810 7302 8876 7318
rect 9002 7352 9068 7368
rect 9116 7364 9146 7390
rect 9212 7368 9242 7390
rect 9002 7318 9018 7352
rect 9052 7318 9068 7352
rect 9002 7302 9068 7318
rect 9194 7352 9260 7368
rect 9308 7364 9338 7390
rect 9404 7368 9434 7390
rect 9194 7318 9210 7352
rect 9244 7318 9260 7352
rect 9194 7302 9260 7318
rect 9386 7352 9452 7368
rect 9500 7364 9530 7390
rect 9386 7318 9402 7352
rect 9436 7318 9452 7352
rect 9386 7302 9452 7318
rect 7658 7244 7724 7260
rect 7658 7210 7674 7244
rect 7708 7210 7724 7244
rect 7658 7194 7724 7210
rect 7850 7244 7916 7260
rect 7850 7210 7866 7244
rect 7900 7210 7916 7244
rect 7676 7172 7706 7194
rect 7772 7172 7802 7198
rect 7850 7194 7916 7210
rect 8042 7244 8108 7260
rect 8042 7210 8058 7244
rect 8092 7210 8108 7244
rect 7868 7172 7898 7194
rect 7964 7172 7994 7198
rect 8042 7194 8108 7210
rect 8234 7244 8300 7260
rect 8234 7210 8250 7244
rect 8284 7210 8300 7244
rect 8060 7172 8090 7194
rect 8156 7172 8186 7198
rect 8234 7194 8300 7210
rect 8426 7244 8492 7260
rect 8426 7210 8442 7244
rect 8476 7210 8492 7244
rect 8252 7172 8282 7194
rect 8348 7172 8378 7198
rect 8426 7194 8492 7210
rect 8618 7244 8684 7260
rect 8618 7210 8634 7244
rect 8668 7210 8684 7244
rect 8444 7172 8474 7194
rect 8540 7172 8570 7198
rect 8618 7194 8684 7210
rect 8810 7244 8876 7260
rect 8810 7210 8826 7244
rect 8860 7210 8876 7244
rect 8636 7172 8666 7194
rect 8732 7172 8762 7198
rect 8810 7194 8876 7210
rect 9002 7244 9068 7260
rect 9002 7210 9018 7244
rect 9052 7210 9068 7244
rect 8828 7172 8858 7194
rect 8924 7172 8954 7198
rect 9002 7194 9068 7210
rect 9194 7244 9260 7260
rect 9194 7210 9210 7244
rect 9244 7210 9260 7244
rect 9020 7172 9050 7194
rect 9116 7172 9146 7198
rect 9194 7194 9260 7210
rect 9386 7244 9452 7260
rect 9386 7210 9402 7244
rect 9436 7210 9452 7244
rect 9212 7172 9242 7194
rect 9308 7172 9338 7198
rect 9386 7194 9452 7210
rect 9404 7172 9434 7194
rect 9500 7172 9530 7198
rect 7676 6746 7706 6772
rect 7772 6750 7802 6772
rect 7754 6734 7820 6750
rect 7868 6746 7898 6772
rect 7964 6750 7994 6772
rect 7754 6700 7770 6734
rect 7804 6700 7820 6734
rect 7754 6684 7820 6700
rect 7946 6734 8012 6750
rect 8060 6746 8090 6772
rect 8156 6750 8186 6772
rect 7946 6700 7962 6734
rect 7996 6700 8012 6734
rect 7946 6684 8012 6700
rect 8138 6734 8204 6750
rect 8252 6746 8282 6772
rect 8348 6750 8378 6772
rect 8138 6700 8154 6734
rect 8188 6700 8204 6734
rect 8138 6684 8204 6700
rect 8330 6734 8396 6750
rect 8444 6746 8474 6772
rect 8540 6750 8570 6772
rect 8330 6700 8346 6734
rect 8380 6700 8396 6734
rect 8330 6684 8396 6700
rect 8522 6734 8588 6750
rect 8636 6746 8666 6772
rect 8732 6750 8762 6772
rect 8522 6700 8538 6734
rect 8572 6700 8588 6734
rect 8522 6684 8588 6700
rect 8714 6734 8780 6750
rect 8828 6746 8858 6772
rect 8924 6750 8954 6772
rect 8714 6700 8730 6734
rect 8764 6700 8780 6734
rect 8714 6684 8780 6700
rect 8906 6734 8972 6750
rect 9020 6746 9050 6772
rect 9116 6750 9146 6772
rect 8906 6700 8922 6734
rect 8956 6700 8972 6734
rect 8906 6684 8972 6700
rect 9098 6734 9164 6750
rect 9212 6746 9242 6772
rect 9308 6750 9338 6772
rect 9098 6700 9114 6734
rect 9148 6700 9164 6734
rect 9098 6684 9164 6700
rect 9290 6734 9356 6750
rect 9404 6746 9434 6772
rect 9500 6750 9530 6772
rect 9290 6700 9306 6734
rect 9340 6700 9356 6734
rect 9290 6684 9356 6700
rect 9482 6734 9548 6750
rect 9482 6700 9498 6734
rect 9532 6700 9548 6734
rect 9482 6684 9548 6700
rect 7754 6626 7820 6642
rect 7754 6592 7770 6626
rect 7804 6592 7820 6626
rect 7676 6554 7706 6580
rect 7754 6576 7820 6592
rect 7946 6626 8012 6642
rect 7946 6592 7962 6626
rect 7996 6592 8012 6626
rect 7772 6554 7802 6576
rect 7868 6554 7898 6580
rect 7946 6576 8012 6592
rect 8138 6626 8204 6642
rect 8138 6592 8154 6626
rect 8188 6592 8204 6626
rect 7964 6554 7994 6576
rect 8060 6554 8090 6580
rect 8138 6576 8204 6592
rect 8330 6626 8396 6642
rect 8330 6592 8346 6626
rect 8380 6592 8396 6626
rect 8156 6554 8186 6576
rect 8252 6554 8282 6580
rect 8330 6576 8396 6592
rect 8522 6626 8588 6642
rect 8522 6592 8538 6626
rect 8572 6592 8588 6626
rect 8348 6554 8378 6576
rect 8444 6554 8474 6580
rect 8522 6576 8588 6592
rect 8714 6626 8780 6642
rect 8714 6592 8730 6626
rect 8764 6592 8780 6626
rect 8540 6554 8570 6576
rect 8636 6554 8666 6580
rect 8714 6576 8780 6592
rect 8906 6626 8972 6642
rect 8906 6592 8922 6626
rect 8956 6592 8972 6626
rect 8732 6554 8762 6576
rect 8828 6554 8858 6580
rect 8906 6576 8972 6592
rect 9098 6626 9164 6642
rect 9098 6592 9114 6626
rect 9148 6592 9164 6626
rect 8924 6554 8954 6576
rect 9020 6554 9050 6580
rect 9098 6576 9164 6592
rect 9290 6626 9356 6642
rect 9290 6592 9306 6626
rect 9340 6592 9356 6626
rect 9116 6554 9146 6576
rect 9212 6554 9242 6580
rect 9290 6576 9356 6592
rect 9482 6626 9548 6642
rect 9482 6592 9498 6626
rect 9532 6592 9548 6626
rect 9308 6554 9338 6576
rect 9404 6554 9434 6580
rect 9482 6576 9548 6592
rect 9500 6554 9530 6576
rect 7676 6132 7706 6154
rect 7658 6116 7724 6132
rect 7772 6128 7802 6154
rect 7868 6132 7898 6154
rect 7658 6082 7674 6116
rect 7708 6082 7724 6116
rect 7658 6066 7724 6082
rect 7850 6116 7916 6132
rect 7964 6128 7994 6154
rect 8060 6132 8090 6154
rect 7850 6082 7866 6116
rect 7900 6082 7916 6116
rect 7850 6066 7916 6082
rect 8042 6116 8108 6132
rect 8156 6128 8186 6154
rect 8252 6132 8282 6154
rect 8042 6082 8058 6116
rect 8092 6082 8108 6116
rect 8042 6066 8108 6082
rect 8234 6116 8300 6132
rect 8348 6128 8378 6154
rect 8444 6132 8474 6154
rect 8234 6082 8250 6116
rect 8284 6082 8300 6116
rect 8234 6066 8300 6082
rect 8426 6116 8492 6132
rect 8540 6128 8570 6154
rect 8636 6132 8666 6154
rect 8426 6082 8442 6116
rect 8476 6082 8492 6116
rect 8426 6066 8492 6082
rect 8618 6116 8684 6132
rect 8732 6128 8762 6154
rect 8828 6132 8858 6154
rect 8618 6082 8634 6116
rect 8668 6082 8684 6116
rect 8618 6066 8684 6082
rect 8810 6116 8876 6132
rect 8924 6128 8954 6154
rect 9020 6132 9050 6154
rect 8810 6082 8826 6116
rect 8860 6082 8876 6116
rect 8810 6066 8876 6082
rect 9002 6116 9068 6132
rect 9116 6128 9146 6154
rect 9212 6132 9242 6154
rect 9002 6082 9018 6116
rect 9052 6082 9068 6116
rect 9002 6066 9068 6082
rect 9194 6116 9260 6132
rect 9308 6128 9338 6154
rect 9404 6132 9434 6154
rect 9194 6082 9210 6116
rect 9244 6082 9260 6116
rect 9194 6066 9260 6082
rect 9386 6116 9452 6132
rect 9500 6128 9530 6154
rect 9386 6082 9402 6116
rect 9436 6082 9452 6116
rect 9386 6066 9452 6082
rect 7658 6008 7724 6024
rect 7658 5974 7674 6008
rect 7708 5974 7724 6008
rect 7658 5958 7724 5974
rect 7850 6008 7916 6024
rect 7850 5974 7866 6008
rect 7900 5974 7916 6008
rect 7676 5936 7706 5958
rect 7772 5936 7802 5962
rect 7850 5958 7916 5974
rect 8042 6008 8108 6024
rect 8042 5974 8058 6008
rect 8092 5974 8108 6008
rect 7868 5936 7898 5958
rect 7964 5936 7994 5962
rect 8042 5958 8108 5974
rect 8234 6008 8300 6024
rect 8234 5974 8250 6008
rect 8284 5974 8300 6008
rect 8060 5936 8090 5958
rect 8156 5936 8186 5962
rect 8234 5958 8300 5974
rect 8426 6008 8492 6024
rect 8426 5974 8442 6008
rect 8476 5974 8492 6008
rect 8252 5936 8282 5958
rect 8348 5936 8378 5962
rect 8426 5958 8492 5974
rect 8618 6008 8684 6024
rect 8618 5974 8634 6008
rect 8668 5974 8684 6008
rect 8444 5936 8474 5958
rect 8540 5936 8570 5962
rect 8618 5958 8684 5974
rect 8810 6008 8876 6024
rect 8810 5974 8826 6008
rect 8860 5974 8876 6008
rect 8636 5936 8666 5958
rect 8732 5936 8762 5962
rect 8810 5958 8876 5974
rect 9002 6008 9068 6024
rect 9002 5974 9018 6008
rect 9052 5974 9068 6008
rect 8828 5936 8858 5958
rect 8924 5936 8954 5962
rect 9002 5958 9068 5974
rect 9194 6008 9260 6024
rect 9194 5974 9210 6008
rect 9244 5974 9260 6008
rect 9020 5936 9050 5958
rect 9116 5936 9146 5962
rect 9194 5958 9260 5974
rect 9386 6008 9452 6024
rect 9386 5974 9402 6008
rect 9436 5974 9452 6008
rect 9212 5936 9242 5958
rect 9308 5936 9338 5962
rect 9386 5958 9452 5974
rect 9404 5936 9434 5958
rect 9500 5936 9530 5962
rect 7676 5510 7706 5536
rect 7772 5514 7802 5536
rect 7754 5498 7820 5514
rect 7868 5510 7898 5536
rect 7964 5514 7994 5536
rect 7754 5464 7770 5498
rect 7804 5464 7820 5498
rect 7754 5448 7820 5464
rect 7946 5498 8012 5514
rect 8060 5510 8090 5536
rect 8156 5514 8186 5536
rect 7946 5464 7962 5498
rect 7996 5464 8012 5498
rect 7946 5448 8012 5464
rect 8138 5498 8204 5514
rect 8252 5510 8282 5536
rect 8348 5514 8378 5536
rect 8138 5464 8154 5498
rect 8188 5464 8204 5498
rect 8138 5448 8204 5464
rect 8330 5498 8396 5514
rect 8444 5510 8474 5536
rect 8540 5514 8570 5536
rect 8330 5464 8346 5498
rect 8380 5464 8396 5498
rect 8330 5448 8396 5464
rect 8522 5498 8588 5514
rect 8636 5510 8666 5536
rect 8732 5514 8762 5536
rect 8522 5464 8538 5498
rect 8572 5464 8588 5498
rect 8522 5448 8588 5464
rect 8714 5498 8780 5514
rect 8828 5510 8858 5536
rect 8924 5514 8954 5536
rect 8714 5464 8730 5498
rect 8764 5464 8780 5498
rect 8714 5448 8780 5464
rect 8906 5498 8972 5514
rect 9020 5510 9050 5536
rect 9116 5514 9146 5536
rect 8906 5464 8922 5498
rect 8956 5464 8972 5498
rect 8906 5448 8972 5464
rect 9098 5498 9164 5514
rect 9212 5510 9242 5536
rect 9308 5514 9338 5536
rect 9098 5464 9114 5498
rect 9148 5464 9164 5498
rect 9098 5448 9164 5464
rect 9290 5498 9356 5514
rect 9404 5510 9434 5536
rect 9500 5514 9530 5536
rect 9290 5464 9306 5498
rect 9340 5464 9356 5498
rect 9290 5448 9356 5464
rect 9482 5498 9548 5514
rect 9482 5464 9498 5498
rect 9532 5464 9548 5498
rect 9482 5448 9548 5464
rect 7754 5390 7820 5406
rect 7754 5356 7770 5390
rect 7804 5356 7820 5390
rect 7676 5318 7706 5344
rect 7754 5340 7820 5356
rect 7946 5390 8012 5406
rect 7946 5356 7962 5390
rect 7996 5356 8012 5390
rect 7772 5318 7802 5340
rect 7868 5318 7898 5344
rect 7946 5340 8012 5356
rect 8138 5390 8204 5406
rect 8138 5356 8154 5390
rect 8188 5356 8204 5390
rect 7964 5318 7994 5340
rect 8060 5318 8090 5344
rect 8138 5340 8204 5356
rect 8330 5390 8396 5406
rect 8330 5356 8346 5390
rect 8380 5356 8396 5390
rect 8156 5318 8186 5340
rect 8252 5318 8282 5344
rect 8330 5340 8396 5356
rect 8522 5390 8588 5406
rect 8522 5356 8538 5390
rect 8572 5356 8588 5390
rect 8348 5318 8378 5340
rect 8444 5318 8474 5344
rect 8522 5340 8588 5356
rect 8714 5390 8780 5406
rect 8714 5356 8730 5390
rect 8764 5356 8780 5390
rect 8540 5318 8570 5340
rect 8636 5318 8666 5344
rect 8714 5340 8780 5356
rect 8906 5390 8972 5406
rect 8906 5356 8922 5390
rect 8956 5356 8972 5390
rect 8732 5318 8762 5340
rect 8828 5318 8858 5344
rect 8906 5340 8972 5356
rect 9098 5390 9164 5406
rect 9098 5356 9114 5390
rect 9148 5356 9164 5390
rect 8924 5318 8954 5340
rect 9020 5318 9050 5344
rect 9098 5340 9164 5356
rect 9290 5390 9356 5406
rect 9290 5356 9306 5390
rect 9340 5356 9356 5390
rect 9116 5318 9146 5340
rect 9212 5318 9242 5344
rect 9290 5340 9356 5356
rect 9482 5390 9548 5406
rect 9482 5356 9498 5390
rect 9532 5356 9548 5390
rect 9308 5318 9338 5340
rect 9404 5318 9434 5344
rect 9482 5340 9548 5356
rect 9500 5318 9530 5340
rect 7676 4896 7706 4918
rect 7658 4880 7724 4896
rect 7772 4892 7802 4918
rect 7868 4896 7898 4918
rect 7658 4846 7674 4880
rect 7708 4846 7724 4880
rect 7658 4830 7724 4846
rect 7850 4880 7916 4896
rect 7964 4892 7994 4918
rect 8060 4896 8090 4918
rect 7850 4846 7866 4880
rect 7900 4846 7916 4880
rect 7850 4830 7916 4846
rect 8042 4880 8108 4896
rect 8156 4892 8186 4918
rect 8252 4896 8282 4918
rect 8042 4846 8058 4880
rect 8092 4846 8108 4880
rect 8042 4830 8108 4846
rect 8234 4880 8300 4896
rect 8348 4892 8378 4918
rect 8444 4896 8474 4918
rect 8234 4846 8250 4880
rect 8284 4846 8300 4880
rect 8234 4830 8300 4846
rect 8426 4880 8492 4896
rect 8540 4892 8570 4918
rect 8636 4896 8666 4918
rect 8426 4846 8442 4880
rect 8476 4846 8492 4880
rect 8426 4830 8492 4846
rect 8618 4880 8684 4896
rect 8732 4892 8762 4918
rect 8828 4896 8858 4918
rect 8618 4846 8634 4880
rect 8668 4846 8684 4880
rect 8618 4830 8684 4846
rect 8810 4880 8876 4896
rect 8924 4892 8954 4918
rect 9020 4896 9050 4918
rect 8810 4846 8826 4880
rect 8860 4846 8876 4880
rect 8810 4830 8876 4846
rect 9002 4880 9068 4896
rect 9116 4892 9146 4918
rect 9212 4896 9242 4918
rect 9002 4846 9018 4880
rect 9052 4846 9068 4880
rect 9002 4830 9068 4846
rect 9194 4880 9260 4896
rect 9308 4892 9338 4918
rect 9404 4896 9434 4918
rect 9194 4846 9210 4880
rect 9244 4846 9260 4880
rect 9194 4830 9260 4846
rect 9386 4880 9452 4896
rect 9500 4892 9530 4918
rect 9386 4846 9402 4880
rect 9436 4846 9452 4880
rect 9386 4830 9452 4846
rect 16218 8802 16284 8818
rect 16218 8768 16234 8802
rect 16268 8768 16284 8802
rect 16140 8730 16170 8756
rect 16218 8752 16284 8768
rect 16410 8802 16476 8818
rect 16410 8768 16426 8802
rect 16460 8768 16476 8802
rect 16236 8730 16266 8752
rect 16332 8730 16362 8756
rect 16410 8752 16476 8768
rect 16602 8802 16668 8818
rect 16602 8768 16618 8802
rect 16652 8768 16668 8802
rect 16428 8730 16458 8752
rect 16524 8730 16554 8756
rect 16602 8752 16668 8768
rect 16794 8802 16860 8818
rect 16794 8768 16810 8802
rect 16844 8768 16860 8802
rect 16620 8730 16650 8752
rect 16716 8730 16746 8756
rect 16794 8752 16860 8768
rect 16986 8802 17052 8818
rect 16986 8768 17002 8802
rect 17036 8768 17052 8802
rect 16812 8730 16842 8752
rect 16908 8730 16938 8756
rect 16986 8752 17052 8768
rect 17178 8802 17244 8818
rect 17178 8768 17194 8802
rect 17228 8768 17244 8802
rect 17004 8730 17034 8752
rect 17100 8730 17130 8756
rect 17178 8752 17244 8768
rect 17370 8802 17436 8818
rect 17370 8768 17386 8802
rect 17420 8768 17436 8802
rect 17196 8730 17226 8752
rect 17292 8730 17322 8756
rect 17370 8752 17436 8768
rect 17562 8802 17628 8818
rect 17562 8768 17578 8802
rect 17612 8768 17628 8802
rect 17388 8730 17418 8752
rect 17484 8730 17514 8756
rect 17562 8752 17628 8768
rect 17754 8802 17820 8818
rect 17754 8768 17770 8802
rect 17804 8768 17820 8802
rect 17580 8730 17610 8752
rect 17676 8730 17706 8756
rect 17754 8752 17820 8768
rect 17946 8802 18012 8818
rect 17946 8768 17962 8802
rect 17996 8768 18012 8802
rect 17772 8730 17802 8752
rect 17868 8730 17898 8756
rect 17946 8752 18012 8768
rect 17964 8730 17994 8752
rect 16140 8308 16170 8330
rect 16122 8292 16188 8308
rect 16236 8304 16266 8330
rect 16332 8308 16362 8330
rect 16122 8258 16138 8292
rect 16172 8258 16188 8292
rect 16122 8242 16188 8258
rect 16314 8292 16380 8308
rect 16428 8304 16458 8330
rect 16524 8308 16554 8330
rect 16314 8258 16330 8292
rect 16364 8258 16380 8292
rect 16314 8242 16380 8258
rect 16506 8292 16572 8308
rect 16620 8304 16650 8330
rect 16716 8308 16746 8330
rect 16506 8258 16522 8292
rect 16556 8258 16572 8292
rect 16506 8242 16572 8258
rect 16698 8292 16764 8308
rect 16812 8304 16842 8330
rect 16908 8308 16938 8330
rect 16698 8258 16714 8292
rect 16748 8258 16764 8292
rect 16698 8242 16764 8258
rect 16890 8292 16956 8308
rect 17004 8304 17034 8330
rect 17100 8308 17130 8330
rect 16890 8258 16906 8292
rect 16940 8258 16956 8292
rect 16890 8242 16956 8258
rect 17082 8292 17148 8308
rect 17196 8304 17226 8330
rect 17292 8308 17322 8330
rect 17082 8258 17098 8292
rect 17132 8258 17148 8292
rect 17082 8242 17148 8258
rect 17274 8292 17340 8308
rect 17388 8304 17418 8330
rect 17484 8308 17514 8330
rect 17274 8258 17290 8292
rect 17324 8258 17340 8292
rect 17274 8242 17340 8258
rect 17466 8292 17532 8308
rect 17580 8304 17610 8330
rect 17676 8308 17706 8330
rect 17466 8258 17482 8292
rect 17516 8258 17532 8292
rect 17466 8242 17532 8258
rect 17658 8292 17724 8308
rect 17772 8304 17802 8330
rect 17868 8308 17898 8330
rect 17658 8258 17674 8292
rect 17708 8258 17724 8292
rect 17658 8242 17724 8258
rect 17850 8292 17916 8308
rect 17964 8304 17994 8330
rect 17850 8258 17866 8292
rect 17900 8258 17916 8292
rect 17850 8242 17916 8258
rect 16218 7982 16284 7998
rect 16218 7948 16234 7982
rect 16268 7948 16284 7982
rect 16140 7910 16170 7936
rect 16218 7932 16284 7948
rect 16410 7982 16476 7998
rect 16410 7948 16426 7982
rect 16460 7948 16476 7982
rect 16236 7910 16266 7932
rect 16332 7910 16362 7936
rect 16410 7932 16476 7948
rect 16602 7982 16668 7998
rect 16602 7948 16618 7982
rect 16652 7948 16668 7982
rect 16428 7910 16458 7932
rect 16524 7910 16554 7936
rect 16602 7932 16668 7948
rect 16794 7982 16860 7998
rect 16794 7948 16810 7982
rect 16844 7948 16860 7982
rect 16620 7910 16650 7932
rect 16716 7910 16746 7936
rect 16794 7932 16860 7948
rect 16986 7982 17052 7998
rect 16986 7948 17002 7982
rect 17036 7948 17052 7982
rect 16812 7910 16842 7932
rect 16908 7910 16938 7936
rect 16986 7932 17052 7948
rect 17178 7982 17244 7998
rect 17178 7948 17194 7982
rect 17228 7948 17244 7982
rect 17004 7910 17034 7932
rect 17100 7910 17130 7936
rect 17178 7932 17244 7948
rect 17370 7982 17436 7998
rect 17370 7948 17386 7982
rect 17420 7948 17436 7982
rect 17196 7910 17226 7932
rect 17292 7910 17322 7936
rect 17370 7932 17436 7948
rect 17562 7982 17628 7998
rect 17562 7948 17578 7982
rect 17612 7948 17628 7982
rect 17388 7910 17418 7932
rect 17484 7910 17514 7936
rect 17562 7932 17628 7948
rect 17754 7982 17820 7998
rect 17754 7948 17770 7982
rect 17804 7948 17820 7982
rect 17580 7910 17610 7932
rect 17676 7910 17706 7936
rect 17754 7932 17820 7948
rect 17946 7982 18012 7998
rect 17946 7948 17962 7982
rect 17996 7948 18012 7982
rect 17772 7910 17802 7932
rect 17868 7910 17898 7936
rect 17946 7932 18012 7948
rect 17964 7910 17994 7932
rect 16140 7488 16170 7510
rect 16122 7472 16188 7488
rect 16236 7484 16266 7510
rect 16332 7488 16362 7510
rect 16122 7438 16138 7472
rect 16172 7438 16188 7472
rect 16122 7422 16188 7438
rect 16314 7472 16380 7488
rect 16428 7484 16458 7510
rect 16524 7488 16554 7510
rect 16314 7438 16330 7472
rect 16364 7438 16380 7472
rect 16314 7422 16380 7438
rect 16506 7472 16572 7488
rect 16620 7484 16650 7510
rect 16716 7488 16746 7510
rect 16506 7438 16522 7472
rect 16556 7438 16572 7472
rect 16506 7422 16572 7438
rect 16698 7472 16764 7488
rect 16812 7484 16842 7510
rect 16908 7488 16938 7510
rect 16698 7438 16714 7472
rect 16748 7438 16764 7472
rect 16698 7422 16764 7438
rect 16890 7472 16956 7488
rect 17004 7484 17034 7510
rect 17100 7488 17130 7510
rect 16890 7438 16906 7472
rect 16940 7438 16956 7472
rect 16890 7422 16956 7438
rect 17082 7472 17148 7488
rect 17196 7484 17226 7510
rect 17292 7488 17322 7510
rect 17082 7438 17098 7472
rect 17132 7438 17148 7472
rect 17082 7422 17148 7438
rect 17274 7472 17340 7488
rect 17388 7484 17418 7510
rect 17484 7488 17514 7510
rect 17274 7438 17290 7472
rect 17324 7438 17340 7472
rect 17274 7422 17340 7438
rect 17466 7472 17532 7488
rect 17580 7484 17610 7510
rect 17676 7488 17706 7510
rect 17466 7438 17482 7472
rect 17516 7438 17532 7472
rect 17466 7422 17532 7438
rect 17658 7472 17724 7488
rect 17772 7484 17802 7510
rect 17868 7488 17898 7510
rect 17658 7438 17674 7472
rect 17708 7438 17724 7472
rect 17658 7422 17724 7438
rect 17850 7472 17916 7488
rect 17964 7484 17994 7510
rect 17850 7438 17866 7472
rect 17900 7438 17916 7472
rect 17850 7422 17916 7438
rect 16218 7162 16284 7178
rect 16218 7128 16234 7162
rect 16268 7128 16284 7162
rect 16140 7090 16170 7116
rect 16218 7112 16284 7128
rect 16410 7162 16476 7178
rect 16410 7128 16426 7162
rect 16460 7128 16476 7162
rect 16236 7090 16266 7112
rect 16332 7090 16362 7116
rect 16410 7112 16476 7128
rect 16602 7162 16668 7178
rect 16602 7128 16618 7162
rect 16652 7128 16668 7162
rect 16428 7090 16458 7112
rect 16524 7090 16554 7116
rect 16602 7112 16668 7128
rect 16794 7162 16860 7178
rect 16794 7128 16810 7162
rect 16844 7128 16860 7162
rect 16620 7090 16650 7112
rect 16716 7090 16746 7116
rect 16794 7112 16860 7128
rect 16986 7162 17052 7178
rect 16986 7128 17002 7162
rect 17036 7128 17052 7162
rect 16812 7090 16842 7112
rect 16908 7090 16938 7116
rect 16986 7112 17052 7128
rect 17178 7162 17244 7178
rect 17178 7128 17194 7162
rect 17228 7128 17244 7162
rect 17004 7090 17034 7112
rect 17100 7090 17130 7116
rect 17178 7112 17244 7128
rect 17370 7162 17436 7178
rect 17370 7128 17386 7162
rect 17420 7128 17436 7162
rect 17196 7090 17226 7112
rect 17292 7090 17322 7116
rect 17370 7112 17436 7128
rect 17562 7162 17628 7178
rect 17562 7128 17578 7162
rect 17612 7128 17628 7162
rect 17388 7090 17418 7112
rect 17484 7090 17514 7116
rect 17562 7112 17628 7128
rect 17754 7162 17820 7178
rect 17754 7128 17770 7162
rect 17804 7128 17820 7162
rect 17580 7090 17610 7112
rect 17676 7090 17706 7116
rect 17754 7112 17820 7128
rect 17946 7162 18012 7178
rect 17946 7128 17962 7162
rect 17996 7128 18012 7162
rect 17772 7090 17802 7112
rect 17868 7090 17898 7116
rect 17946 7112 18012 7128
rect 17964 7090 17994 7112
rect 16140 6668 16170 6690
rect 16122 6652 16188 6668
rect 16236 6664 16266 6690
rect 16332 6668 16362 6690
rect 16122 6618 16138 6652
rect 16172 6618 16188 6652
rect 16122 6602 16188 6618
rect 16314 6652 16380 6668
rect 16428 6664 16458 6690
rect 16524 6668 16554 6690
rect 16314 6618 16330 6652
rect 16364 6618 16380 6652
rect 16314 6602 16380 6618
rect 16506 6652 16572 6668
rect 16620 6664 16650 6690
rect 16716 6668 16746 6690
rect 16506 6618 16522 6652
rect 16556 6618 16572 6652
rect 16506 6602 16572 6618
rect 16698 6652 16764 6668
rect 16812 6664 16842 6690
rect 16908 6668 16938 6690
rect 16698 6618 16714 6652
rect 16748 6618 16764 6652
rect 16698 6602 16764 6618
rect 16890 6652 16956 6668
rect 17004 6664 17034 6690
rect 17100 6668 17130 6690
rect 16890 6618 16906 6652
rect 16940 6618 16956 6652
rect 16890 6602 16956 6618
rect 17082 6652 17148 6668
rect 17196 6664 17226 6690
rect 17292 6668 17322 6690
rect 17082 6618 17098 6652
rect 17132 6618 17148 6652
rect 17082 6602 17148 6618
rect 17274 6652 17340 6668
rect 17388 6664 17418 6690
rect 17484 6668 17514 6690
rect 17274 6618 17290 6652
rect 17324 6618 17340 6652
rect 17274 6602 17340 6618
rect 17466 6652 17532 6668
rect 17580 6664 17610 6690
rect 17676 6668 17706 6690
rect 17466 6618 17482 6652
rect 17516 6618 17532 6652
rect 17466 6602 17532 6618
rect 17658 6652 17724 6668
rect 17772 6664 17802 6690
rect 17868 6668 17898 6690
rect 17658 6618 17674 6652
rect 17708 6618 17724 6652
rect 17658 6602 17724 6618
rect 17850 6652 17916 6668
rect 17964 6664 17994 6690
rect 17850 6618 17866 6652
rect 17900 6618 17916 6652
rect 17850 6602 17916 6618
rect 19558 10364 19624 10380
rect 19558 10330 19574 10364
rect 19608 10330 19624 10364
rect 19558 10314 19624 10330
rect 19750 10364 19816 10380
rect 19750 10330 19766 10364
rect 19800 10330 19816 10364
rect 19750 10314 19816 10330
rect 19942 10364 20008 10380
rect 19942 10330 19958 10364
rect 19992 10330 20008 10364
rect 19942 10314 20008 10330
rect 20134 10364 20200 10380
rect 20134 10330 20150 10364
rect 20184 10330 20200 10364
rect 20134 10314 20200 10330
rect 20326 10364 20392 10380
rect 20326 10330 20342 10364
rect 20376 10330 20392 10364
rect 20326 10314 20392 10330
rect 20518 10364 20584 10380
rect 20518 10330 20534 10364
rect 20568 10330 20584 10364
rect 20518 10314 20584 10330
rect 20710 10364 20776 10380
rect 20710 10330 20726 10364
rect 20760 10330 20776 10364
rect 20710 10314 20776 10330
rect 20902 10364 20968 10380
rect 20902 10330 20918 10364
rect 20952 10330 20968 10364
rect 20902 10314 20968 10330
rect 21094 10364 21160 10380
rect 21094 10330 21110 10364
rect 21144 10330 21160 10364
rect 21094 10314 21160 10330
rect 21286 10364 21352 10380
rect 21286 10330 21302 10364
rect 21336 10330 21352 10364
rect 21286 10314 21352 10330
rect 19576 10283 19606 10314
rect 19672 10283 19702 10309
rect 19768 10283 19798 10314
rect 19864 10283 19894 10309
rect 19960 10283 19990 10314
rect 20056 10283 20086 10309
rect 20152 10283 20182 10314
rect 20248 10283 20278 10309
rect 20344 10283 20374 10314
rect 20440 10283 20470 10309
rect 20536 10283 20566 10314
rect 20632 10283 20662 10309
rect 20728 10283 20758 10314
rect 20824 10283 20854 10309
rect 20920 10283 20950 10314
rect 21016 10283 21046 10309
rect 21112 10283 21142 10314
rect 21208 10283 21238 10309
rect 21304 10283 21334 10314
rect 21400 10283 21430 10309
rect 19576 9857 19606 9883
rect 19672 9852 19702 9883
rect 19768 9857 19798 9883
rect 19864 9852 19894 9883
rect 19960 9857 19990 9883
rect 20056 9852 20086 9883
rect 20152 9857 20182 9883
rect 20248 9852 20278 9883
rect 20344 9857 20374 9883
rect 20440 9852 20470 9883
rect 20536 9857 20566 9883
rect 20632 9852 20662 9883
rect 20728 9857 20758 9883
rect 20824 9852 20854 9883
rect 20920 9857 20950 9883
rect 21016 9852 21046 9883
rect 21112 9857 21142 9883
rect 21208 9852 21238 9883
rect 21304 9857 21334 9883
rect 21400 9852 21430 9883
rect 19654 9836 19720 9852
rect 19654 9802 19670 9836
rect 19704 9802 19720 9836
rect 19654 9786 19720 9802
rect 19846 9836 19912 9852
rect 19846 9802 19862 9836
rect 19896 9802 19912 9836
rect 19846 9786 19912 9802
rect 20038 9836 20104 9852
rect 20038 9802 20054 9836
rect 20088 9802 20104 9836
rect 20038 9786 20104 9802
rect 20230 9836 20296 9852
rect 20230 9802 20246 9836
rect 20280 9802 20296 9836
rect 20230 9786 20296 9802
rect 20422 9836 20488 9852
rect 20422 9802 20438 9836
rect 20472 9802 20488 9836
rect 20422 9786 20488 9802
rect 20614 9836 20680 9852
rect 20614 9802 20630 9836
rect 20664 9802 20680 9836
rect 20614 9786 20680 9802
rect 20806 9836 20872 9852
rect 20806 9802 20822 9836
rect 20856 9802 20872 9836
rect 20806 9786 20872 9802
rect 20998 9836 21064 9852
rect 20998 9802 21014 9836
rect 21048 9802 21064 9836
rect 20998 9786 21064 9802
rect 21190 9836 21256 9852
rect 21190 9802 21206 9836
rect 21240 9802 21256 9836
rect 21190 9786 21256 9802
rect 21382 9836 21448 9852
rect 21382 9802 21398 9836
rect 21432 9802 21448 9836
rect 21382 9786 21448 9802
rect 19654 9728 19720 9744
rect 19654 9694 19670 9728
rect 19704 9694 19720 9728
rect 19654 9678 19720 9694
rect 19846 9728 19912 9744
rect 19846 9694 19862 9728
rect 19896 9694 19912 9728
rect 19846 9678 19912 9694
rect 20038 9728 20104 9744
rect 20038 9694 20054 9728
rect 20088 9694 20104 9728
rect 20038 9678 20104 9694
rect 20230 9728 20296 9744
rect 20230 9694 20246 9728
rect 20280 9694 20296 9728
rect 20230 9678 20296 9694
rect 20422 9728 20488 9744
rect 20422 9694 20438 9728
rect 20472 9694 20488 9728
rect 20422 9678 20488 9694
rect 20614 9728 20680 9744
rect 20614 9694 20630 9728
rect 20664 9694 20680 9728
rect 20614 9678 20680 9694
rect 20806 9728 20872 9744
rect 20806 9694 20822 9728
rect 20856 9694 20872 9728
rect 20806 9678 20872 9694
rect 20998 9728 21064 9744
rect 20998 9694 21014 9728
rect 21048 9694 21064 9728
rect 20998 9678 21064 9694
rect 21190 9728 21256 9744
rect 21190 9694 21206 9728
rect 21240 9694 21256 9728
rect 21190 9678 21256 9694
rect 21382 9728 21448 9744
rect 21382 9694 21398 9728
rect 21432 9694 21448 9728
rect 21382 9678 21448 9694
rect 19576 9647 19606 9673
rect 19672 9647 19702 9678
rect 19768 9647 19798 9673
rect 19864 9647 19894 9678
rect 19960 9647 19990 9673
rect 20056 9647 20086 9678
rect 20152 9647 20182 9673
rect 20248 9647 20278 9678
rect 20344 9647 20374 9673
rect 20440 9647 20470 9678
rect 20536 9647 20566 9673
rect 20632 9647 20662 9678
rect 20728 9647 20758 9673
rect 20824 9647 20854 9678
rect 20920 9647 20950 9673
rect 21016 9647 21046 9678
rect 21112 9647 21142 9673
rect 21208 9647 21238 9678
rect 21304 9647 21334 9673
rect 21400 9647 21430 9678
rect 19576 9216 19606 9247
rect 19672 9221 19702 9247
rect 19768 9216 19798 9247
rect 19864 9221 19894 9247
rect 19960 9216 19990 9247
rect 20056 9221 20086 9247
rect 20152 9216 20182 9247
rect 20248 9221 20278 9247
rect 20344 9216 20374 9247
rect 20440 9221 20470 9247
rect 20536 9216 20566 9247
rect 20632 9221 20662 9247
rect 20728 9216 20758 9247
rect 20824 9221 20854 9247
rect 20920 9216 20950 9247
rect 21016 9221 21046 9247
rect 21112 9216 21142 9247
rect 21208 9221 21238 9247
rect 21304 9216 21334 9247
rect 21400 9221 21430 9247
rect 19558 9200 19624 9216
rect 19558 9166 19574 9200
rect 19608 9166 19624 9200
rect 19558 9150 19624 9166
rect 19750 9200 19816 9216
rect 19750 9166 19766 9200
rect 19800 9166 19816 9200
rect 19750 9150 19816 9166
rect 19942 9200 20008 9216
rect 19942 9166 19958 9200
rect 19992 9166 20008 9200
rect 19942 9150 20008 9166
rect 20134 9200 20200 9216
rect 20134 9166 20150 9200
rect 20184 9166 20200 9200
rect 20134 9150 20200 9166
rect 20326 9200 20392 9216
rect 20326 9166 20342 9200
rect 20376 9166 20392 9200
rect 20326 9150 20392 9166
rect 20518 9200 20584 9216
rect 20518 9166 20534 9200
rect 20568 9166 20584 9200
rect 20518 9150 20584 9166
rect 20710 9200 20776 9216
rect 20710 9166 20726 9200
rect 20760 9166 20776 9200
rect 20710 9150 20776 9166
rect 20902 9200 20968 9216
rect 20902 9166 20918 9200
rect 20952 9166 20968 9200
rect 20902 9150 20968 9166
rect 21094 9200 21160 9216
rect 21094 9166 21110 9200
rect 21144 9166 21160 9200
rect 21094 9150 21160 9166
rect 21286 9200 21352 9216
rect 21286 9166 21302 9200
rect 21336 9166 21352 9200
rect 21286 9150 21352 9166
rect 19558 8768 19624 8784
rect 19558 8734 19574 8768
rect 19608 8734 19624 8768
rect 19558 8718 19624 8734
rect 19750 8768 19816 8784
rect 19750 8734 19766 8768
rect 19800 8734 19816 8768
rect 19576 8696 19606 8718
rect 19672 8696 19702 8722
rect 19750 8718 19816 8734
rect 19942 8768 20008 8784
rect 19942 8734 19958 8768
rect 19992 8734 20008 8768
rect 19768 8696 19798 8718
rect 19864 8696 19894 8722
rect 19942 8718 20008 8734
rect 20134 8768 20200 8784
rect 20134 8734 20150 8768
rect 20184 8734 20200 8768
rect 19960 8696 19990 8718
rect 20056 8696 20086 8722
rect 20134 8718 20200 8734
rect 20326 8768 20392 8784
rect 20326 8734 20342 8768
rect 20376 8734 20392 8768
rect 20152 8696 20182 8718
rect 20248 8696 20278 8722
rect 20326 8718 20392 8734
rect 20518 8768 20584 8784
rect 20518 8734 20534 8768
rect 20568 8734 20584 8768
rect 20344 8696 20374 8718
rect 20440 8696 20470 8722
rect 20518 8718 20584 8734
rect 20710 8768 20776 8784
rect 20710 8734 20726 8768
rect 20760 8734 20776 8768
rect 20536 8696 20566 8718
rect 20632 8696 20662 8722
rect 20710 8718 20776 8734
rect 20902 8768 20968 8784
rect 20902 8734 20918 8768
rect 20952 8734 20968 8768
rect 20728 8696 20758 8718
rect 20824 8696 20854 8722
rect 20902 8718 20968 8734
rect 21094 8768 21160 8784
rect 21094 8734 21110 8768
rect 21144 8734 21160 8768
rect 20920 8696 20950 8718
rect 21016 8696 21046 8722
rect 21094 8718 21160 8734
rect 21286 8768 21352 8784
rect 21286 8734 21302 8768
rect 21336 8734 21352 8768
rect 21112 8696 21142 8718
rect 21208 8696 21238 8722
rect 21286 8718 21352 8734
rect 21304 8696 21334 8718
rect 21400 8696 21430 8722
rect 19576 8270 19606 8296
rect 19672 8274 19702 8296
rect 19654 8258 19720 8274
rect 19768 8270 19798 8296
rect 19864 8274 19894 8296
rect 19654 8224 19670 8258
rect 19704 8224 19720 8258
rect 19654 8208 19720 8224
rect 19846 8258 19912 8274
rect 19960 8270 19990 8296
rect 20056 8274 20086 8296
rect 19846 8224 19862 8258
rect 19896 8224 19912 8258
rect 19846 8208 19912 8224
rect 20038 8258 20104 8274
rect 20152 8270 20182 8296
rect 20248 8274 20278 8296
rect 20038 8224 20054 8258
rect 20088 8224 20104 8258
rect 20038 8208 20104 8224
rect 20230 8258 20296 8274
rect 20344 8270 20374 8296
rect 20440 8274 20470 8296
rect 20230 8224 20246 8258
rect 20280 8224 20296 8258
rect 20230 8208 20296 8224
rect 20422 8258 20488 8274
rect 20536 8270 20566 8296
rect 20632 8274 20662 8296
rect 20422 8224 20438 8258
rect 20472 8224 20488 8258
rect 20422 8208 20488 8224
rect 20614 8258 20680 8274
rect 20728 8270 20758 8296
rect 20824 8274 20854 8296
rect 20614 8224 20630 8258
rect 20664 8224 20680 8258
rect 20614 8208 20680 8224
rect 20806 8258 20872 8274
rect 20920 8270 20950 8296
rect 21016 8274 21046 8296
rect 20806 8224 20822 8258
rect 20856 8224 20872 8258
rect 20806 8208 20872 8224
rect 20998 8258 21064 8274
rect 21112 8270 21142 8296
rect 21208 8274 21238 8296
rect 20998 8224 21014 8258
rect 21048 8224 21064 8258
rect 20998 8208 21064 8224
rect 21190 8258 21256 8274
rect 21304 8270 21334 8296
rect 21400 8274 21430 8296
rect 21190 8224 21206 8258
rect 21240 8224 21256 8258
rect 21190 8208 21256 8224
rect 21382 8258 21448 8274
rect 21382 8224 21398 8258
rect 21432 8224 21448 8258
rect 21382 8208 21448 8224
rect 19654 8150 19720 8166
rect 19654 8116 19670 8150
rect 19704 8116 19720 8150
rect 19576 8078 19606 8104
rect 19654 8100 19720 8116
rect 19846 8150 19912 8166
rect 19846 8116 19862 8150
rect 19896 8116 19912 8150
rect 19672 8078 19702 8100
rect 19768 8078 19798 8104
rect 19846 8100 19912 8116
rect 20038 8150 20104 8166
rect 20038 8116 20054 8150
rect 20088 8116 20104 8150
rect 19864 8078 19894 8100
rect 19960 8078 19990 8104
rect 20038 8100 20104 8116
rect 20230 8150 20296 8166
rect 20230 8116 20246 8150
rect 20280 8116 20296 8150
rect 20056 8078 20086 8100
rect 20152 8078 20182 8104
rect 20230 8100 20296 8116
rect 20422 8150 20488 8166
rect 20422 8116 20438 8150
rect 20472 8116 20488 8150
rect 20248 8078 20278 8100
rect 20344 8078 20374 8104
rect 20422 8100 20488 8116
rect 20614 8150 20680 8166
rect 20614 8116 20630 8150
rect 20664 8116 20680 8150
rect 20440 8078 20470 8100
rect 20536 8078 20566 8104
rect 20614 8100 20680 8116
rect 20806 8150 20872 8166
rect 20806 8116 20822 8150
rect 20856 8116 20872 8150
rect 20632 8078 20662 8100
rect 20728 8078 20758 8104
rect 20806 8100 20872 8116
rect 20998 8150 21064 8166
rect 20998 8116 21014 8150
rect 21048 8116 21064 8150
rect 20824 8078 20854 8100
rect 20920 8078 20950 8104
rect 20998 8100 21064 8116
rect 21190 8150 21256 8166
rect 21190 8116 21206 8150
rect 21240 8116 21256 8150
rect 21016 8078 21046 8100
rect 21112 8078 21142 8104
rect 21190 8100 21256 8116
rect 21382 8150 21448 8166
rect 21382 8116 21398 8150
rect 21432 8116 21448 8150
rect 21208 8078 21238 8100
rect 21304 8078 21334 8104
rect 21382 8100 21448 8116
rect 21400 8078 21430 8100
rect 19576 7656 19606 7678
rect 19558 7640 19624 7656
rect 19672 7652 19702 7678
rect 19768 7656 19798 7678
rect 19558 7606 19574 7640
rect 19608 7606 19624 7640
rect 19558 7590 19624 7606
rect 19750 7640 19816 7656
rect 19864 7652 19894 7678
rect 19960 7656 19990 7678
rect 19750 7606 19766 7640
rect 19800 7606 19816 7640
rect 19750 7590 19816 7606
rect 19942 7640 20008 7656
rect 20056 7652 20086 7678
rect 20152 7656 20182 7678
rect 19942 7606 19958 7640
rect 19992 7606 20008 7640
rect 19942 7590 20008 7606
rect 20134 7640 20200 7656
rect 20248 7652 20278 7678
rect 20344 7656 20374 7678
rect 20134 7606 20150 7640
rect 20184 7606 20200 7640
rect 20134 7590 20200 7606
rect 20326 7640 20392 7656
rect 20440 7652 20470 7678
rect 20536 7656 20566 7678
rect 20326 7606 20342 7640
rect 20376 7606 20392 7640
rect 20326 7590 20392 7606
rect 20518 7640 20584 7656
rect 20632 7652 20662 7678
rect 20728 7656 20758 7678
rect 20518 7606 20534 7640
rect 20568 7606 20584 7640
rect 20518 7590 20584 7606
rect 20710 7640 20776 7656
rect 20824 7652 20854 7678
rect 20920 7656 20950 7678
rect 20710 7606 20726 7640
rect 20760 7606 20776 7640
rect 20710 7590 20776 7606
rect 20902 7640 20968 7656
rect 21016 7652 21046 7678
rect 21112 7656 21142 7678
rect 20902 7606 20918 7640
rect 20952 7606 20968 7640
rect 20902 7590 20968 7606
rect 21094 7640 21160 7656
rect 21208 7652 21238 7678
rect 21304 7656 21334 7678
rect 21094 7606 21110 7640
rect 21144 7606 21160 7640
rect 21094 7590 21160 7606
rect 21286 7640 21352 7656
rect 21400 7652 21430 7678
rect 21286 7606 21302 7640
rect 21336 7606 21352 7640
rect 21286 7590 21352 7606
rect 14754 5946 14820 5962
rect 14754 5912 14770 5946
rect 14804 5912 14820 5946
rect 14676 5874 14706 5900
rect 14754 5896 14820 5912
rect 14946 5946 15012 5962
rect 14946 5912 14962 5946
rect 14996 5912 15012 5946
rect 14772 5874 14802 5896
rect 14868 5874 14898 5900
rect 14946 5896 15012 5912
rect 15138 5946 15204 5962
rect 15138 5912 15154 5946
rect 15188 5912 15204 5946
rect 14964 5874 14994 5896
rect 15060 5874 15090 5900
rect 15138 5896 15204 5912
rect 15330 5946 15396 5962
rect 15330 5912 15346 5946
rect 15380 5912 15396 5946
rect 15156 5874 15186 5896
rect 15252 5874 15282 5900
rect 15330 5896 15396 5912
rect 15522 5946 15588 5962
rect 15522 5912 15538 5946
rect 15572 5912 15588 5946
rect 15348 5874 15378 5896
rect 15444 5874 15474 5900
rect 15522 5896 15588 5912
rect 15540 5874 15570 5896
rect 14676 5452 14706 5474
rect 14658 5436 14724 5452
rect 14772 5448 14802 5474
rect 14868 5452 14898 5474
rect 14658 5402 14674 5436
rect 14708 5402 14724 5436
rect 14658 5386 14724 5402
rect 14850 5436 14916 5452
rect 14964 5448 14994 5474
rect 15060 5452 15090 5474
rect 14850 5402 14866 5436
rect 14900 5402 14916 5436
rect 14850 5386 14916 5402
rect 15042 5436 15108 5452
rect 15156 5448 15186 5474
rect 15252 5452 15282 5474
rect 15042 5402 15058 5436
rect 15092 5402 15108 5436
rect 15042 5386 15108 5402
rect 15234 5436 15300 5452
rect 15348 5448 15378 5474
rect 15444 5452 15474 5474
rect 15234 5402 15250 5436
rect 15284 5402 15300 5436
rect 15234 5386 15300 5402
rect 15426 5436 15492 5452
rect 15540 5448 15570 5474
rect 15426 5402 15442 5436
rect 15476 5402 15492 5436
rect 15426 5386 15492 5402
rect 14658 5328 14724 5344
rect 14658 5294 14674 5328
rect 14708 5294 14724 5328
rect 14658 5278 14724 5294
rect 14850 5328 14916 5344
rect 14850 5294 14866 5328
rect 14900 5294 14916 5328
rect 14676 5256 14706 5278
rect 14772 5256 14802 5282
rect 14850 5278 14916 5294
rect 15042 5328 15108 5344
rect 15042 5294 15058 5328
rect 15092 5294 15108 5328
rect 14868 5256 14898 5278
rect 14964 5256 14994 5282
rect 15042 5278 15108 5294
rect 15234 5328 15300 5344
rect 15234 5294 15250 5328
rect 15284 5294 15300 5328
rect 15060 5256 15090 5278
rect 15156 5256 15186 5282
rect 15234 5278 15300 5294
rect 15426 5328 15492 5344
rect 15426 5294 15442 5328
rect 15476 5294 15492 5328
rect 15252 5256 15282 5278
rect 15348 5256 15378 5282
rect 15426 5278 15492 5294
rect 15444 5256 15474 5278
rect 15540 5256 15570 5282
rect 14676 4830 14706 4856
rect 14772 4834 14802 4856
rect 14754 4818 14820 4834
rect 14868 4830 14898 4856
rect 14964 4834 14994 4856
rect 14754 4784 14770 4818
rect 14804 4784 14820 4818
rect 14754 4768 14820 4784
rect 14946 4818 15012 4834
rect 15060 4830 15090 4856
rect 15156 4834 15186 4856
rect 14946 4784 14962 4818
rect 14996 4784 15012 4818
rect 14946 4768 15012 4784
rect 15138 4818 15204 4834
rect 15252 4830 15282 4856
rect 15348 4834 15378 4856
rect 15138 4784 15154 4818
rect 15188 4784 15204 4818
rect 15138 4768 15204 4784
rect 15330 4818 15396 4834
rect 15444 4830 15474 4856
rect 15540 4834 15570 4856
rect 15330 4784 15346 4818
rect 15380 4784 15396 4818
rect 15330 4768 15396 4784
rect 15522 4818 15588 4834
rect 15522 4784 15538 4818
rect 15572 4784 15588 4818
rect 15522 4768 15588 4784
rect 14754 4710 14820 4726
rect 14754 4676 14770 4710
rect 14804 4676 14820 4710
rect 14676 4638 14706 4664
rect 14754 4660 14820 4676
rect 14946 4710 15012 4726
rect 14946 4676 14962 4710
rect 14996 4676 15012 4710
rect 14772 4638 14802 4660
rect 14868 4638 14898 4664
rect 14946 4660 15012 4676
rect 15138 4710 15204 4726
rect 15138 4676 15154 4710
rect 15188 4676 15204 4710
rect 14964 4638 14994 4660
rect 15060 4638 15090 4664
rect 15138 4660 15204 4676
rect 15330 4710 15396 4726
rect 15330 4676 15346 4710
rect 15380 4676 15396 4710
rect 15156 4638 15186 4660
rect 15252 4638 15282 4664
rect 15330 4660 15396 4676
rect 15522 4710 15588 4726
rect 15522 4676 15538 4710
rect 15572 4676 15588 4710
rect 15348 4638 15378 4660
rect 15444 4638 15474 4664
rect 15522 4660 15588 4676
rect 15540 4638 15570 4660
rect 14676 4216 14706 4238
rect 14658 4200 14724 4216
rect 14772 4212 14802 4238
rect 14868 4216 14898 4238
rect 14658 4166 14674 4200
rect 14708 4166 14724 4200
rect 14658 4150 14724 4166
rect 14850 4200 14916 4216
rect 14964 4212 14994 4238
rect 15060 4216 15090 4238
rect 14850 4166 14866 4200
rect 14900 4166 14916 4200
rect 14850 4150 14916 4166
rect 15042 4200 15108 4216
rect 15156 4212 15186 4238
rect 15252 4216 15282 4238
rect 15042 4166 15058 4200
rect 15092 4166 15108 4200
rect 15042 4150 15108 4166
rect 15234 4200 15300 4216
rect 15348 4212 15378 4238
rect 15444 4216 15474 4238
rect 15234 4166 15250 4200
rect 15284 4166 15300 4200
rect 15234 4150 15300 4166
rect 15426 4200 15492 4216
rect 15540 4212 15570 4238
rect 15426 4166 15442 4200
rect 15476 4166 15492 4200
rect 15426 4150 15492 4166
rect 16554 5946 16620 5962
rect 16554 5912 16570 5946
rect 16604 5912 16620 5946
rect 16476 5874 16506 5900
rect 16554 5896 16620 5912
rect 16746 5946 16812 5962
rect 16746 5912 16762 5946
rect 16796 5912 16812 5946
rect 16572 5874 16602 5896
rect 16668 5874 16698 5900
rect 16746 5896 16812 5912
rect 16938 5946 17004 5962
rect 16938 5912 16954 5946
rect 16988 5912 17004 5946
rect 16764 5874 16794 5896
rect 16860 5874 16890 5900
rect 16938 5896 17004 5912
rect 17130 5946 17196 5962
rect 17130 5912 17146 5946
rect 17180 5912 17196 5946
rect 16956 5874 16986 5896
rect 17052 5874 17082 5900
rect 17130 5896 17196 5912
rect 17322 5946 17388 5962
rect 17322 5912 17338 5946
rect 17372 5912 17388 5946
rect 17148 5874 17178 5896
rect 17244 5874 17274 5900
rect 17322 5896 17388 5912
rect 17340 5874 17370 5896
rect 16476 5452 16506 5474
rect 16458 5436 16524 5452
rect 16572 5448 16602 5474
rect 16668 5452 16698 5474
rect 16458 5402 16474 5436
rect 16508 5402 16524 5436
rect 16458 5386 16524 5402
rect 16650 5436 16716 5452
rect 16764 5448 16794 5474
rect 16860 5452 16890 5474
rect 16650 5402 16666 5436
rect 16700 5402 16716 5436
rect 16650 5386 16716 5402
rect 16842 5436 16908 5452
rect 16956 5448 16986 5474
rect 17052 5452 17082 5474
rect 16842 5402 16858 5436
rect 16892 5402 16908 5436
rect 16842 5386 16908 5402
rect 17034 5436 17100 5452
rect 17148 5448 17178 5474
rect 17244 5452 17274 5474
rect 17034 5402 17050 5436
rect 17084 5402 17100 5436
rect 17034 5386 17100 5402
rect 17226 5436 17292 5452
rect 17340 5448 17370 5474
rect 17226 5402 17242 5436
rect 17276 5402 17292 5436
rect 17226 5386 17292 5402
rect 16458 5328 16524 5344
rect 16458 5294 16474 5328
rect 16508 5294 16524 5328
rect 16458 5278 16524 5294
rect 16650 5328 16716 5344
rect 16650 5294 16666 5328
rect 16700 5294 16716 5328
rect 16476 5256 16506 5278
rect 16572 5256 16602 5282
rect 16650 5278 16716 5294
rect 16842 5328 16908 5344
rect 16842 5294 16858 5328
rect 16892 5294 16908 5328
rect 16668 5256 16698 5278
rect 16764 5256 16794 5282
rect 16842 5278 16908 5294
rect 17034 5328 17100 5344
rect 17034 5294 17050 5328
rect 17084 5294 17100 5328
rect 16860 5256 16890 5278
rect 16956 5256 16986 5282
rect 17034 5278 17100 5294
rect 17226 5328 17292 5344
rect 17226 5294 17242 5328
rect 17276 5294 17292 5328
rect 17052 5256 17082 5278
rect 17148 5256 17178 5282
rect 17226 5278 17292 5294
rect 17244 5256 17274 5278
rect 17340 5256 17370 5282
rect 16476 4830 16506 4856
rect 16572 4834 16602 4856
rect 16554 4818 16620 4834
rect 16668 4830 16698 4856
rect 16764 4834 16794 4856
rect 16554 4784 16570 4818
rect 16604 4784 16620 4818
rect 16554 4768 16620 4784
rect 16746 4818 16812 4834
rect 16860 4830 16890 4856
rect 16956 4834 16986 4856
rect 16746 4784 16762 4818
rect 16796 4784 16812 4818
rect 16746 4768 16812 4784
rect 16938 4818 17004 4834
rect 17052 4830 17082 4856
rect 17148 4834 17178 4856
rect 16938 4784 16954 4818
rect 16988 4784 17004 4818
rect 16938 4768 17004 4784
rect 17130 4818 17196 4834
rect 17244 4830 17274 4856
rect 17340 4834 17370 4856
rect 17130 4784 17146 4818
rect 17180 4784 17196 4818
rect 17130 4768 17196 4784
rect 17322 4818 17388 4834
rect 17322 4784 17338 4818
rect 17372 4784 17388 4818
rect 17322 4768 17388 4784
rect 16554 4710 16620 4726
rect 16554 4676 16570 4710
rect 16604 4676 16620 4710
rect 16476 4638 16506 4664
rect 16554 4660 16620 4676
rect 16746 4710 16812 4726
rect 16746 4676 16762 4710
rect 16796 4676 16812 4710
rect 16572 4638 16602 4660
rect 16668 4638 16698 4664
rect 16746 4660 16812 4676
rect 16938 4710 17004 4726
rect 16938 4676 16954 4710
rect 16988 4676 17004 4710
rect 16764 4638 16794 4660
rect 16860 4638 16890 4664
rect 16938 4660 17004 4676
rect 17130 4710 17196 4726
rect 17130 4676 17146 4710
rect 17180 4676 17196 4710
rect 16956 4638 16986 4660
rect 17052 4638 17082 4664
rect 17130 4660 17196 4676
rect 17322 4710 17388 4726
rect 17322 4676 17338 4710
rect 17372 4676 17388 4710
rect 17148 4638 17178 4660
rect 17244 4638 17274 4664
rect 17322 4660 17388 4676
rect 17340 4638 17370 4660
rect 16476 4216 16506 4238
rect 16458 4200 16524 4216
rect 16572 4212 16602 4238
rect 16668 4216 16698 4238
rect 16458 4166 16474 4200
rect 16508 4166 16524 4200
rect 16458 4150 16524 4166
rect 16650 4200 16716 4216
rect 16764 4212 16794 4238
rect 16860 4216 16890 4238
rect 16650 4166 16666 4200
rect 16700 4166 16716 4200
rect 16650 4150 16716 4166
rect 16842 4200 16908 4216
rect 16956 4212 16986 4238
rect 17052 4216 17082 4238
rect 16842 4166 16858 4200
rect 16892 4166 16908 4200
rect 16842 4150 16908 4166
rect 17034 4200 17100 4216
rect 17148 4212 17178 4238
rect 17244 4216 17274 4238
rect 17034 4166 17050 4200
rect 17084 4166 17100 4200
rect 17034 4150 17100 4166
rect 17226 4200 17292 4216
rect 17340 4212 17370 4238
rect 17226 4166 17242 4200
rect 17276 4166 17292 4200
rect 17226 4150 17292 4166
rect 18354 5946 18420 5962
rect 18354 5912 18370 5946
rect 18404 5912 18420 5946
rect 18276 5874 18306 5900
rect 18354 5896 18420 5912
rect 18546 5946 18612 5962
rect 18546 5912 18562 5946
rect 18596 5912 18612 5946
rect 18372 5874 18402 5896
rect 18468 5874 18498 5900
rect 18546 5896 18612 5912
rect 18738 5946 18804 5962
rect 18738 5912 18754 5946
rect 18788 5912 18804 5946
rect 18564 5874 18594 5896
rect 18660 5874 18690 5900
rect 18738 5896 18804 5912
rect 18930 5946 18996 5962
rect 18930 5912 18946 5946
rect 18980 5912 18996 5946
rect 18756 5874 18786 5896
rect 18852 5874 18882 5900
rect 18930 5896 18996 5912
rect 19122 5946 19188 5962
rect 19122 5912 19138 5946
rect 19172 5912 19188 5946
rect 18948 5874 18978 5896
rect 19044 5874 19074 5900
rect 19122 5896 19188 5912
rect 19140 5874 19170 5896
rect 18276 5452 18306 5474
rect 18258 5436 18324 5452
rect 18372 5448 18402 5474
rect 18468 5452 18498 5474
rect 18258 5402 18274 5436
rect 18308 5402 18324 5436
rect 18258 5386 18324 5402
rect 18450 5436 18516 5452
rect 18564 5448 18594 5474
rect 18660 5452 18690 5474
rect 18450 5402 18466 5436
rect 18500 5402 18516 5436
rect 18450 5386 18516 5402
rect 18642 5436 18708 5452
rect 18756 5448 18786 5474
rect 18852 5452 18882 5474
rect 18642 5402 18658 5436
rect 18692 5402 18708 5436
rect 18642 5386 18708 5402
rect 18834 5436 18900 5452
rect 18948 5448 18978 5474
rect 19044 5452 19074 5474
rect 18834 5402 18850 5436
rect 18884 5402 18900 5436
rect 18834 5386 18900 5402
rect 19026 5436 19092 5452
rect 19140 5448 19170 5474
rect 19026 5402 19042 5436
rect 19076 5402 19092 5436
rect 19026 5386 19092 5402
rect 18258 5328 18324 5344
rect 18258 5294 18274 5328
rect 18308 5294 18324 5328
rect 18258 5278 18324 5294
rect 18450 5328 18516 5344
rect 18450 5294 18466 5328
rect 18500 5294 18516 5328
rect 18276 5256 18306 5278
rect 18372 5256 18402 5282
rect 18450 5278 18516 5294
rect 18642 5328 18708 5344
rect 18642 5294 18658 5328
rect 18692 5294 18708 5328
rect 18468 5256 18498 5278
rect 18564 5256 18594 5282
rect 18642 5278 18708 5294
rect 18834 5328 18900 5344
rect 18834 5294 18850 5328
rect 18884 5294 18900 5328
rect 18660 5256 18690 5278
rect 18756 5256 18786 5282
rect 18834 5278 18900 5294
rect 19026 5328 19092 5344
rect 19026 5294 19042 5328
rect 19076 5294 19092 5328
rect 18852 5256 18882 5278
rect 18948 5256 18978 5282
rect 19026 5278 19092 5294
rect 19044 5256 19074 5278
rect 19140 5256 19170 5282
rect 18276 4830 18306 4856
rect 18372 4834 18402 4856
rect 18354 4818 18420 4834
rect 18468 4830 18498 4856
rect 18564 4834 18594 4856
rect 18354 4784 18370 4818
rect 18404 4784 18420 4818
rect 18354 4768 18420 4784
rect 18546 4818 18612 4834
rect 18660 4830 18690 4856
rect 18756 4834 18786 4856
rect 18546 4784 18562 4818
rect 18596 4784 18612 4818
rect 18546 4768 18612 4784
rect 18738 4818 18804 4834
rect 18852 4830 18882 4856
rect 18948 4834 18978 4856
rect 18738 4784 18754 4818
rect 18788 4784 18804 4818
rect 18738 4768 18804 4784
rect 18930 4818 18996 4834
rect 19044 4830 19074 4856
rect 19140 4834 19170 4856
rect 18930 4784 18946 4818
rect 18980 4784 18996 4818
rect 18930 4768 18996 4784
rect 19122 4818 19188 4834
rect 19122 4784 19138 4818
rect 19172 4784 19188 4818
rect 19122 4768 19188 4784
rect 18354 4710 18420 4726
rect 18354 4676 18370 4710
rect 18404 4676 18420 4710
rect 18276 4638 18306 4664
rect 18354 4660 18420 4676
rect 18546 4710 18612 4726
rect 18546 4676 18562 4710
rect 18596 4676 18612 4710
rect 18372 4638 18402 4660
rect 18468 4638 18498 4664
rect 18546 4660 18612 4676
rect 18738 4710 18804 4726
rect 18738 4676 18754 4710
rect 18788 4676 18804 4710
rect 18564 4638 18594 4660
rect 18660 4638 18690 4664
rect 18738 4660 18804 4676
rect 18930 4710 18996 4726
rect 18930 4676 18946 4710
rect 18980 4676 18996 4710
rect 18756 4638 18786 4660
rect 18852 4638 18882 4664
rect 18930 4660 18996 4676
rect 19122 4710 19188 4726
rect 19122 4676 19138 4710
rect 19172 4676 19188 4710
rect 18948 4638 18978 4660
rect 19044 4638 19074 4664
rect 19122 4660 19188 4676
rect 19140 4638 19170 4660
rect 18276 4216 18306 4238
rect 18258 4200 18324 4216
rect 18372 4212 18402 4238
rect 18468 4216 18498 4238
rect 18258 4166 18274 4200
rect 18308 4166 18324 4200
rect 18258 4150 18324 4166
rect 18450 4200 18516 4216
rect 18564 4212 18594 4238
rect 18660 4216 18690 4238
rect 18450 4166 18466 4200
rect 18500 4166 18516 4200
rect 18450 4150 18516 4166
rect 18642 4200 18708 4216
rect 18756 4212 18786 4238
rect 18852 4216 18882 4238
rect 18642 4166 18658 4200
rect 18692 4166 18708 4200
rect 18642 4150 18708 4166
rect 18834 4200 18900 4216
rect 18948 4212 18978 4238
rect 19044 4216 19074 4238
rect 18834 4166 18850 4200
rect 18884 4166 18900 4200
rect 18834 4150 18900 4166
rect 19026 4200 19092 4216
rect 19140 4212 19170 4238
rect 19026 4166 19042 4200
rect 19076 4166 19092 4200
rect 19026 4150 19092 4166
rect 20154 5946 20220 5962
rect 20154 5912 20170 5946
rect 20204 5912 20220 5946
rect 20076 5874 20106 5900
rect 20154 5896 20220 5912
rect 20346 5946 20412 5962
rect 20346 5912 20362 5946
rect 20396 5912 20412 5946
rect 20172 5874 20202 5896
rect 20268 5874 20298 5900
rect 20346 5896 20412 5912
rect 20538 5946 20604 5962
rect 20538 5912 20554 5946
rect 20588 5912 20604 5946
rect 20364 5874 20394 5896
rect 20460 5874 20490 5900
rect 20538 5896 20604 5912
rect 20730 5946 20796 5962
rect 20730 5912 20746 5946
rect 20780 5912 20796 5946
rect 20556 5874 20586 5896
rect 20652 5874 20682 5900
rect 20730 5896 20796 5912
rect 20922 5946 20988 5962
rect 20922 5912 20938 5946
rect 20972 5912 20988 5946
rect 20748 5874 20778 5896
rect 20844 5874 20874 5900
rect 20922 5896 20988 5912
rect 20940 5874 20970 5896
rect 20076 5452 20106 5474
rect 20058 5436 20124 5452
rect 20172 5448 20202 5474
rect 20268 5452 20298 5474
rect 20058 5402 20074 5436
rect 20108 5402 20124 5436
rect 20058 5386 20124 5402
rect 20250 5436 20316 5452
rect 20364 5448 20394 5474
rect 20460 5452 20490 5474
rect 20250 5402 20266 5436
rect 20300 5402 20316 5436
rect 20250 5386 20316 5402
rect 20442 5436 20508 5452
rect 20556 5448 20586 5474
rect 20652 5452 20682 5474
rect 20442 5402 20458 5436
rect 20492 5402 20508 5436
rect 20442 5386 20508 5402
rect 20634 5436 20700 5452
rect 20748 5448 20778 5474
rect 20844 5452 20874 5474
rect 20634 5402 20650 5436
rect 20684 5402 20700 5436
rect 20634 5386 20700 5402
rect 20826 5436 20892 5452
rect 20940 5448 20970 5474
rect 20826 5402 20842 5436
rect 20876 5402 20892 5436
rect 20826 5386 20892 5402
rect 20058 5328 20124 5344
rect 20058 5294 20074 5328
rect 20108 5294 20124 5328
rect 20058 5278 20124 5294
rect 20250 5328 20316 5344
rect 20250 5294 20266 5328
rect 20300 5294 20316 5328
rect 20076 5256 20106 5278
rect 20172 5256 20202 5282
rect 20250 5278 20316 5294
rect 20442 5328 20508 5344
rect 20442 5294 20458 5328
rect 20492 5294 20508 5328
rect 20268 5256 20298 5278
rect 20364 5256 20394 5282
rect 20442 5278 20508 5294
rect 20634 5328 20700 5344
rect 20634 5294 20650 5328
rect 20684 5294 20700 5328
rect 20460 5256 20490 5278
rect 20556 5256 20586 5282
rect 20634 5278 20700 5294
rect 20826 5328 20892 5344
rect 20826 5294 20842 5328
rect 20876 5294 20892 5328
rect 20652 5256 20682 5278
rect 20748 5256 20778 5282
rect 20826 5278 20892 5294
rect 20844 5256 20874 5278
rect 20940 5256 20970 5282
rect 20076 4830 20106 4856
rect 20172 4834 20202 4856
rect 20154 4818 20220 4834
rect 20268 4830 20298 4856
rect 20364 4834 20394 4856
rect 20154 4784 20170 4818
rect 20204 4784 20220 4818
rect 20154 4768 20220 4784
rect 20346 4818 20412 4834
rect 20460 4830 20490 4856
rect 20556 4834 20586 4856
rect 20346 4784 20362 4818
rect 20396 4784 20412 4818
rect 20346 4768 20412 4784
rect 20538 4818 20604 4834
rect 20652 4830 20682 4856
rect 20748 4834 20778 4856
rect 20538 4784 20554 4818
rect 20588 4784 20604 4818
rect 20538 4768 20604 4784
rect 20730 4818 20796 4834
rect 20844 4830 20874 4856
rect 20940 4834 20970 4856
rect 20730 4784 20746 4818
rect 20780 4784 20796 4818
rect 20730 4768 20796 4784
rect 20922 4818 20988 4834
rect 20922 4784 20938 4818
rect 20972 4784 20988 4818
rect 20922 4768 20988 4784
rect 20154 4710 20220 4726
rect 20154 4676 20170 4710
rect 20204 4676 20220 4710
rect 20076 4638 20106 4664
rect 20154 4660 20220 4676
rect 20346 4710 20412 4726
rect 20346 4676 20362 4710
rect 20396 4676 20412 4710
rect 20172 4638 20202 4660
rect 20268 4638 20298 4664
rect 20346 4660 20412 4676
rect 20538 4710 20604 4726
rect 20538 4676 20554 4710
rect 20588 4676 20604 4710
rect 20364 4638 20394 4660
rect 20460 4638 20490 4664
rect 20538 4660 20604 4676
rect 20730 4710 20796 4726
rect 20730 4676 20746 4710
rect 20780 4676 20796 4710
rect 20556 4638 20586 4660
rect 20652 4638 20682 4664
rect 20730 4660 20796 4676
rect 20922 4710 20988 4726
rect 20922 4676 20938 4710
rect 20972 4676 20988 4710
rect 20748 4638 20778 4660
rect 20844 4638 20874 4664
rect 20922 4660 20988 4676
rect 20940 4638 20970 4660
rect 20076 4216 20106 4238
rect 20058 4200 20124 4216
rect 20172 4212 20202 4238
rect 20268 4216 20298 4238
rect 20058 4166 20074 4200
rect 20108 4166 20124 4200
rect 20058 4150 20124 4166
rect 20250 4200 20316 4216
rect 20364 4212 20394 4238
rect 20460 4216 20490 4238
rect 20250 4166 20266 4200
rect 20300 4166 20316 4200
rect 20250 4150 20316 4166
rect 20442 4200 20508 4216
rect 20556 4212 20586 4238
rect 20652 4216 20682 4238
rect 20442 4166 20458 4200
rect 20492 4166 20508 4200
rect 20442 4150 20508 4166
rect 20634 4200 20700 4216
rect 20748 4212 20778 4238
rect 20844 4216 20874 4238
rect 20634 4166 20650 4200
rect 20684 4166 20700 4200
rect 20634 4150 20700 4166
rect 20826 4200 20892 4216
rect 20940 4212 20970 4238
rect 20826 4166 20842 4200
rect 20876 4166 20892 4200
rect 20826 4150 20892 4166
rect 22154 10334 22220 10350
rect 22154 10300 22170 10334
rect 22204 10300 22220 10334
rect 22076 10262 22106 10288
rect 22154 10284 22220 10300
rect 22346 10334 22412 10350
rect 22346 10300 22362 10334
rect 22396 10300 22412 10334
rect 22172 10262 22202 10284
rect 22268 10262 22298 10288
rect 22346 10284 22412 10300
rect 22538 10334 22604 10350
rect 22538 10300 22554 10334
rect 22588 10300 22604 10334
rect 22364 10262 22394 10284
rect 22460 10262 22490 10288
rect 22538 10284 22604 10300
rect 22730 10334 22796 10350
rect 22730 10300 22746 10334
rect 22780 10300 22796 10334
rect 22556 10262 22586 10284
rect 22652 10262 22682 10288
rect 22730 10284 22796 10300
rect 22922 10334 22988 10350
rect 22922 10300 22938 10334
rect 22972 10300 22988 10334
rect 22748 10262 22778 10284
rect 22844 10262 22874 10288
rect 22922 10284 22988 10300
rect 23114 10334 23180 10350
rect 23114 10300 23130 10334
rect 23164 10300 23180 10334
rect 22940 10262 22970 10284
rect 23036 10262 23066 10288
rect 23114 10284 23180 10300
rect 23306 10334 23372 10350
rect 23306 10300 23322 10334
rect 23356 10300 23372 10334
rect 23132 10262 23162 10284
rect 23228 10262 23258 10288
rect 23306 10284 23372 10300
rect 23498 10334 23564 10350
rect 23498 10300 23514 10334
rect 23548 10300 23564 10334
rect 23324 10262 23354 10284
rect 23420 10262 23450 10288
rect 23498 10284 23564 10300
rect 23690 10334 23756 10350
rect 23690 10300 23706 10334
rect 23740 10300 23756 10334
rect 23516 10262 23546 10284
rect 23612 10262 23642 10288
rect 23690 10284 23756 10300
rect 23882 10334 23948 10350
rect 23882 10300 23898 10334
rect 23932 10300 23948 10334
rect 23708 10262 23738 10284
rect 23804 10262 23834 10288
rect 23882 10284 23948 10300
rect 23900 10262 23930 10284
rect 22076 9840 22106 9862
rect 22058 9824 22124 9840
rect 22172 9836 22202 9862
rect 22268 9840 22298 9862
rect 22058 9790 22074 9824
rect 22108 9790 22124 9824
rect 22058 9774 22124 9790
rect 22250 9824 22316 9840
rect 22364 9836 22394 9862
rect 22460 9840 22490 9862
rect 22250 9790 22266 9824
rect 22300 9790 22316 9824
rect 22250 9774 22316 9790
rect 22442 9824 22508 9840
rect 22556 9836 22586 9862
rect 22652 9840 22682 9862
rect 22442 9790 22458 9824
rect 22492 9790 22508 9824
rect 22442 9774 22508 9790
rect 22634 9824 22700 9840
rect 22748 9836 22778 9862
rect 22844 9840 22874 9862
rect 22634 9790 22650 9824
rect 22684 9790 22700 9824
rect 22634 9774 22700 9790
rect 22826 9824 22892 9840
rect 22940 9836 22970 9862
rect 23036 9840 23066 9862
rect 22826 9790 22842 9824
rect 22876 9790 22892 9824
rect 22826 9774 22892 9790
rect 23018 9824 23084 9840
rect 23132 9836 23162 9862
rect 23228 9840 23258 9862
rect 23018 9790 23034 9824
rect 23068 9790 23084 9824
rect 23018 9774 23084 9790
rect 23210 9824 23276 9840
rect 23324 9836 23354 9862
rect 23420 9840 23450 9862
rect 23210 9790 23226 9824
rect 23260 9790 23276 9824
rect 23210 9774 23276 9790
rect 23402 9824 23468 9840
rect 23516 9836 23546 9862
rect 23612 9840 23642 9862
rect 23402 9790 23418 9824
rect 23452 9790 23468 9824
rect 23402 9774 23468 9790
rect 23594 9824 23660 9840
rect 23708 9836 23738 9862
rect 23804 9840 23834 9862
rect 23594 9790 23610 9824
rect 23644 9790 23660 9824
rect 23594 9774 23660 9790
rect 23786 9824 23852 9840
rect 23900 9836 23930 9862
rect 23786 9790 23802 9824
rect 23836 9790 23852 9824
rect 23786 9774 23852 9790
rect 22058 9716 22124 9732
rect 22058 9682 22074 9716
rect 22108 9682 22124 9716
rect 22058 9666 22124 9682
rect 22250 9716 22316 9732
rect 22250 9682 22266 9716
rect 22300 9682 22316 9716
rect 22076 9644 22106 9666
rect 22172 9644 22202 9670
rect 22250 9666 22316 9682
rect 22442 9716 22508 9732
rect 22442 9682 22458 9716
rect 22492 9682 22508 9716
rect 22268 9644 22298 9666
rect 22364 9644 22394 9670
rect 22442 9666 22508 9682
rect 22634 9716 22700 9732
rect 22634 9682 22650 9716
rect 22684 9682 22700 9716
rect 22460 9644 22490 9666
rect 22556 9644 22586 9670
rect 22634 9666 22700 9682
rect 22826 9716 22892 9732
rect 22826 9682 22842 9716
rect 22876 9682 22892 9716
rect 22652 9644 22682 9666
rect 22748 9644 22778 9670
rect 22826 9666 22892 9682
rect 23018 9716 23084 9732
rect 23018 9682 23034 9716
rect 23068 9682 23084 9716
rect 22844 9644 22874 9666
rect 22940 9644 22970 9670
rect 23018 9666 23084 9682
rect 23210 9716 23276 9732
rect 23210 9682 23226 9716
rect 23260 9682 23276 9716
rect 23036 9644 23066 9666
rect 23132 9644 23162 9670
rect 23210 9666 23276 9682
rect 23402 9716 23468 9732
rect 23402 9682 23418 9716
rect 23452 9682 23468 9716
rect 23228 9644 23258 9666
rect 23324 9644 23354 9670
rect 23402 9666 23468 9682
rect 23594 9716 23660 9732
rect 23594 9682 23610 9716
rect 23644 9682 23660 9716
rect 23420 9644 23450 9666
rect 23516 9644 23546 9670
rect 23594 9666 23660 9682
rect 23786 9716 23852 9732
rect 23786 9682 23802 9716
rect 23836 9682 23852 9716
rect 23612 9644 23642 9666
rect 23708 9644 23738 9670
rect 23786 9666 23852 9682
rect 23804 9644 23834 9666
rect 23900 9644 23930 9670
rect 22076 9218 22106 9244
rect 22172 9222 22202 9244
rect 22154 9206 22220 9222
rect 22268 9218 22298 9244
rect 22364 9222 22394 9244
rect 22154 9172 22170 9206
rect 22204 9172 22220 9206
rect 22154 9156 22220 9172
rect 22346 9206 22412 9222
rect 22460 9218 22490 9244
rect 22556 9222 22586 9244
rect 22346 9172 22362 9206
rect 22396 9172 22412 9206
rect 22346 9156 22412 9172
rect 22538 9206 22604 9222
rect 22652 9218 22682 9244
rect 22748 9222 22778 9244
rect 22538 9172 22554 9206
rect 22588 9172 22604 9206
rect 22538 9156 22604 9172
rect 22730 9206 22796 9222
rect 22844 9218 22874 9244
rect 22940 9222 22970 9244
rect 22730 9172 22746 9206
rect 22780 9172 22796 9206
rect 22730 9156 22796 9172
rect 22922 9206 22988 9222
rect 23036 9218 23066 9244
rect 23132 9222 23162 9244
rect 22922 9172 22938 9206
rect 22972 9172 22988 9206
rect 22922 9156 22988 9172
rect 23114 9206 23180 9222
rect 23228 9218 23258 9244
rect 23324 9222 23354 9244
rect 23114 9172 23130 9206
rect 23164 9172 23180 9206
rect 23114 9156 23180 9172
rect 23306 9206 23372 9222
rect 23420 9218 23450 9244
rect 23516 9222 23546 9244
rect 23306 9172 23322 9206
rect 23356 9172 23372 9206
rect 23306 9156 23372 9172
rect 23498 9206 23564 9222
rect 23612 9218 23642 9244
rect 23708 9222 23738 9244
rect 23498 9172 23514 9206
rect 23548 9172 23564 9206
rect 23498 9156 23564 9172
rect 23690 9206 23756 9222
rect 23804 9218 23834 9244
rect 23900 9222 23930 9244
rect 23690 9172 23706 9206
rect 23740 9172 23756 9206
rect 23690 9156 23756 9172
rect 23882 9206 23948 9222
rect 23882 9172 23898 9206
rect 23932 9172 23948 9206
rect 23882 9156 23948 9172
rect 22154 9098 22220 9114
rect 22154 9064 22170 9098
rect 22204 9064 22220 9098
rect 22076 9026 22106 9052
rect 22154 9048 22220 9064
rect 22346 9098 22412 9114
rect 22346 9064 22362 9098
rect 22396 9064 22412 9098
rect 22172 9026 22202 9048
rect 22268 9026 22298 9052
rect 22346 9048 22412 9064
rect 22538 9098 22604 9114
rect 22538 9064 22554 9098
rect 22588 9064 22604 9098
rect 22364 9026 22394 9048
rect 22460 9026 22490 9052
rect 22538 9048 22604 9064
rect 22730 9098 22796 9114
rect 22730 9064 22746 9098
rect 22780 9064 22796 9098
rect 22556 9026 22586 9048
rect 22652 9026 22682 9052
rect 22730 9048 22796 9064
rect 22922 9098 22988 9114
rect 22922 9064 22938 9098
rect 22972 9064 22988 9098
rect 22748 9026 22778 9048
rect 22844 9026 22874 9052
rect 22922 9048 22988 9064
rect 23114 9098 23180 9114
rect 23114 9064 23130 9098
rect 23164 9064 23180 9098
rect 22940 9026 22970 9048
rect 23036 9026 23066 9052
rect 23114 9048 23180 9064
rect 23306 9098 23372 9114
rect 23306 9064 23322 9098
rect 23356 9064 23372 9098
rect 23132 9026 23162 9048
rect 23228 9026 23258 9052
rect 23306 9048 23372 9064
rect 23498 9098 23564 9114
rect 23498 9064 23514 9098
rect 23548 9064 23564 9098
rect 23324 9026 23354 9048
rect 23420 9026 23450 9052
rect 23498 9048 23564 9064
rect 23690 9098 23756 9114
rect 23690 9064 23706 9098
rect 23740 9064 23756 9098
rect 23516 9026 23546 9048
rect 23612 9026 23642 9052
rect 23690 9048 23756 9064
rect 23882 9098 23948 9114
rect 23882 9064 23898 9098
rect 23932 9064 23948 9098
rect 23708 9026 23738 9048
rect 23804 9026 23834 9052
rect 23882 9048 23948 9064
rect 23900 9026 23930 9048
rect 22076 8604 22106 8626
rect 22058 8588 22124 8604
rect 22172 8600 22202 8626
rect 22268 8604 22298 8626
rect 22058 8554 22074 8588
rect 22108 8554 22124 8588
rect 22058 8538 22124 8554
rect 22250 8588 22316 8604
rect 22364 8600 22394 8626
rect 22460 8604 22490 8626
rect 22250 8554 22266 8588
rect 22300 8554 22316 8588
rect 22250 8538 22316 8554
rect 22442 8588 22508 8604
rect 22556 8600 22586 8626
rect 22652 8604 22682 8626
rect 22442 8554 22458 8588
rect 22492 8554 22508 8588
rect 22442 8538 22508 8554
rect 22634 8588 22700 8604
rect 22748 8600 22778 8626
rect 22844 8604 22874 8626
rect 22634 8554 22650 8588
rect 22684 8554 22700 8588
rect 22634 8538 22700 8554
rect 22826 8588 22892 8604
rect 22940 8600 22970 8626
rect 23036 8604 23066 8626
rect 22826 8554 22842 8588
rect 22876 8554 22892 8588
rect 22826 8538 22892 8554
rect 23018 8588 23084 8604
rect 23132 8600 23162 8626
rect 23228 8604 23258 8626
rect 23018 8554 23034 8588
rect 23068 8554 23084 8588
rect 23018 8538 23084 8554
rect 23210 8588 23276 8604
rect 23324 8600 23354 8626
rect 23420 8604 23450 8626
rect 23210 8554 23226 8588
rect 23260 8554 23276 8588
rect 23210 8538 23276 8554
rect 23402 8588 23468 8604
rect 23516 8600 23546 8626
rect 23612 8604 23642 8626
rect 23402 8554 23418 8588
rect 23452 8554 23468 8588
rect 23402 8538 23468 8554
rect 23594 8588 23660 8604
rect 23708 8600 23738 8626
rect 23804 8604 23834 8626
rect 23594 8554 23610 8588
rect 23644 8554 23660 8588
rect 23594 8538 23660 8554
rect 23786 8588 23852 8604
rect 23900 8600 23930 8626
rect 23786 8554 23802 8588
rect 23836 8554 23852 8588
rect 23786 8538 23852 8554
rect 22058 8480 22124 8496
rect 22058 8446 22074 8480
rect 22108 8446 22124 8480
rect 22058 8430 22124 8446
rect 22250 8480 22316 8496
rect 22250 8446 22266 8480
rect 22300 8446 22316 8480
rect 22076 8408 22106 8430
rect 22172 8408 22202 8434
rect 22250 8430 22316 8446
rect 22442 8480 22508 8496
rect 22442 8446 22458 8480
rect 22492 8446 22508 8480
rect 22268 8408 22298 8430
rect 22364 8408 22394 8434
rect 22442 8430 22508 8446
rect 22634 8480 22700 8496
rect 22634 8446 22650 8480
rect 22684 8446 22700 8480
rect 22460 8408 22490 8430
rect 22556 8408 22586 8434
rect 22634 8430 22700 8446
rect 22826 8480 22892 8496
rect 22826 8446 22842 8480
rect 22876 8446 22892 8480
rect 22652 8408 22682 8430
rect 22748 8408 22778 8434
rect 22826 8430 22892 8446
rect 23018 8480 23084 8496
rect 23018 8446 23034 8480
rect 23068 8446 23084 8480
rect 22844 8408 22874 8430
rect 22940 8408 22970 8434
rect 23018 8430 23084 8446
rect 23210 8480 23276 8496
rect 23210 8446 23226 8480
rect 23260 8446 23276 8480
rect 23036 8408 23066 8430
rect 23132 8408 23162 8434
rect 23210 8430 23276 8446
rect 23402 8480 23468 8496
rect 23402 8446 23418 8480
rect 23452 8446 23468 8480
rect 23228 8408 23258 8430
rect 23324 8408 23354 8434
rect 23402 8430 23468 8446
rect 23594 8480 23660 8496
rect 23594 8446 23610 8480
rect 23644 8446 23660 8480
rect 23420 8408 23450 8430
rect 23516 8408 23546 8434
rect 23594 8430 23660 8446
rect 23786 8480 23852 8496
rect 23786 8446 23802 8480
rect 23836 8446 23852 8480
rect 23612 8408 23642 8430
rect 23708 8408 23738 8434
rect 23786 8430 23852 8446
rect 23804 8408 23834 8430
rect 23900 8408 23930 8434
rect 22076 7982 22106 8008
rect 22172 7986 22202 8008
rect 22154 7970 22220 7986
rect 22268 7982 22298 8008
rect 22364 7986 22394 8008
rect 22154 7936 22170 7970
rect 22204 7936 22220 7970
rect 22154 7920 22220 7936
rect 22346 7970 22412 7986
rect 22460 7982 22490 8008
rect 22556 7986 22586 8008
rect 22346 7936 22362 7970
rect 22396 7936 22412 7970
rect 22346 7920 22412 7936
rect 22538 7970 22604 7986
rect 22652 7982 22682 8008
rect 22748 7986 22778 8008
rect 22538 7936 22554 7970
rect 22588 7936 22604 7970
rect 22538 7920 22604 7936
rect 22730 7970 22796 7986
rect 22844 7982 22874 8008
rect 22940 7986 22970 8008
rect 22730 7936 22746 7970
rect 22780 7936 22796 7970
rect 22730 7920 22796 7936
rect 22922 7970 22988 7986
rect 23036 7982 23066 8008
rect 23132 7986 23162 8008
rect 22922 7936 22938 7970
rect 22972 7936 22988 7970
rect 22922 7920 22988 7936
rect 23114 7970 23180 7986
rect 23228 7982 23258 8008
rect 23324 7986 23354 8008
rect 23114 7936 23130 7970
rect 23164 7936 23180 7970
rect 23114 7920 23180 7936
rect 23306 7970 23372 7986
rect 23420 7982 23450 8008
rect 23516 7986 23546 8008
rect 23306 7936 23322 7970
rect 23356 7936 23372 7970
rect 23306 7920 23372 7936
rect 23498 7970 23564 7986
rect 23612 7982 23642 8008
rect 23708 7986 23738 8008
rect 23498 7936 23514 7970
rect 23548 7936 23564 7970
rect 23498 7920 23564 7936
rect 23690 7970 23756 7986
rect 23804 7982 23834 8008
rect 23900 7986 23930 8008
rect 23690 7936 23706 7970
rect 23740 7936 23756 7970
rect 23690 7920 23756 7936
rect 23882 7970 23948 7986
rect 23882 7936 23898 7970
rect 23932 7936 23948 7970
rect 23882 7920 23948 7936
rect 22154 7862 22220 7878
rect 22154 7828 22170 7862
rect 22204 7828 22220 7862
rect 22076 7790 22106 7816
rect 22154 7812 22220 7828
rect 22346 7862 22412 7878
rect 22346 7828 22362 7862
rect 22396 7828 22412 7862
rect 22172 7790 22202 7812
rect 22268 7790 22298 7816
rect 22346 7812 22412 7828
rect 22538 7862 22604 7878
rect 22538 7828 22554 7862
rect 22588 7828 22604 7862
rect 22364 7790 22394 7812
rect 22460 7790 22490 7816
rect 22538 7812 22604 7828
rect 22730 7862 22796 7878
rect 22730 7828 22746 7862
rect 22780 7828 22796 7862
rect 22556 7790 22586 7812
rect 22652 7790 22682 7816
rect 22730 7812 22796 7828
rect 22922 7862 22988 7878
rect 22922 7828 22938 7862
rect 22972 7828 22988 7862
rect 22748 7790 22778 7812
rect 22844 7790 22874 7816
rect 22922 7812 22988 7828
rect 23114 7862 23180 7878
rect 23114 7828 23130 7862
rect 23164 7828 23180 7862
rect 22940 7790 22970 7812
rect 23036 7790 23066 7816
rect 23114 7812 23180 7828
rect 23306 7862 23372 7878
rect 23306 7828 23322 7862
rect 23356 7828 23372 7862
rect 23132 7790 23162 7812
rect 23228 7790 23258 7816
rect 23306 7812 23372 7828
rect 23498 7862 23564 7878
rect 23498 7828 23514 7862
rect 23548 7828 23564 7862
rect 23324 7790 23354 7812
rect 23420 7790 23450 7816
rect 23498 7812 23564 7828
rect 23690 7862 23756 7878
rect 23690 7828 23706 7862
rect 23740 7828 23756 7862
rect 23516 7790 23546 7812
rect 23612 7790 23642 7816
rect 23690 7812 23756 7828
rect 23882 7862 23948 7878
rect 23882 7828 23898 7862
rect 23932 7828 23948 7862
rect 23708 7790 23738 7812
rect 23804 7790 23834 7816
rect 23882 7812 23948 7828
rect 23900 7790 23930 7812
rect 22076 7368 22106 7390
rect 22058 7352 22124 7368
rect 22172 7364 22202 7390
rect 22268 7368 22298 7390
rect 22058 7318 22074 7352
rect 22108 7318 22124 7352
rect 22058 7302 22124 7318
rect 22250 7352 22316 7368
rect 22364 7364 22394 7390
rect 22460 7368 22490 7390
rect 22250 7318 22266 7352
rect 22300 7318 22316 7352
rect 22250 7302 22316 7318
rect 22442 7352 22508 7368
rect 22556 7364 22586 7390
rect 22652 7368 22682 7390
rect 22442 7318 22458 7352
rect 22492 7318 22508 7352
rect 22442 7302 22508 7318
rect 22634 7352 22700 7368
rect 22748 7364 22778 7390
rect 22844 7368 22874 7390
rect 22634 7318 22650 7352
rect 22684 7318 22700 7352
rect 22634 7302 22700 7318
rect 22826 7352 22892 7368
rect 22940 7364 22970 7390
rect 23036 7368 23066 7390
rect 22826 7318 22842 7352
rect 22876 7318 22892 7352
rect 22826 7302 22892 7318
rect 23018 7352 23084 7368
rect 23132 7364 23162 7390
rect 23228 7368 23258 7390
rect 23018 7318 23034 7352
rect 23068 7318 23084 7352
rect 23018 7302 23084 7318
rect 23210 7352 23276 7368
rect 23324 7364 23354 7390
rect 23420 7368 23450 7390
rect 23210 7318 23226 7352
rect 23260 7318 23276 7352
rect 23210 7302 23276 7318
rect 23402 7352 23468 7368
rect 23516 7364 23546 7390
rect 23612 7368 23642 7390
rect 23402 7318 23418 7352
rect 23452 7318 23468 7352
rect 23402 7302 23468 7318
rect 23594 7352 23660 7368
rect 23708 7364 23738 7390
rect 23804 7368 23834 7390
rect 23594 7318 23610 7352
rect 23644 7318 23660 7352
rect 23594 7302 23660 7318
rect 23786 7352 23852 7368
rect 23900 7364 23930 7390
rect 23786 7318 23802 7352
rect 23836 7318 23852 7352
rect 23786 7302 23852 7318
rect 22058 7244 22124 7260
rect 22058 7210 22074 7244
rect 22108 7210 22124 7244
rect 22058 7194 22124 7210
rect 22250 7244 22316 7260
rect 22250 7210 22266 7244
rect 22300 7210 22316 7244
rect 22076 7172 22106 7194
rect 22172 7172 22202 7198
rect 22250 7194 22316 7210
rect 22442 7244 22508 7260
rect 22442 7210 22458 7244
rect 22492 7210 22508 7244
rect 22268 7172 22298 7194
rect 22364 7172 22394 7198
rect 22442 7194 22508 7210
rect 22634 7244 22700 7260
rect 22634 7210 22650 7244
rect 22684 7210 22700 7244
rect 22460 7172 22490 7194
rect 22556 7172 22586 7198
rect 22634 7194 22700 7210
rect 22826 7244 22892 7260
rect 22826 7210 22842 7244
rect 22876 7210 22892 7244
rect 22652 7172 22682 7194
rect 22748 7172 22778 7198
rect 22826 7194 22892 7210
rect 23018 7244 23084 7260
rect 23018 7210 23034 7244
rect 23068 7210 23084 7244
rect 22844 7172 22874 7194
rect 22940 7172 22970 7198
rect 23018 7194 23084 7210
rect 23210 7244 23276 7260
rect 23210 7210 23226 7244
rect 23260 7210 23276 7244
rect 23036 7172 23066 7194
rect 23132 7172 23162 7198
rect 23210 7194 23276 7210
rect 23402 7244 23468 7260
rect 23402 7210 23418 7244
rect 23452 7210 23468 7244
rect 23228 7172 23258 7194
rect 23324 7172 23354 7198
rect 23402 7194 23468 7210
rect 23594 7244 23660 7260
rect 23594 7210 23610 7244
rect 23644 7210 23660 7244
rect 23420 7172 23450 7194
rect 23516 7172 23546 7198
rect 23594 7194 23660 7210
rect 23786 7244 23852 7260
rect 23786 7210 23802 7244
rect 23836 7210 23852 7244
rect 23612 7172 23642 7194
rect 23708 7172 23738 7198
rect 23786 7194 23852 7210
rect 23804 7172 23834 7194
rect 23900 7172 23930 7198
rect 22076 6746 22106 6772
rect 22172 6750 22202 6772
rect 22154 6734 22220 6750
rect 22268 6746 22298 6772
rect 22364 6750 22394 6772
rect 22154 6700 22170 6734
rect 22204 6700 22220 6734
rect 22154 6684 22220 6700
rect 22346 6734 22412 6750
rect 22460 6746 22490 6772
rect 22556 6750 22586 6772
rect 22346 6700 22362 6734
rect 22396 6700 22412 6734
rect 22346 6684 22412 6700
rect 22538 6734 22604 6750
rect 22652 6746 22682 6772
rect 22748 6750 22778 6772
rect 22538 6700 22554 6734
rect 22588 6700 22604 6734
rect 22538 6684 22604 6700
rect 22730 6734 22796 6750
rect 22844 6746 22874 6772
rect 22940 6750 22970 6772
rect 22730 6700 22746 6734
rect 22780 6700 22796 6734
rect 22730 6684 22796 6700
rect 22922 6734 22988 6750
rect 23036 6746 23066 6772
rect 23132 6750 23162 6772
rect 22922 6700 22938 6734
rect 22972 6700 22988 6734
rect 22922 6684 22988 6700
rect 23114 6734 23180 6750
rect 23228 6746 23258 6772
rect 23324 6750 23354 6772
rect 23114 6700 23130 6734
rect 23164 6700 23180 6734
rect 23114 6684 23180 6700
rect 23306 6734 23372 6750
rect 23420 6746 23450 6772
rect 23516 6750 23546 6772
rect 23306 6700 23322 6734
rect 23356 6700 23372 6734
rect 23306 6684 23372 6700
rect 23498 6734 23564 6750
rect 23612 6746 23642 6772
rect 23708 6750 23738 6772
rect 23498 6700 23514 6734
rect 23548 6700 23564 6734
rect 23498 6684 23564 6700
rect 23690 6734 23756 6750
rect 23804 6746 23834 6772
rect 23900 6750 23930 6772
rect 23690 6700 23706 6734
rect 23740 6700 23756 6734
rect 23690 6684 23756 6700
rect 23882 6734 23948 6750
rect 23882 6700 23898 6734
rect 23932 6700 23948 6734
rect 23882 6684 23948 6700
rect 22154 6626 22220 6642
rect 22154 6592 22170 6626
rect 22204 6592 22220 6626
rect 22076 6554 22106 6580
rect 22154 6576 22220 6592
rect 22346 6626 22412 6642
rect 22346 6592 22362 6626
rect 22396 6592 22412 6626
rect 22172 6554 22202 6576
rect 22268 6554 22298 6580
rect 22346 6576 22412 6592
rect 22538 6626 22604 6642
rect 22538 6592 22554 6626
rect 22588 6592 22604 6626
rect 22364 6554 22394 6576
rect 22460 6554 22490 6580
rect 22538 6576 22604 6592
rect 22730 6626 22796 6642
rect 22730 6592 22746 6626
rect 22780 6592 22796 6626
rect 22556 6554 22586 6576
rect 22652 6554 22682 6580
rect 22730 6576 22796 6592
rect 22922 6626 22988 6642
rect 22922 6592 22938 6626
rect 22972 6592 22988 6626
rect 22748 6554 22778 6576
rect 22844 6554 22874 6580
rect 22922 6576 22988 6592
rect 23114 6626 23180 6642
rect 23114 6592 23130 6626
rect 23164 6592 23180 6626
rect 22940 6554 22970 6576
rect 23036 6554 23066 6580
rect 23114 6576 23180 6592
rect 23306 6626 23372 6642
rect 23306 6592 23322 6626
rect 23356 6592 23372 6626
rect 23132 6554 23162 6576
rect 23228 6554 23258 6580
rect 23306 6576 23372 6592
rect 23498 6626 23564 6642
rect 23498 6592 23514 6626
rect 23548 6592 23564 6626
rect 23324 6554 23354 6576
rect 23420 6554 23450 6580
rect 23498 6576 23564 6592
rect 23690 6626 23756 6642
rect 23690 6592 23706 6626
rect 23740 6592 23756 6626
rect 23516 6554 23546 6576
rect 23612 6554 23642 6580
rect 23690 6576 23756 6592
rect 23882 6626 23948 6642
rect 23882 6592 23898 6626
rect 23932 6592 23948 6626
rect 23708 6554 23738 6576
rect 23804 6554 23834 6580
rect 23882 6576 23948 6592
rect 23900 6554 23930 6576
rect 22076 6132 22106 6154
rect 22058 6116 22124 6132
rect 22172 6128 22202 6154
rect 22268 6132 22298 6154
rect 22058 6082 22074 6116
rect 22108 6082 22124 6116
rect 22058 6066 22124 6082
rect 22250 6116 22316 6132
rect 22364 6128 22394 6154
rect 22460 6132 22490 6154
rect 22250 6082 22266 6116
rect 22300 6082 22316 6116
rect 22250 6066 22316 6082
rect 22442 6116 22508 6132
rect 22556 6128 22586 6154
rect 22652 6132 22682 6154
rect 22442 6082 22458 6116
rect 22492 6082 22508 6116
rect 22442 6066 22508 6082
rect 22634 6116 22700 6132
rect 22748 6128 22778 6154
rect 22844 6132 22874 6154
rect 22634 6082 22650 6116
rect 22684 6082 22700 6116
rect 22634 6066 22700 6082
rect 22826 6116 22892 6132
rect 22940 6128 22970 6154
rect 23036 6132 23066 6154
rect 22826 6082 22842 6116
rect 22876 6082 22892 6116
rect 22826 6066 22892 6082
rect 23018 6116 23084 6132
rect 23132 6128 23162 6154
rect 23228 6132 23258 6154
rect 23018 6082 23034 6116
rect 23068 6082 23084 6116
rect 23018 6066 23084 6082
rect 23210 6116 23276 6132
rect 23324 6128 23354 6154
rect 23420 6132 23450 6154
rect 23210 6082 23226 6116
rect 23260 6082 23276 6116
rect 23210 6066 23276 6082
rect 23402 6116 23468 6132
rect 23516 6128 23546 6154
rect 23612 6132 23642 6154
rect 23402 6082 23418 6116
rect 23452 6082 23468 6116
rect 23402 6066 23468 6082
rect 23594 6116 23660 6132
rect 23708 6128 23738 6154
rect 23804 6132 23834 6154
rect 23594 6082 23610 6116
rect 23644 6082 23660 6116
rect 23594 6066 23660 6082
rect 23786 6116 23852 6132
rect 23900 6128 23930 6154
rect 23786 6082 23802 6116
rect 23836 6082 23852 6116
rect 23786 6066 23852 6082
rect 22058 6008 22124 6024
rect 22058 5974 22074 6008
rect 22108 5974 22124 6008
rect 22058 5958 22124 5974
rect 22250 6008 22316 6024
rect 22250 5974 22266 6008
rect 22300 5974 22316 6008
rect 22076 5936 22106 5958
rect 22172 5936 22202 5962
rect 22250 5958 22316 5974
rect 22442 6008 22508 6024
rect 22442 5974 22458 6008
rect 22492 5974 22508 6008
rect 22268 5936 22298 5958
rect 22364 5936 22394 5962
rect 22442 5958 22508 5974
rect 22634 6008 22700 6024
rect 22634 5974 22650 6008
rect 22684 5974 22700 6008
rect 22460 5936 22490 5958
rect 22556 5936 22586 5962
rect 22634 5958 22700 5974
rect 22826 6008 22892 6024
rect 22826 5974 22842 6008
rect 22876 5974 22892 6008
rect 22652 5936 22682 5958
rect 22748 5936 22778 5962
rect 22826 5958 22892 5974
rect 23018 6008 23084 6024
rect 23018 5974 23034 6008
rect 23068 5974 23084 6008
rect 22844 5936 22874 5958
rect 22940 5936 22970 5962
rect 23018 5958 23084 5974
rect 23210 6008 23276 6024
rect 23210 5974 23226 6008
rect 23260 5974 23276 6008
rect 23036 5936 23066 5958
rect 23132 5936 23162 5962
rect 23210 5958 23276 5974
rect 23402 6008 23468 6024
rect 23402 5974 23418 6008
rect 23452 5974 23468 6008
rect 23228 5936 23258 5958
rect 23324 5936 23354 5962
rect 23402 5958 23468 5974
rect 23594 6008 23660 6024
rect 23594 5974 23610 6008
rect 23644 5974 23660 6008
rect 23420 5936 23450 5958
rect 23516 5936 23546 5962
rect 23594 5958 23660 5974
rect 23786 6008 23852 6024
rect 23786 5974 23802 6008
rect 23836 5974 23852 6008
rect 23612 5936 23642 5958
rect 23708 5936 23738 5962
rect 23786 5958 23852 5974
rect 23804 5936 23834 5958
rect 23900 5936 23930 5962
rect 22076 5510 22106 5536
rect 22172 5514 22202 5536
rect 22154 5498 22220 5514
rect 22268 5510 22298 5536
rect 22364 5514 22394 5536
rect 22154 5464 22170 5498
rect 22204 5464 22220 5498
rect 22154 5448 22220 5464
rect 22346 5498 22412 5514
rect 22460 5510 22490 5536
rect 22556 5514 22586 5536
rect 22346 5464 22362 5498
rect 22396 5464 22412 5498
rect 22346 5448 22412 5464
rect 22538 5498 22604 5514
rect 22652 5510 22682 5536
rect 22748 5514 22778 5536
rect 22538 5464 22554 5498
rect 22588 5464 22604 5498
rect 22538 5448 22604 5464
rect 22730 5498 22796 5514
rect 22844 5510 22874 5536
rect 22940 5514 22970 5536
rect 22730 5464 22746 5498
rect 22780 5464 22796 5498
rect 22730 5448 22796 5464
rect 22922 5498 22988 5514
rect 23036 5510 23066 5536
rect 23132 5514 23162 5536
rect 22922 5464 22938 5498
rect 22972 5464 22988 5498
rect 22922 5448 22988 5464
rect 23114 5498 23180 5514
rect 23228 5510 23258 5536
rect 23324 5514 23354 5536
rect 23114 5464 23130 5498
rect 23164 5464 23180 5498
rect 23114 5448 23180 5464
rect 23306 5498 23372 5514
rect 23420 5510 23450 5536
rect 23516 5514 23546 5536
rect 23306 5464 23322 5498
rect 23356 5464 23372 5498
rect 23306 5448 23372 5464
rect 23498 5498 23564 5514
rect 23612 5510 23642 5536
rect 23708 5514 23738 5536
rect 23498 5464 23514 5498
rect 23548 5464 23564 5498
rect 23498 5448 23564 5464
rect 23690 5498 23756 5514
rect 23804 5510 23834 5536
rect 23900 5514 23930 5536
rect 23690 5464 23706 5498
rect 23740 5464 23756 5498
rect 23690 5448 23756 5464
rect 23882 5498 23948 5514
rect 23882 5464 23898 5498
rect 23932 5464 23948 5498
rect 23882 5448 23948 5464
rect 22154 5390 22220 5406
rect 22154 5356 22170 5390
rect 22204 5356 22220 5390
rect 22076 5318 22106 5344
rect 22154 5340 22220 5356
rect 22346 5390 22412 5406
rect 22346 5356 22362 5390
rect 22396 5356 22412 5390
rect 22172 5318 22202 5340
rect 22268 5318 22298 5344
rect 22346 5340 22412 5356
rect 22538 5390 22604 5406
rect 22538 5356 22554 5390
rect 22588 5356 22604 5390
rect 22364 5318 22394 5340
rect 22460 5318 22490 5344
rect 22538 5340 22604 5356
rect 22730 5390 22796 5406
rect 22730 5356 22746 5390
rect 22780 5356 22796 5390
rect 22556 5318 22586 5340
rect 22652 5318 22682 5344
rect 22730 5340 22796 5356
rect 22922 5390 22988 5406
rect 22922 5356 22938 5390
rect 22972 5356 22988 5390
rect 22748 5318 22778 5340
rect 22844 5318 22874 5344
rect 22922 5340 22988 5356
rect 23114 5390 23180 5406
rect 23114 5356 23130 5390
rect 23164 5356 23180 5390
rect 22940 5318 22970 5340
rect 23036 5318 23066 5344
rect 23114 5340 23180 5356
rect 23306 5390 23372 5406
rect 23306 5356 23322 5390
rect 23356 5356 23372 5390
rect 23132 5318 23162 5340
rect 23228 5318 23258 5344
rect 23306 5340 23372 5356
rect 23498 5390 23564 5406
rect 23498 5356 23514 5390
rect 23548 5356 23564 5390
rect 23324 5318 23354 5340
rect 23420 5318 23450 5344
rect 23498 5340 23564 5356
rect 23690 5390 23756 5406
rect 23690 5356 23706 5390
rect 23740 5356 23756 5390
rect 23516 5318 23546 5340
rect 23612 5318 23642 5344
rect 23690 5340 23756 5356
rect 23882 5390 23948 5406
rect 23882 5356 23898 5390
rect 23932 5356 23948 5390
rect 23708 5318 23738 5340
rect 23804 5318 23834 5344
rect 23882 5340 23948 5356
rect 23900 5318 23930 5340
rect 22076 4896 22106 4918
rect 22058 4880 22124 4896
rect 22172 4892 22202 4918
rect 22268 4896 22298 4918
rect 22058 4846 22074 4880
rect 22108 4846 22124 4880
rect 22058 4830 22124 4846
rect 22250 4880 22316 4896
rect 22364 4892 22394 4918
rect 22460 4896 22490 4918
rect 22250 4846 22266 4880
rect 22300 4846 22316 4880
rect 22250 4830 22316 4846
rect 22442 4880 22508 4896
rect 22556 4892 22586 4918
rect 22652 4896 22682 4918
rect 22442 4846 22458 4880
rect 22492 4846 22508 4880
rect 22442 4830 22508 4846
rect 22634 4880 22700 4896
rect 22748 4892 22778 4918
rect 22844 4896 22874 4918
rect 22634 4846 22650 4880
rect 22684 4846 22700 4880
rect 22634 4830 22700 4846
rect 22826 4880 22892 4896
rect 22940 4892 22970 4918
rect 23036 4896 23066 4918
rect 22826 4846 22842 4880
rect 22876 4846 22892 4880
rect 22826 4830 22892 4846
rect 23018 4880 23084 4896
rect 23132 4892 23162 4918
rect 23228 4896 23258 4918
rect 23018 4846 23034 4880
rect 23068 4846 23084 4880
rect 23018 4830 23084 4846
rect 23210 4880 23276 4896
rect 23324 4892 23354 4918
rect 23420 4896 23450 4918
rect 23210 4846 23226 4880
rect 23260 4846 23276 4880
rect 23210 4830 23276 4846
rect 23402 4880 23468 4896
rect 23516 4892 23546 4918
rect 23612 4896 23642 4918
rect 23402 4846 23418 4880
rect 23452 4846 23468 4880
rect 23402 4830 23468 4846
rect 23594 4880 23660 4896
rect 23708 4892 23738 4918
rect 23804 4896 23834 4918
rect 23594 4846 23610 4880
rect 23644 4846 23660 4880
rect 23594 4830 23660 4846
rect 23786 4880 23852 4896
rect 23900 4892 23930 4918
rect 23786 4846 23802 4880
rect 23836 4846 23852 4880
rect 23786 4830 23852 4846
rect 272 3800 472 3816
rect 272 3766 288 3800
rect 456 3766 472 3800
rect 272 3728 472 3766
rect 530 3800 730 3816
rect 530 3766 546 3800
rect 714 3766 730 3800
rect 530 3728 730 3766
rect 788 3800 988 3816
rect 788 3766 804 3800
rect 972 3766 988 3800
rect 788 3728 988 3766
rect 1046 3800 1246 3816
rect 1046 3766 1062 3800
rect 1230 3766 1246 3800
rect 1046 3728 1246 3766
rect 1304 3800 1504 3816
rect 1304 3766 1320 3800
rect 1488 3766 1504 3800
rect 1304 3728 1504 3766
rect 272 3290 472 3328
rect 272 3256 288 3290
rect 456 3256 472 3290
rect 272 3240 472 3256
rect 530 3290 730 3328
rect 530 3256 546 3290
rect 714 3256 730 3290
rect 530 3240 730 3256
rect 788 3290 988 3328
rect 788 3256 804 3290
rect 972 3256 988 3290
rect 788 3240 988 3256
rect 1046 3290 1246 3328
rect 1046 3256 1062 3290
rect 1230 3256 1246 3290
rect 1046 3240 1246 3256
rect 1304 3290 1504 3328
rect 1304 3256 1320 3290
rect 1488 3256 1504 3290
rect 1304 3240 1504 3256
rect 272 3182 472 3198
rect 272 3148 288 3182
rect 456 3148 472 3182
rect 272 3110 472 3148
rect 530 3182 730 3198
rect 530 3148 546 3182
rect 714 3148 730 3182
rect 530 3110 730 3148
rect 788 3182 988 3198
rect 788 3148 804 3182
rect 972 3148 988 3182
rect 788 3110 988 3148
rect 1046 3182 1246 3198
rect 1046 3148 1062 3182
rect 1230 3148 1246 3182
rect 1046 3110 1246 3148
rect 1304 3182 1504 3198
rect 1304 3148 1320 3182
rect 1488 3148 1504 3182
rect 1304 3110 1504 3148
rect 272 2672 472 2710
rect 272 2638 288 2672
rect 456 2638 472 2672
rect 272 2622 472 2638
rect 530 2672 730 2710
rect 530 2638 546 2672
rect 714 2638 730 2672
rect 530 2622 730 2638
rect 788 2672 988 2710
rect 788 2638 804 2672
rect 972 2638 988 2672
rect 788 2622 988 2638
rect 1046 2672 1246 2710
rect 1046 2638 1062 2672
rect 1230 2638 1246 2672
rect 1046 2622 1246 2638
rect 1304 2672 1504 2710
rect 1304 2638 1320 2672
rect 1488 2638 1504 2672
rect 1304 2622 1504 2638
rect 272 2564 472 2580
rect 272 2530 288 2564
rect 456 2530 472 2564
rect 272 2492 472 2530
rect 530 2564 730 2580
rect 530 2530 546 2564
rect 714 2530 730 2564
rect 530 2492 730 2530
rect 788 2564 988 2580
rect 788 2530 804 2564
rect 972 2530 988 2564
rect 788 2492 988 2530
rect 1046 2564 1246 2580
rect 1046 2530 1062 2564
rect 1230 2530 1246 2564
rect 1046 2492 1246 2530
rect 1304 2564 1504 2580
rect 1304 2530 1320 2564
rect 1488 2530 1504 2564
rect 1304 2492 1504 2530
rect 272 2054 472 2092
rect 272 2020 288 2054
rect 456 2020 472 2054
rect 272 2004 472 2020
rect 530 2054 730 2092
rect 530 2020 546 2054
rect 714 2020 730 2054
rect 530 2004 730 2020
rect 788 2054 988 2092
rect 788 2020 804 2054
rect 972 2020 988 2054
rect 788 2004 988 2020
rect 1046 2054 1246 2092
rect 1046 2020 1062 2054
rect 1230 2020 1246 2054
rect 1046 2004 1246 2020
rect 1304 2054 1504 2092
rect 1304 2020 1320 2054
rect 1488 2020 1504 2054
rect 1304 2004 1504 2020
rect 272 1946 472 1962
rect 272 1912 288 1946
rect 456 1912 472 1946
rect 272 1874 472 1912
rect 530 1946 730 1962
rect 530 1912 546 1946
rect 714 1912 730 1946
rect 530 1874 730 1912
rect 788 1946 988 1962
rect 788 1912 804 1946
rect 972 1912 988 1946
rect 788 1874 988 1912
rect 1046 1946 1246 1962
rect 1046 1912 1062 1946
rect 1230 1912 1246 1946
rect 1046 1874 1246 1912
rect 1304 1946 1504 1962
rect 1304 1912 1320 1946
rect 1488 1912 1504 1946
rect 1304 1874 1504 1912
rect 272 1436 472 1474
rect 272 1402 288 1436
rect 456 1402 472 1436
rect 272 1386 472 1402
rect 530 1436 730 1474
rect 530 1402 546 1436
rect 714 1402 730 1436
rect 530 1386 730 1402
rect 788 1436 988 1474
rect 788 1402 804 1436
rect 972 1402 988 1436
rect 788 1386 988 1402
rect 1046 1436 1246 1474
rect 1046 1402 1062 1436
rect 1230 1402 1246 1436
rect 1046 1386 1246 1402
rect 1304 1436 1504 1474
rect 1304 1402 1320 1436
rect 1488 1402 1504 1436
rect 1304 1386 1504 1402
rect 272 1328 472 1344
rect 272 1294 288 1328
rect 456 1294 472 1328
rect 272 1256 472 1294
rect 530 1328 730 1344
rect 530 1294 546 1328
rect 714 1294 730 1328
rect 530 1256 730 1294
rect 788 1328 988 1344
rect 788 1294 804 1328
rect 972 1294 988 1328
rect 788 1256 988 1294
rect 1046 1328 1246 1344
rect 1046 1294 1062 1328
rect 1230 1294 1246 1328
rect 1046 1256 1246 1294
rect 1304 1328 1504 1344
rect 1304 1294 1320 1328
rect 1488 1294 1504 1328
rect 1304 1256 1504 1294
rect 272 818 472 856
rect 272 784 288 818
rect 456 784 472 818
rect 272 768 472 784
rect 530 818 730 856
rect 530 784 546 818
rect 714 784 730 818
rect 530 768 730 784
rect 788 818 988 856
rect 788 784 804 818
rect 972 784 988 818
rect 788 768 988 784
rect 1046 818 1246 856
rect 1046 784 1062 818
rect 1230 784 1246 818
rect 1046 768 1246 784
rect 1304 818 1504 856
rect 1304 784 1320 818
rect 1488 784 1504 818
rect 1304 768 1504 784
rect 272 710 472 726
rect 272 676 288 710
rect 456 676 472 710
rect 272 638 472 676
rect 530 710 730 726
rect 530 676 546 710
rect 714 676 730 710
rect 530 638 730 676
rect 788 710 988 726
rect 788 676 804 710
rect 972 676 988 710
rect 788 638 988 676
rect 1046 710 1246 726
rect 1046 676 1062 710
rect 1230 676 1246 710
rect 1046 638 1246 676
rect 1304 710 1504 726
rect 1304 676 1320 710
rect 1488 676 1504 710
rect 1304 638 1504 676
rect 272 200 472 238
rect 272 166 288 200
rect 456 166 472 200
rect 272 150 472 166
rect 530 200 730 238
rect 530 166 546 200
rect 714 166 730 200
rect 530 150 730 166
rect 788 200 988 238
rect 788 166 804 200
rect 972 166 988 200
rect 788 150 988 166
rect 1046 200 1246 238
rect 1046 166 1062 200
rect 1230 166 1246 200
rect 1046 150 1246 166
rect 1304 200 1504 238
rect 1304 166 1320 200
rect 1488 166 1504 200
rect 1304 150 1504 166
rect 2072 3800 2272 3816
rect 2072 3766 2088 3800
rect 2256 3766 2272 3800
rect 2072 3728 2272 3766
rect 2330 3800 2530 3816
rect 2330 3766 2346 3800
rect 2514 3766 2530 3800
rect 2330 3728 2530 3766
rect 2588 3800 2788 3816
rect 2588 3766 2604 3800
rect 2772 3766 2788 3800
rect 2588 3728 2788 3766
rect 2846 3800 3046 3816
rect 2846 3766 2862 3800
rect 3030 3766 3046 3800
rect 2846 3728 3046 3766
rect 3104 3800 3304 3816
rect 3104 3766 3120 3800
rect 3288 3766 3304 3800
rect 3104 3728 3304 3766
rect 2072 3290 2272 3328
rect 2072 3256 2088 3290
rect 2256 3256 2272 3290
rect 2072 3240 2272 3256
rect 2330 3290 2530 3328
rect 2330 3256 2346 3290
rect 2514 3256 2530 3290
rect 2330 3240 2530 3256
rect 2588 3290 2788 3328
rect 2588 3256 2604 3290
rect 2772 3256 2788 3290
rect 2588 3240 2788 3256
rect 2846 3290 3046 3328
rect 2846 3256 2862 3290
rect 3030 3256 3046 3290
rect 2846 3240 3046 3256
rect 3104 3290 3304 3328
rect 3104 3256 3120 3290
rect 3288 3256 3304 3290
rect 3104 3240 3304 3256
rect 2072 3182 2272 3198
rect 2072 3148 2088 3182
rect 2256 3148 2272 3182
rect 2072 3110 2272 3148
rect 2330 3182 2530 3198
rect 2330 3148 2346 3182
rect 2514 3148 2530 3182
rect 2330 3110 2530 3148
rect 2588 3182 2788 3198
rect 2588 3148 2604 3182
rect 2772 3148 2788 3182
rect 2588 3110 2788 3148
rect 2846 3182 3046 3198
rect 2846 3148 2862 3182
rect 3030 3148 3046 3182
rect 2846 3110 3046 3148
rect 3104 3182 3304 3198
rect 3104 3148 3120 3182
rect 3288 3148 3304 3182
rect 3104 3110 3304 3148
rect 2072 2672 2272 2710
rect 2072 2638 2088 2672
rect 2256 2638 2272 2672
rect 2072 2622 2272 2638
rect 2330 2672 2530 2710
rect 2330 2638 2346 2672
rect 2514 2638 2530 2672
rect 2330 2622 2530 2638
rect 2588 2672 2788 2710
rect 2588 2638 2604 2672
rect 2772 2638 2788 2672
rect 2588 2622 2788 2638
rect 2846 2672 3046 2710
rect 2846 2638 2862 2672
rect 3030 2638 3046 2672
rect 2846 2622 3046 2638
rect 3104 2672 3304 2710
rect 3104 2638 3120 2672
rect 3288 2638 3304 2672
rect 3104 2622 3304 2638
rect 2072 2564 2272 2580
rect 2072 2530 2088 2564
rect 2256 2530 2272 2564
rect 2072 2492 2272 2530
rect 2330 2564 2530 2580
rect 2330 2530 2346 2564
rect 2514 2530 2530 2564
rect 2330 2492 2530 2530
rect 2588 2564 2788 2580
rect 2588 2530 2604 2564
rect 2772 2530 2788 2564
rect 2588 2492 2788 2530
rect 2846 2564 3046 2580
rect 2846 2530 2862 2564
rect 3030 2530 3046 2564
rect 2846 2492 3046 2530
rect 3104 2564 3304 2580
rect 3104 2530 3120 2564
rect 3288 2530 3304 2564
rect 3104 2492 3304 2530
rect 2072 2054 2272 2092
rect 2072 2020 2088 2054
rect 2256 2020 2272 2054
rect 2072 2004 2272 2020
rect 2330 2054 2530 2092
rect 2330 2020 2346 2054
rect 2514 2020 2530 2054
rect 2330 2004 2530 2020
rect 2588 2054 2788 2092
rect 2588 2020 2604 2054
rect 2772 2020 2788 2054
rect 2588 2004 2788 2020
rect 2846 2054 3046 2092
rect 2846 2020 2862 2054
rect 3030 2020 3046 2054
rect 2846 2004 3046 2020
rect 3104 2054 3304 2092
rect 3104 2020 3120 2054
rect 3288 2020 3304 2054
rect 3104 2004 3304 2020
rect 2072 1946 2272 1962
rect 2072 1912 2088 1946
rect 2256 1912 2272 1946
rect 2072 1874 2272 1912
rect 2330 1946 2530 1962
rect 2330 1912 2346 1946
rect 2514 1912 2530 1946
rect 2330 1874 2530 1912
rect 2588 1946 2788 1962
rect 2588 1912 2604 1946
rect 2772 1912 2788 1946
rect 2588 1874 2788 1912
rect 2846 1946 3046 1962
rect 2846 1912 2862 1946
rect 3030 1912 3046 1946
rect 2846 1874 3046 1912
rect 3104 1946 3304 1962
rect 3104 1912 3120 1946
rect 3288 1912 3304 1946
rect 3104 1874 3304 1912
rect 2072 1436 2272 1474
rect 2072 1402 2088 1436
rect 2256 1402 2272 1436
rect 2072 1386 2272 1402
rect 2330 1436 2530 1474
rect 2330 1402 2346 1436
rect 2514 1402 2530 1436
rect 2330 1386 2530 1402
rect 2588 1436 2788 1474
rect 2588 1402 2604 1436
rect 2772 1402 2788 1436
rect 2588 1386 2788 1402
rect 2846 1436 3046 1474
rect 2846 1402 2862 1436
rect 3030 1402 3046 1436
rect 2846 1386 3046 1402
rect 3104 1436 3304 1474
rect 3104 1402 3120 1436
rect 3288 1402 3304 1436
rect 3104 1386 3304 1402
rect 2072 1328 2272 1344
rect 2072 1294 2088 1328
rect 2256 1294 2272 1328
rect 2072 1256 2272 1294
rect 2330 1328 2530 1344
rect 2330 1294 2346 1328
rect 2514 1294 2530 1328
rect 2330 1256 2530 1294
rect 2588 1328 2788 1344
rect 2588 1294 2604 1328
rect 2772 1294 2788 1328
rect 2588 1256 2788 1294
rect 2846 1328 3046 1344
rect 2846 1294 2862 1328
rect 3030 1294 3046 1328
rect 2846 1256 3046 1294
rect 3104 1328 3304 1344
rect 3104 1294 3120 1328
rect 3288 1294 3304 1328
rect 3104 1256 3304 1294
rect 2072 818 2272 856
rect 2072 784 2088 818
rect 2256 784 2272 818
rect 2072 768 2272 784
rect 2330 818 2530 856
rect 2330 784 2346 818
rect 2514 784 2530 818
rect 2330 768 2530 784
rect 2588 818 2788 856
rect 2588 784 2604 818
rect 2772 784 2788 818
rect 2588 768 2788 784
rect 2846 818 3046 856
rect 2846 784 2862 818
rect 3030 784 3046 818
rect 2846 768 3046 784
rect 3104 818 3304 856
rect 3104 784 3120 818
rect 3288 784 3304 818
rect 3104 768 3304 784
rect 2072 710 2272 726
rect 2072 676 2088 710
rect 2256 676 2272 710
rect 2072 638 2272 676
rect 2330 710 2530 726
rect 2330 676 2346 710
rect 2514 676 2530 710
rect 2330 638 2530 676
rect 2588 710 2788 726
rect 2588 676 2604 710
rect 2772 676 2788 710
rect 2588 638 2788 676
rect 2846 710 3046 726
rect 2846 676 2862 710
rect 3030 676 3046 710
rect 2846 638 3046 676
rect 3104 710 3304 726
rect 3104 676 3120 710
rect 3288 676 3304 710
rect 3104 638 3304 676
rect 2072 200 2272 238
rect 2072 166 2088 200
rect 2256 166 2272 200
rect 2072 150 2272 166
rect 2330 200 2530 238
rect 2330 166 2346 200
rect 2514 166 2530 200
rect 2330 150 2530 166
rect 2588 200 2788 238
rect 2588 166 2604 200
rect 2772 166 2788 200
rect 2588 150 2788 166
rect 2846 200 3046 238
rect 2846 166 2862 200
rect 3030 166 3046 200
rect 2846 150 3046 166
rect 3104 200 3304 238
rect 3104 166 3120 200
rect 3288 166 3304 200
rect 3104 150 3304 166
rect 3872 3800 4072 3816
rect 3872 3766 3888 3800
rect 4056 3766 4072 3800
rect 3872 3728 4072 3766
rect 4130 3800 4330 3816
rect 4130 3766 4146 3800
rect 4314 3766 4330 3800
rect 4130 3728 4330 3766
rect 4388 3800 4588 3816
rect 4388 3766 4404 3800
rect 4572 3766 4588 3800
rect 4388 3728 4588 3766
rect 4646 3800 4846 3816
rect 4646 3766 4662 3800
rect 4830 3766 4846 3800
rect 4646 3728 4846 3766
rect 4904 3800 5104 3816
rect 4904 3766 4920 3800
rect 5088 3766 5104 3800
rect 4904 3728 5104 3766
rect 3872 3290 4072 3328
rect 3872 3256 3888 3290
rect 4056 3256 4072 3290
rect 3872 3240 4072 3256
rect 4130 3290 4330 3328
rect 4130 3256 4146 3290
rect 4314 3256 4330 3290
rect 4130 3240 4330 3256
rect 4388 3290 4588 3328
rect 4388 3256 4404 3290
rect 4572 3256 4588 3290
rect 4388 3240 4588 3256
rect 4646 3290 4846 3328
rect 4646 3256 4662 3290
rect 4830 3256 4846 3290
rect 4646 3240 4846 3256
rect 4904 3290 5104 3328
rect 4904 3256 4920 3290
rect 5088 3256 5104 3290
rect 4904 3240 5104 3256
rect 3872 3182 4072 3198
rect 3872 3148 3888 3182
rect 4056 3148 4072 3182
rect 3872 3110 4072 3148
rect 4130 3182 4330 3198
rect 4130 3148 4146 3182
rect 4314 3148 4330 3182
rect 4130 3110 4330 3148
rect 4388 3182 4588 3198
rect 4388 3148 4404 3182
rect 4572 3148 4588 3182
rect 4388 3110 4588 3148
rect 4646 3182 4846 3198
rect 4646 3148 4662 3182
rect 4830 3148 4846 3182
rect 4646 3110 4846 3148
rect 4904 3182 5104 3198
rect 4904 3148 4920 3182
rect 5088 3148 5104 3182
rect 4904 3110 5104 3148
rect 3872 2672 4072 2710
rect 3872 2638 3888 2672
rect 4056 2638 4072 2672
rect 3872 2622 4072 2638
rect 4130 2672 4330 2710
rect 4130 2638 4146 2672
rect 4314 2638 4330 2672
rect 4130 2622 4330 2638
rect 4388 2672 4588 2710
rect 4388 2638 4404 2672
rect 4572 2638 4588 2672
rect 4388 2622 4588 2638
rect 4646 2672 4846 2710
rect 4646 2638 4662 2672
rect 4830 2638 4846 2672
rect 4646 2622 4846 2638
rect 4904 2672 5104 2710
rect 4904 2638 4920 2672
rect 5088 2638 5104 2672
rect 4904 2622 5104 2638
rect 3872 2564 4072 2580
rect 3872 2530 3888 2564
rect 4056 2530 4072 2564
rect 3872 2492 4072 2530
rect 4130 2564 4330 2580
rect 4130 2530 4146 2564
rect 4314 2530 4330 2564
rect 4130 2492 4330 2530
rect 4388 2564 4588 2580
rect 4388 2530 4404 2564
rect 4572 2530 4588 2564
rect 4388 2492 4588 2530
rect 4646 2564 4846 2580
rect 4646 2530 4662 2564
rect 4830 2530 4846 2564
rect 4646 2492 4846 2530
rect 4904 2564 5104 2580
rect 4904 2530 4920 2564
rect 5088 2530 5104 2564
rect 4904 2492 5104 2530
rect 3872 2054 4072 2092
rect 3872 2020 3888 2054
rect 4056 2020 4072 2054
rect 3872 2004 4072 2020
rect 4130 2054 4330 2092
rect 4130 2020 4146 2054
rect 4314 2020 4330 2054
rect 4130 2004 4330 2020
rect 4388 2054 4588 2092
rect 4388 2020 4404 2054
rect 4572 2020 4588 2054
rect 4388 2004 4588 2020
rect 4646 2054 4846 2092
rect 4646 2020 4662 2054
rect 4830 2020 4846 2054
rect 4646 2004 4846 2020
rect 4904 2054 5104 2092
rect 4904 2020 4920 2054
rect 5088 2020 5104 2054
rect 4904 2004 5104 2020
rect 3872 1946 4072 1962
rect 3872 1912 3888 1946
rect 4056 1912 4072 1946
rect 3872 1874 4072 1912
rect 4130 1946 4330 1962
rect 4130 1912 4146 1946
rect 4314 1912 4330 1946
rect 4130 1874 4330 1912
rect 4388 1946 4588 1962
rect 4388 1912 4404 1946
rect 4572 1912 4588 1946
rect 4388 1874 4588 1912
rect 4646 1946 4846 1962
rect 4646 1912 4662 1946
rect 4830 1912 4846 1946
rect 4646 1874 4846 1912
rect 4904 1946 5104 1962
rect 4904 1912 4920 1946
rect 5088 1912 5104 1946
rect 4904 1874 5104 1912
rect 3872 1436 4072 1474
rect 3872 1402 3888 1436
rect 4056 1402 4072 1436
rect 3872 1386 4072 1402
rect 4130 1436 4330 1474
rect 4130 1402 4146 1436
rect 4314 1402 4330 1436
rect 4130 1386 4330 1402
rect 4388 1436 4588 1474
rect 4388 1402 4404 1436
rect 4572 1402 4588 1436
rect 4388 1386 4588 1402
rect 4646 1436 4846 1474
rect 4646 1402 4662 1436
rect 4830 1402 4846 1436
rect 4646 1386 4846 1402
rect 4904 1436 5104 1474
rect 4904 1402 4920 1436
rect 5088 1402 5104 1436
rect 4904 1386 5104 1402
rect 3872 1328 4072 1344
rect 3872 1294 3888 1328
rect 4056 1294 4072 1328
rect 3872 1256 4072 1294
rect 4130 1328 4330 1344
rect 4130 1294 4146 1328
rect 4314 1294 4330 1328
rect 4130 1256 4330 1294
rect 4388 1328 4588 1344
rect 4388 1294 4404 1328
rect 4572 1294 4588 1328
rect 4388 1256 4588 1294
rect 4646 1328 4846 1344
rect 4646 1294 4662 1328
rect 4830 1294 4846 1328
rect 4646 1256 4846 1294
rect 4904 1328 5104 1344
rect 4904 1294 4920 1328
rect 5088 1294 5104 1328
rect 4904 1256 5104 1294
rect 3872 818 4072 856
rect 3872 784 3888 818
rect 4056 784 4072 818
rect 3872 768 4072 784
rect 4130 818 4330 856
rect 4130 784 4146 818
rect 4314 784 4330 818
rect 4130 768 4330 784
rect 4388 818 4588 856
rect 4388 784 4404 818
rect 4572 784 4588 818
rect 4388 768 4588 784
rect 4646 818 4846 856
rect 4646 784 4662 818
rect 4830 784 4846 818
rect 4646 768 4846 784
rect 4904 818 5104 856
rect 4904 784 4920 818
rect 5088 784 5104 818
rect 4904 768 5104 784
rect 3872 710 4072 726
rect 3872 676 3888 710
rect 4056 676 4072 710
rect 3872 638 4072 676
rect 4130 710 4330 726
rect 4130 676 4146 710
rect 4314 676 4330 710
rect 4130 638 4330 676
rect 4388 710 4588 726
rect 4388 676 4404 710
rect 4572 676 4588 710
rect 4388 638 4588 676
rect 4646 710 4846 726
rect 4646 676 4662 710
rect 4830 676 4846 710
rect 4646 638 4846 676
rect 4904 710 5104 726
rect 4904 676 4920 710
rect 5088 676 5104 710
rect 4904 638 5104 676
rect 3872 200 4072 238
rect 3872 166 3888 200
rect 4056 166 4072 200
rect 3872 150 4072 166
rect 4130 200 4330 238
rect 4130 166 4146 200
rect 4314 166 4330 200
rect 4130 150 4330 166
rect 4388 200 4588 238
rect 4388 166 4404 200
rect 4572 166 4588 200
rect 4388 150 4588 166
rect 4646 200 4846 238
rect 4646 166 4662 200
rect 4830 166 4846 200
rect 4646 150 4846 166
rect 4904 200 5104 238
rect 4904 166 4920 200
rect 5088 166 5104 200
rect 4904 150 5104 166
rect 5672 3800 5872 3816
rect 5672 3766 5688 3800
rect 5856 3766 5872 3800
rect 5672 3728 5872 3766
rect 5930 3800 6130 3816
rect 5930 3766 5946 3800
rect 6114 3766 6130 3800
rect 5930 3728 6130 3766
rect 6188 3800 6388 3816
rect 6188 3766 6204 3800
rect 6372 3766 6388 3800
rect 6188 3728 6388 3766
rect 6446 3800 6646 3816
rect 6446 3766 6462 3800
rect 6630 3766 6646 3800
rect 6446 3728 6646 3766
rect 6704 3800 6904 3816
rect 6704 3766 6720 3800
rect 6888 3766 6904 3800
rect 6704 3728 6904 3766
rect 5672 3290 5872 3328
rect 5672 3256 5688 3290
rect 5856 3256 5872 3290
rect 5672 3240 5872 3256
rect 5930 3290 6130 3328
rect 5930 3256 5946 3290
rect 6114 3256 6130 3290
rect 5930 3240 6130 3256
rect 6188 3290 6388 3328
rect 6188 3256 6204 3290
rect 6372 3256 6388 3290
rect 6188 3240 6388 3256
rect 6446 3290 6646 3328
rect 6446 3256 6462 3290
rect 6630 3256 6646 3290
rect 6446 3240 6646 3256
rect 6704 3290 6904 3328
rect 6704 3256 6720 3290
rect 6888 3256 6904 3290
rect 6704 3240 6904 3256
rect 5672 3182 5872 3198
rect 5672 3148 5688 3182
rect 5856 3148 5872 3182
rect 5672 3110 5872 3148
rect 5930 3182 6130 3198
rect 5930 3148 5946 3182
rect 6114 3148 6130 3182
rect 5930 3110 6130 3148
rect 6188 3182 6388 3198
rect 6188 3148 6204 3182
rect 6372 3148 6388 3182
rect 6188 3110 6388 3148
rect 6446 3182 6646 3198
rect 6446 3148 6462 3182
rect 6630 3148 6646 3182
rect 6446 3110 6646 3148
rect 6704 3182 6904 3198
rect 6704 3148 6720 3182
rect 6888 3148 6904 3182
rect 6704 3110 6904 3148
rect 5672 2672 5872 2710
rect 5672 2638 5688 2672
rect 5856 2638 5872 2672
rect 5672 2622 5872 2638
rect 5930 2672 6130 2710
rect 5930 2638 5946 2672
rect 6114 2638 6130 2672
rect 5930 2622 6130 2638
rect 6188 2672 6388 2710
rect 6188 2638 6204 2672
rect 6372 2638 6388 2672
rect 6188 2622 6388 2638
rect 6446 2672 6646 2710
rect 6446 2638 6462 2672
rect 6630 2638 6646 2672
rect 6446 2622 6646 2638
rect 6704 2672 6904 2710
rect 6704 2638 6720 2672
rect 6888 2638 6904 2672
rect 6704 2622 6904 2638
rect 5672 2564 5872 2580
rect 5672 2530 5688 2564
rect 5856 2530 5872 2564
rect 5672 2492 5872 2530
rect 5930 2564 6130 2580
rect 5930 2530 5946 2564
rect 6114 2530 6130 2564
rect 5930 2492 6130 2530
rect 6188 2564 6388 2580
rect 6188 2530 6204 2564
rect 6372 2530 6388 2564
rect 6188 2492 6388 2530
rect 6446 2564 6646 2580
rect 6446 2530 6462 2564
rect 6630 2530 6646 2564
rect 6446 2492 6646 2530
rect 6704 2564 6904 2580
rect 6704 2530 6720 2564
rect 6888 2530 6904 2564
rect 6704 2492 6904 2530
rect 5672 2054 5872 2092
rect 5672 2020 5688 2054
rect 5856 2020 5872 2054
rect 5672 2004 5872 2020
rect 5930 2054 6130 2092
rect 5930 2020 5946 2054
rect 6114 2020 6130 2054
rect 5930 2004 6130 2020
rect 6188 2054 6388 2092
rect 6188 2020 6204 2054
rect 6372 2020 6388 2054
rect 6188 2004 6388 2020
rect 6446 2054 6646 2092
rect 6446 2020 6462 2054
rect 6630 2020 6646 2054
rect 6446 2004 6646 2020
rect 6704 2054 6904 2092
rect 6704 2020 6720 2054
rect 6888 2020 6904 2054
rect 6704 2004 6904 2020
rect 5672 1946 5872 1962
rect 5672 1912 5688 1946
rect 5856 1912 5872 1946
rect 5672 1874 5872 1912
rect 5930 1946 6130 1962
rect 5930 1912 5946 1946
rect 6114 1912 6130 1946
rect 5930 1874 6130 1912
rect 6188 1946 6388 1962
rect 6188 1912 6204 1946
rect 6372 1912 6388 1946
rect 6188 1874 6388 1912
rect 6446 1946 6646 1962
rect 6446 1912 6462 1946
rect 6630 1912 6646 1946
rect 6446 1874 6646 1912
rect 6704 1946 6904 1962
rect 6704 1912 6720 1946
rect 6888 1912 6904 1946
rect 6704 1874 6904 1912
rect 5672 1436 5872 1474
rect 5672 1402 5688 1436
rect 5856 1402 5872 1436
rect 5672 1386 5872 1402
rect 5930 1436 6130 1474
rect 5930 1402 5946 1436
rect 6114 1402 6130 1436
rect 5930 1386 6130 1402
rect 6188 1436 6388 1474
rect 6188 1402 6204 1436
rect 6372 1402 6388 1436
rect 6188 1386 6388 1402
rect 6446 1436 6646 1474
rect 6446 1402 6462 1436
rect 6630 1402 6646 1436
rect 6446 1386 6646 1402
rect 6704 1436 6904 1474
rect 6704 1402 6720 1436
rect 6888 1402 6904 1436
rect 6704 1386 6904 1402
rect 5672 1328 5872 1344
rect 5672 1294 5688 1328
rect 5856 1294 5872 1328
rect 5672 1256 5872 1294
rect 5930 1328 6130 1344
rect 5930 1294 5946 1328
rect 6114 1294 6130 1328
rect 5930 1256 6130 1294
rect 6188 1328 6388 1344
rect 6188 1294 6204 1328
rect 6372 1294 6388 1328
rect 6188 1256 6388 1294
rect 6446 1328 6646 1344
rect 6446 1294 6462 1328
rect 6630 1294 6646 1328
rect 6446 1256 6646 1294
rect 6704 1328 6904 1344
rect 6704 1294 6720 1328
rect 6888 1294 6904 1328
rect 6704 1256 6904 1294
rect 5672 818 5872 856
rect 5672 784 5688 818
rect 5856 784 5872 818
rect 5672 768 5872 784
rect 5930 818 6130 856
rect 5930 784 5946 818
rect 6114 784 6130 818
rect 5930 768 6130 784
rect 6188 818 6388 856
rect 6188 784 6204 818
rect 6372 784 6388 818
rect 6188 768 6388 784
rect 6446 818 6646 856
rect 6446 784 6462 818
rect 6630 784 6646 818
rect 6446 768 6646 784
rect 6704 818 6904 856
rect 6704 784 6720 818
rect 6888 784 6904 818
rect 6704 768 6904 784
rect 5672 710 5872 726
rect 5672 676 5688 710
rect 5856 676 5872 710
rect 5672 638 5872 676
rect 5930 710 6130 726
rect 5930 676 5946 710
rect 6114 676 6130 710
rect 5930 638 6130 676
rect 6188 710 6388 726
rect 6188 676 6204 710
rect 6372 676 6388 710
rect 6188 638 6388 676
rect 6446 710 6646 726
rect 6446 676 6462 710
rect 6630 676 6646 710
rect 6446 638 6646 676
rect 6704 710 6904 726
rect 6704 676 6720 710
rect 6888 676 6904 710
rect 6704 638 6904 676
rect 5672 200 5872 238
rect 5672 166 5688 200
rect 5856 166 5872 200
rect 5672 150 5872 166
rect 5930 200 6130 238
rect 5930 166 5946 200
rect 6114 166 6130 200
rect 5930 150 6130 166
rect 6188 200 6388 238
rect 6188 166 6204 200
rect 6372 166 6388 200
rect 6188 150 6388 166
rect 6446 200 6646 238
rect 6446 166 6462 200
rect 6630 166 6646 200
rect 6446 150 6646 166
rect 6704 200 6904 238
rect 6704 166 6720 200
rect 6888 166 6904 200
rect 6704 150 6904 166
rect 14672 3800 14872 3816
rect 14672 3766 14688 3800
rect 14856 3766 14872 3800
rect 14672 3728 14872 3766
rect 14930 3800 15130 3816
rect 14930 3766 14946 3800
rect 15114 3766 15130 3800
rect 14930 3728 15130 3766
rect 15188 3800 15388 3816
rect 15188 3766 15204 3800
rect 15372 3766 15388 3800
rect 15188 3728 15388 3766
rect 15446 3800 15646 3816
rect 15446 3766 15462 3800
rect 15630 3766 15646 3800
rect 15446 3728 15646 3766
rect 15704 3800 15904 3816
rect 15704 3766 15720 3800
rect 15888 3766 15904 3800
rect 15704 3728 15904 3766
rect 14672 3290 14872 3328
rect 14672 3256 14688 3290
rect 14856 3256 14872 3290
rect 14672 3240 14872 3256
rect 14930 3290 15130 3328
rect 14930 3256 14946 3290
rect 15114 3256 15130 3290
rect 14930 3240 15130 3256
rect 15188 3290 15388 3328
rect 15188 3256 15204 3290
rect 15372 3256 15388 3290
rect 15188 3240 15388 3256
rect 15446 3290 15646 3328
rect 15446 3256 15462 3290
rect 15630 3256 15646 3290
rect 15446 3240 15646 3256
rect 15704 3290 15904 3328
rect 15704 3256 15720 3290
rect 15888 3256 15904 3290
rect 15704 3240 15904 3256
rect 14672 3182 14872 3198
rect 14672 3148 14688 3182
rect 14856 3148 14872 3182
rect 14672 3110 14872 3148
rect 14930 3182 15130 3198
rect 14930 3148 14946 3182
rect 15114 3148 15130 3182
rect 14930 3110 15130 3148
rect 15188 3182 15388 3198
rect 15188 3148 15204 3182
rect 15372 3148 15388 3182
rect 15188 3110 15388 3148
rect 15446 3182 15646 3198
rect 15446 3148 15462 3182
rect 15630 3148 15646 3182
rect 15446 3110 15646 3148
rect 15704 3182 15904 3198
rect 15704 3148 15720 3182
rect 15888 3148 15904 3182
rect 15704 3110 15904 3148
rect 14672 2672 14872 2710
rect 14672 2638 14688 2672
rect 14856 2638 14872 2672
rect 14672 2622 14872 2638
rect 14930 2672 15130 2710
rect 14930 2638 14946 2672
rect 15114 2638 15130 2672
rect 14930 2622 15130 2638
rect 15188 2672 15388 2710
rect 15188 2638 15204 2672
rect 15372 2638 15388 2672
rect 15188 2622 15388 2638
rect 15446 2672 15646 2710
rect 15446 2638 15462 2672
rect 15630 2638 15646 2672
rect 15446 2622 15646 2638
rect 15704 2672 15904 2710
rect 15704 2638 15720 2672
rect 15888 2638 15904 2672
rect 15704 2622 15904 2638
rect 14672 2564 14872 2580
rect 14672 2530 14688 2564
rect 14856 2530 14872 2564
rect 14672 2492 14872 2530
rect 14930 2564 15130 2580
rect 14930 2530 14946 2564
rect 15114 2530 15130 2564
rect 14930 2492 15130 2530
rect 15188 2564 15388 2580
rect 15188 2530 15204 2564
rect 15372 2530 15388 2564
rect 15188 2492 15388 2530
rect 15446 2564 15646 2580
rect 15446 2530 15462 2564
rect 15630 2530 15646 2564
rect 15446 2492 15646 2530
rect 15704 2564 15904 2580
rect 15704 2530 15720 2564
rect 15888 2530 15904 2564
rect 15704 2492 15904 2530
rect 14672 2054 14872 2092
rect 14672 2020 14688 2054
rect 14856 2020 14872 2054
rect 14672 2004 14872 2020
rect 14930 2054 15130 2092
rect 14930 2020 14946 2054
rect 15114 2020 15130 2054
rect 14930 2004 15130 2020
rect 15188 2054 15388 2092
rect 15188 2020 15204 2054
rect 15372 2020 15388 2054
rect 15188 2004 15388 2020
rect 15446 2054 15646 2092
rect 15446 2020 15462 2054
rect 15630 2020 15646 2054
rect 15446 2004 15646 2020
rect 15704 2054 15904 2092
rect 15704 2020 15720 2054
rect 15888 2020 15904 2054
rect 15704 2004 15904 2020
rect 14672 1946 14872 1962
rect 14672 1912 14688 1946
rect 14856 1912 14872 1946
rect 14672 1874 14872 1912
rect 14930 1946 15130 1962
rect 14930 1912 14946 1946
rect 15114 1912 15130 1946
rect 14930 1874 15130 1912
rect 15188 1946 15388 1962
rect 15188 1912 15204 1946
rect 15372 1912 15388 1946
rect 15188 1874 15388 1912
rect 15446 1946 15646 1962
rect 15446 1912 15462 1946
rect 15630 1912 15646 1946
rect 15446 1874 15646 1912
rect 15704 1946 15904 1962
rect 15704 1912 15720 1946
rect 15888 1912 15904 1946
rect 15704 1874 15904 1912
rect 14672 1436 14872 1474
rect 14672 1402 14688 1436
rect 14856 1402 14872 1436
rect 14672 1386 14872 1402
rect 14930 1436 15130 1474
rect 14930 1402 14946 1436
rect 15114 1402 15130 1436
rect 14930 1386 15130 1402
rect 15188 1436 15388 1474
rect 15188 1402 15204 1436
rect 15372 1402 15388 1436
rect 15188 1386 15388 1402
rect 15446 1436 15646 1474
rect 15446 1402 15462 1436
rect 15630 1402 15646 1436
rect 15446 1386 15646 1402
rect 15704 1436 15904 1474
rect 15704 1402 15720 1436
rect 15888 1402 15904 1436
rect 15704 1386 15904 1402
rect 14672 1328 14872 1344
rect 14672 1294 14688 1328
rect 14856 1294 14872 1328
rect 14672 1256 14872 1294
rect 14930 1328 15130 1344
rect 14930 1294 14946 1328
rect 15114 1294 15130 1328
rect 14930 1256 15130 1294
rect 15188 1328 15388 1344
rect 15188 1294 15204 1328
rect 15372 1294 15388 1328
rect 15188 1256 15388 1294
rect 15446 1328 15646 1344
rect 15446 1294 15462 1328
rect 15630 1294 15646 1328
rect 15446 1256 15646 1294
rect 15704 1328 15904 1344
rect 15704 1294 15720 1328
rect 15888 1294 15904 1328
rect 15704 1256 15904 1294
rect 14672 818 14872 856
rect 14672 784 14688 818
rect 14856 784 14872 818
rect 14672 768 14872 784
rect 14930 818 15130 856
rect 14930 784 14946 818
rect 15114 784 15130 818
rect 14930 768 15130 784
rect 15188 818 15388 856
rect 15188 784 15204 818
rect 15372 784 15388 818
rect 15188 768 15388 784
rect 15446 818 15646 856
rect 15446 784 15462 818
rect 15630 784 15646 818
rect 15446 768 15646 784
rect 15704 818 15904 856
rect 15704 784 15720 818
rect 15888 784 15904 818
rect 15704 768 15904 784
rect 14672 710 14872 726
rect 14672 676 14688 710
rect 14856 676 14872 710
rect 14672 638 14872 676
rect 14930 710 15130 726
rect 14930 676 14946 710
rect 15114 676 15130 710
rect 14930 638 15130 676
rect 15188 710 15388 726
rect 15188 676 15204 710
rect 15372 676 15388 710
rect 15188 638 15388 676
rect 15446 710 15646 726
rect 15446 676 15462 710
rect 15630 676 15646 710
rect 15446 638 15646 676
rect 15704 710 15904 726
rect 15704 676 15720 710
rect 15888 676 15904 710
rect 15704 638 15904 676
rect 14672 200 14872 238
rect 14672 166 14688 200
rect 14856 166 14872 200
rect 14672 150 14872 166
rect 14930 200 15130 238
rect 14930 166 14946 200
rect 15114 166 15130 200
rect 14930 150 15130 166
rect 15188 200 15388 238
rect 15188 166 15204 200
rect 15372 166 15388 200
rect 15188 150 15388 166
rect 15446 200 15646 238
rect 15446 166 15462 200
rect 15630 166 15646 200
rect 15446 150 15646 166
rect 15704 200 15904 238
rect 15704 166 15720 200
rect 15888 166 15904 200
rect 15704 150 15904 166
rect 16472 3800 16672 3816
rect 16472 3766 16488 3800
rect 16656 3766 16672 3800
rect 16472 3728 16672 3766
rect 16730 3800 16930 3816
rect 16730 3766 16746 3800
rect 16914 3766 16930 3800
rect 16730 3728 16930 3766
rect 16988 3800 17188 3816
rect 16988 3766 17004 3800
rect 17172 3766 17188 3800
rect 16988 3728 17188 3766
rect 17246 3800 17446 3816
rect 17246 3766 17262 3800
rect 17430 3766 17446 3800
rect 17246 3728 17446 3766
rect 17504 3800 17704 3816
rect 17504 3766 17520 3800
rect 17688 3766 17704 3800
rect 17504 3728 17704 3766
rect 16472 3290 16672 3328
rect 16472 3256 16488 3290
rect 16656 3256 16672 3290
rect 16472 3240 16672 3256
rect 16730 3290 16930 3328
rect 16730 3256 16746 3290
rect 16914 3256 16930 3290
rect 16730 3240 16930 3256
rect 16988 3290 17188 3328
rect 16988 3256 17004 3290
rect 17172 3256 17188 3290
rect 16988 3240 17188 3256
rect 17246 3290 17446 3328
rect 17246 3256 17262 3290
rect 17430 3256 17446 3290
rect 17246 3240 17446 3256
rect 17504 3290 17704 3328
rect 17504 3256 17520 3290
rect 17688 3256 17704 3290
rect 17504 3240 17704 3256
rect 16472 3182 16672 3198
rect 16472 3148 16488 3182
rect 16656 3148 16672 3182
rect 16472 3110 16672 3148
rect 16730 3182 16930 3198
rect 16730 3148 16746 3182
rect 16914 3148 16930 3182
rect 16730 3110 16930 3148
rect 16988 3182 17188 3198
rect 16988 3148 17004 3182
rect 17172 3148 17188 3182
rect 16988 3110 17188 3148
rect 17246 3182 17446 3198
rect 17246 3148 17262 3182
rect 17430 3148 17446 3182
rect 17246 3110 17446 3148
rect 17504 3182 17704 3198
rect 17504 3148 17520 3182
rect 17688 3148 17704 3182
rect 17504 3110 17704 3148
rect 16472 2672 16672 2710
rect 16472 2638 16488 2672
rect 16656 2638 16672 2672
rect 16472 2622 16672 2638
rect 16730 2672 16930 2710
rect 16730 2638 16746 2672
rect 16914 2638 16930 2672
rect 16730 2622 16930 2638
rect 16988 2672 17188 2710
rect 16988 2638 17004 2672
rect 17172 2638 17188 2672
rect 16988 2622 17188 2638
rect 17246 2672 17446 2710
rect 17246 2638 17262 2672
rect 17430 2638 17446 2672
rect 17246 2622 17446 2638
rect 17504 2672 17704 2710
rect 17504 2638 17520 2672
rect 17688 2638 17704 2672
rect 17504 2622 17704 2638
rect 16472 2564 16672 2580
rect 16472 2530 16488 2564
rect 16656 2530 16672 2564
rect 16472 2492 16672 2530
rect 16730 2564 16930 2580
rect 16730 2530 16746 2564
rect 16914 2530 16930 2564
rect 16730 2492 16930 2530
rect 16988 2564 17188 2580
rect 16988 2530 17004 2564
rect 17172 2530 17188 2564
rect 16988 2492 17188 2530
rect 17246 2564 17446 2580
rect 17246 2530 17262 2564
rect 17430 2530 17446 2564
rect 17246 2492 17446 2530
rect 17504 2564 17704 2580
rect 17504 2530 17520 2564
rect 17688 2530 17704 2564
rect 17504 2492 17704 2530
rect 16472 2054 16672 2092
rect 16472 2020 16488 2054
rect 16656 2020 16672 2054
rect 16472 2004 16672 2020
rect 16730 2054 16930 2092
rect 16730 2020 16746 2054
rect 16914 2020 16930 2054
rect 16730 2004 16930 2020
rect 16988 2054 17188 2092
rect 16988 2020 17004 2054
rect 17172 2020 17188 2054
rect 16988 2004 17188 2020
rect 17246 2054 17446 2092
rect 17246 2020 17262 2054
rect 17430 2020 17446 2054
rect 17246 2004 17446 2020
rect 17504 2054 17704 2092
rect 17504 2020 17520 2054
rect 17688 2020 17704 2054
rect 17504 2004 17704 2020
rect 16472 1946 16672 1962
rect 16472 1912 16488 1946
rect 16656 1912 16672 1946
rect 16472 1874 16672 1912
rect 16730 1946 16930 1962
rect 16730 1912 16746 1946
rect 16914 1912 16930 1946
rect 16730 1874 16930 1912
rect 16988 1946 17188 1962
rect 16988 1912 17004 1946
rect 17172 1912 17188 1946
rect 16988 1874 17188 1912
rect 17246 1946 17446 1962
rect 17246 1912 17262 1946
rect 17430 1912 17446 1946
rect 17246 1874 17446 1912
rect 17504 1946 17704 1962
rect 17504 1912 17520 1946
rect 17688 1912 17704 1946
rect 17504 1874 17704 1912
rect 16472 1436 16672 1474
rect 16472 1402 16488 1436
rect 16656 1402 16672 1436
rect 16472 1386 16672 1402
rect 16730 1436 16930 1474
rect 16730 1402 16746 1436
rect 16914 1402 16930 1436
rect 16730 1386 16930 1402
rect 16988 1436 17188 1474
rect 16988 1402 17004 1436
rect 17172 1402 17188 1436
rect 16988 1386 17188 1402
rect 17246 1436 17446 1474
rect 17246 1402 17262 1436
rect 17430 1402 17446 1436
rect 17246 1386 17446 1402
rect 17504 1436 17704 1474
rect 17504 1402 17520 1436
rect 17688 1402 17704 1436
rect 17504 1386 17704 1402
rect 16472 1328 16672 1344
rect 16472 1294 16488 1328
rect 16656 1294 16672 1328
rect 16472 1256 16672 1294
rect 16730 1328 16930 1344
rect 16730 1294 16746 1328
rect 16914 1294 16930 1328
rect 16730 1256 16930 1294
rect 16988 1328 17188 1344
rect 16988 1294 17004 1328
rect 17172 1294 17188 1328
rect 16988 1256 17188 1294
rect 17246 1328 17446 1344
rect 17246 1294 17262 1328
rect 17430 1294 17446 1328
rect 17246 1256 17446 1294
rect 17504 1328 17704 1344
rect 17504 1294 17520 1328
rect 17688 1294 17704 1328
rect 17504 1256 17704 1294
rect 16472 818 16672 856
rect 16472 784 16488 818
rect 16656 784 16672 818
rect 16472 768 16672 784
rect 16730 818 16930 856
rect 16730 784 16746 818
rect 16914 784 16930 818
rect 16730 768 16930 784
rect 16988 818 17188 856
rect 16988 784 17004 818
rect 17172 784 17188 818
rect 16988 768 17188 784
rect 17246 818 17446 856
rect 17246 784 17262 818
rect 17430 784 17446 818
rect 17246 768 17446 784
rect 17504 818 17704 856
rect 17504 784 17520 818
rect 17688 784 17704 818
rect 17504 768 17704 784
rect 16472 710 16672 726
rect 16472 676 16488 710
rect 16656 676 16672 710
rect 16472 638 16672 676
rect 16730 710 16930 726
rect 16730 676 16746 710
rect 16914 676 16930 710
rect 16730 638 16930 676
rect 16988 710 17188 726
rect 16988 676 17004 710
rect 17172 676 17188 710
rect 16988 638 17188 676
rect 17246 710 17446 726
rect 17246 676 17262 710
rect 17430 676 17446 710
rect 17246 638 17446 676
rect 17504 710 17704 726
rect 17504 676 17520 710
rect 17688 676 17704 710
rect 17504 638 17704 676
rect 16472 200 16672 238
rect 16472 166 16488 200
rect 16656 166 16672 200
rect 16472 150 16672 166
rect 16730 200 16930 238
rect 16730 166 16746 200
rect 16914 166 16930 200
rect 16730 150 16930 166
rect 16988 200 17188 238
rect 16988 166 17004 200
rect 17172 166 17188 200
rect 16988 150 17188 166
rect 17246 200 17446 238
rect 17246 166 17262 200
rect 17430 166 17446 200
rect 17246 150 17446 166
rect 17504 200 17704 238
rect 17504 166 17520 200
rect 17688 166 17704 200
rect 17504 150 17704 166
rect 18272 3800 18472 3816
rect 18272 3766 18288 3800
rect 18456 3766 18472 3800
rect 18272 3728 18472 3766
rect 18530 3800 18730 3816
rect 18530 3766 18546 3800
rect 18714 3766 18730 3800
rect 18530 3728 18730 3766
rect 18788 3800 18988 3816
rect 18788 3766 18804 3800
rect 18972 3766 18988 3800
rect 18788 3728 18988 3766
rect 19046 3800 19246 3816
rect 19046 3766 19062 3800
rect 19230 3766 19246 3800
rect 19046 3728 19246 3766
rect 19304 3800 19504 3816
rect 19304 3766 19320 3800
rect 19488 3766 19504 3800
rect 19304 3728 19504 3766
rect 18272 3290 18472 3328
rect 18272 3256 18288 3290
rect 18456 3256 18472 3290
rect 18272 3240 18472 3256
rect 18530 3290 18730 3328
rect 18530 3256 18546 3290
rect 18714 3256 18730 3290
rect 18530 3240 18730 3256
rect 18788 3290 18988 3328
rect 18788 3256 18804 3290
rect 18972 3256 18988 3290
rect 18788 3240 18988 3256
rect 19046 3290 19246 3328
rect 19046 3256 19062 3290
rect 19230 3256 19246 3290
rect 19046 3240 19246 3256
rect 19304 3290 19504 3328
rect 19304 3256 19320 3290
rect 19488 3256 19504 3290
rect 19304 3240 19504 3256
rect 18272 3182 18472 3198
rect 18272 3148 18288 3182
rect 18456 3148 18472 3182
rect 18272 3110 18472 3148
rect 18530 3182 18730 3198
rect 18530 3148 18546 3182
rect 18714 3148 18730 3182
rect 18530 3110 18730 3148
rect 18788 3182 18988 3198
rect 18788 3148 18804 3182
rect 18972 3148 18988 3182
rect 18788 3110 18988 3148
rect 19046 3182 19246 3198
rect 19046 3148 19062 3182
rect 19230 3148 19246 3182
rect 19046 3110 19246 3148
rect 19304 3182 19504 3198
rect 19304 3148 19320 3182
rect 19488 3148 19504 3182
rect 19304 3110 19504 3148
rect 18272 2672 18472 2710
rect 18272 2638 18288 2672
rect 18456 2638 18472 2672
rect 18272 2622 18472 2638
rect 18530 2672 18730 2710
rect 18530 2638 18546 2672
rect 18714 2638 18730 2672
rect 18530 2622 18730 2638
rect 18788 2672 18988 2710
rect 18788 2638 18804 2672
rect 18972 2638 18988 2672
rect 18788 2622 18988 2638
rect 19046 2672 19246 2710
rect 19046 2638 19062 2672
rect 19230 2638 19246 2672
rect 19046 2622 19246 2638
rect 19304 2672 19504 2710
rect 19304 2638 19320 2672
rect 19488 2638 19504 2672
rect 19304 2622 19504 2638
rect 18272 2564 18472 2580
rect 18272 2530 18288 2564
rect 18456 2530 18472 2564
rect 18272 2492 18472 2530
rect 18530 2564 18730 2580
rect 18530 2530 18546 2564
rect 18714 2530 18730 2564
rect 18530 2492 18730 2530
rect 18788 2564 18988 2580
rect 18788 2530 18804 2564
rect 18972 2530 18988 2564
rect 18788 2492 18988 2530
rect 19046 2564 19246 2580
rect 19046 2530 19062 2564
rect 19230 2530 19246 2564
rect 19046 2492 19246 2530
rect 19304 2564 19504 2580
rect 19304 2530 19320 2564
rect 19488 2530 19504 2564
rect 19304 2492 19504 2530
rect 18272 2054 18472 2092
rect 18272 2020 18288 2054
rect 18456 2020 18472 2054
rect 18272 2004 18472 2020
rect 18530 2054 18730 2092
rect 18530 2020 18546 2054
rect 18714 2020 18730 2054
rect 18530 2004 18730 2020
rect 18788 2054 18988 2092
rect 18788 2020 18804 2054
rect 18972 2020 18988 2054
rect 18788 2004 18988 2020
rect 19046 2054 19246 2092
rect 19046 2020 19062 2054
rect 19230 2020 19246 2054
rect 19046 2004 19246 2020
rect 19304 2054 19504 2092
rect 19304 2020 19320 2054
rect 19488 2020 19504 2054
rect 19304 2004 19504 2020
rect 18272 1946 18472 1962
rect 18272 1912 18288 1946
rect 18456 1912 18472 1946
rect 18272 1874 18472 1912
rect 18530 1946 18730 1962
rect 18530 1912 18546 1946
rect 18714 1912 18730 1946
rect 18530 1874 18730 1912
rect 18788 1946 18988 1962
rect 18788 1912 18804 1946
rect 18972 1912 18988 1946
rect 18788 1874 18988 1912
rect 19046 1946 19246 1962
rect 19046 1912 19062 1946
rect 19230 1912 19246 1946
rect 19046 1874 19246 1912
rect 19304 1946 19504 1962
rect 19304 1912 19320 1946
rect 19488 1912 19504 1946
rect 19304 1874 19504 1912
rect 18272 1436 18472 1474
rect 18272 1402 18288 1436
rect 18456 1402 18472 1436
rect 18272 1386 18472 1402
rect 18530 1436 18730 1474
rect 18530 1402 18546 1436
rect 18714 1402 18730 1436
rect 18530 1386 18730 1402
rect 18788 1436 18988 1474
rect 18788 1402 18804 1436
rect 18972 1402 18988 1436
rect 18788 1386 18988 1402
rect 19046 1436 19246 1474
rect 19046 1402 19062 1436
rect 19230 1402 19246 1436
rect 19046 1386 19246 1402
rect 19304 1436 19504 1474
rect 19304 1402 19320 1436
rect 19488 1402 19504 1436
rect 19304 1386 19504 1402
rect 18272 1328 18472 1344
rect 18272 1294 18288 1328
rect 18456 1294 18472 1328
rect 18272 1256 18472 1294
rect 18530 1328 18730 1344
rect 18530 1294 18546 1328
rect 18714 1294 18730 1328
rect 18530 1256 18730 1294
rect 18788 1328 18988 1344
rect 18788 1294 18804 1328
rect 18972 1294 18988 1328
rect 18788 1256 18988 1294
rect 19046 1328 19246 1344
rect 19046 1294 19062 1328
rect 19230 1294 19246 1328
rect 19046 1256 19246 1294
rect 19304 1328 19504 1344
rect 19304 1294 19320 1328
rect 19488 1294 19504 1328
rect 19304 1256 19504 1294
rect 18272 818 18472 856
rect 18272 784 18288 818
rect 18456 784 18472 818
rect 18272 768 18472 784
rect 18530 818 18730 856
rect 18530 784 18546 818
rect 18714 784 18730 818
rect 18530 768 18730 784
rect 18788 818 18988 856
rect 18788 784 18804 818
rect 18972 784 18988 818
rect 18788 768 18988 784
rect 19046 818 19246 856
rect 19046 784 19062 818
rect 19230 784 19246 818
rect 19046 768 19246 784
rect 19304 818 19504 856
rect 19304 784 19320 818
rect 19488 784 19504 818
rect 19304 768 19504 784
rect 18272 710 18472 726
rect 18272 676 18288 710
rect 18456 676 18472 710
rect 18272 638 18472 676
rect 18530 710 18730 726
rect 18530 676 18546 710
rect 18714 676 18730 710
rect 18530 638 18730 676
rect 18788 710 18988 726
rect 18788 676 18804 710
rect 18972 676 18988 710
rect 18788 638 18988 676
rect 19046 710 19246 726
rect 19046 676 19062 710
rect 19230 676 19246 710
rect 19046 638 19246 676
rect 19304 710 19504 726
rect 19304 676 19320 710
rect 19488 676 19504 710
rect 19304 638 19504 676
rect 18272 200 18472 238
rect 18272 166 18288 200
rect 18456 166 18472 200
rect 18272 150 18472 166
rect 18530 200 18730 238
rect 18530 166 18546 200
rect 18714 166 18730 200
rect 18530 150 18730 166
rect 18788 200 18988 238
rect 18788 166 18804 200
rect 18972 166 18988 200
rect 18788 150 18988 166
rect 19046 200 19246 238
rect 19046 166 19062 200
rect 19230 166 19246 200
rect 19046 150 19246 166
rect 19304 200 19504 238
rect 19304 166 19320 200
rect 19488 166 19504 200
rect 19304 150 19504 166
rect 20072 3800 20272 3816
rect 20072 3766 20088 3800
rect 20256 3766 20272 3800
rect 20072 3728 20272 3766
rect 20330 3800 20530 3816
rect 20330 3766 20346 3800
rect 20514 3766 20530 3800
rect 20330 3728 20530 3766
rect 20588 3800 20788 3816
rect 20588 3766 20604 3800
rect 20772 3766 20788 3800
rect 20588 3728 20788 3766
rect 20846 3800 21046 3816
rect 20846 3766 20862 3800
rect 21030 3766 21046 3800
rect 20846 3728 21046 3766
rect 21104 3800 21304 3816
rect 21104 3766 21120 3800
rect 21288 3766 21304 3800
rect 21104 3728 21304 3766
rect 20072 3290 20272 3328
rect 20072 3256 20088 3290
rect 20256 3256 20272 3290
rect 20072 3240 20272 3256
rect 20330 3290 20530 3328
rect 20330 3256 20346 3290
rect 20514 3256 20530 3290
rect 20330 3240 20530 3256
rect 20588 3290 20788 3328
rect 20588 3256 20604 3290
rect 20772 3256 20788 3290
rect 20588 3240 20788 3256
rect 20846 3290 21046 3328
rect 20846 3256 20862 3290
rect 21030 3256 21046 3290
rect 20846 3240 21046 3256
rect 21104 3290 21304 3328
rect 21104 3256 21120 3290
rect 21288 3256 21304 3290
rect 21104 3240 21304 3256
rect 20072 3182 20272 3198
rect 20072 3148 20088 3182
rect 20256 3148 20272 3182
rect 20072 3110 20272 3148
rect 20330 3182 20530 3198
rect 20330 3148 20346 3182
rect 20514 3148 20530 3182
rect 20330 3110 20530 3148
rect 20588 3182 20788 3198
rect 20588 3148 20604 3182
rect 20772 3148 20788 3182
rect 20588 3110 20788 3148
rect 20846 3182 21046 3198
rect 20846 3148 20862 3182
rect 21030 3148 21046 3182
rect 20846 3110 21046 3148
rect 21104 3182 21304 3198
rect 21104 3148 21120 3182
rect 21288 3148 21304 3182
rect 21104 3110 21304 3148
rect 20072 2672 20272 2710
rect 20072 2638 20088 2672
rect 20256 2638 20272 2672
rect 20072 2622 20272 2638
rect 20330 2672 20530 2710
rect 20330 2638 20346 2672
rect 20514 2638 20530 2672
rect 20330 2622 20530 2638
rect 20588 2672 20788 2710
rect 20588 2638 20604 2672
rect 20772 2638 20788 2672
rect 20588 2622 20788 2638
rect 20846 2672 21046 2710
rect 20846 2638 20862 2672
rect 21030 2638 21046 2672
rect 20846 2622 21046 2638
rect 21104 2672 21304 2710
rect 21104 2638 21120 2672
rect 21288 2638 21304 2672
rect 21104 2622 21304 2638
rect 20072 2564 20272 2580
rect 20072 2530 20088 2564
rect 20256 2530 20272 2564
rect 20072 2492 20272 2530
rect 20330 2564 20530 2580
rect 20330 2530 20346 2564
rect 20514 2530 20530 2564
rect 20330 2492 20530 2530
rect 20588 2564 20788 2580
rect 20588 2530 20604 2564
rect 20772 2530 20788 2564
rect 20588 2492 20788 2530
rect 20846 2564 21046 2580
rect 20846 2530 20862 2564
rect 21030 2530 21046 2564
rect 20846 2492 21046 2530
rect 21104 2564 21304 2580
rect 21104 2530 21120 2564
rect 21288 2530 21304 2564
rect 21104 2492 21304 2530
rect 20072 2054 20272 2092
rect 20072 2020 20088 2054
rect 20256 2020 20272 2054
rect 20072 2004 20272 2020
rect 20330 2054 20530 2092
rect 20330 2020 20346 2054
rect 20514 2020 20530 2054
rect 20330 2004 20530 2020
rect 20588 2054 20788 2092
rect 20588 2020 20604 2054
rect 20772 2020 20788 2054
rect 20588 2004 20788 2020
rect 20846 2054 21046 2092
rect 20846 2020 20862 2054
rect 21030 2020 21046 2054
rect 20846 2004 21046 2020
rect 21104 2054 21304 2092
rect 21104 2020 21120 2054
rect 21288 2020 21304 2054
rect 21104 2004 21304 2020
rect 20072 1946 20272 1962
rect 20072 1912 20088 1946
rect 20256 1912 20272 1946
rect 20072 1874 20272 1912
rect 20330 1946 20530 1962
rect 20330 1912 20346 1946
rect 20514 1912 20530 1946
rect 20330 1874 20530 1912
rect 20588 1946 20788 1962
rect 20588 1912 20604 1946
rect 20772 1912 20788 1946
rect 20588 1874 20788 1912
rect 20846 1946 21046 1962
rect 20846 1912 20862 1946
rect 21030 1912 21046 1946
rect 20846 1874 21046 1912
rect 21104 1946 21304 1962
rect 21104 1912 21120 1946
rect 21288 1912 21304 1946
rect 21104 1874 21304 1912
rect 20072 1436 20272 1474
rect 20072 1402 20088 1436
rect 20256 1402 20272 1436
rect 20072 1386 20272 1402
rect 20330 1436 20530 1474
rect 20330 1402 20346 1436
rect 20514 1402 20530 1436
rect 20330 1386 20530 1402
rect 20588 1436 20788 1474
rect 20588 1402 20604 1436
rect 20772 1402 20788 1436
rect 20588 1386 20788 1402
rect 20846 1436 21046 1474
rect 20846 1402 20862 1436
rect 21030 1402 21046 1436
rect 20846 1386 21046 1402
rect 21104 1436 21304 1474
rect 21104 1402 21120 1436
rect 21288 1402 21304 1436
rect 21104 1386 21304 1402
rect 20072 1328 20272 1344
rect 20072 1294 20088 1328
rect 20256 1294 20272 1328
rect 20072 1256 20272 1294
rect 20330 1328 20530 1344
rect 20330 1294 20346 1328
rect 20514 1294 20530 1328
rect 20330 1256 20530 1294
rect 20588 1328 20788 1344
rect 20588 1294 20604 1328
rect 20772 1294 20788 1328
rect 20588 1256 20788 1294
rect 20846 1328 21046 1344
rect 20846 1294 20862 1328
rect 21030 1294 21046 1328
rect 20846 1256 21046 1294
rect 21104 1328 21304 1344
rect 21104 1294 21120 1328
rect 21288 1294 21304 1328
rect 21104 1256 21304 1294
rect 20072 818 20272 856
rect 20072 784 20088 818
rect 20256 784 20272 818
rect 20072 768 20272 784
rect 20330 818 20530 856
rect 20330 784 20346 818
rect 20514 784 20530 818
rect 20330 768 20530 784
rect 20588 818 20788 856
rect 20588 784 20604 818
rect 20772 784 20788 818
rect 20588 768 20788 784
rect 20846 818 21046 856
rect 20846 784 20862 818
rect 21030 784 21046 818
rect 20846 768 21046 784
rect 21104 818 21304 856
rect 21104 784 21120 818
rect 21288 784 21304 818
rect 21104 768 21304 784
rect 20072 710 20272 726
rect 20072 676 20088 710
rect 20256 676 20272 710
rect 20072 638 20272 676
rect 20330 710 20530 726
rect 20330 676 20346 710
rect 20514 676 20530 710
rect 20330 638 20530 676
rect 20588 710 20788 726
rect 20588 676 20604 710
rect 20772 676 20788 710
rect 20588 638 20788 676
rect 20846 710 21046 726
rect 20846 676 20862 710
rect 21030 676 21046 710
rect 20846 638 21046 676
rect 21104 710 21304 726
rect 21104 676 21120 710
rect 21288 676 21304 710
rect 21104 638 21304 676
rect 20072 200 20272 238
rect 20072 166 20088 200
rect 20256 166 20272 200
rect 20072 150 20272 166
rect 20330 200 20530 238
rect 20330 166 20346 200
rect 20514 166 20530 200
rect 20330 150 20530 166
rect 20588 200 20788 238
rect 20588 166 20604 200
rect 20772 166 20788 200
rect 20588 150 20788 166
rect 20846 200 21046 238
rect 20846 166 20862 200
rect 21030 166 21046 200
rect 20846 150 21046 166
rect 21104 200 21304 238
rect 21104 166 21120 200
rect 21288 166 21304 200
rect 21104 150 21304 166
<< polycont >>
rect 6552 27134 6620 27168
rect 6710 27134 6778 27168
rect 6868 27134 6936 27168
rect 7026 27134 7094 27168
rect 7184 27134 7252 27168
rect 7342 27134 7410 27168
rect 7500 27134 7568 27168
rect 7658 27134 7726 27168
rect 7816 27134 7884 27168
rect 7974 27134 8042 27168
rect 6552 26606 6620 26640
rect 6710 26606 6778 26640
rect 6868 26606 6936 26640
rect 7026 26606 7094 26640
rect 7184 26606 7252 26640
rect 7342 26606 7410 26640
rect 7500 26606 7568 26640
rect 7658 26606 7726 26640
rect 7816 26606 7884 26640
rect 7974 26606 8042 26640
rect 6552 26498 6620 26532
rect 6710 26498 6778 26532
rect 6868 26498 6936 26532
rect 7026 26498 7094 26532
rect 7184 26498 7252 26532
rect 7342 26498 7410 26532
rect 7500 26498 7568 26532
rect 7658 26498 7726 26532
rect 7816 26498 7884 26532
rect 7974 26498 8042 26532
rect 6552 25970 6620 26004
rect 6710 25970 6778 26004
rect 6868 25970 6936 26004
rect 7026 25970 7094 26004
rect 7184 25970 7252 26004
rect 7342 25970 7410 26004
rect 7500 25970 7568 26004
rect 7658 25970 7726 26004
rect 7816 25970 7884 26004
rect 7974 25970 8042 26004
rect 6552 25862 6620 25896
rect 6710 25862 6778 25896
rect 6868 25862 6936 25896
rect 7026 25862 7094 25896
rect 7184 25862 7252 25896
rect 7342 25862 7410 25896
rect 7500 25862 7568 25896
rect 7658 25862 7726 25896
rect 7816 25862 7884 25896
rect 7974 25862 8042 25896
rect 6552 25334 6620 25368
rect 6710 25334 6778 25368
rect 6868 25334 6936 25368
rect 7026 25334 7094 25368
rect 7184 25334 7252 25368
rect 7342 25334 7410 25368
rect 7500 25334 7568 25368
rect 7658 25334 7726 25368
rect 7816 25334 7884 25368
rect 7974 25334 8042 25368
rect 8772 27134 8840 27168
rect 8930 27134 8998 27168
rect 9088 27134 9156 27168
rect 9246 27134 9314 27168
rect 9404 27134 9472 27168
rect 9562 27134 9630 27168
rect 9720 27134 9788 27168
rect 9878 27134 9946 27168
rect 10036 27134 10104 27168
rect 10194 27134 10262 27168
rect 8772 26606 8840 26640
rect 8930 26606 8998 26640
rect 9088 26606 9156 26640
rect 9246 26606 9314 26640
rect 9404 26606 9472 26640
rect 9562 26606 9630 26640
rect 9720 26606 9788 26640
rect 9878 26606 9946 26640
rect 10036 26606 10104 26640
rect 10194 26606 10262 26640
rect 8772 26498 8840 26532
rect 8930 26498 8998 26532
rect 9088 26498 9156 26532
rect 9246 26498 9314 26532
rect 9404 26498 9472 26532
rect 9562 26498 9630 26532
rect 9720 26498 9788 26532
rect 9878 26498 9946 26532
rect 10036 26498 10104 26532
rect 10194 26498 10262 26532
rect 8772 25970 8840 26004
rect 8930 25970 8998 26004
rect 9088 25970 9156 26004
rect 9246 25970 9314 26004
rect 9404 25970 9472 26004
rect 9562 25970 9630 26004
rect 9720 25970 9788 26004
rect 9878 25970 9946 26004
rect 10036 25970 10104 26004
rect 10194 25970 10262 26004
rect 8772 25862 8840 25896
rect 8930 25862 8998 25896
rect 9088 25862 9156 25896
rect 9246 25862 9314 25896
rect 9404 25862 9472 25896
rect 9562 25862 9630 25896
rect 9720 25862 9788 25896
rect 9878 25862 9946 25896
rect 10036 25862 10104 25896
rect 10194 25862 10262 25896
rect 8772 25334 8840 25368
rect 8930 25334 8998 25368
rect 9088 25334 9156 25368
rect 9246 25334 9314 25368
rect 9404 25334 9472 25368
rect 9562 25334 9630 25368
rect 9720 25334 9788 25368
rect 9878 25334 9946 25368
rect 10036 25334 10104 25368
rect 10194 25334 10262 25368
rect 10952 27134 11020 27168
rect 11110 27134 11178 27168
rect 11268 27134 11336 27168
rect 11426 27134 11494 27168
rect 11584 27134 11652 27168
rect 11742 27134 11810 27168
rect 11900 27134 11968 27168
rect 12058 27134 12126 27168
rect 12216 27134 12284 27168
rect 12374 27134 12442 27168
rect 10952 26606 11020 26640
rect 11110 26606 11178 26640
rect 11268 26606 11336 26640
rect 11426 26606 11494 26640
rect 11584 26606 11652 26640
rect 11742 26606 11810 26640
rect 11900 26606 11968 26640
rect 12058 26606 12126 26640
rect 12216 26606 12284 26640
rect 12374 26606 12442 26640
rect 10952 26498 11020 26532
rect 11110 26498 11178 26532
rect 11268 26498 11336 26532
rect 11426 26498 11494 26532
rect 11584 26498 11652 26532
rect 11742 26498 11810 26532
rect 11900 26498 11968 26532
rect 12058 26498 12126 26532
rect 12216 26498 12284 26532
rect 12374 26498 12442 26532
rect 10952 25970 11020 26004
rect 11110 25970 11178 26004
rect 11268 25970 11336 26004
rect 11426 25970 11494 26004
rect 11584 25970 11652 26004
rect 11742 25970 11810 26004
rect 11900 25970 11968 26004
rect 12058 25970 12126 26004
rect 12216 25970 12284 26004
rect 12374 25970 12442 26004
rect 10952 25862 11020 25896
rect 11110 25862 11178 25896
rect 11268 25862 11336 25896
rect 11426 25862 11494 25896
rect 11584 25862 11652 25896
rect 11742 25862 11810 25896
rect 11900 25862 11968 25896
rect 12058 25862 12126 25896
rect 12216 25862 12284 25896
rect 12374 25862 12442 25896
rect 10952 25334 11020 25368
rect 11110 25334 11178 25368
rect 11268 25334 11336 25368
rect 11426 25334 11494 25368
rect 11584 25334 11652 25368
rect 11742 25334 11810 25368
rect 11900 25334 11968 25368
rect 12058 25334 12126 25368
rect 12216 25334 12284 25368
rect 12374 25334 12442 25368
rect 13132 27134 13200 27168
rect 13290 27134 13358 27168
rect 13448 27134 13516 27168
rect 13606 27134 13674 27168
rect 13764 27134 13832 27168
rect 13922 27134 13990 27168
rect 14080 27134 14148 27168
rect 14238 27134 14306 27168
rect 14396 27134 14464 27168
rect 14554 27134 14622 27168
rect 13132 26606 13200 26640
rect 13290 26606 13358 26640
rect 13448 26606 13516 26640
rect 13606 26606 13674 26640
rect 13764 26606 13832 26640
rect 13922 26606 13990 26640
rect 14080 26606 14148 26640
rect 14238 26606 14306 26640
rect 14396 26606 14464 26640
rect 14554 26606 14622 26640
rect 13132 26498 13200 26532
rect 13290 26498 13358 26532
rect 13448 26498 13516 26532
rect 13606 26498 13674 26532
rect 13764 26498 13832 26532
rect 13922 26498 13990 26532
rect 14080 26498 14148 26532
rect 14238 26498 14306 26532
rect 14396 26498 14464 26532
rect 14554 26498 14622 26532
rect 13132 25970 13200 26004
rect 13290 25970 13358 26004
rect 13448 25970 13516 26004
rect 13606 25970 13674 26004
rect 13764 25970 13832 26004
rect 13922 25970 13990 26004
rect 14080 25970 14148 26004
rect 14238 25970 14306 26004
rect 14396 25970 14464 26004
rect 14554 25970 14622 26004
rect 13132 25862 13200 25896
rect 13290 25862 13358 25896
rect 13448 25862 13516 25896
rect 13606 25862 13674 25896
rect 13764 25862 13832 25896
rect 13922 25862 13990 25896
rect 14080 25862 14148 25896
rect 14238 25862 14306 25896
rect 14396 25862 14464 25896
rect 14554 25862 14622 25896
rect 13132 25334 13200 25368
rect 13290 25334 13358 25368
rect 13448 25334 13516 25368
rect 13606 25334 13674 25368
rect 13764 25334 13832 25368
rect 13922 25334 13990 25368
rect 14080 25334 14148 25368
rect 14238 25334 14306 25368
rect 14396 25334 14464 25368
rect 14554 25334 14622 25368
rect 15332 27134 15400 27168
rect 15490 27134 15558 27168
rect 15648 27134 15716 27168
rect 15806 27134 15874 27168
rect 15964 27134 16032 27168
rect 16122 27134 16190 27168
rect 16280 27134 16348 27168
rect 16438 27134 16506 27168
rect 16596 27134 16664 27168
rect 16754 27134 16822 27168
rect 15332 26606 15400 26640
rect 15490 26606 15558 26640
rect 15648 26606 15716 26640
rect 15806 26606 15874 26640
rect 15964 26606 16032 26640
rect 16122 26606 16190 26640
rect 16280 26606 16348 26640
rect 16438 26606 16506 26640
rect 16596 26606 16664 26640
rect 16754 26606 16822 26640
rect 15332 26498 15400 26532
rect 15490 26498 15558 26532
rect 15648 26498 15716 26532
rect 15806 26498 15874 26532
rect 15964 26498 16032 26532
rect 16122 26498 16190 26532
rect 16280 26498 16348 26532
rect 16438 26498 16506 26532
rect 16596 26498 16664 26532
rect 16754 26498 16822 26532
rect 15332 25970 15400 26004
rect 15490 25970 15558 26004
rect 15648 25970 15716 26004
rect 15806 25970 15874 26004
rect 15964 25970 16032 26004
rect 16122 25970 16190 26004
rect 16280 25970 16348 26004
rect 16438 25970 16506 26004
rect 16596 25970 16664 26004
rect 16754 25970 16822 26004
rect 15332 25862 15400 25896
rect 15490 25862 15558 25896
rect 15648 25862 15716 25896
rect 15806 25862 15874 25896
rect 15964 25862 16032 25896
rect 16122 25862 16190 25896
rect 16280 25862 16348 25896
rect 16438 25862 16506 25896
rect 16596 25862 16664 25896
rect 16754 25862 16822 25896
rect 15332 25334 15400 25368
rect 15490 25334 15558 25368
rect 15648 25334 15716 25368
rect 15806 25334 15874 25368
rect 15964 25334 16032 25368
rect 16122 25334 16190 25368
rect 16280 25334 16348 25368
rect 16438 25334 16506 25368
rect 16596 25334 16664 25368
rect 16754 25334 16822 25368
rect 6538 25038 6572 25072
rect 6730 25038 6764 25072
rect 6922 25038 6956 25072
rect 7114 25038 7148 25072
rect 7306 25038 7340 25072
rect 7498 25038 7532 25072
rect 7690 25038 7724 25072
rect 7882 25038 7916 25072
rect 6634 24510 6668 24544
rect 6826 24510 6860 24544
rect 7018 24510 7052 24544
rect 7210 24510 7244 24544
rect 7402 24510 7436 24544
rect 7594 24510 7628 24544
rect 7786 24510 7820 24544
rect 6634 24402 6668 24436
rect 6826 24402 6860 24436
rect 7018 24402 7052 24436
rect 7210 24402 7244 24436
rect 7402 24402 7436 24436
rect 7594 24402 7628 24436
rect 7786 24402 7820 24436
rect 6538 23874 6572 23908
rect 6730 23874 6764 23908
rect 6922 23874 6956 23908
rect 7114 23874 7148 23908
rect 7306 23874 7340 23908
rect 7498 23874 7532 23908
rect 7690 23874 7724 23908
rect 7882 23874 7916 23908
rect 8758 25038 8792 25072
rect 8950 25038 8984 25072
rect 9142 25038 9176 25072
rect 9334 25038 9368 25072
rect 9526 25038 9560 25072
rect 9718 25038 9752 25072
rect 9910 25038 9944 25072
rect 10102 25038 10136 25072
rect 8854 24510 8888 24544
rect 9046 24510 9080 24544
rect 9238 24510 9272 24544
rect 9430 24510 9464 24544
rect 9622 24510 9656 24544
rect 9814 24510 9848 24544
rect 10006 24510 10040 24544
rect 8854 24402 8888 24436
rect 9046 24402 9080 24436
rect 9238 24402 9272 24436
rect 9430 24402 9464 24436
rect 9622 24402 9656 24436
rect 9814 24402 9848 24436
rect 10006 24402 10040 24436
rect 8758 23874 8792 23908
rect 8950 23874 8984 23908
rect 9142 23874 9176 23908
rect 9334 23874 9368 23908
rect 9526 23874 9560 23908
rect 9718 23874 9752 23908
rect 9910 23874 9944 23908
rect 10102 23874 10136 23908
rect 10938 25038 10972 25072
rect 11130 25038 11164 25072
rect 11322 25038 11356 25072
rect 11514 25038 11548 25072
rect 11706 25038 11740 25072
rect 11898 25038 11932 25072
rect 12090 25038 12124 25072
rect 12282 25038 12316 25072
rect 11034 24510 11068 24544
rect 11226 24510 11260 24544
rect 11418 24510 11452 24544
rect 11610 24510 11644 24544
rect 11802 24510 11836 24544
rect 11994 24510 12028 24544
rect 12186 24510 12220 24544
rect 11034 24402 11068 24436
rect 11226 24402 11260 24436
rect 11418 24402 11452 24436
rect 11610 24402 11644 24436
rect 11802 24402 11836 24436
rect 11994 24402 12028 24436
rect 12186 24402 12220 24436
rect 10938 23874 10972 23908
rect 11130 23874 11164 23908
rect 11322 23874 11356 23908
rect 11514 23874 11548 23908
rect 11706 23874 11740 23908
rect 11898 23874 11932 23908
rect 12090 23874 12124 23908
rect 12282 23874 12316 23908
rect 13118 25038 13152 25072
rect 13310 25038 13344 25072
rect 13502 25038 13536 25072
rect 13694 25038 13728 25072
rect 13886 25038 13920 25072
rect 14078 25038 14112 25072
rect 14270 25038 14304 25072
rect 14462 25038 14496 25072
rect 13214 24510 13248 24544
rect 13406 24510 13440 24544
rect 13598 24510 13632 24544
rect 13790 24510 13824 24544
rect 13982 24510 14016 24544
rect 14174 24510 14208 24544
rect 14366 24510 14400 24544
rect 13214 24402 13248 24436
rect 13406 24402 13440 24436
rect 13598 24402 13632 24436
rect 13790 24402 13824 24436
rect 13982 24402 14016 24436
rect 14174 24402 14208 24436
rect 14366 24402 14400 24436
rect 13118 23874 13152 23908
rect 13310 23874 13344 23908
rect 13502 23874 13536 23908
rect 13694 23874 13728 23908
rect 13886 23874 13920 23908
rect 14078 23874 14112 23908
rect 14270 23874 14304 23908
rect 14462 23874 14496 23908
rect 15318 25038 15352 25072
rect 15510 25038 15544 25072
rect 15702 25038 15736 25072
rect 15894 25038 15928 25072
rect 16086 25038 16120 25072
rect 16278 25038 16312 25072
rect 16470 25038 16504 25072
rect 16662 25038 16696 25072
rect 15414 24510 15448 24544
rect 15606 24510 15640 24544
rect 15798 24510 15832 24544
rect 15990 24510 16024 24544
rect 16182 24510 16216 24544
rect 16374 24510 16408 24544
rect 16566 24510 16600 24544
rect 15414 24402 15448 24436
rect 15606 24402 15640 24436
rect 15798 24402 15832 24436
rect 15990 24402 16024 24436
rect 16182 24402 16216 24436
rect 16374 24402 16408 24436
rect 16566 24402 16600 24436
rect 15318 23874 15352 23908
rect 15510 23874 15544 23908
rect 15702 23874 15736 23908
rect 15894 23874 15928 23908
rect 16086 23874 16120 23908
rect 16278 23874 16312 23908
rect 16470 23874 16504 23908
rect 16662 23874 16696 23908
rect 6754 23460 6788 23494
rect 6946 23460 6980 23494
rect 7138 23460 7172 23494
rect 7330 23460 7364 23494
rect 7522 23460 7556 23494
rect 6658 22950 6692 22984
rect 6850 22950 6884 22984
rect 7042 22950 7076 22984
rect 7234 22950 7268 22984
rect 7426 22950 7460 22984
rect 6658 22842 6692 22876
rect 6850 22842 6884 22876
rect 7042 22842 7076 22876
rect 7234 22842 7268 22876
rect 7426 22842 7460 22876
rect 6754 22332 6788 22366
rect 6946 22332 6980 22366
rect 7138 22332 7172 22366
rect 7330 22332 7364 22366
rect 7522 22332 7556 22366
rect 6754 22224 6788 22258
rect 6946 22224 6980 22258
rect 7138 22224 7172 22258
rect 7330 22224 7364 22258
rect 7522 22224 7556 22258
rect 6658 21714 6692 21748
rect 6850 21714 6884 21748
rect 7042 21714 7076 21748
rect 7234 21714 7268 21748
rect 7426 21714 7460 21748
rect 8474 23460 8508 23494
rect 8666 23460 8700 23494
rect 8858 23460 8892 23494
rect 9050 23460 9084 23494
rect 9242 23460 9276 23494
rect 8378 22950 8412 22984
rect 8570 22950 8604 22984
rect 8762 22950 8796 22984
rect 8954 22950 8988 22984
rect 9146 22950 9180 22984
rect 8378 22842 8412 22876
rect 8570 22842 8604 22876
rect 8762 22842 8796 22876
rect 8954 22842 8988 22876
rect 9146 22842 9180 22876
rect 8474 22332 8508 22366
rect 8666 22332 8700 22366
rect 8858 22332 8892 22366
rect 9050 22332 9084 22366
rect 9242 22332 9276 22366
rect 8474 22224 8508 22258
rect 8666 22224 8700 22258
rect 8858 22224 8892 22258
rect 9050 22224 9084 22258
rect 9242 22224 9276 22258
rect 8378 21714 8412 21748
rect 8570 21714 8604 21748
rect 8762 21714 8796 21748
rect 8954 21714 8988 21748
rect 9146 21714 9180 21748
rect 18958 23452 18992 25020
rect 19286 23452 19320 25020
rect 18454 23070 18488 23104
rect 18646 23070 18680 23104
rect 18838 23070 18872 23104
rect 19030 23070 19064 23104
rect 19222 23070 19256 23104
rect 18358 22542 18392 22576
rect 18550 22542 18584 22576
rect 18742 22542 18776 22576
rect 18934 22542 18968 22576
rect 19126 22542 19160 22576
rect 6672 21314 6840 21348
rect 6930 21314 7098 21348
rect 7188 21314 7356 21348
rect 7446 21314 7614 21348
rect 7704 21314 7872 21348
rect 6672 20804 6840 20838
rect 6930 20804 7098 20838
rect 7188 20804 7356 20838
rect 7446 20804 7614 20838
rect 7704 20804 7872 20838
rect 6672 20696 6840 20730
rect 6930 20696 7098 20730
rect 7188 20696 7356 20730
rect 7446 20696 7614 20730
rect 7704 20696 7872 20730
rect 6672 20186 6840 20220
rect 6930 20186 7098 20220
rect 7188 20186 7356 20220
rect 7446 20186 7614 20220
rect 7704 20186 7872 20220
rect 6672 20078 6840 20112
rect 6930 20078 7098 20112
rect 7188 20078 7356 20112
rect 7446 20078 7614 20112
rect 7704 20078 7872 20112
rect 6672 19568 6840 19602
rect 6930 19568 7098 19602
rect 7188 19568 7356 19602
rect 7446 19568 7614 19602
rect 7704 19568 7872 19602
rect 6672 19460 6840 19494
rect 6930 19460 7098 19494
rect 7188 19460 7356 19494
rect 7446 19460 7614 19494
rect 7704 19460 7872 19494
rect 6672 18950 6840 18984
rect 6930 18950 7098 18984
rect 7188 18950 7356 18984
rect 7446 18950 7614 18984
rect 7704 18950 7872 18984
rect 6672 18842 6840 18876
rect 6930 18842 7098 18876
rect 7188 18842 7356 18876
rect 7446 18842 7614 18876
rect 7704 18842 7872 18876
rect 6672 18332 6840 18366
rect 6930 18332 7098 18366
rect 7188 18332 7356 18366
rect 7446 18332 7614 18366
rect 7704 18332 7872 18366
rect 6672 18224 6840 18258
rect 6930 18224 7098 18258
rect 7188 18224 7356 18258
rect 7446 18224 7614 18258
rect 7704 18224 7872 18258
rect 6672 17714 6840 17748
rect 6930 17714 7098 17748
rect 7188 17714 7356 17748
rect 7446 17714 7614 17748
rect 7704 17714 7872 17748
rect 8392 21314 8560 21348
rect 8650 21314 8818 21348
rect 8908 21314 9076 21348
rect 9166 21314 9334 21348
rect 9424 21314 9592 21348
rect 8392 20804 8560 20838
rect 8650 20804 8818 20838
rect 8908 20804 9076 20838
rect 9166 20804 9334 20838
rect 9424 20804 9592 20838
rect 8392 20696 8560 20730
rect 8650 20696 8818 20730
rect 8908 20696 9076 20730
rect 9166 20696 9334 20730
rect 9424 20696 9592 20730
rect 8392 20186 8560 20220
rect 8650 20186 8818 20220
rect 8908 20186 9076 20220
rect 9166 20186 9334 20220
rect 9424 20186 9592 20220
rect 8392 20078 8560 20112
rect 8650 20078 8818 20112
rect 8908 20078 9076 20112
rect 9166 20078 9334 20112
rect 9424 20078 9592 20112
rect 8392 19568 8560 19602
rect 8650 19568 8818 19602
rect 8908 19568 9076 19602
rect 9166 19568 9334 19602
rect 9424 19568 9592 19602
rect 8392 19460 8560 19494
rect 8650 19460 8818 19494
rect 8908 19460 9076 19494
rect 9166 19460 9334 19494
rect 9424 19460 9592 19494
rect 8392 18950 8560 18984
rect 8650 18950 8818 18984
rect 8908 18950 9076 18984
rect 9166 18950 9334 18984
rect 9424 18950 9592 18984
rect 8392 18842 8560 18876
rect 8650 18842 8818 18876
rect 8908 18842 9076 18876
rect 9166 18842 9334 18876
rect 9424 18842 9592 18876
rect 8392 18332 8560 18366
rect 8650 18332 8818 18366
rect 8908 18332 9076 18366
rect 9166 18332 9334 18366
rect 9424 18332 9592 18366
rect 8392 18224 8560 18258
rect 8650 18224 8818 18258
rect 8908 18224 9076 18258
rect 9166 18224 9334 18258
rect 9424 18224 9592 18258
rect 8392 17714 8560 17748
rect 8650 17714 8818 17748
rect 8908 17714 9076 17748
rect 9166 17714 9334 17748
rect 9424 17714 9592 17748
rect 18454 22202 18488 22236
rect 18646 22202 18680 22236
rect 18838 22202 18872 22236
rect 19030 22202 19064 22236
rect 19222 22202 19256 22236
rect 18358 21692 18392 21726
rect 18550 21692 18584 21726
rect 18742 21692 18776 21726
rect 18934 21692 18968 21726
rect 19126 21692 19160 21726
rect 18358 21584 18392 21618
rect 18550 21584 18584 21618
rect 18742 21584 18776 21618
rect 18934 21584 18968 21618
rect 19126 21584 19160 21618
rect 18454 21074 18488 21108
rect 18646 21074 18680 21108
rect 18838 21074 18872 21108
rect 19030 21074 19064 21108
rect 19222 21074 19256 21108
rect 10314 19764 10348 19798
rect 10506 19764 10540 19798
rect 10698 19764 10732 19798
rect 10218 19254 10252 19288
rect 10410 19254 10444 19288
rect 10602 19254 10636 19288
rect 10794 19254 10828 19288
rect 10218 18842 10252 18876
rect 10410 18842 10444 18876
rect 10602 18842 10636 18876
rect 10794 18842 10828 18876
rect 10986 18842 11020 18876
rect 10314 18332 10348 18366
rect 10506 18332 10540 18366
rect 10698 18332 10732 18366
rect 10890 18332 10924 18366
rect 11082 18332 11116 18366
rect 10314 18224 10348 18258
rect 10506 18224 10540 18258
rect 10698 18224 10732 18258
rect 10890 18224 10924 18258
rect 11082 18224 11116 18258
rect 10218 17714 10252 17748
rect 10410 17714 10444 17748
rect 10602 17714 10636 17748
rect 10794 17714 10828 17748
rect 10986 17714 11020 17748
rect 18372 20718 18540 20752
rect 18630 20718 18798 20752
rect 18888 20718 19056 20752
rect 19146 20718 19314 20752
rect 19404 20718 19572 20752
rect 18372 20208 18540 20242
rect 18630 20208 18798 20242
rect 18888 20208 19056 20242
rect 19146 20208 19314 20242
rect 19404 20208 19572 20242
rect 18372 20100 18540 20134
rect 18630 20100 18798 20134
rect 18888 20100 19056 20134
rect 19146 20100 19314 20134
rect 19404 20100 19572 20134
rect 18372 19590 18540 19624
rect 18630 19590 18798 19624
rect 18888 19590 19056 19624
rect 19146 19590 19314 19624
rect 19404 19590 19572 19624
rect 18372 19482 18540 19516
rect 18630 19482 18798 19516
rect 18888 19482 19056 19516
rect 19146 19482 19314 19516
rect 19404 19482 19572 19516
rect 18372 18972 18540 19006
rect 18630 18972 18798 19006
rect 18888 18972 19056 19006
rect 19146 18972 19314 19006
rect 19404 18972 19572 19006
rect 18372 18864 18540 18898
rect 18630 18864 18798 18898
rect 18888 18864 19056 18898
rect 19146 18864 19314 18898
rect 19404 18864 19572 18898
rect 18372 18354 18540 18388
rect 18630 18354 18798 18388
rect 18888 18354 19056 18388
rect 19146 18354 19314 18388
rect 19404 18354 19572 18388
rect -9906 8272 -9872 8306
rect -9714 8272 -9680 8306
rect -9522 8272 -9488 8306
rect -9330 8272 -9296 8306
rect -9138 8272 -9104 8306
rect -10002 7762 -9968 7796
rect -9810 7762 -9776 7796
rect -9618 7762 -9584 7796
rect -9426 7762 -9392 7796
rect -9234 7762 -9200 7796
rect -10002 7654 -9968 7688
rect -9810 7654 -9776 7688
rect -9618 7654 -9584 7688
rect -9426 7654 -9392 7688
rect -9234 7654 -9200 7688
rect -9906 7144 -9872 7178
rect -9714 7144 -9680 7178
rect -9522 7144 -9488 7178
rect -9330 7144 -9296 7178
rect -9138 7144 -9104 7178
rect -9906 7036 -9872 7070
rect -9714 7036 -9680 7070
rect -9522 7036 -9488 7070
rect -9330 7036 -9296 7070
rect -9138 7036 -9104 7070
rect -10002 6526 -9968 6560
rect -9810 6526 -9776 6560
rect -9618 6526 -9584 6560
rect -9426 6526 -9392 6560
rect -9234 6526 -9200 6560
rect -8742 6600 -8708 8168
rect -8432 6600 -8398 8168
rect -9906 6192 -9872 6226
rect -9714 6192 -9680 6226
rect -9522 6192 -9488 6226
rect -9330 6192 -9296 6226
rect -9138 6192 -9104 6226
rect -10002 5682 -9968 5716
rect -9810 5682 -9776 5716
rect -9618 5682 -9584 5716
rect -9426 5682 -9392 5716
rect -9234 5682 -9200 5716
rect -10002 5574 -9968 5608
rect -9810 5574 -9776 5608
rect -9618 5574 -9584 5608
rect -9426 5574 -9392 5608
rect -9234 5574 -9200 5608
rect -9906 5064 -9872 5098
rect -9714 5064 -9680 5098
rect -9522 5064 -9488 5098
rect -9330 5064 -9296 5098
rect -9138 5064 -9104 5098
rect -9906 4956 -9872 4990
rect -9714 4956 -9680 4990
rect -9522 4956 -9488 4990
rect -9330 4956 -9296 4990
rect -9138 4956 -9104 4990
rect -10002 4446 -9968 4480
rect -9810 4446 -9776 4480
rect -9618 4446 -9584 4480
rect -9426 4446 -9392 4480
rect -9234 4446 -9200 4480
rect 1834 8768 1868 8802
rect 2026 8768 2060 8802
rect 2218 8768 2252 8802
rect 2410 8768 2444 8802
rect 2602 8768 2636 8802
rect 2794 8768 2828 8802
rect 2986 8768 3020 8802
rect 3178 8768 3212 8802
rect 3370 8768 3404 8802
rect 3562 8768 3596 8802
rect 1738 8258 1772 8292
rect 1930 8258 1964 8292
rect 2122 8258 2156 8292
rect 2314 8258 2348 8292
rect 2506 8258 2540 8292
rect 2698 8258 2732 8292
rect 2890 8258 2924 8292
rect 3082 8258 3116 8292
rect 3274 8258 3308 8292
rect 3466 8258 3500 8292
rect 1834 7948 1868 7982
rect 2026 7948 2060 7982
rect 2218 7948 2252 7982
rect 2410 7948 2444 7982
rect 2602 7948 2636 7982
rect 2794 7948 2828 7982
rect 2986 7948 3020 7982
rect 3178 7948 3212 7982
rect 3370 7948 3404 7982
rect 3562 7948 3596 7982
rect 1738 7438 1772 7472
rect 1930 7438 1964 7472
rect 2122 7438 2156 7472
rect 2314 7438 2348 7472
rect 2506 7438 2540 7472
rect 2698 7438 2732 7472
rect 2890 7438 2924 7472
rect 3082 7438 3116 7472
rect 3274 7438 3308 7472
rect 3466 7438 3500 7472
rect 1834 7128 1868 7162
rect 2026 7128 2060 7162
rect 2218 7128 2252 7162
rect 2410 7128 2444 7162
rect 2602 7128 2636 7162
rect 2794 7128 2828 7162
rect 2986 7128 3020 7162
rect 3178 7128 3212 7162
rect 3370 7128 3404 7162
rect 3562 7128 3596 7162
rect 1738 6618 1772 6652
rect 1930 6618 1964 6652
rect 2122 6618 2156 6652
rect 2314 6618 2348 6652
rect 2506 6618 2540 6652
rect 2698 6618 2732 6652
rect 2890 6618 2924 6652
rect 3082 6618 3116 6652
rect 3274 6618 3308 6652
rect 3466 6618 3500 6652
rect 5174 10330 5208 10364
rect 5366 10330 5400 10364
rect 5558 10330 5592 10364
rect 5750 10330 5784 10364
rect 5942 10330 5976 10364
rect 6134 10330 6168 10364
rect 6326 10330 6360 10364
rect 6518 10330 6552 10364
rect 6710 10330 6744 10364
rect 6902 10330 6936 10364
rect 5270 9802 5304 9836
rect 5462 9802 5496 9836
rect 5654 9802 5688 9836
rect 5846 9802 5880 9836
rect 6038 9802 6072 9836
rect 6230 9802 6264 9836
rect 6422 9802 6456 9836
rect 6614 9802 6648 9836
rect 6806 9802 6840 9836
rect 6998 9802 7032 9836
rect 5270 9694 5304 9728
rect 5462 9694 5496 9728
rect 5654 9694 5688 9728
rect 5846 9694 5880 9728
rect 6038 9694 6072 9728
rect 6230 9694 6264 9728
rect 6422 9694 6456 9728
rect 6614 9694 6648 9728
rect 6806 9694 6840 9728
rect 6998 9694 7032 9728
rect 5174 9166 5208 9200
rect 5366 9166 5400 9200
rect 5558 9166 5592 9200
rect 5750 9166 5784 9200
rect 5942 9166 5976 9200
rect 6134 9166 6168 9200
rect 6326 9166 6360 9200
rect 6518 9166 6552 9200
rect 6710 9166 6744 9200
rect 6902 9166 6936 9200
rect 5174 8734 5208 8768
rect 5366 8734 5400 8768
rect 5558 8734 5592 8768
rect 5750 8734 5784 8768
rect 5942 8734 5976 8768
rect 6134 8734 6168 8768
rect 6326 8734 6360 8768
rect 6518 8734 6552 8768
rect 6710 8734 6744 8768
rect 6902 8734 6936 8768
rect 5270 8224 5304 8258
rect 5462 8224 5496 8258
rect 5654 8224 5688 8258
rect 5846 8224 5880 8258
rect 6038 8224 6072 8258
rect 6230 8224 6264 8258
rect 6422 8224 6456 8258
rect 6614 8224 6648 8258
rect 6806 8224 6840 8258
rect 6998 8224 7032 8258
rect 5270 8116 5304 8150
rect 5462 8116 5496 8150
rect 5654 8116 5688 8150
rect 5846 8116 5880 8150
rect 6038 8116 6072 8150
rect 6230 8116 6264 8150
rect 6422 8116 6456 8150
rect 6614 8116 6648 8150
rect 6806 8116 6840 8150
rect 6998 8116 7032 8150
rect 5174 7606 5208 7640
rect 5366 7606 5400 7640
rect 5558 7606 5592 7640
rect 5750 7606 5784 7640
rect 5942 7606 5976 7640
rect 6134 7606 6168 7640
rect 6326 7606 6360 7640
rect 6518 7606 6552 7640
rect 6710 7606 6744 7640
rect 6902 7606 6936 7640
rect -9988 4046 -9820 4080
rect -9730 4046 -9562 4080
rect -9472 4046 -9304 4080
rect -9214 4046 -9046 4080
rect -8956 4046 -8788 4080
rect -9988 3536 -9820 3570
rect -9730 3536 -9562 3570
rect -9472 3536 -9304 3570
rect -9214 3536 -9046 3570
rect -8956 3536 -8788 3570
rect -9988 3428 -9820 3462
rect -9730 3428 -9562 3462
rect -9472 3428 -9304 3462
rect -9214 3428 -9046 3462
rect -8956 3428 -8788 3462
rect -9988 2918 -9820 2952
rect -9730 2918 -9562 2952
rect -9472 2918 -9304 2952
rect -9214 2918 -9046 2952
rect -8956 2918 -8788 2952
rect -9988 2810 -9820 2844
rect -9730 2810 -9562 2844
rect -9472 2810 -9304 2844
rect -9214 2810 -9046 2844
rect -8956 2810 -8788 2844
rect -9988 2300 -9820 2334
rect -9730 2300 -9562 2334
rect -9472 2300 -9304 2334
rect -9214 2300 -9046 2334
rect -8956 2300 -8788 2334
rect -9988 2192 -9820 2226
rect -9730 2192 -9562 2226
rect -9472 2192 -9304 2226
rect -9214 2192 -9046 2226
rect -8956 2192 -8788 2226
rect -9988 1682 -9820 1716
rect -9730 1682 -9562 1716
rect -9472 1682 -9304 1716
rect -9214 1682 -9046 1716
rect -8956 1682 -8788 1716
rect -9988 1574 -9820 1608
rect -9730 1574 -9562 1608
rect -9472 1574 -9304 1608
rect -9214 1574 -9046 1608
rect -8956 1574 -8788 1608
rect -9988 1064 -9820 1098
rect -9730 1064 -9562 1098
rect -9472 1064 -9304 1098
rect -9214 1064 -9046 1098
rect -8956 1064 -8788 1098
rect -9988 956 -9820 990
rect -9730 956 -9562 990
rect -9472 956 -9304 990
rect -9214 956 -9046 990
rect -8956 956 -8788 990
rect -9988 446 -9820 480
rect -9730 446 -9562 480
rect -9472 446 -9304 480
rect -9214 446 -9046 480
rect -8956 446 -8788 480
rect 370 5912 404 5946
rect 562 5912 596 5946
rect 754 5912 788 5946
rect 946 5912 980 5946
rect 1138 5912 1172 5946
rect 274 5402 308 5436
rect 466 5402 500 5436
rect 658 5402 692 5436
rect 850 5402 884 5436
rect 1042 5402 1076 5436
rect 274 5294 308 5328
rect 466 5294 500 5328
rect 658 5294 692 5328
rect 850 5294 884 5328
rect 1042 5294 1076 5328
rect 370 4784 404 4818
rect 562 4784 596 4818
rect 754 4784 788 4818
rect 946 4784 980 4818
rect 1138 4784 1172 4818
rect 370 4676 404 4710
rect 562 4676 596 4710
rect 754 4676 788 4710
rect 946 4676 980 4710
rect 1138 4676 1172 4710
rect 274 4166 308 4200
rect 466 4166 500 4200
rect 658 4166 692 4200
rect 850 4166 884 4200
rect 1042 4166 1076 4200
rect 2170 5912 2204 5946
rect 2362 5912 2396 5946
rect 2554 5912 2588 5946
rect 2746 5912 2780 5946
rect 2938 5912 2972 5946
rect 2074 5402 2108 5436
rect 2266 5402 2300 5436
rect 2458 5402 2492 5436
rect 2650 5402 2684 5436
rect 2842 5402 2876 5436
rect 2074 5294 2108 5328
rect 2266 5294 2300 5328
rect 2458 5294 2492 5328
rect 2650 5294 2684 5328
rect 2842 5294 2876 5328
rect 2170 4784 2204 4818
rect 2362 4784 2396 4818
rect 2554 4784 2588 4818
rect 2746 4784 2780 4818
rect 2938 4784 2972 4818
rect 2170 4676 2204 4710
rect 2362 4676 2396 4710
rect 2554 4676 2588 4710
rect 2746 4676 2780 4710
rect 2938 4676 2972 4710
rect 2074 4166 2108 4200
rect 2266 4166 2300 4200
rect 2458 4166 2492 4200
rect 2650 4166 2684 4200
rect 2842 4166 2876 4200
rect 3970 5912 4004 5946
rect 4162 5912 4196 5946
rect 4354 5912 4388 5946
rect 4546 5912 4580 5946
rect 4738 5912 4772 5946
rect 3874 5402 3908 5436
rect 4066 5402 4100 5436
rect 4258 5402 4292 5436
rect 4450 5402 4484 5436
rect 4642 5402 4676 5436
rect 3874 5294 3908 5328
rect 4066 5294 4100 5328
rect 4258 5294 4292 5328
rect 4450 5294 4484 5328
rect 4642 5294 4676 5328
rect 3970 4784 4004 4818
rect 4162 4784 4196 4818
rect 4354 4784 4388 4818
rect 4546 4784 4580 4818
rect 4738 4784 4772 4818
rect 3970 4676 4004 4710
rect 4162 4676 4196 4710
rect 4354 4676 4388 4710
rect 4546 4676 4580 4710
rect 4738 4676 4772 4710
rect 3874 4166 3908 4200
rect 4066 4166 4100 4200
rect 4258 4166 4292 4200
rect 4450 4166 4484 4200
rect 4642 4166 4676 4200
rect 5770 5912 5804 5946
rect 5962 5912 5996 5946
rect 6154 5912 6188 5946
rect 6346 5912 6380 5946
rect 6538 5912 6572 5946
rect 5674 5402 5708 5436
rect 5866 5402 5900 5436
rect 6058 5402 6092 5436
rect 6250 5402 6284 5436
rect 6442 5402 6476 5436
rect 5674 5294 5708 5328
rect 5866 5294 5900 5328
rect 6058 5294 6092 5328
rect 6250 5294 6284 5328
rect 6442 5294 6476 5328
rect 5770 4784 5804 4818
rect 5962 4784 5996 4818
rect 6154 4784 6188 4818
rect 6346 4784 6380 4818
rect 6538 4784 6572 4818
rect 5770 4676 5804 4710
rect 5962 4676 5996 4710
rect 6154 4676 6188 4710
rect 6346 4676 6380 4710
rect 6538 4676 6572 4710
rect 5674 4166 5708 4200
rect 5866 4166 5900 4200
rect 6058 4166 6092 4200
rect 6250 4166 6284 4200
rect 6442 4166 6476 4200
rect 7770 10300 7804 10334
rect 7962 10300 7996 10334
rect 8154 10300 8188 10334
rect 8346 10300 8380 10334
rect 8538 10300 8572 10334
rect 8730 10300 8764 10334
rect 8922 10300 8956 10334
rect 9114 10300 9148 10334
rect 9306 10300 9340 10334
rect 9498 10300 9532 10334
rect 7674 9790 7708 9824
rect 7866 9790 7900 9824
rect 8058 9790 8092 9824
rect 8250 9790 8284 9824
rect 8442 9790 8476 9824
rect 8634 9790 8668 9824
rect 8826 9790 8860 9824
rect 9018 9790 9052 9824
rect 9210 9790 9244 9824
rect 9402 9790 9436 9824
rect 7674 9682 7708 9716
rect 7866 9682 7900 9716
rect 8058 9682 8092 9716
rect 8250 9682 8284 9716
rect 8442 9682 8476 9716
rect 8634 9682 8668 9716
rect 8826 9682 8860 9716
rect 9018 9682 9052 9716
rect 9210 9682 9244 9716
rect 9402 9682 9436 9716
rect 7770 9172 7804 9206
rect 7962 9172 7996 9206
rect 8154 9172 8188 9206
rect 8346 9172 8380 9206
rect 8538 9172 8572 9206
rect 8730 9172 8764 9206
rect 8922 9172 8956 9206
rect 9114 9172 9148 9206
rect 9306 9172 9340 9206
rect 9498 9172 9532 9206
rect 7770 9064 7804 9098
rect 7962 9064 7996 9098
rect 8154 9064 8188 9098
rect 8346 9064 8380 9098
rect 8538 9064 8572 9098
rect 8730 9064 8764 9098
rect 8922 9064 8956 9098
rect 9114 9064 9148 9098
rect 9306 9064 9340 9098
rect 9498 9064 9532 9098
rect 7674 8554 7708 8588
rect 7866 8554 7900 8588
rect 8058 8554 8092 8588
rect 8250 8554 8284 8588
rect 8442 8554 8476 8588
rect 8634 8554 8668 8588
rect 8826 8554 8860 8588
rect 9018 8554 9052 8588
rect 9210 8554 9244 8588
rect 9402 8554 9436 8588
rect 7674 8446 7708 8480
rect 7866 8446 7900 8480
rect 8058 8446 8092 8480
rect 8250 8446 8284 8480
rect 8442 8446 8476 8480
rect 8634 8446 8668 8480
rect 8826 8446 8860 8480
rect 9018 8446 9052 8480
rect 9210 8446 9244 8480
rect 9402 8446 9436 8480
rect 7770 7936 7804 7970
rect 7962 7936 7996 7970
rect 8154 7936 8188 7970
rect 8346 7936 8380 7970
rect 8538 7936 8572 7970
rect 8730 7936 8764 7970
rect 8922 7936 8956 7970
rect 9114 7936 9148 7970
rect 9306 7936 9340 7970
rect 9498 7936 9532 7970
rect 7770 7828 7804 7862
rect 7962 7828 7996 7862
rect 8154 7828 8188 7862
rect 8346 7828 8380 7862
rect 8538 7828 8572 7862
rect 8730 7828 8764 7862
rect 8922 7828 8956 7862
rect 9114 7828 9148 7862
rect 9306 7828 9340 7862
rect 9498 7828 9532 7862
rect 7674 7318 7708 7352
rect 7866 7318 7900 7352
rect 8058 7318 8092 7352
rect 8250 7318 8284 7352
rect 8442 7318 8476 7352
rect 8634 7318 8668 7352
rect 8826 7318 8860 7352
rect 9018 7318 9052 7352
rect 9210 7318 9244 7352
rect 9402 7318 9436 7352
rect 7674 7210 7708 7244
rect 7866 7210 7900 7244
rect 8058 7210 8092 7244
rect 8250 7210 8284 7244
rect 8442 7210 8476 7244
rect 8634 7210 8668 7244
rect 8826 7210 8860 7244
rect 9018 7210 9052 7244
rect 9210 7210 9244 7244
rect 9402 7210 9436 7244
rect 7770 6700 7804 6734
rect 7962 6700 7996 6734
rect 8154 6700 8188 6734
rect 8346 6700 8380 6734
rect 8538 6700 8572 6734
rect 8730 6700 8764 6734
rect 8922 6700 8956 6734
rect 9114 6700 9148 6734
rect 9306 6700 9340 6734
rect 9498 6700 9532 6734
rect 7770 6592 7804 6626
rect 7962 6592 7996 6626
rect 8154 6592 8188 6626
rect 8346 6592 8380 6626
rect 8538 6592 8572 6626
rect 8730 6592 8764 6626
rect 8922 6592 8956 6626
rect 9114 6592 9148 6626
rect 9306 6592 9340 6626
rect 9498 6592 9532 6626
rect 7674 6082 7708 6116
rect 7866 6082 7900 6116
rect 8058 6082 8092 6116
rect 8250 6082 8284 6116
rect 8442 6082 8476 6116
rect 8634 6082 8668 6116
rect 8826 6082 8860 6116
rect 9018 6082 9052 6116
rect 9210 6082 9244 6116
rect 9402 6082 9436 6116
rect 7674 5974 7708 6008
rect 7866 5974 7900 6008
rect 8058 5974 8092 6008
rect 8250 5974 8284 6008
rect 8442 5974 8476 6008
rect 8634 5974 8668 6008
rect 8826 5974 8860 6008
rect 9018 5974 9052 6008
rect 9210 5974 9244 6008
rect 9402 5974 9436 6008
rect 7770 5464 7804 5498
rect 7962 5464 7996 5498
rect 8154 5464 8188 5498
rect 8346 5464 8380 5498
rect 8538 5464 8572 5498
rect 8730 5464 8764 5498
rect 8922 5464 8956 5498
rect 9114 5464 9148 5498
rect 9306 5464 9340 5498
rect 9498 5464 9532 5498
rect 7770 5356 7804 5390
rect 7962 5356 7996 5390
rect 8154 5356 8188 5390
rect 8346 5356 8380 5390
rect 8538 5356 8572 5390
rect 8730 5356 8764 5390
rect 8922 5356 8956 5390
rect 9114 5356 9148 5390
rect 9306 5356 9340 5390
rect 9498 5356 9532 5390
rect 7674 4846 7708 4880
rect 7866 4846 7900 4880
rect 8058 4846 8092 4880
rect 8250 4846 8284 4880
rect 8442 4846 8476 4880
rect 8634 4846 8668 4880
rect 8826 4846 8860 4880
rect 9018 4846 9052 4880
rect 9210 4846 9244 4880
rect 9402 4846 9436 4880
rect 16234 8768 16268 8802
rect 16426 8768 16460 8802
rect 16618 8768 16652 8802
rect 16810 8768 16844 8802
rect 17002 8768 17036 8802
rect 17194 8768 17228 8802
rect 17386 8768 17420 8802
rect 17578 8768 17612 8802
rect 17770 8768 17804 8802
rect 17962 8768 17996 8802
rect 16138 8258 16172 8292
rect 16330 8258 16364 8292
rect 16522 8258 16556 8292
rect 16714 8258 16748 8292
rect 16906 8258 16940 8292
rect 17098 8258 17132 8292
rect 17290 8258 17324 8292
rect 17482 8258 17516 8292
rect 17674 8258 17708 8292
rect 17866 8258 17900 8292
rect 16234 7948 16268 7982
rect 16426 7948 16460 7982
rect 16618 7948 16652 7982
rect 16810 7948 16844 7982
rect 17002 7948 17036 7982
rect 17194 7948 17228 7982
rect 17386 7948 17420 7982
rect 17578 7948 17612 7982
rect 17770 7948 17804 7982
rect 17962 7948 17996 7982
rect 16138 7438 16172 7472
rect 16330 7438 16364 7472
rect 16522 7438 16556 7472
rect 16714 7438 16748 7472
rect 16906 7438 16940 7472
rect 17098 7438 17132 7472
rect 17290 7438 17324 7472
rect 17482 7438 17516 7472
rect 17674 7438 17708 7472
rect 17866 7438 17900 7472
rect 16234 7128 16268 7162
rect 16426 7128 16460 7162
rect 16618 7128 16652 7162
rect 16810 7128 16844 7162
rect 17002 7128 17036 7162
rect 17194 7128 17228 7162
rect 17386 7128 17420 7162
rect 17578 7128 17612 7162
rect 17770 7128 17804 7162
rect 17962 7128 17996 7162
rect 16138 6618 16172 6652
rect 16330 6618 16364 6652
rect 16522 6618 16556 6652
rect 16714 6618 16748 6652
rect 16906 6618 16940 6652
rect 17098 6618 17132 6652
rect 17290 6618 17324 6652
rect 17482 6618 17516 6652
rect 17674 6618 17708 6652
rect 17866 6618 17900 6652
rect 19574 10330 19608 10364
rect 19766 10330 19800 10364
rect 19958 10330 19992 10364
rect 20150 10330 20184 10364
rect 20342 10330 20376 10364
rect 20534 10330 20568 10364
rect 20726 10330 20760 10364
rect 20918 10330 20952 10364
rect 21110 10330 21144 10364
rect 21302 10330 21336 10364
rect 19670 9802 19704 9836
rect 19862 9802 19896 9836
rect 20054 9802 20088 9836
rect 20246 9802 20280 9836
rect 20438 9802 20472 9836
rect 20630 9802 20664 9836
rect 20822 9802 20856 9836
rect 21014 9802 21048 9836
rect 21206 9802 21240 9836
rect 21398 9802 21432 9836
rect 19670 9694 19704 9728
rect 19862 9694 19896 9728
rect 20054 9694 20088 9728
rect 20246 9694 20280 9728
rect 20438 9694 20472 9728
rect 20630 9694 20664 9728
rect 20822 9694 20856 9728
rect 21014 9694 21048 9728
rect 21206 9694 21240 9728
rect 21398 9694 21432 9728
rect 19574 9166 19608 9200
rect 19766 9166 19800 9200
rect 19958 9166 19992 9200
rect 20150 9166 20184 9200
rect 20342 9166 20376 9200
rect 20534 9166 20568 9200
rect 20726 9166 20760 9200
rect 20918 9166 20952 9200
rect 21110 9166 21144 9200
rect 21302 9166 21336 9200
rect 19574 8734 19608 8768
rect 19766 8734 19800 8768
rect 19958 8734 19992 8768
rect 20150 8734 20184 8768
rect 20342 8734 20376 8768
rect 20534 8734 20568 8768
rect 20726 8734 20760 8768
rect 20918 8734 20952 8768
rect 21110 8734 21144 8768
rect 21302 8734 21336 8768
rect 19670 8224 19704 8258
rect 19862 8224 19896 8258
rect 20054 8224 20088 8258
rect 20246 8224 20280 8258
rect 20438 8224 20472 8258
rect 20630 8224 20664 8258
rect 20822 8224 20856 8258
rect 21014 8224 21048 8258
rect 21206 8224 21240 8258
rect 21398 8224 21432 8258
rect 19670 8116 19704 8150
rect 19862 8116 19896 8150
rect 20054 8116 20088 8150
rect 20246 8116 20280 8150
rect 20438 8116 20472 8150
rect 20630 8116 20664 8150
rect 20822 8116 20856 8150
rect 21014 8116 21048 8150
rect 21206 8116 21240 8150
rect 21398 8116 21432 8150
rect 19574 7606 19608 7640
rect 19766 7606 19800 7640
rect 19958 7606 19992 7640
rect 20150 7606 20184 7640
rect 20342 7606 20376 7640
rect 20534 7606 20568 7640
rect 20726 7606 20760 7640
rect 20918 7606 20952 7640
rect 21110 7606 21144 7640
rect 21302 7606 21336 7640
rect 14770 5912 14804 5946
rect 14962 5912 14996 5946
rect 15154 5912 15188 5946
rect 15346 5912 15380 5946
rect 15538 5912 15572 5946
rect 14674 5402 14708 5436
rect 14866 5402 14900 5436
rect 15058 5402 15092 5436
rect 15250 5402 15284 5436
rect 15442 5402 15476 5436
rect 14674 5294 14708 5328
rect 14866 5294 14900 5328
rect 15058 5294 15092 5328
rect 15250 5294 15284 5328
rect 15442 5294 15476 5328
rect 14770 4784 14804 4818
rect 14962 4784 14996 4818
rect 15154 4784 15188 4818
rect 15346 4784 15380 4818
rect 15538 4784 15572 4818
rect 14770 4676 14804 4710
rect 14962 4676 14996 4710
rect 15154 4676 15188 4710
rect 15346 4676 15380 4710
rect 15538 4676 15572 4710
rect 14674 4166 14708 4200
rect 14866 4166 14900 4200
rect 15058 4166 15092 4200
rect 15250 4166 15284 4200
rect 15442 4166 15476 4200
rect 16570 5912 16604 5946
rect 16762 5912 16796 5946
rect 16954 5912 16988 5946
rect 17146 5912 17180 5946
rect 17338 5912 17372 5946
rect 16474 5402 16508 5436
rect 16666 5402 16700 5436
rect 16858 5402 16892 5436
rect 17050 5402 17084 5436
rect 17242 5402 17276 5436
rect 16474 5294 16508 5328
rect 16666 5294 16700 5328
rect 16858 5294 16892 5328
rect 17050 5294 17084 5328
rect 17242 5294 17276 5328
rect 16570 4784 16604 4818
rect 16762 4784 16796 4818
rect 16954 4784 16988 4818
rect 17146 4784 17180 4818
rect 17338 4784 17372 4818
rect 16570 4676 16604 4710
rect 16762 4676 16796 4710
rect 16954 4676 16988 4710
rect 17146 4676 17180 4710
rect 17338 4676 17372 4710
rect 16474 4166 16508 4200
rect 16666 4166 16700 4200
rect 16858 4166 16892 4200
rect 17050 4166 17084 4200
rect 17242 4166 17276 4200
rect 18370 5912 18404 5946
rect 18562 5912 18596 5946
rect 18754 5912 18788 5946
rect 18946 5912 18980 5946
rect 19138 5912 19172 5946
rect 18274 5402 18308 5436
rect 18466 5402 18500 5436
rect 18658 5402 18692 5436
rect 18850 5402 18884 5436
rect 19042 5402 19076 5436
rect 18274 5294 18308 5328
rect 18466 5294 18500 5328
rect 18658 5294 18692 5328
rect 18850 5294 18884 5328
rect 19042 5294 19076 5328
rect 18370 4784 18404 4818
rect 18562 4784 18596 4818
rect 18754 4784 18788 4818
rect 18946 4784 18980 4818
rect 19138 4784 19172 4818
rect 18370 4676 18404 4710
rect 18562 4676 18596 4710
rect 18754 4676 18788 4710
rect 18946 4676 18980 4710
rect 19138 4676 19172 4710
rect 18274 4166 18308 4200
rect 18466 4166 18500 4200
rect 18658 4166 18692 4200
rect 18850 4166 18884 4200
rect 19042 4166 19076 4200
rect 20170 5912 20204 5946
rect 20362 5912 20396 5946
rect 20554 5912 20588 5946
rect 20746 5912 20780 5946
rect 20938 5912 20972 5946
rect 20074 5402 20108 5436
rect 20266 5402 20300 5436
rect 20458 5402 20492 5436
rect 20650 5402 20684 5436
rect 20842 5402 20876 5436
rect 20074 5294 20108 5328
rect 20266 5294 20300 5328
rect 20458 5294 20492 5328
rect 20650 5294 20684 5328
rect 20842 5294 20876 5328
rect 20170 4784 20204 4818
rect 20362 4784 20396 4818
rect 20554 4784 20588 4818
rect 20746 4784 20780 4818
rect 20938 4784 20972 4818
rect 20170 4676 20204 4710
rect 20362 4676 20396 4710
rect 20554 4676 20588 4710
rect 20746 4676 20780 4710
rect 20938 4676 20972 4710
rect 20074 4166 20108 4200
rect 20266 4166 20300 4200
rect 20458 4166 20492 4200
rect 20650 4166 20684 4200
rect 20842 4166 20876 4200
rect 22170 10300 22204 10334
rect 22362 10300 22396 10334
rect 22554 10300 22588 10334
rect 22746 10300 22780 10334
rect 22938 10300 22972 10334
rect 23130 10300 23164 10334
rect 23322 10300 23356 10334
rect 23514 10300 23548 10334
rect 23706 10300 23740 10334
rect 23898 10300 23932 10334
rect 22074 9790 22108 9824
rect 22266 9790 22300 9824
rect 22458 9790 22492 9824
rect 22650 9790 22684 9824
rect 22842 9790 22876 9824
rect 23034 9790 23068 9824
rect 23226 9790 23260 9824
rect 23418 9790 23452 9824
rect 23610 9790 23644 9824
rect 23802 9790 23836 9824
rect 22074 9682 22108 9716
rect 22266 9682 22300 9716
rect 22458 9682 22492 9716
rect 22650 9682 22684 9716
rect 22842 9682 22876 9716
rect 23034 9682 23068 9716
rect 23226 9682 23260 9716
rect 23418 9682 23452 9716
rect 23610 9682 23644 9716
rect 23802 9682 23836 9716
rect 22170 9172 22204 9206
rect 22362 9172 22396 9206
rect 22554 9172 22588 9206
rect 22746 9172 22780 9206
rect 22938 9172 22972 9206
rect 23130 9172 23164 9206
rect 23322 9172 23356 9206
rect 23514 9172 23548 9206
rect 23706 9172 23740 9206
rect 23898 9172 23932 9206
rect 22170 9064 22204 9098
rect 22362 9064 22396 9098
rect 22554 9064 22588 9098
rect 22746 9064 22780 9098
rect 22938 9064 22972 9098
rect 23130 9064 23164 9098
rect 23322 9064 23356 9098
rect 23514 9064 23548 9098
rect 23706 9064 23740 9098
rect 23898 9064 23932 9098
rect 22074 8554 22108 8588
rect 22266 8554 22300 8588
rect 22458 8554 22492 8588
rect 22650 8554 22684 8588
rect 22842 8554 22876 8588
rect 23034 8554 23068 8588
rect 23226 8554 23260 8588
rect 23418 8554 23452 8588
rect 23610 8554 23644 8588
rect 23802 8554 23836 8588
rect 22074 8446 22108 8480
rect 22266 8446 22300 8480
rect 22458 8446 22492 8480
rect 22650 8446 22684 8480
rect 22842 8446 22876 8480
rect 23034 8446 23068 8480
rect 23226 8446 23260 8480
rect 23418 8446 23452 8480
rect 23610 8446 23644 8480
rect 23802 8446 23836 8480
rect 22170 7936 22204 7970
rect 22362 7936 22396 7970
rect 22554 7936 22588 7970
rect 22746 7936 22780 7970
rect 22938 7936 22972 7970
rect 23130 7936 23164 7970
rect 23322 7936 23356 7970
rect 23514 7936 23548 7970
rect 23706 7936 23740 7970
rect 23898 7936 23932 7970
rect 22170 7828 22204 7862
rect 22362 7828 22396 7862
rect 22554 7828 22588 7862
rect 22746 7828 22780 7862
rect 22938 7828 22972 7862
rect 23130 7828 23164 7862
rect 23322 7828 23356 7862
rect 23514 7828 23548 7862
rect 23706 7828 23740 7862
rect 23898 7828 23932 7862
rect 22074 7318 22108 7352
rect 22266 7318 22300 7352
rect 22458 7318 22492 7352
rect 22650 7318 22684 7352
rect 22842 7318 22876 7352
rect 23034 7318 23068 7352
rect 23226 7318 23260 7352
rect 23418 7318 23452 7352
rect 23610 7318 23644 7352
rect 23802 7318 23836 7352
rect 22074 7210 22108 7244
rect 22266 7210 22300 7244
rect 22458 7210 22492 7244
rect 22650 7210 22684 7244
rect 22842 7210 22876 7244
rect 23034 7210 23068 7244
rect 23226 7210 23260 7244
rect 23418 7210 23452 7244
rect 23610 7210 23644 7244
rect 23802 7210 23836 7244
rect 22170 6700 22204 6734
rect 22362 6700 22396 6734
rect 22554 6700 22588 6734
rect 22746 6700 22780 6734
rect 22938 6700 22972 6734
rect 23130 6700 23164 6734
rect 23322 6700 23356 6734
rect 23514 6700 23548 6734
rect 23706 6700 23740 6734
rect 23898 6700 23932 6734
rect 22170 6592 22204 6626
rect 22362 6592 22396 6626
rect 22554 6592 22588 6626
rect 22746 6592 22780 6626
rect 22938 6592 22972 6626
rect 23130 6592 23164 6626
rect 23322 6592 23356 6626
rect 23514 6592 23548 6626
rect 23706 6592 23740 6626
rect 23898 6592 23932 6626
rect 22074 6082 22108 6116
rect 22266 6082 22300 6116
rect 22458 6082 22492 6116
rect 22650 6082 22684 6116
rect 22842 6082 22876 6116
rect 23034 6082 23068 6116
rect 23226 6082 23260 6116
rect 23418 6082 23452 6116
rect 23610 6082 23644 6116
rect 23802 6082 23836 6116
rect 22074 5974 22108 6008
rect 22266 5974 22300 6008
rect 22458 5974 22492 6008
rect 22650 5974 22684 6008
rect 22842 5974 22876 6008
rect 23034 5974 23068 6008
rect 23226 5974 23260 6008
rect 23418 5974 23452 6008
rect 23610 5974 23644 6008
rect 23802 5974 23836 6008
rect 22170 5464 22204 5498
rect 22362 5464 22396 5498
rect 22554 5464 22588 5498
rect 22746 5464 22780 5498
rect 22938 5464 22972 5498
rect 23130 5464 23164 5498
rect 23322 5464 23356 5498
rect 23514 5464 23548 5498
rect 23706 5464 23740 5498
rect 23898 5464 23932 5498
rect 22170 5356 22204 5390
rect 22362 5356 22396 5390
rect 22554 5356 22588 5390
rect 22746 5356 22780 5390
rect 22938 5356 22972 5390
rect 23130 5356 23164 5390
rect 23322 5356 23356 5390
rect 23514 5356 23548 5390
rect 23706 5356 23740 5390
rect 23898 5356 23932 5390
rect 22074 4846 22108 4880
rect 22266 4846 22300 4880
rect 22458 4846 22492 4880
rect 22650 4846 22684 4880
rect 22842 4846 22876 4880
rect 23034 4846 23068 4880
rect 23226 4846 23260 4880
rect 23418 4846 23452 4880
rect 23610 4846 23644 4880
rect 23802 4846 23836 4880
rect 288 3766 456 3800
rect 546 3766 714 3800
rect 804 3766 972 3800
rect 1062 3766 1230 3800
rect 1320 3766 1488 3800
rect 288 3256 456 3290
rect 546 3256 714 3290
rect 804 3256 972 3290
rect 1062 3256 1230 3290
rect 1320 3256 1488 3290
rect 288 3148 456 3182
rect 546 3148 714 3182
rect 804 3148 972 3182
rect 1062 3148 1230 3182
rect 1320 3148 1488 3182
rect 288 2638 456 2672
rect 546 2638 714 2672
rect 804 2638 972 2672
rect 1062 2638 1230 2672
rect 1320 2638 1488 2672
rect 288 2530 456 2564
rect 546 2530 714 2564
rect 804 2530 972 2564
rect 1062 2530 1230 2564
rect 1320 2530 1488 2564
rect 288 2020 456 2054
rect 546 2020 714 2054
rect 804 2020 972 2054
rect 1062 2020 1230 2054
rect 1320 2020 1488 2054
rect 288 1912 456 1946
rect 546 1912 714 1946
rect 804 1912 972 1946
rect 1062 1912 1230 1946
rect 1320 1912 1488 1946
rect 288 1402 456 1436
rect 546 1402 714 1436
rect 804 1402 972 1436
rect 1062 1402 1230 1436
rect 1320 1402 1488 1436
rect 288 1294 456 1328
rect 546 1294 714 1328
rect 804 1294 972 1328
rect 1062 1294 1230 1328
rect 1320 1294 1488 1328
rect 288 784 456 818
rect 546 784 714 818
rect 804 784 972 818
rect 1062 784 1230 818
rect 1320 784 1488 818
rect 288 676 456 710
rect 546 676 714 710
rect 804 676 972 710
rect 1062 676 1230 710
rect 1320 676 1488 710
rect 288 166 456 200
rect 546 166 714 200
rect 804 166 972 200
rect 1062 166 1230 200
rect 1320 166 1488 200
rect 2088 3766 2256 3800
rect 2346 3766 2514 3800
rect 2604 3766 2772 3800
rect 2862 3766 3030 3800
rect 3120 3766 3288 3800
rect 2088 3256 2256 3290
rect 2346 3256 2514 3290
rect 2604 3256 2772 3290
rect 2862 3256 3030 3290
rect 3120 3256 3288 3290
rect 2088 3148 2256 3182
rect 2346 3148 2514 3182
rect 2604 3148 2772 3182
rect 2862 3148 3030 3182
rect 3120 3148 3288 3182
rect 2088 2638 2256 2672
rect 2346 2638 2514 2672
rect 2604 2638 2772 2672
rect 2862 2638 3030 2672
rect 3120 2638 3288 2672
rect 2088 2530 2256 2564
rect 2346 2530 2514 2564
rect 2604 2530 2772 2564
rect 2862 2530 3030 2564
rect 3120 2530 3288 2564
rect 2088 2020 2256 2054
rect 2346 2020 2514 2054
rect 2604 2020 2772 2054
rect 2862 2020 3030 2054
rect 3120 2020 3288 2054
rect 2088 1912 2256 1946
rect 2346 1912 2514 1946
rect 2604 1912 2772 1946
rect 2862 1912 3030 1946
rect 3120 1912 3288 1946
rect 2088 1402 2256 1436
rect 2346 1402 2514 1436
rect 2604 1402 2772 1436
rect 2862 1402 3030 1436
rect 3120 1402 3288 1436
rect 2088 1294 2256 1328
rect 2346 1294 2514 1328
rect 2604 1294 2772 1328
rect 2862 1294 3030 1328
rect 3120 1294 3288 1328
rect 2088 784 2256 818
rect 2346 784 2514 818
rect 2604 784 2772 818
rect 2862 784 3030 818
rect 3120 784 3288 818
rect 2088 676 2256 710
rect 2346 676 2514 710
rect 2604 676 2772 710
rect 2862 676 3030 710
rect 3120 676 3288 710
rect 2088 166 2256 200
rect 2346 166 2514 200
rect 2604 166 2772 200
rect 2862 166 3030 200
rect 3120 166 3288 200
rect 3888 3766 4056 3800
rect 4146 3766 4314 3800
rect 4404 3766 4572 3800
rect 4662 3766 4830 3800
rect 4920 3766 5088 3800
rect 3888 3256 4056 3290
rect 4146 3256 4314 3290
rect 4404 3256 4572 3290
rect 4662 3256 4830 3290
rect 4920 3256 5088 3290
rect 3888 3148 4056 3182
rect 4146 3148 4314 3182
rect 4404 3148 4572 3182
rect 4662 3148 4830 3182
rect 4920 3148 5088 3182
rect 3888 2638 4056 2672
rect 4146 2638 4314 2672
rect 4404 2638 4572 2672
rect 4662 2638 4830 2672
rect 4920 2638 5088 2672
rect 3888 2530 4056 2564
rect 4146 2530 4314 2564
rect 4404 2530 4572 2564
rect 4662 2530 4830 2564
rect 4920 2530 5088 2564
rect 3888 2020 4056 2054
rect 4146 2020 4314 2054
rect 4404 2020 4572 2054
rect 4662 2020 4830 2054
rect 4920 2020 5088 2054
rect 3888 1912 4056 1946
rect 4146 1912 4314 1946
rect 4404 1912 4572 1946
rect 4662 1912 4830 1946
rect 4920 1912 5088 1946
rect 3888 1402 4056 1436
rect 4146 1402 4314 1436
rect 4404 1402 4572 1436
rect 4662 1402 4830 1436
rect 4920 1402 5088 1436
rect 3888 1294 4056 1328
rect 4146 1294 4314 1328
rect 4404 1294 4572 1328
rect 4662 1294 4830 1328
rect 4920 1294 5088 1328
rect 3888 784 4056 818
rect 4146 784 4314 818
rect 4404 784 4572 818
rect 4662 784 4830 818
rect 4920 784 5088 818
rect 3888 676 4056 710
rect 4146 676 4314 710
rect 4404 676 4572 710
rect 4662 676 4830 710
rect 4920 676 5088 710
rect 3888 166 4056 200
rect 4146 166 4314 200
rect 4404 166 4572 200
rect 4662 166 4830 200
rect 4920 166 5088 200
rect 5688 3766 5856 3800
rect 5946 3766 6114 3800
rect 6204 3766 6372 3800
rect 6462 3766 6630 3800
rect 6720 3766 6888 3800
rect 5688 3256 5856 3290
rect 5946 3256 6114 3290
rect 6204 3256 6372 3290
rect 6462 3256 6630 3290
rect 6720 3256 6888 3290
rect 5688 3148 5856 3182
rect 5946 3148 6114 3182
rect 6204 3148 6372 3182
rect 6462 3148 6630 3182
rect 6720 3148 6888 3182
rect 5688 2638 5856 2672
rect 5946 2638 6114 2672
rect 6204 2638 6372 2672
rect 6462 2638 6630 2672
rect 6720 2638 6888 2672
rect 5688 2530 5856 2564
rect 5946 2530 6114 2564
rect 6204 2530 6372 2564
rect 6462 2530 6630 2564
rect 6720 2530 6888 2564
rect 5688 2020 5856 2054
rect 5946 2020 6114 2054
rect 6204 2020 6372 2054
rect 6462 2020 6630 2054
rect 6720 2020 6888 2054
rect 5688 1912 5856 1946
rect 5946 1912 6114 1946
rect 6204 1912 6372 1946
rect 6462 1912 6630 1946
rect 6720 1912 6888 1946
rect 5688 1402 5856 1436
rect 5946 1402 6114 1436
rect 6204 1402 6372 1436
rect 6462 1402 6630 1436
rect 6720 1402 6888 1436
rect 5688 1294 5856 1328
rect 5946 1294 6114 1328
rect 6204 1294 6372 1328
rect 6462 1294 6630 1328
rect 6720 1294 6888 1328
rect 5688 784 5856 818
rect 5946 784 6114 818
rect 6204 784 6372 818
rect 6462 784 6630 818
rect 6720 784 6888 818
rect 5688 676 5856 710
rect 5946 676 6114 710
rect 6204 676 6372 710
rect 6462 676 6630 710
rect 6720 676 6888 710
rect 5688 166 5856 200
rect 5946 166 6114 200
rect 6204 166 6372 200
rect 6462 166 6630 200
rect 6720 166 6888 200
rect 14688 3766 14856 3800
rect 14946 3766 15114 3800
rect 15204 3766 15372 3800
rect 15462 3766 15630 3800
rect 15720 3766 15888 3800
rect 14688 3256 14856 3290
rect 14946 3256 15114 3290
rect 15204 3256 15372 3290
rect 15462 3256 15630 3290
rect 15720 3256 15888 3290
rect 14688 3148 14856 3182
rect 14946 3148 15114 3182
rect 15204 3148 15372 3182
rect 15462 3148 15630 3182
rect 15720 3148 15888 3182
rect 14688 2638 14856 2672
rect 14946 2638 15114 2672
rect 15204 2638 15372 2672
rect 15462 2638 15630 2672
rect 15720 2638 15888 2672
rect 14688 2530 14856 2564
rect 14946 2530 15114 2564
rect 15204 2530 15372 2564
rect 15462 2530 15630 2564
rect 15720 2530 15888 2564
rect 14688 2020 14856 2054
rect 14946 2020 15114 2054
rect 15204 2020 15372 2054
rect 15462 2020 15630 2054
rect 15720 2020 15888 2054
rect 14688 1912 14856 1946
rect 14946 1912 15114 1946
rect 15204 1912 15372 1946
rect 15462 1912 15630 1946
rect 15720 1912 15888 1946
rect 14688 1402 14856 1436
rect 14946 1402 15114 1436
rect 15204 1402 15372 1436
rect 15462 1402 15630 1436
rect 15720 1402 15888 1436
rect 14688 1294 14856 1328
rect 14946 1294 15114 1328
rect 15204 1294 15372 1328
rect 15462 1294 15630 1328
rect 15720 1294 15888 1328
rect 14688 784 14856 818
rect 14946 784 15114 818
rect 15204 784 15372 818
rect 15462 784 15630 818
rect 15720 784 15888 818
rect 14688 676 14856 710
rect 14946 676 15114 710
rect 15204 676 15372 710
rect 15462 676 15630 710
rect 15720 676 15888 710
rect 14688 166 14856 200
rect 14946 166 15114 200
rect 15204 166 15372 200
rect 15462 166 15630 200
rect 15720 166 15888 200
rect 16488 3766 16656 3800
rect 16746 3766 16914 3800
rect 17004 3766 17172 3800
rect 17262 3766 17430 3800
rect 17520 3766 17688 3800
rect 16488 3256 16656 3290
rect 16746 3256 16914 3290
rect 17004 3256 17172 3290
rect 17262 3256 17430 3290
rect 17520 3256 17688 3290
rect 16488 3148 16656 3182
rect 16746 3148 16914 3182
rect 17004 3148 17172 3182
rect 17262 3148 17430 3182
rect 17520 3148 17688 3182
rect 16488 2638 16656 2672
rect 16746 2638 16914 2672
rect 17004 2638 17172 2672
rect 17262 2638 17430 2672
rect 17520 2638 17688 2672
rect 16488 2530 16656 2564
rect 16746 2530 16914 2564
rect 17004 2530 17172 2564
rect 17262 2530 17430 2564
rect 17520 2530 17688 2564
rect 16488 2020 16656 2054
rect 16746 2020 16914 2054
rect 17004 2020 17172 2054
rect 17262 2020 17430 2054
rect 17520 2020 17688 2054
rect 16488 1912 16656 1946
rect 16746 1912 16914 1946
rect 17004 1912 17172 1946
rect 17262 1912 17430 1946
rect 17520 1912 17688 1946
rect 16488 1402 16656 1436
rect 16746 1402 16914 1436
rect 17004 1402 17172 1436
rect 17262 1402 17430 1436
rect 17520 1402 17688 1436
rect 16488 1294 16656 1328
rect 16746 1294 16914 1328
rect 17004 1294 17172 1328
rect 17262 1294 17430 1328
rect 17520 1294 17688 1328
rect 16488 784 16656 818
rect 16746 784 16914 818
rect 17004 784 17172 818
rect 17262 784 17430 818
rect 17520 784 17688 818
rect 16488 676 16656 710
rect 16746 676 16914 710
rect 17004 676 17172 710
rect 17262 676 17430 710
rect 17520 676 17688 710
rect 16488 166 16656 200
rect 16746 166 16914 200
rect 17004 166 17172 200
rect 17262 166 17430 200
rect 17520 166 17688 200
rect 18288 3766 18456 3800
rect 18546 3766 18714 3800
rect 18804 3766 18972 3800
rect 19062 3766 19230 3800
rect 19320 3766 19488 3800
rect 18288 3256 18456 3290
rect 18546 3256 18714 3290
rect 18804 3256 18972 3290
rect 19062 3256 19230 3290
rect 19320 3256 19488 3290
rect 18288 3148 18456 3182
rect 18546 3148 18714 3182
rect 18804 3148 18972 3182
rect 19062 3148 19230 3182
rect 19320 3148 19488 3182
rect 18288 2638 18456 2672
rect 18546 2638 18714 2672
rect 18804 2638 18972 2672
rect 19062 2638 19230 2672
rect 19320 2638 19488 2672
rect 18288 2530 18456 2564
rect 18546 2530 18714 2564
rect 18804 2530 18972 2564
rect 19062 2530 19230 2564
rect 19320 2530 19488 2564
rect 18288 2020 18456 2054
rect 18546 2020 18714 2054
rect 18804 2020 18972 2054
rect 19062 2020 19230 2054
rect 19320 2020 19488 2054
rect 18288 1912 18456 1946
rect 18546 1912 18714 1946
rect 18804 1912 18972 1946
rect 19062 1912 19230 1946
rect 19320 1912 19488 1946
rect 18288 1402 18456 1436
rect 18546 1402 18714 1436
rect 18804 1402 18972 1436
rect 19062 1402 19230 1436
rect 19320 1402 19488 1436
rect 18288 1294 18456 1328
rect 18546 1294 18714 1328
rect 18804 1294 18972 1328
rect 19062 1294 19230 1328
rect 19320 1294 19488 1328
rect 18288 784 18456 818
rect 18546 784 18714 818
rect 18804 784 18972 818
rect 19062 784 19230 818
rect 19320 784 19488 818
rect 18288 676 18456 710
rect 18546 676 18714 710
rect 18804 676 18972 710
rect 19062 676 19230 710
rect 19320 676 19488 710
rect 18288 166 18456 200
rect 18546 166 18714 200
rect 18804 166 18972 200
rect 19062 166 19230 200
rect 19320 166 19488 200
rect 20088 3766 20256 3800
rect 20346 3766 20514 3800
rect 20604 3766 20772 3800
rect 20862 3766 21030 3800
rect 21120 3766 21288 3800
rect 20088 3256 20256 3290
rect 20346 3256 20514 3290
rect 20604 3256 20772 3290
rect 20862 3256 21030 3290
rect 21120 3256 21288 3290
rect 20088 3148 20256 3182
rect 20346 3148 20514 3182
rect 20604 3148 20772 3182
rect 20862 3148 21030 3182
rect 21120 3148 21288 3182
rect 20088 2638 20256 2672
rect 20346 2638 20514 2672
rect 20604 2638 20772 2672
rect 20862 2638 21030 2672
rect 21120 2638 21288 2672
rect 20088 2530 20256 2564
rect 20346 2530 20514 2564
rect 20604 2530 20772 2564
rect 20862 2530 21030 2564
rect 21120 2530 21288 2564
rect 20088 2020 20256 2054
rect 20346 2020 20514 2054
rect 20604 2020 20772 2054
rect 20862 2020 21030 2054
rect 21120 2020 21288 2054
rect 20088 1912 20256 1946
rect 20346 1912 20514 1946
rect 20604 1912 20772 1946
rect 20862 1912 21030 1946
rect 21120 1912 21288 1946
rect 20088 1402 20256 1436
rect 20346 1402 20514 1436
rect 20604 1402 20772 1436
rect 20862 1402 21030 1436
rect 21120 1402 21288 1436
rect 20088 1294 20256 1328
rect 20346 1294 20514 1328
rect 20604 1294 20772 1328
rect 20862 1294 21030 1328
rect 21120 1294 21288 1328
rect 20088 784 20256 818
rect 20346 784 20514 818
rect 20604 784 20772 818
rect 20862 784 21030 818
rect 21120 784 21288 818
rect 20088 676 20256 710
rect 20346 676 20514 710
rect 20604 676 20772 710
rect 20862 676 21030 710
rect 21120 676 21288 710
rect 20088 166 20256 200
rect 20346 166 20514 200
rect 20604 166 20772 200
rect 20862 166 21030 200
rect 21120 166 21288 200
<< xpolycontact >>
rect 18326 24654 18608 25086
rect 18326 23422 18608 23854
rect 2602 10686 2884 11118
rect 2602 9454 2884 9886
rect 2980 10686 3262 11118
rect 2980 9454 3262 9886
rect 3358 10686 3640 11118
rect 3358 9454 3640 9886
rect 3736 10686 4018 11118
rect 3736 9454 4018 9886
rect 4114 10686 4396 11118
rect 4114 9454 4396 9886
rect 4492 10686 4774 11118
rect 4492 9454 4774 9886
rect 17002 10686 17284 11118
rect 17002 9454 17284 9886
rect 17380 10686 17662 11118
rect 17380 9454 17662 9886
rect 17758 10686 18040 11118
rect 17758 9454 18040 9886
rect 18136 10686 18418 11118
rect 18136 9454 18418 9886
rect 18514 10686 18796 11118
rect 18514 9454 18796 9886
rect 18892 10686 19174 11118
rect 18892 9454 19174 9886
<< xpolyres >>
rect 18326 23854 18608 24654
rect 2602 9886 2884 10686
rect 2980 9886 3262 10686
rect 3358 9886 3640 10686
rect 3736 9886 4018 10686
rect 4114 9886 4396 10686
rect 4492 9886 4774 10686
rect 17002 9886 17284 10686
rect 17380 9886 17662 10686
rect 17758 9886 18040 10686
rect 18136 9886 18418 10686
rect 18514 9886 18796 10686
rect 18892 9886 19174 10686
<< locali >>
rect 7440 27270 7540 27336
rect 6376 27236 6472 27270
rect 8122 27256 8218 27270
rect 8596 27256 8692 27270
rect 8122 27236 8692 27256
rect 10342 27256 10438 27270
rect 10776 27256 10872 27270
rect 10342 27236 10872 27256
rect 12522 27236 12618 27270
rect 6376 27174 6410 27236
rect 8184 27176 8630 27236
rect 8184 27174 8218 27176
rect 6536 27134 6552 27168
rect 6620 27134 6636 27168
rect 6694 27134 6710 27168
rect 6778 27134 6794 27168
rect 6852 27134 6868 27168
rect 6936 27134 6952 27168
rect 7010 27134 7026 27168
rect 7094 27134 7110 27168
rect 7168 27134 7184 27168
rect 7252 27134 7268 27168
rect 7326 27134 7342 27168
rect 7410 27134 7426 27168
rect 7484 27134 7500 27168
rect 7568 27134 7584 27168
rect 7642 27134 7658 27168
rect 7726 27134 7742 27168
rect 7800 27134 7816 27168
rect 7884 27134 7900 27168
rect 7958 27134 7974 27168
rect 8042 27134 8058 27168
rect 6490 27075 6524 27091
rect 6490 26683 6524 26699
rect 6648 27075 6682 27091
rect 6648 26683 6682 26699
rect 6806 27075 6840 27091
rect 6806 26683 6840 26699
rect 6964 27075 6998 27091
rect 6964 26683 6998 26699
rect 7122 27075 7156 27091
rect 7122 26683 7156 26699
rect 7280 27075 7314 27091
rect 7280 26683 7314 26699
rect 7438 27075 7472 27091
rect 7438 26683 7472 26699
rect 7596 27075 7630 27091
rect 7596 26683 7630 26699
rect 7754 27075 7788 27091
rect 7754 26683 7788 26699
rect 7912 27075 7946 27091
rect 7912 26683 7946 26699
rect 8070 27075 8104 27091
rect 8070 26683 8104 26699
rect 6536 26606 6552 26640
rect 6620 26606 6636 26640
rect 6694 26606 6710 26640
rect 6778 26606 6794 26640
rect 6852 26606 6868 26640
rect 6936 26606 6952 26640
rect 7010 26606 7026 26640
rect 7094 26606 7110 26640
rect 7168 26606 7184 26640
rect 7252 26606 7268 26640
rect 7326 26606 7342 26640
rect 7410 26606 7426 26640
rect 7484 26606 7500 26640
rect 7568 26606 7584 26640
rect 7642 26606 7658 26640
rect 7726 26606 7742 26640
rect 7800 26606 7816 26640
rect 7884 26606 7900 26640
rect 7958 26606 7974 26640
rect 8042 26606 8058 26640
rect 6536 26498 6552 26532
rect 6620 26498 6636 26532
rect 6694 26498 6710 26532
rect 6778 26498 6794 26532
rect 6852 26498 6868 26532
rect 6936 26498 6952 26532
rect 7010 26498 7026 26532
rect 7094 26498 7110 26532
rect 7168 26498 7184 26532
rect 7252 26498 7268 26532
rect 7326 26498 7342 26532
rect 7410 26498 7426 26532
rect 7484 26498 7500 26532
rect 7568 26498 7584 26532
rect 7642 26498 7658 26532
rect 7726 26498 7742 26532
rect 7800 26498 7816 26532
rect 7884 26498 7900 26532
rect 7958 26498 7974 26532
rect 8042 26498 8058 26532
rect 6490 26439 6524 26455
rect 6490 26047 6524 26063
rect 6648 26439 6682 26455
rect 6648 26047 6682 26063
rect 6806 26439 6840 26455
rect 6806 26047 6840 26063
rect 6964 26439 6998 26455
rect 6964 26047 6998 26063
rect 7122 26439 7156 26455
rect 7122 26047 7156 26063
rect 7280 26439 7314 26455
rect 7280 26047 7314 26063
rect 7438 26439 7472 26455
rect 7438 26047 7472 26063
rect 7596 26439 7630 26455
rect 7596 26047 7630 26063
rect 7754 26439 7788 26455
rect 7754 26047 7788 26063
rect 7912 26439 7946 26455
rect 7912 26047 7946 26063
rect 8070 26439 8104 26455
rect 8070 26047 8104 26063
rect 6536 25970 6552 26004
rect 6620 25970 6636 26004
rect 6694 25970 6710 26004
rect 6778 25970 6794 26004
rect 6852 25970 6868 26004
rect 6936 25970 6952 26004
rect 7010 25970 7026 26004
rect 7094 25970 7110 26004
rect 7168 25970 7184 26004
rect 7252 25970 7268 26004
rect 7326 25970 7342 26004
rect 7410 25970 7426 26004
rect 7484 25970 7500 26004
rect 7568 25970 7584 26004
rect 7642 25970 7658 26004
rect 7726 25970 7742 26004
rect 7800 25970 7816 26004
rect 7884 25970 7900 26004
rect 7958 25970 7974 26004
rect 8042 25970 8058 26004
rect 6536 25862 6552 25896
rect 6620 25862 6636 25896
rect 6694 25862 6710 25896
rect 6778 25862 6794 25896
rect 6852 25862 6868 25896
rect 6936 25862 6952 25896
rect 7010 25862 7026 25896
rect 7094 25862 7110 25896
rect 7168 25862 7184 25896
rect 7252 25862 7268 25896
rect 7326 25862 7342 25896
rect 7410 25862 7426 25896
rect 7484 25862 7500 25896
rect 7568 25862 7584 25896
rect 7642 25862 7658 25896
rect 7726 25862 7742 25896
rect 7800 25862 7816 25896
rect 7884 25862 7900 25896
rect 7958 25862 7974 25896
rect 8042 25862 8058 25896
rect 6490 25803 6524 25819
rect 6490 25411 6524 25427
rect 6648 25803 6682 25819
rect 6648 25411 6682 25427
rect 6806 25803 6840 25819
rect 6806 25411 6840 25427
rect 6964 25803 6998 25819
rect 6964 25411 6998 25427
rect 7122 25803 7156 25819
rect 7122 25411 7156 25427
rect 7280 25803 7314 25819
rect 7280 25411 7314 25427
rect 7438 25803 7472 25819
rect 7438 25411 7472 25427
rect 7596 25803 7630 25819
rect 7596 25411 7630 25427
rect 7754 25803 7788 25819
rect 7754 25411 7788 25427
rect 7912 25803 7946 25819
rect 7912 25411 7946 25427
rect 8070 25803 8104 25819
rect 8070 25411 8104 25427
rect 6536 25334 6552 25368
rect 6620 25334 6636 25368
rect 6694 25334 6710 25368
rect 6778 25334 6794 25368
rect 6852 25334 6868 25368
rect 6936 25334 6952 25368
rect 7010 25334 7026 25368
rect 7094 25334 7110 25368
rect 7168 25334 7184 25368
rect 7252 25334 7268 25368
rect 7326 25334 7342 25368
rect 7410 25334 7426 25368
rect 7484 25334 7500 25368
rect 7568 25334 7584 25368
rect 7642 25334 7658 25368
rect 7726 25334 7742 25368
rect 7800 25334 7816 25368
rect 7884 25334 7900 25368
rect 7958 25334 7974 25368
rect 8042 25334 8058 25368
rect 6376 25266 6410 25328
rect 8184 25266 8218 25328
rect 6376 25232 6472 25266
rect 8122 25232 8218 25266
rect 8596 27174 8630 27176
rect 10404 27174 10810 27236
rect 8756 27134 8772 27168
rect 8840 27134 8856 27168
rect 8914 27134 8930 27168
rect 8998 27134 9014 27168
rect 9072 27134 9088 27168
rect 9156 27134 9172 27168
rect 9230 27134 9246 27168
rect 9314 27134 9330 27168
rect 9388 27134 9404 27168
rect 9472 27134 9488 27168
rect 9546 27134 9562 27168
rect 9630 27134 9646 27168
rect 9704 27134 9720 27168
rect 9788 27134 9804 27168
rect 9862 27134 9878 27168
rect 9946 27134 9962 27168
rect 10020 27134 10036 27168
rect 10104 27134 10120 27168
rect 10178 27134 10194 27168
rect 10262 27134 10278 27168
rect 8710 27075 8744 27091
rect 8710 26683 8744 26699
rect 8868 27075 8902 27091
rect 8868 26683 8902 26699
rect 9026 27075 9060 27091
rect 9026 26683 9060 26699
rect 9184 27075 9218 27091
rect 9184 26683 9218 26699
rect 9342 27075 9376 27091
rect 9342 26683 9376 26699
rect 9500 27075 9534 27091
rect 9500 26683 9534 26699
rect 9658 27075 9692 27091
rect 9658 26683 9692 26699
rect 9816 27075 9850 27091
rect 9816 26683 9850 26699
rect 9974 27075 10008 27091
rect 9974 26683 10008 26699
rect 10132 27075 10166 27091
rect 10132 26683 10166 26699
rect 10290 27075 10324 27091
rect 10290 26683 10324 26699
rect 8756 26606 8772 26640
rect 8840 26606 8856 26640
rect 8914 26606 8930 26640
rect 8998 26606 9014 26640
rect 9072 26606 9088 26640
rect 9156 26606 9172 26640
rect 9230 26606 9246 26640
rect 9314 26606 9330 26640
rect 9388 26606 9404 26640
rect 9472 26606 9488 26640
rect 9546 26606 9562 26640
rect 9630 26606 9646 26640
rect 9704 26606 9720 26640
rect 9788 26606 9804 26640
rect 9862 26606 9878 26640
rect 9946 26606 9962 26640
rect 10020 26606 10036 26640
rect 10104 26606 10120 26640
rect 10178 26606 10194 26640
rect 10262 26606 10278 26640
rect 8756 26498 8772 26532
rect 8840 26498 8856 26532
rect 8914 26498 8930 26532
rect 8998 26498 9014 26532
rect 9072 26498 9088 26532
rect 9156 26498 9172 26532
rect 9230 26498 9246 26532
rect 9314 26498 9330 26532
rect 9388 26498 9404 26532
rect 9472 26498 9488 26532
rect 9546 26498 9562 26532
rect 9630 26498 9646 26532
rect 9704 26498 9720 26532
rect 9788 26498 9804 26532
rect 9862 26498 9878 26532
rect 9946 26498 9962 26532
rect 10020 26498 10036 26532
rect 10104 26498 10120 26532
rect 10178 26498 10194 26532
rect 10262 26498 10278 26532
rect 8710 26439 8744 26455
rect 8710 26047 8744 26063
rect 8868 26439 8902 26455
rect 8868 26047 8902 26063
rect 9026 26439 9060 26455
rect 9026 26047 9060 26063
rect 9184 26439 9218 26455
rect 9184 26047 9218 26063
rect 9342 26439 9376 26455
rect 9342 26047 9376 26063
rect 9500 26439 9534 26455
rect 9500 26047 9534 26063
rect 9658 26439 9692 26455
rect 9658 26047 9692 26063
rect 9816 26439 9850 26455
rect 9816 26047 9850 26063
rect 9974 26439 10008 26455
rect 9974 26047 10008 26063
rect 10132 26439 10166 26455
rect 10132 26047 10166 26063
rect 10290 26439 10324 26455
rect 10290 26047 10324 26063
rect 8756 25970 8772 26004
rect 8840 25970 8856 26004
rect 8914 25970 8930 26004
rect 8998 25970 9014 26004
rect 9072 25970 9088 26004
rect 9156 25970 9172 26004
rect 9230 25970 9246 26004
rect 9314 25970 9330 26004
rect 9388 25970 9404 26004
rect 9472 25970 9488 26004
rect 9546 25970 9562 26004
rect 9630 25970 9646 26004
rect 9704 25970 9720 26004
rect 9788 25970 9804 26004
rect 9862 25970 9878 26004
rect 9946 25970 9962 26004
rect 10020 25970 10036 26004
rect 10104 25970 10120 26004
rect 10178 25970 10194 26004
rect 10262 25970 10278 26004
rect 8756 25862 8772 25896
rect 8840 25862 8856 25896
rect 8914 25862 8930 25896
rect 8998 25862 9014 25896
rect 9072 25862 9088 25896
rect 9156 25862 9172 25896
rect 9230 25862 9246 25896
rect 9314 25862 9330 25896
rect 9388 25862 9404 25896
rect 9472 25862 9488 25896
rect 9546 25862 9562 25896
rect 9630 25862 9646 25896
rect 9704 25862 9720 25896
rect 9788 25862 9804 25896
rect 9862 25862 9878 25896
rect 9946 25862 9962 25896
rect 10020 25862 10036 25896
rect 10104 25862 10120 25896
rect 10178 25862 10194 25896
rect 10262 25862 10278 25896
rect 8710 25803 8744 25819
rect 8710 25411 8744 25427
rect 8868 25803 8902 25819
rect 8868 25411 8902 25427
rect 9026 25803 9060 25819
rect 9026 25411 9060 25427
rect 9184 25803 9218 25819
rect 9184 25411 9218 25427
rect 9342 25803 9376 25819
rect 9342 25411 9376 25427
rect 9500 25803 9534 25819
rect 9500 25411 9534 25427
rect 9658 25803 9692 25819
rect 9658 25411 9692 25427
rect 9816 25803 9850 25819
rect 9816 25411 9850 25427
rect 9974 25803 10008 25819
rect 9974 25411 10008 25427
rect 10132 25803 10166 25819
rect 10132 25411 10166 25427
rect 10290 25803 10324 25819
rect 10290 25411 10324 25427
rect 8756 25334 8772 25368
rect 8840 25334 8856 25368
rect 8914 25334 8930 25368
rect 8998 25334 9014 25368
rect 9072 25334 9088 25368
rect 9156 25334 9172 25368
rect 9230 25334 9246 25368
rect 9314 25334 9330 25368
rect 9388 25334 9404 25368
rect 9472 25334 9488 25368
rect 9546 25334 9562 25368
rect 9630 25334 9646 25368
rect 9704 25334 9720 25368
rect 9788 25334 9804 25368
rect 9862 25334 9878 25368
rect 9946 25334 9962 25368
rect 10020 25334 10036 25368
rect 10104 25334 10120 25368
rect 10178 25334 10194 25368
rect 10262 25334 10278 25368
rect 8596 25266 8630 25328
rect 10438 27156 10776 27174
rect 10404 25266 10438 25328
rect 8596 25232 8692 25266
rect 10342 25232 10438 25266
rect 12584 27216 12618 27236
rect 12956 27236 13052 27270
rect 14702 27236 14798 27270
rect 15156 27236 15252 27270
rect 16902 27236 16998 27270
rect 12956 27216 12990 27236
rect 12584 27174 12990 27216
rect 10936 27134 10952 27168
rect 11020 27134 11036 27168
rect 11094 27134 11110 27168
rect 11178 27134 11194 27168
rect 11252 27134 11268 27168
rect 11336 27134 11352 27168
rect 11410 27134 11426 27168
rect 11494 27134 11510 27168
rect 11568 27134 11584 27168
rect 11652 27134 11668 27168
rect 11726 27134 11742 27168
rect 11810 27134 11826 27168
rect 11884 27134 11900 27168
rect 11968 27134 11984 27168
rect 12042 27134 12058 27168
rect 12126 27134 12142 27168
rect 12200 27134 12216 27168
rect 12284 27134 12300 27168
rect 12358 27134 12374 27168
rect 12442 27134 12458 27168
rect 10890 27075 10924 27091
rect 10890 26683 10924 26699
rect 11048 27075 11082 27091
rect 11048 26683 11082 26699
rect 11206 27075 11240 27091
rect 11206 26683 11240 26699
rect 11364 27075 11398 27091
rect 11364 26683 11398 26699
rect 11522 27075 11556 27091
rect 11522 26683 11556 26699
rect 11680 27075 11714 27091
rect 11680 26683 11714 26699
rect 11838 27075 11872 27091
rect 11838 26683 11872 26699
rect 11996 27075 12030 27091
rect 11996 26683 12030 26699
rect 12154 27075 12188 27091
rect 12154 26683 12188 26699
rect 12312 27075 12346 27091
rect 12312 26683 12346 26699
rect 12470 27075 12504 27091
rect 12470 26683 12504 26699
rect 10936 26606 10952 26640
rect 11020 26606 11036 26640
rect 11094 26606 11110 26640
rect 11178 26606 11194 26640
rect 11252 26606 11268 26640
rect 11336 26606 11352 26640
rect 11410 26606 11426 26640
rect 11494 26606 11510 26640
rect 11568 26606 11584 26640
rect 11652 26606 11668 26640
rect 11726 26606 11742 26640
rect 11810 26606 11826 26640
rect 11884 26606 11900 26640
rect 11968 26606 11984 26640
rect 12042 26606 12058 26640
rect 12126 26606 12142 26640
rect 12200 26606 12216 26640
rect 12284 26606 12300 26640
rect 12358 26606 12374 26640
rect 12442 26606 12458 26640
rect 10936 26498 10952 26532
rect 11020 26498 11036 26532
rect 11094 26498 11110 26532
rect 11178 26498 11194 26532
rect 11252 26498 11268 26532
rect 11336 26498 11352 26532
rect 11410 26498 11426 26532
rect 11494 26498 11510 26532
rect 11568 26498 11584 26532
rect 11652 26498 11668 26532
rect 11726 26498 11742 26532
rect 11810 26498 11826 26532
rect 11884 26498 11900 26532
rect 11968 26498 11984 26532
rect 12042 26498 12058 26532
rect 12126 26498 12142 26532
rect 12200 26498 12216 26532
rect 12284 26498 12300 26532
rect 12358 26498 12374 26532
rect 12442 26498 12458 26532
rect 10890 26439 10924 26455
rect 10890 26047 10924 26063
rect 11048 26439 11082 26455
rect 11048 26047 11082 26063
rect 11206 26439 11240 26455
rect 11206 26047 11240 26063
rect 11364 26439 11398 26455
rect 11364 26047 11398 26063
rect 11522 26439 11556 26455
rect 11522 26047 11556 26063
rect 11680 26439 11714 26455
rect 11680 26047 11714 26063
rect 11838 26439 11872 26455
rect 11838 26047 11872 26063
rect 11996 26439 12030 26455
rect 11996 26047 12030 26063
rect 12154 26439 12188 26455
rect 12154 26047 12188 26063
rect 12312 26439 12346 26455
rect 12312 26047 12346 26063
rect 12470 26439 12504 26455
rect 12470 26047 12504 26063
rect 10936 25970 10952 26004
rect 11020 25970 11036 26004
rect 11094 25970 11110 26004
rect 11178 25970 11194 26004
rect 11252 25970 11268 26004
rect 11336 25970 11352 26004
rect 11410 25970 11426 26004
rect 11494 25970 11510 26004
rect 11568 25970 11584 26004
rect 11652 25970 11668 26004
rect 11726 25970 11742 26004
rect 11810 25970 11826 26004
rect 11884 25970 11900 26004
rect 11968 25970 11984 26004
rect 12042 25970 12058 26004
rect 12126 25970 12142 26004
rect 12200 25970 12216 26004
rect 12284 25970 12300 26004
rect 12358 25970 12374 26004
rect 12442 25970 12458 26004
rect 10936 25862 10952 25896
rect 11020 25862 11036 25896
rect 11094 25862 11110 25896
rect 11178 25862 11194 25896
rect 11252 25862 11268 25896
rect 11336 25862 11352 25896
rect 11410 25862 11426 25896
rect 11494 25862 11510 25896
rect 11568 25862 11584 25896
rect 11652 25862 11668 25896
rect 11726 25862 11742 25896
rect 11810 25862 11826 25896
rect 11884 25862 11900 25896
rect 11968 25862 11984 25896
rect 12042 25862 12058 25896
rect 12126 25862 12142 25896
rect 12200 25862 12216 25896
rect 12284 25862 12300 25896
rect 12358 25862 12374 25896
rect 12442 25862 12458 25896
rect 10890 25803 10924 25819
rect 10890 25411 10924 25427
rect 11048 25803 11082 25819
rect 11048 25411 11082 25427
rect 11206 25803 11240 25819
rect 11206 25411 11240 25427
rect 11364 25803 11398 25819
rect 11364 25411 11398 25427
rect 11522 25803 11556 25819
rect 11522 25411 11556 25427
rect 11680 25803 11714 25819
rect 11680 25411 11714 25427
rect 11838 25803 11872 25819
rect 11838 25411 11872 25427
rect 11996 25803 12030 25819
rect 11996 25411 12030 25427
rect 12154 25803 12188 25819
rect 12154 25411 12188 25427
rect 12312 25803 12346 25819
rect 12312 25411 12346 25427
rect 12470 25803 12504 25819
rect 12470 25411 12504 25427
rect 10936 25334 10952 25368
rect 11020 25334 11036 25368
rect 11094 25334 11110 25368
rect 11178 25334 11194 25368
rect 11252 25334 11268 25368
rect 11336 25334 11352 25368
rect 11410 25334 11426 25368
rect 11494 25334 11510 25368
rect 11568 25334 11584 25368
rect 11652 25334 11668 25368
rect 11726 25334 11742 25368
rect 11810 25334 11826 25368
rect 11884 25334 11900 25368
rect 11968 25334 11984 25368
rect 12042 25334 12058 25368
rect 12126 25334 12142 25368
rect 12200 25334 12216 25368
rect 12284 25334 12300 25368
rect 12358 25334 12374 25368
rect 12442 25334 12458 25368
rect 10776 25266 10810 25328
rect 12618 27116 12956 27174
rect 12584 25266 12618 25328
rect 10776 25232 10872 25266
rect 12522 25232 12618 25266
rect 14764 27174 15190 27236
rect 13116 27134 13132 27168
rect 13200 27134 13216 27168
rect 13274 27134 13290 27168
rect 13358 27134 13374 27168
rect 13432 27134 13448 27168
rect 13516 27134 13532 27168
rect 13590 27134 13606 27168
rect 13674 27134 13690 27168
rect 13748 27134 13764 27168
rect 13832 27134 13848 27168
rect 13906 27134 13922 27168
rect 13990 27134 14006 27168
rect 14064 27134 14080 27168
rect 14148 27134 14164 27168
rect 14222 27134 14238 27168
rect 14306 27134 14322 27168
rect 14380 27134 14396 27168
rect 14464 27134 14480 27168
rect 14538 27134 14554 27168
rect 14622 27134 14638 27168
rect 13070 27075 13104 27091
rect 13070 26683 13104 26699
rect 13228 27075 13262 27091
rect 13228 26683 13262 26699
rect 13386 27075 13420 27091
rect 13386 26683 13420 26699
rect 13544 27075 13578 27091
rect 13544 26683 13578 26699
rect 13702 27075 13736 27091
rect 13702 26683 13736 26699
rect 13860 27075 13894 27091
rect 13860 26683 13894 26699
rect 14018 27075 14052 27091
rect 14018 26683 14052 26699
rect 14176 27075 14210 27091
rect 14176 26683 14210 26699
rect 14334 27075 14368 27091
rect 14334 26683 14368 26699
rect 14492 27075 14526 27091
rect 14492 26683 14526 26699
rect 14650 27075 14684 27091
rect 14650 26683 14684 26699
rect 13116 26606 13132 26640
rect 13200 26606 13216 26640
rect 13274 26606 13290 26640
rect 13358 26606 13374 26640
rect 13432 26606 13448 26640
rect 13516 26606 13532 26640
rect 13590 26606 13606 26640
rect 13674 26606 13690 26640
rect 13748 26606 13764 26640
rect 13832 26606 13848 26640
rect 13906 26606 13922 26640
rect 13990 26606 14006 26640
rect 14064 26606 14080 26640
rect 14148 26606 14164 26640
rect 14222 26606 14238 26640
rect 14306 26606 14322 26640
rect 14380 26606 14396 26640
rect 14464 26606 14480 26640
rect 14538 26606 14554 26640
rect 14622 26606 14638 26640
rect 13116 26498 13132 26532
rect 13200 26498 13216 26532
rect 13274 26498 13290 26532
rect 13358 26498 13374 26532
rect 13432 26498 13448 26532
rect 13516 26498 13532 26532
rect 13590 26498 13606 26532
rect 13674 26498 13690 26532
rect 13748 26498 13764 26532
rect 13832 26498 13848 26532
rect 13906 26498 13922 26532
rect 13990 26498 14006 26532
rect 14064 26498 14080 26532
rect 14148 26498 14164 26532
rect 14222 26498 14238 26532
rect 14306 26498 14322 26532
rect 14380 26498 14396 26532
rect 14464 26498 14480 26532
rect 14538 26498 14554 26532
rect 14622 26498 14638 26532
rect 13070 26439 13104 26455
rect 13070 26047 13104 26063
rect 13228 26439 13262 26455
rect 13228 26047 13262 26063
rect 13386 26439 13420 26455
rect 13386 26047 13420 26063
rect 13544 26439 13578 26455
rect 13544 26047 13578 26063
rect 13702 26439 13736 26455
rect 13702 26047 13736 26063
rect 13860 26439 13894 26455
rect 13860 26047 13894 26063
rect 14018 26439 14052 26455
rect 14018 26047 14052 26063
rect 14176 26439 14210 26455
rect 14176 26047 14210 26063
rect 14334 26439 14368 26455
rect 14334 26047 14368 26063
rect 14492 26439 14526 26455
rect 14492 26047 14526 26063
rect 14650 26439 14684 26455
rect 14650 26047 14684 26063
rect 13116 25970 13132 26004
rect 13200 25970 13216 26004
rect 13274 25970 13290 26004
rect 13358 25970 13374 26004
rect 13432 25970 13448 26004
rect 13516 25970 13532 26004
rect 13590 25970 13606 26004
rect 13674 25970 13690 26004
rect 13748 25970 13764 26004
rect 13832 25970 13848 26004
rect 13906 25970 13922 26004
rect 13990 25970 14006 26004
rect 14064 25970 14080 26004
rect 14148 25970 14164 26004
rect 14222 25970 14238 26004
rect 14306 25970 14322 26004
rect 14380 25970 14396 26004
rect 14464 25970 14480 26004
rect 14538 25970 14554 26004
rect 14622 25970 14638 26004
rect 13116 25862 13132 25896
rect 13200 25862 13216 25896
rect 13274 25862 13290 25896
rect 13358 25862 13374 25896
rect 13432 25862 13448 25896
rect 13516 25862 13532 25896
rect 13590 25862 13606 25896
rect 13674 25862 13690 25896
rect 13748 25862 13764 25896
rect 13832 25862 13848 25896
rect 13906 25862 13922 25896
rect 13990 25862 14006 25896
rect 14064 25862 14080 25896
rect 14148 25862 14164 25896
rect 14222 25862 14238 25896
rect 14306 25862 14322 25896
rect 14380 25862 14396 25896
rect 14464 25862 14480 25896
rect 14538 25862 14554 25896
rect 14622 25862 14638 25896
rect 13070 25803 13104 25819
rect 13070 25411 13104 25427
rect 13228 25803 13262 25819
rect 13228 25411 13262 25427
rect 13386 25803 13420 25819
rect 13386 25411 13420 25427
rect 13544 25803 13578 25819
rect 13544 25411 13578 25427
rect 13702 25803 13736 25819
rect 13702 25411 13736 25427
rect 13860 25803 13894 25819
rect 13860 25411 13894 25427
rect 14018 25803 14052 25819
rect 14018 25411 14052 25427
rect 14176 25803 14210 25819
rect 14176 25411 14210 25427
rect 14334 25803 14368 25819
rect 14334 25411 14368 25427
rect 14492 25803 14526 25819
rect 14492 25411 14526 25427
rect 14650 25803 14684 25819
rect 14650 25411 14684 25427
rect 13116 25334 13132 25368
rect 13200 25334 13216 25368
rect 13274 25334 13290 25368
rect 13358 25334 13374 25368
rect 13432 25334 13448 25368
rect 13516 25334 13532 25368
rect 13590 25334 13606 25368
rect 13674 25334 13690 25368
rect 13748 25334 13764 25368
rect 13832 25334 13848 25368
rect 13906 25334 13922 25368
rect 13990 25334 14006 25368
rect 14064 25334 14080 25368
rect 14148 25334 14164 25368
rect 14222 25334 14238 25368
rect 14306 25334 14322 25368
rect 14380 25334 14396 25368
rect 14464 25334 14480 25368
rect 14538 25334 14554 25368
rect 14622 25334 14638 25368
rect 12956 25266 12990 25328
rect 14798 27136 15156 27174
rect 14764 25266 14798 25328
rect 12956 25232 13052 25266
rect 14702 25232 14798 25266
rect 16964 27174 16998 27236
rect 15316 27134 15332 27168
rect 15400 27134 15416 27168
rect 15474 27134 15490 27168
rect 15558 27134 15574 27168
rect 15632 27134 15648 27168
rect 15716 27134 15732 27168
rect 15790 27134 15806 27168
rect 15874 27134 15890 27168
rect 15948 27134 15964 27168
rect 16032 27134 16048 27168
rect 16106 27134 16122 27168
rect 16190 27134 16206 27168
rect 16264 27134 16280 27168
rect 16348 27134 16364 27168
rect 16422 27134 16438 27168
rect 16506 27134 16522 27168
rect 16580 27134 16596 27168
rect 16664 27134 16680 27168
rect 16738 27134 16754 27168
rect 16822 27134 16838 27168
rect 15270 27075 15304 27091
rect 15270 26683 15304 26699
rect 15428 27075 15462 27091
rect 15428 26683 15462 26699
rect 15586 27075 15620 27091
rect 15586 26683 15620 26699
rect 15744 27075 15778 27091
rect 15744 26683 15778 26699
rect 15902 27075 15936 27091
rect 15902 26683 15936 26699
rect 16060 27075 16094 27091
rect 16060 26683 16094 26699
rect 16218 27075 16252 27091
rect 16218 26683 16252 26699
rect 16376 27075 16410 27091
rect 16376 26683 16410 26699
rect 16534 27075 16568 27091
rect 16534 26683 16568 26699
rect 16692 27075 16726 27091
rect 16692 26683 16726 26699
rect 16850 27075 16884 27091
rect 16850 26683 16884 26699
rect 15316 26606 15332 26640
rect 15400 26606 15416 26640
rect 15474 26606 15490 26640
rect 15558 26606 15574 26640
rect 15632 26606 15648 26640
rect 15716 26606 15732 26640
rect 15790 26606 15806 26640
rect 15874 26606 15890 26640
rect 15948 26606 15964 26640
rect 16032 26606 16048 26640
rect 16106 26606 16122 26640
rect 16190 26606 16206 26640
rect 16264 26606 16280 26640
rect 16348 26606 16364 26640
rect 16422 26606 16438 26640
rect 16506 26606 16522 26640
rect 16580 26606 16596 26640
rect 16664 26606 16680 26640
rect 16738 26606 16754 26640
rect 16822 26606 16838 26640
rect 15316 26498 15332 26532
rect 15400 26498 15416 26532
rect 15474 26498 15490 26532
rect 15558 26498 15574 26532
rect 15632 26498 15648 26532
rect 15716 26498 15732 26532
rect 15790 26498 15806 26532
rect 15874 26498 15890 26532
rect 15948 26498 15964 26532
rect 16032 26498 16048 26532
rect 16106 26498 16122 26532
rect 16190 26498 16206 26532
rect 16264 26498 16280 26532
rect 16348 26498 16364 26532
rect 16422 26498 16438 26532
rect 16506 26498 16522 26532
rect 16580 26498 16596 26532
rect 16664 26498 16680 26532
rect 16738 26498 16754 26532
rect 16822 26498 16838 26532
rect 15270 26439 15304 26455
rect 15270 26047 15304 26063
rect 15428 26439 15462 26455
rect 15428 26047 15462 26063
rect 15586 26439 15620 26455
rect 15586 26047 15620 26063
rect 15744 26439 15778 26455
rect 15744 26047 15778 26063
rect 15902 26439 15936 26455
rect 15902 26047 15936 26063
rect 16060 26439 16094 26455
rect 16060 26047 16094 26063
rect 16218 26439 16252 26455
rect 16218 26047 16252 26063
rect 16376 26439 16410 26455
rect 16376 26047 16410 26063
rect 16534 26439 16568 26455
rect 16534 26047 16568 26063
rect 16692 26439 16726 26455
rect 16692 26047 16726 26063
rect 16850 26439 16884 26455
rect 16850 26047 16884 26063
rect 15316 25970 15332 26004
rect 15400 25970 15416 26004
rect 15474 25970 15490 26004
rect 15558 25970 15574 26004
rect 15632 25970 15648 26004
rect 15716 25970 15732 26004
rect 15790 25970 15806 26004
rect 15874 25970 15890 26004
rect 15948 25970 15964 26004
rect 16032 25970 16048 26004
rect 16106 25970 16122 26004
rect 16190 25970 16206 26004
rect 16264 25970 16280 26004
rect 16348 25970 16364 26004
rect 16422 25970 16438 26004
rect 16506 25970 16522 26004
rect 16580 25970 16596 26004
rect 16664 25970 16680 26004
rect 16738 25970 16754 26004
rect 16822 25970 16838 26004
rect 15316 25862 15332 25896
rect 15400 25862 15416 25896
rect 15474 25862 15490 25896
rect 15558 25862 15574 25896
rect 15632 25862 15648 25896
rect 15716 25862 15732 25896
rect 15790 25862 15806 25896
rect 15874 25862 15890 25896
rect 15948 25862 15964 25896
rect 16032 25862 16048 25896
rect 16106 25862 16122 25896
rect 16190 25862 16206 25896
rect 16264 25862 16280 25896
rect 16348 25862 16364 25896
rect 16422 25862 16438 25896
rect 16506 25862 16522 25896
rect 16580 25862 16596 25896
rect 16664 25862 16680 25896
rect 16738 25862 16754 25896
rect 16822 25862 16838 25896
rect 15270 25803 15304 25819
rect 15270 25411 15304 25427
rect 15428 25803 15462 25819
rect 15428 25411 15462 25427
rect 15586 25803 15620 25819
rect 15586 25411 15620 25427
rect 15744 25803 15778 25819
rect 15744 25411 15778 25427
rect 15902 25803 15936 25819
rect 15902 25411 15936 25427
rect 16060 25803 16094 25819
rect 16060 25411 16094 25427
rect 16218 25803 16252 25819
rect 16218 25411 16252 25427
rect 16376 25803 16410 25819
rect 16376 25411 16410 25427
rect 16534 25803 16568 25819
rect 16534 25411 16568 25427
rect 16692 25803 16726 25819
rect 16692 25411 16726 25427
rect 16850 25803 16884 25819
rect 16850 25411 16884 25427
rect 15316 25334 15332 25368
rect 15400 25334 15416 25368
rect 15474 25334 15490 25368
rect 15558 25334 15574 25368
rect 15632 25334 15648 25368
rect 15716 25334 15732 25368
rect 15790 25334 15806 25368
rect 15874 25334 15890 25368
rect 15948 25334 15964 25368
rect 16032 25334 16048 25368
rect 16106 25334 16122 25368
rect 16190 25334 16206 25368
rect 16264 25334 16280 25368
rect 16348 25334 16364 25368
rect 16422 25334 16438 25368
rect 16506 25334 16522 25368
rect 16580 25334 16596 25368
rect 16664 25334 16680 25368
rect 16738 25334 16754 25368
rect 16822 25334 16838 25368
rect 15156 25266 15190 25328
rect 16964 25266 16998 25328
rect 15156 25232 15252 25266
rect 16902 25232 16998 25266
rect 7340 25174 7440 25232
rect 9000 25174 9100 25232
rect 11140 25174 11240 25232
rect 13140 25174 13240 25232
rect 15300 25174 15400 25232
rect 18196 25182 18292 25216
rect 18642 25182 18738 25216
rect 19060 25196 19220 25296
rect 6376 25140 6472 25174
rect 7982 25140 8078 25174
rect 6376 25078 6410 25140
rect 8044 25078 8078 25140
rect 6522 25038 6538 25072
rect 6572 25038 6588 25072
rect 6714 25038 6730 25072
rect 6764 25038 6780 25072
rect 6906 25038 6922 25072
rect 6956 25038 6972 25072
rect 7098 25038 7114 25072
rect 7148 25038 7164 25072
rect 7290 25038 7306 25072
rect 7340 25038 7356 25072
rect 7482 25038 7498 25072
rect 7532 25038 7548 25072
rect 7674 25038 7690 25072
rect 7724 25038 7740 25072
rect 7866 25038 7882 25072
rect 7916 25038 7932 25072
rect 6490 24979 6524 24995
rect 6490 24587 6524 24603
rect 6586 24979 6620 24995
rect 6586 24587 6620 24603
rect 6682 24979 6716 24995
rect 6682 24587 6716 24603
rect 6778 24979 6812 24995
rect 6778 24587 6812 24603
rect 6874 24979 6908 24995
rect 6874 24587 6908 24603
rect 6970 24979 7004 24995
rect 6970 24587 7004 24603
rect 7066 24979 7100 24995
rect 7066 24587 7100 24603
rect 7162 24979 7196 24995
rect 7162 24587 7196 24603
rect 7258 24979 7292 24995
rect 7258 24587 7292 24603
rect 7354 24979 7388 24995
rect 7354 24587 7388 24603
rect 7450 24979 7484 24995
rect 7450 24587 7484 24603
rect 7546 24979 7580 24995
rect 7546 24587 7580 24603
rect 7642 24979 7676 24995
rect 7642 24587 7676 24603
rect 7738 24979 7772 24995
rect 7738 24587 7772 24603
rect 7834 24979 7868 24995
rect 7834 24587 7868 24603
rect 7930 24979 7964 24995
rect 7930 24587 7964 24603
rect 6618 24510 6634 24544
rect 6668 24510 6684 24544
rect 6810 24510 6826 24544
rect 6860 24510 6876 24544
rect 7002 24510 7018 24544
rect 7052 24510 7068 24544
rect 7194 24510 7210 24544
rect 7244 24510 7260 24544
rect 7386 24510 7402 24544
rect 7436 24510 7452 24544
rect 7578 24510 7594 24544
rect 7628 24510 7644 24544
rect 7770 24510 7786 24544
rect 7820 24510 7836 24544
rect 6618 24402 6634 24436
rect 6668 24402 6684 24436
rect 6810 24402 6826 24436
rect 6860 24402 6876 24436
rect 7002 24402 7018 24436
rect 7052 24402 7068 24436
rect 7194 24402 7210 24436
rect 7244 24402 7260 24436
rect 7386 24402 7402 24436
rect 7436 24402 7452 24436
rect 7578 24402 7594 24436
rect 7628 24402 7644 24436
rect 7770 24402 7786 24436
rect 7820 24402 7836 24436
rect 6490 24343 6524 24359
rect 6490 23951 6524 23967
rect 6586 24343 6620 24359
rect 6586 23951 6620 23967
rect 6682 24343 6716 24359
rect 6682 23951 6716 23967
rect 6778 24343 6812 24359
rect 6778 23951 6812 23967
rect 6874 24343 6908 24359
rect 6874 23951 6908 23967
rect 6970 24343 7004 24359
rect 6970 23951 7004 23967
rect 7066 24343 7100 24359
rect 7066 23951 7100 23967
rect 7162 24343 7196 24359
rect 7162 23951 7196 23967
rect 7258 24343 7292 24359
rect 7258 23951 7292 23967
rect 7354 24343 7388 24359
rect 7354 23951 7388 23967
rect 7450 24343 7484 24359
rect 7450 23951 7484 23967
rect 7546 24343 7580 24359
rect 7546 23951 7580 23967
rect 7642 24343 7676 24359
rect 7642 23951 7676 23967
rect 7738 24343 7772 24359
rect 7738 23951 7772 23967
rect 7834 24343 7868 24359
rect 7834 23951 7868 23967
rect 7930 24343 7964 24359
rect 7930 23951 7964 23967
rect 6522 23874 6538 23908
rect 6572 23874 6588 23908
rect 6714 23874 6730 23908
rect 6764 23874 6780 23908
rect 6906 23874 6922 23908
rect 6956 23874 6972 23908
rect 7098 23874 7114 23908
rect 7148 23874 7164 23908
rect 7290 23874 7306 23908
rect 7340 23874 7356 23908
rect 7482 23874 7498 23908
rect 7532 23874 7548 23908
rect 7674 23874 7690 23908
rect 7724 23874 7740 23908
rect 7866 23874 7882 23908
rect 7916 23874 7932 23908
rect 6376 23806 6410 23868
rect 8044 23806 8078 23868
rect 6376 23772 6472 23806
rect 7982 23772 8078 23806
rect 8596 25140 8692 25174
rect 10202 25140 10298 25174
rect 8596 25078 8630 25140
rect 10264 25078 10298 25140
rect 8742 25038 8758 25072
rect 8792 25038 8808 25072
rect 8934 25038 8950 25072
rect 8984 25038 9000 25072
rect 9126 25038 9142 25072
rect 9176 25038 9192 25072
rect 9318 25038 9334 25072
rect 9368 25038 9384 25072
rect 9510 25038 9526 25072
rect 9560 25038 9576 25072
rect 9702 25038 9718 25072
rect 9752 25038 9768 25072
rect 9894 25038 9910 25072
rect 9944 25038 9960 25072
rect 10086 25038 10102 25072
rect 10136 25038 10152 25072
rect 8710 24979 8744 24995
rect 8710 24587 8744 24603
rect 8806 24979 8840 24995
rect 8806 24587 8840 24603
rect 8902 24979 8936 24995
rect 8902 24587 8936 24603
rect 8998 24979 9032 24995
rect 8998 24587 9032 24603
rect 9094 24979 9128 24995
rect 9094 24587 9128 24603
rect 9190 24979 9224 24995
rect 9190 24587 9224 24603
rect 9286 24979 9320 24995
rect 9286 24587 9320 24603
rect 9382 24979 9416 24995
rect 9382 24587 9416 24603
rect 9478 24979 9512 24995
rect 9478 24587 9512 24603
rect 9574 24979 9608 24995
rect 9574 24587 9608 24603
rect 9670 24979 9704 24995
rect 9670 24587 9704 24603
rect 9766 24979 9800 24995
rect 9766 24587 9800 24603
rect 9862 24979 9896 24995
rect 9862 24587 9896 24603
rect 9958 24979 9992 24995
rect 9958 24587 9992 24603
rect 10054 24979 10088 24995
rect 10054 24587 10088 24603
rect 10150 24979 10184 24995
rect 10150 24587 10184 24603
rect 8838 24510 8854 24544
rect 8888 24510 8904 24544
rect 9030 24510 9046 24544
rect 9080 24510 9096 24544
rect 9222 24510 9238 24544
rect 9272 24510 9288 24544
rect 9414 24510 9430 24544
rect 9464 24510 9480 24544
rect 9606 24510 9622 24544
rect 9656 24510 9672 24544
rect 9798 24510 9814 24544
rect 9848 24510 9864 24544
rect 9990 24510 10006 24544
rect 10040 24510 10056 24544
rect 8838 24402 8854 24436
rect 8888 24402 8904 24436
rect 9030 24402 9046 24436
rect 9080 24402 9096 24436
rect 9222 24402 9238 24436
rect 9272 24402 9288 24436
rect 9414 24402 9430 24436
rect 9464 24402 9480 24436
rect 9606 24402 9622 24436
rect 9656 24402 9672 24436
rect 9798 24402 9814 24436
rect 9848 24402 9864 24436
rect 9990 24402 10006 24436
rect 10040 24402 10056 24436
rect 8710 24343 8744 24359
rect 8710 23951 8744 23967
rect 8806 24343 8840 24359
rect 8806 23951 8840 23967
rect 8902 24343 8936 24359
rect 8902 23951 8936 23967
rect 8998 24343 9032 24359
rect 8998 23951 9032 23967
rect 9094 24343 9128 24359
rect 9094 23951 9128 23967
rect 9190 24343 9224 24359
rect 9190 23951 9224 23967
rect 9286 24343 9320 24359
rect 9286 23951 9320 23967
rect 9382 24343 9416 24359
rect 9382 23951 9416 23967
rect 9478 24343 9512 24359
rect 9478 23951 9512 23967
rect 9574 24343 9608 24359
rect 9574 23951 9608 23967
rect 9670 24343 9704 24359
rect 9670 23951 9704 23967
rect 9766 24343 9800 24359
rect 9766 23951 9800 23967
rect 9862 24343 9896 24359
rect 9862 23951 9896 23967
rect 9958 24343 9992 24359
rect 9958 23951 9992 23967
rect 10054 24343 10088 24359
rect 10054 23951 10088 23967
rect 10150 24343 10184 24359
rect 10150 23951 10184 23967
rect 8742 23874 8758 23908
rect 8792 23874 8808 23908
rect 8934 23874 8950 23908
rect 8984 23874 9000 23908
rect 9126 23874 9142 23908
rect 9176 23874 9192 23908
rect 9318 23874 9334 23908
rect 9368 23874 9384 23908
rect 9510 23874 9526 23908
rect 9560 23874 9576 23908
rect 9702 23874 9718 23908
rect 9752 23874 9768 23908
rect 9894 23874 9910 23908
rect 9944 23874 9960 23908
rect 10086 23874 10102 23908
rect 10136 23874 10152 23908
rect 8596 23806 8630 23868
rect 10264 23806 10298 23868
rect 8596 23772 8692 23806
rect 10202 23772 10298 23806
rect 10776 25140 10872 25174
rect 12382 25140 12478 25174
rect 10776 25078 10810 25140
rect 12444 25078 12478 25140
rect 10922 25038 10938 25072
rect 10972 25038 10988 25072
rect 11114 25038 11130 25072
rect 11164 25038 11180 25072
rect 11306 25038 11322 25072
rect 11356 25038 11372 25072
rect 11498 25038 11514 25072
rect 11548 25038 11564 25072
rect 11690 25038 11706 25072
rect 11740 25038 11756 25072
rect 11882 25038 11898 25072
rect 11932 25038 11948 25072
rect 12074 25038 12090 25072
rect 12124 25038 12140 25072
rect 12266 25038 12282 25072
rect 12316 25038 12332 25072
rect 10890 24979 10924 24995
rect 10890 24587 10924 24603
rect 10986 24979 11020 24995
rect 10986 24587 11020 24603
rect 11082 24979 11116 24995
rect 11082 24587 11116 24603
rect 11178 24979 11212 24995
rect 11178 24587 11212 24603
rect 11274 24979 11308 24995
rect 11274 24587 11308 24603
rect 11370 24979 11404 24995
rect 11370 24587 11404 24603
rect 11466 24979 11500 24995
rect 11466 24587 11500 24603
rect 11562 24979 11596 24995
rect 11562 24587 11596 24603
rect 11658 24979 11692 24995
rect 11658 24587 11692 24603
rect 11754 24979 11788 24995
rect 11754 24587 11788 24603
rect 11850 24979 11884 24995
rect 11850 24587 11884 24603
rect 11946 24979 11980 24995
rect 11946 24587 11980 24603
rect 12042 24979 12076 24995
rect 12042 24587 12076 24603
rect 12138 24979 12172 24995
rect 12138 24587 12172 24603
rect 12234 24979 12268 24995
rect 12234 24587 12268 24603
rect 12330 24979 12364 24995
rect 12330 24587 12364 24603
rect 11018 24510 11034 24544
rect 11068 24510 11084 24544
rect 11210 24510 11226 24544
rect 11260 24510 11276 24544
rect 11402 24510 11418 24544
rect 11452 24510 11468 24544
rect 11594 24510 11610 24544
rect 11644 24510 11660 24544
rect 11786 24510 11802 24544
rect 11836 24510 11852 24544
rect 11978 24510 11994 24544
rect 12028 24510 12044 24544
rect 12170 24510 12186 24544
rect 12220 24510 12236 24544
rect 11018 24402 11034 24436
rect 11068 24402 11084 24436
rect 11210 24402 11226 24436
rect 11260 24402 11276 24436
rect 11402 24402 11418 24436
rect 11452 24402 11468 24436
rect 11594 24402 11610 24436
rect 11644 24402 11660 24436
rect 11786 24402 11802 24436
rect 11836 24402 11852 24436
rect 11978 24402 11994 24436
rect 12028 24402 12044 24436
rect 12170 24402 12186 24436
rect 12220 24402 12236 24436
rect 10890 24343 10924 24359
rect 10890 23951 10924 23967
rect 10986 24343 11020 24359
rect 10986 23951 11020 23967
rect 11082 24343 11116 24359
rect 11082 23951 11116 23967
rect 11178 24343 11212 24359
rect 11178 23951 11212 23967
rect 11274 24343 11308 24359
rect 11274 23951 11308 23967
rect 11370 24343 11404 24359
rect 11370 23951 11404 23967
rect 11466 24343 11500 24359
rect 11466 23951 11500 23967
rect 11562 24343 11596 24359
rect 11562 23951 11596 23967
rect 11658 24343 11692 24359
rect 11658 23951 11692 23967
rect 11754 24343 11788 24359
rect 11754 23951 11788 23967
rect 11850 24343 11884 24359
rect 11850 23951 11884 23967
rect 11946 24343 11980 24359
rect 11946 23951 11980 23967
rect 12042 24343 12076 24359
rect 12042 23951 12076 23967
rect 12138 24343 12172 24359
rect 12138 23951 12172 23967
rect 12234 24343 12268 24359
rect 12234 23951 12268 23967
rect 12330 24343 12364 24359
rect 12330 23951 12364 23967
rect 10922 23874 10938 23908
rect 10972 23874 10988 23908
rect 11114 23874 11130 23908
rect 11164 23874 11180 23908
rect 11306 23874 11322 23908
rect 11356 23874 11372 23908
rect 11498 23874 11514 23908
rect 11548 23874 11564 23908
rect 11690 23874 11706 23908
rect 11740 23874 11756 23908
rect 11882 23874 11898 23908
rect 11932 23874 11948 23908
rect 12074 23874 12090 23908
rect 12124 23874 12140 23908
rect 12266 23874 12282 23908
rect 12316 23874 12332 23908
rect 10776 23806 10810 23868
rect 12444 23806 12478 23868
rect 10776 23772 10872 23806
rect 12382 23772 12478 23806
rect 12956 25140 13052 25174
rect 14562 25140 14658 25174
rect 12956 25078 12990 25140
rect 14624 25078 14658 25140
rect 13102 25038 13118 25072
rect 13152 25038 13168 25072
rect 13294 25038 13310 25072
rect 13344 25038 13360 25072
rect 13486 25038 13502 25072
rect 13536 25038 13552 25072
rect 13678 25038 13694 25072
rect 13728 25038 13744 25072
rect 13870 25038 13886 25072
rect 13920 25038 13936 25072
rect 14062 25038 14078 25072
rect 14112 25038 14128 25072
rect 14254 25038 14270 25072
rect 14304 25038 14320 25072
rect 14446 25038 14462 25072
rect 14496 25038 14512 25072
rect 13070 24979 13104 24995
rect 13070 24587 13104 24603
rect 13166 24979 13200 24995
rect 13166 24587 13200 24603
rect 13262 24979 13296 24995
rect 13262 24587 13296 24603
rect 13358 24979 13392 24995
rect 13358 24587 13392 24603
rect 13454 24979 13488 24995
rect 13454 24587 13488 24603
rect 13550 24979 13584 24995
rect 13550 24587 13584 24603
rect 13646 24979 13680 24995
rect 13646 24587 13680 24603
rect 13742 24979 13776 24995
rect 13742 24587 13776 24603
rect 13838 24979 13872 24995
rect 13838 24587 13872 24603
rect 13934 24979 13968 24995
rect 13934 24587 13968 24603
rect 14030 24979 14064 24995
rect 14030 24587 14064 24603
rect 14126 24979 14160 24995
rect 14126 24587 14160 24603
rect 14222 24979 14256 24995
rect 14222 24587 14256 24603
rect 14318 24979 14352 24995
rect 14318 24587 14352 24603
rect 14414 24979 14448 24995
rect 14414 24587 14448 24603
rect 14510 24979 14544 24995
rect 14510 24587 14544 24603
rect 13198 24510 13214 24544
rect 13248 24510 13264 24544
rect 13390 24510 13406 24544
rect 13440 24510 13456 24544
rect 13582 24510 13598 24544
rect 13632 24510 13648 24544
rect 13774 24510 13790 24544
rect 13824 24510 13840 24544
rect 13966 24510 13982 24544
rect 14016 24510 14032 24544
rect 14158 24510 14174 24544
rect 14208 24510 14224 24544
rect 14350 24510 14366 24544
rect 14400 24510 14416 24544
rect 13198 24402 13214 24436
rect 13248 24402 13264 24436
rect 13390 24402 13406 24436
rect 13440 24402 13456 24436
rect 13582 24402 13598 24436
rect 13632 24402 13648 24436
rect 13774 24402 13790 24436
rect 13824 24402 13840 24436
rect 13966 24402 13982 24436
rect 14016 24402 14032 24436
rect 14158 24402 14174 24436
rect 14208 24402 14224 24436
rect 14350 24402 14366 24436
rect 14400 24402 14416 24436
rect 13070 24343 13104 24359
rect 13070 23951 13104 23967
rect 13166 24343 13200 24359
rect 13166 23951 13200 23967
rect 13262 24343 13296 24359
rect 13262 23951 13296 23967
rect 13358 24343 13392 24359
rect 13358 23951 13392 23967
rect 13454 24343 13488 24359
rect 13454 23951 13488 23967
rect 13550 24343 13584 24359
rect 13550 23951 13584 23967
rect 13646 24343 13680 24359
rect 13646 23951 13680 23967
rect 13742 24343 13776 24359
rect 13742 23951 13776 23967
rect 13838 24343 13872 24359
rect 13838 23951 13872 23967
rect 13934 24343 13968 24359
rect 13934 23951 13968 23967
rect 14030 24343 14064 24359
rect 14030 23951 14064 23967
rect 14126 24343 14160 24359
rect 14126 23951 14160 23967
rect 14222 24343 14256 24359
rect 14222 23951 14256 23967
rect 14318 24343 14352 24359
rect 14318 23951 14352 23967
rect 14414 24343 14448 24359
rect 14414 23951 14448 23967
rect 14510 24343 14544 24359
rect 14510 23951 14544 23967
rect 13102 23874 13118 23908
rect 13152 23874 13168 23908
rect 13294 23874 13310 23908
rect 13344 23874 13360 23908
rect 13486 23874 13502 23908
rect 13536 23874 13552 23908
rect 13678 23874 13694 23908
rect 13728 23874 13744 23908
rect 13870 23874 13886 23908
rect 13920 23874 13936 23908
rect 14062 23874 14078 23908
rect 14112 23874 14128 23908
rect 14254 23874 14270 23908
rect 14304 23874 14320 23908
rect 14446 23874 14462 23908
rect 14496 23874 14512 23908
rect 12956 23806 12990 23868
rect 14624 23806 14658 23868
rect 12956 23772 13052 23806
rect 14562 23772 14658 23806
rect 15156 25140 15252 25174
rect 16762 25140 16858 25174
rect 15156 25078 15190 25140
rect 16824 25078 16858 25140
rect 15302 25038 15318 25072
rect 15352 25038 15368 25072
rect 15494 25038 15510 25072
rect 15544 25038 15560 25072
rect 15686 25038 15702 25072
rect 15736 25038 15752 25072
rect 15878 25038 15894 25072
rect 15928 25038 15944 25072
rect 16070 25038 16086 25072
rect 16120 25038 16136 25072
rect 16262 25038 16278 25072
rect 16312 25038 16328 25072
rect 16454 25038 16470 25072
rect 16504 25038 16520 25072
rect 16646 25038 16662 25072
rect 16696 25038 16712 25072
rect 15270 24979 15304 24995
rect 15270 24587 15304 24603
rect 15366 24979 15400 24995
rect 15366 24587 15400 24603
rect 15462 24979 15496 24995
rect 15462 24587 15496 24603
rect 15558 24979 15592 24995
rect 15558 24587 15592 24603
rect 15654 24979 15688 24995
rect 15654 24587 15688 24603
rect 15750 24979 15784 24995
rect 15750 24587 15784 24603
rect 15846 24979 15880 24995
rect 15846 24587 15880 24603
rect 15942 24979 15976 24995
rect 15942 24587 15976 24603
rect 16038 24979 16072 24995
rect 16038 24587 16072 24603
rect 16134 24979 16168 24995
rect 16134 24587 16168 24603
rect 16230 24979 16264 24995
rect 16230 24587 16264 24603
rect 16326 24979 16360 24995
rect 16326 24587 16360 24603
rect 16422 24979 16456 24995
rect 16422 24587 16456 24603
rect 16518 24979 16552 24995
rect 16518 24587 16552 24603
rect 16614 24979 16648 24995
rect 16614 24587 16648 24603
rect 16710 24979 16744 24995
rect 16710 24587 16744 24603
rect 15398 24510 15414 24544
rect 15448 24510 15464 24544
rect 15590 24510 15606 24544
rect 15640 24510 15656 24544
rect 15782 24510 15798 24544
rect 15832 24510 15848 24544
rect 15974 24510 15990 24544
rect 16024 24510 16040 24544
rect 16166 24510 16182 24544
rect 16216 24510 16232 24544
rect 16358 24510 16374 24544
rect 16408 24510 16424 24544
rect 16550 24510 16566 24544
rect 16600 24510 16616 24544
rect 15398 24402 15414 24436
rect 15448 24402 15464 24436
rect 15590 24402 15606 24436
rect 15640 24402 15656 24436
rect 15782 24402 15798 24436
rect 15832 24402 15848 24436
rect 15974 24402 15990 24436
rect 16024 24402 16040 24436
rect 16166 24402 16182 24436
rect 16216 24402 16232 24436
rect 16358 24402 16374 24436
rect 16408 24402 16424 24436
rect 16550 24402 16566 24436
rect 16600 24402 16616 24436
rect 15270 24343 15304 24359
rect 15270 23951 15304 23967
rect 15366 24343 15400 24359
rect 15366 23951 15400 23967
rect 15462 24343 15496 24359
rect 15462 23951 15496 23967
rect 15558 24343 15592 24359
rect 15558 23951 15592 23967
rect 15654 24343 15688 24359
rect 15654 23951 15688 23967
rect 15750 24343 15784 24359
rect 15750 23951 15784 23967
rect 15846 24343 15880 24359
rect 15846 23951 15880 23967
rect 15942 24343 15976 24359
rect 15942 23951 15976 23967
rect 16038 24343 16072 24359
rect 16038 23951 16072 23967
rect 16134 24343 16168 24359
rect 16134 23951 16168 23967
rect 16230 24343 16264 24359
rect 16230 23951 16264 23967
rect 16326 24343 16360 24359
rect 16326 23951 16360 23967
rect 16422 24343 16456 24359
rect 16422 23951 16456 23967
rect 16518 24343 16552 24359
rect 16518 23951 16552 23967
rect 16614 24343 16648 24359
rect 16614 23951 16648 23967
rect 16710 24343 16744 24359
rect 16710 23951 16744 23967
rect 15302 23874 15318 23908
rect 15352 23874 15368 23908
rect 15494 23874 15510 23908
rect 15544 23874 15560 23908
rect 15686 23874 15702 23908
rect 15736 23874 15752 23908
rect 15878 23874 15894 23908
rect 15928 23874 15944 23908
rect 16070 23874 16086 23908
rect 16120 23874 16136 23908
rect 16262 23874 16278 23908
rect 16312 23874 16328 23908
rect 16454 23874 16470 23908
rect 16504 23874 16520 23908
rect 16646 23874 16662 23908
rect 16696 23874 16712 23908
rect 15156 23806 15190 23868
rect 16824 23806 16858 23868
rect 15156 23772 15252 23806
rect 16762 23772 16858 23806
rect 18196 25120 18230 25182
rect 6496 23562 6592 23596
rect 7622 23562 7718 23596
rect 6496 23500 6530 23562
rect 7684 23500 7718 23562
rect 6738 23460 6754 23494
rect 6788 23460 6804 23494
rect 6930 23460 6946 23494
rect 6980 23460 6996 23494
rect 7122 23460 7138 23494
rect 7172 23460 7188 23494
rect 7314 23460 7330 23494
rect 7364 23460 7380 23494
rect 7506 23460 7522 23494
rect 7556 23460 7572 23494
rect 6610 23410 6644 23426
rect 6610 23018 6644 23034
rect 6706 23410 6740 23426
rect 6706 23018 6740 23034
rect 6802 23410 6836 23426
rect 6802 23018 6836 23034
rect 6898 23410 6932 23426
rect 6898 23018 6932 23034
rect 6994 23410 7028 23426
rect 6994 23018 7028 23034
rect 7090 23410 7124 23426
rect 7090 23018 7124 23034
rect 7186 23410 7220 23426
rect 7186 23018 7220 23034
rect 7282 23410 7316 23426
rect 7282 23018 7316 23034
rect 7378 23410 7412 23426
rect 7378 23018 7412 23034
rect 7474 23410 7508 23426
rect 7474 23018 7508 23034
rect 7570 23410 7604 23426
rect 7570 23018 7604 23034
rect 6642 22950 6658 22984
rect 6692 22950 6708 22984
rect 6834 22950 6850 22984
rect 6884 22950 6900 22984
rect 7026 22950 7042 22984
rect 7076 22950 7092 22984
rect 7218 22950 7234 22984
rect 7268 22950 7284 22984
rect 7410 22950 7426 22984
rect 7460 22950 7476 22984
rect 6642 22842 6658 22876
rect 6692 22842 6708 22876
rect 6834 22842 6850 22876
rect 6884 22842 6900 22876
rect 7026 22842 7042 22876
rect 7076 22842 7092 22876
rect 7218 22842 7234 22876
rect 7268 22842 7284 22876
rect 7410 22842 7426 22876
rect 7460 22842 7476 22876
rect 6610 22792 6644 22808
rect 6610 22400 6644 22416
rect 6706 22792 6740 22808
rect 6706 22400 6740 22416
rect 6802 22792 6836 22808
rect 6802 22400 6836 22416
rect 6898 22792 6932 22808
rect 6898 22400 6932 22416
rect 6994 22792 7028 22808
rect 6994 22400 7028 22416
rect 7090 22792 7124 22808
rect 7090 22400 7124 22416
rect 7186 22792 7220 22808
rect 7186 22400 7220 22416
rect 7282 22792 7316 22808
rect 7282 22400 7316 22416
rect 7378 22792 7412 22808
rect 7378 22400 7412 22416
rect 7474 22792 7508 22808
rect 7474 22400 7508 22416
rect 7570 22792 7604 22808
rect 7570 22400 7604 22416
rect 6738 22332 6754 22366
rect 6788 22332 6804 22366
rect 6930 22332 6946 22366
rect 6980 22332 6996 22366
rect 7122 22332 7138 22366
rect 7172 22332 7188 22366
rect 7314 22332 7330 22366
rect 7364 22332 7380 22366
rect 7506 22332 7522 22366
rect 7556 22332 7572 22366
rect 6738 22224 6754 22258
rect 6788 22224 6804 22258
rect 6930 22224 6946 22258
rect 6980 22224 6996 22258
rect 7122 22224 7138 22258
rect 7172 22224 7188 22258
rect 7314 22224 7330 22258
rect 7364 22224 7380 22258
rect 7506 22224 7522 22258
rect 7556 22224 7572 22258
rect 6610 22174 6644 22190
rect 6610 21782 6644 21798
rect 6706 22174 6740 22190
rect 6706 21782 6740 21798
rect 6802 22174 6836 22190
rect 6802 21782 6836 21798
rect 6898 22174 6932 22190
rect 6898 21782 6932 21798
rect 6994 22174 7028 22190
rect 6994 21782 7028 21798
rect 7090 22174 7124 22190
rect 7090 21782 7124 21798
rect 7186 22174 7220 22190
rect 7186 21782 7220 21798
rect 7282 22174 7316 22190
rect 7282 21782 7316 21798
rect 7378 22174 7412 22190
rect 7378 21782 7412 21798
rect 7474 22174 7508 22190
rect 7474 21782 7508 21798
rect 7570 22174 7604 22190
rect 7570 21782 7604 21798
rect 6642 21714 6658 21748
rect 6692 21714 6708 21748
rect 6834 21714 6850 21748
rect 6884 21714 6900 21748
rect 7026 21714 7042 21748
rect 7076 21714 7092 21748
rect 7218 21714 7234 21748
rect 7268 21714 7284 21748
rect 7410 21714 7426 21748
rect 7460 21714 7476 21748
rect 6496 21646 6530 21708
rect 7684 21646 7718 21708
rect 6496 21612 6592 21646
rect 7622 21612 7718 21646
rect 8216 23562 8312 23596
rect 9342 23562 9438 23596
rect 8216 23500 8250 23562
rect 9404 23500 9438 23562
rect 8458 23460 8474 23494
rect 8508 23460 8524 23494
rect 8650 23460 8666 23494
rect 8700 23460 8716 23494
rect 8842 23460 8858 23494
rect 8892 23460 8908 23494
rect 9034 23460 9050 23494
rect 9084 23460 9100 23494
rect 9226 23460 9242 23494
rect 9276 23460 9292 23494
rect 8330 23410 8364 23426
rect 8330 23018 8364 23034
rect 8426 23410 8460 23426
rect 8426 23018 8460 23034
rect 8522 23410 8556 23426
rect 8522 23018 8556 23034
rect 8618 23410 8652 23426
rect 8618 23018 8652 23034
rect 8714 23410 8748 23426
rect 8714 23018 8748 23034
rect 8810 23410 8844 23426
rect 8810 23018 8844 23034
rect 8906 23410 8940 23426
rect 8906 23018 8940 23034
rect 9002 23410 9036 23426
rect 9002 23018 9036 23034
rect 9098 23410 9132 23426
rect 9098 23018 9132 23034
rect 9194 23410 9228 23426
rect 9194 23018 9228 23034
rect 9290 23410 9324 23426
rect 9290 23018 9324 23034
rect 8362 22950 8378 22984
rect 8412 22950 8428 22984
rect 8554 22950 8570 22984
rect 8604 22950 8620 22984
rect 8746 22950 8762 22984
rect 8796 22950 8812 22984
rect 8938 22950 8954 22984
rect 8988 22950 9004 22984
rect 9130 22950 9146 22984
rect 9180 22950 9196 22984
rect 8362 22842 8378 22876
rect 8412 22842 8428 22876
rect 8554 22842 8570 22876
rect 8604 22842 8620 22876
rect 8746 22842 8762 22876
rect 8796 22842 8812 22876
rect 8938 22842 8954 22876
rect 8988 22842 9004 22876
rect 9130 22842 9146 22876
rect 9180 22842 9196 22876
rect 8330 22792 8364 22808
rect 8330 22400 8364 22416
rect 8426 22792 8460 22808
rect 8426 22400 8460 22416
rect 8522 22792 8556 22808
rect 8522 22400 8556 22416
rect 8618 22792 8652 22808
rect 8618 22400 8652 22416
rect 8714 22792 8748 22808
rect 8714 22400 8748 22416
rect 8810 22792 8844 22808
rect 8810 22400 8844 22416
rect 8906 22792 8940 22808
rect 8906 22400 8940 22416
rect 9002 22792 9036 22808
rect 9002 22400 9036 22416
rect 9098 22792 9132 22808
rect 9098 22400 9132 22416
rect 9194 22792 9228 22808
rect 9194 22400 9228 22416
rect 9290 22792 9324 22808
rect 9290 22400 9324 22416
rect 8458 22332 8474 22366
rect 8508 22332 8524 22366
rect 8650 22332 8666 22366
rect 8700 22332 8716 22366
rect 8842 22332 8858 22366
rect 8892 22332 8908 22366
rect 9034 22332 9050 22366
rect 9084 22332 9100 22366
rect 9226 22332 9242 22366
rect 9276 22332 9292 22366
rect 8458 22224 8474 22258
rect 8508 22224 8524 22258
rect 8650 22224 8666 22258
rect 8700 22224 8716 22258
rect 8842 22224 8858 22258
rect 8892 22224 8908 22258
rect 9034 22224 9050 22258
rect 9084 22224 9100 22258
rect 9226 22224 9242 22258
rect 9276 22224 9292 22258
rect 8330 22174 8364 22190
rect 8330 21782 8364 21798
rect 8426 22174 8460 22190
rect 8426 21782 8460 21798
rect 8522 22174 8556 22190
rect 8522 21782 8556 21798
rect 8618 22174 8652 22190
rect 8618 21782 8652 21798
rect 8714 22174 8748 22190
rect 8714 21782 8748 21798
rect 8810 22174 8844 22190
rect 8810 21782 8844 21798
rect 8906 22174 8940 22190
rect 8906 21782 8940 21798
rect 9002 22174 9036 22190
rect 9002 21782 9036 21798
rect 9098 22174 9132 22190
rect 9098 21782 9132 21798
rect 9194 22174 9228 22190
rect 9194 21782 9228 21798
rect 9290 22174 9324 22190
rect 9290 21782 9324 21798
rect 8362 21714 8378 21748
rect 8412 21714 8428 21748
rect 8554 21714 8570 21748
rect 8604 21714 8620 21748
rect 8746 21714 8762 21748
rect 8796 21714 8812 21748
rect 8938 21714 8954 21748
rect 8988 21714 9004 21748
rect 9130 21714 9146 21748
rect 9180 21714 9196 21748
rect 8216 21646 8250 21708
rect 18060 23388 18196 23396
rect 18704 25120 18738 25182
rect 18060 23326 18230 23388
rect 18704 23326 18738 23388
rect 18060 23296 18292 23326
rect 18060 22376 18140 23296
rect 18196 23292 18292 23296
rect 18642 23292 18738 23326
rect 18856 25162 18952 25196
rect 19326 25162 19422 25196
rect 18856 25100 18890 25162
rect 19388 25100 19422 25162
rect 19035 25048 19051 25082
rect 19227 25048 19243 25082
rect 18958 25020 18992 25036
rect 18958 23436 18992 23452
rect 19286 25020 19320 25036
rect 19286 23436 19320 23452
rect 19035 23390 19051 23424
rect 19227 23390 19243 23424
rect 18856 23310 18890 23372
rect 19388 23310 19422 23372
rect 18856 23276 18952 23310
rect 19326 23276 19422 23310
rect 19080 23206 19200 23276
rect 18196 23172 18292 23206
rect 19322 23172 19418 23206
rect 18196 23110 18230 23172
rect 19384 23110 19418 23172
rect 18438 23070 18454 23104
rect 18488 23070 18504 23104
rect 18630 23070 18646 23104
rect 18680 23070 18696 23104
rect 18822 23070 18838 23104
rect 18872 23070 18888 23104
rect 19014 23070 19030 23104
rect 19064 23070 19080 23104
rect 19206 23070 19222 23104
rect 19256 23070 19272 23104
rect 18310 23011 18344 23027
rect 18310 22619 18344 22635
rect 18406 23011 18440 23027
rect 18406 22619 18440 22635
rect 18502 23011 18536 23027
rect 18502 22619 18536 22635
rect 18598 23011 18632 23027
rect 18598 22619 18632 22635
rect 18694 23011 18728 23027
rect 18694 22619 18728 22635
rect 18790 23011 18824 23027
rect 18790 22619 18824 22635
rect 18886 23011 18920 23027
rect 18886 22619 18920 22635
rect 18982 23011 19016 23027
rect 18982 22619 19016 22635
rect 19078 23011 19112 23027
rect 19078 22619 19112 22635
rect 19174 23011 19208 23027
rect 19174 22619 19208 22635
rect 19270 23011 19304 23027
rect 19270 22619 19304 22635
rect 18342 22542 18358 22576
rect 18392 22542 18408 22576
rect 18534 22542 18550 22576
rect 18584 22542 18600 22576
rect 18726 22542 18742 22576
rect 18776 22542 18792 22576
rect 18918 22542 18934 22576
rect 18968 22542 18984 22576
rect 19110 22542 19126 22576
rect 19160 22542 19176 22576
rect 18196 22474 18230 22536
rect 19384 22474 19418 22536
rect 18196 22440 18292 22474
rect 19322 22440 19418 22474
rect 18060 22338 18200 22376
rect 18060 22304 18292 22338
rect 19322 22304 19418 22338
rect 18060 22242 18230 22304
rect 18060 22176 18196 22242
rect 9404 21646 9438 21708
rect 8216 21612 8312 21646
rect 9342 21612 9438 21646
rect 6500 21450 6660 21612
rect 8220 21450 8380 21612
rect 6496 21416 6592 21450
rect 7952 21416 8048 21450
rect 6496 21354 6530 21416
rect 8014 21354 8048 21416
rect 6656 21314 6672 21348
rect 6840 21314 6856 21348
rect 6914 21314 6930 21348
rect 7098 21314 7114 21348
rect 7172 21314 7188 21348
rect 7356 21314 7372 21348
rect 7430 21314 7446 21348
rect 7614 21314 7630 21348
rect 7688 21314 7704 21348
rect 7872 21314 7888 21348
rect 6610 21264 6644 21280
rect 6610 20872 6644 20888
rect 6868 21264 6902 21280
rect 6868 20872 6902 20888
rect 7126 21264 7160 21280
rect 7126 20872 7160 20888
rect 7384 21264 7418 21280
rect 7384 20872 7418 20888
rect 7642 21264 7676 21280
rect 7642 20872 7676 20888
rect 7900 21264 7934 21280
rect 7900 20872 7934 20888
rect 6656 20804 6672 20838
rect 6840 20804 6856 20838
rect 6914 20804 6930 20838
rect 7098 20804 7114 20838
rect 7172 20804 7188 20838
rect 7356 20804 7372 20838
rect 7430 20804 7446 20838
rect 7614 20804 7630 20838
rect 7688 20804 7704 20838
rect 7872 20804 7888 20838
rect 6656 20696 6672 20730
rect 6840 20696 6856 20730
rect 6914 20696 6930 20730
rect 7098 20696 7114 20730
rect 7172 20696 7188 20730
rect 7356 20696 7372 20730
rect 7430 20696 7446 20730
rect 7614 20696 7630 20730
rect 7688 20696 7704 20730
rect 7872 20696 7888 20730
rect 6610 20646 6644 20662
rect 6610 20254 6644 20270
rect 6868 20646 6902 20662
rect 6868 20254 6902 20270
rect 7126 20646 7160 20662
rect 7126 20254 7160 20270
rect 7384 20646 7418 20662
rect 7384 20254 7418 20270
rect 7642 20646 7676 20662
rect 7642 20254 7676 20270
rect 7900 20646 7934 20662
rect 7900 20254 7934 20270
rect 6656 20186 6672 20220
rect 6840 20186 6856 20220
rect 6914 20186 6930 20220
rect 7098 20186 7114 20220
rect 7172 20186 7188 20220
rect 7356 20186 7372 20220
rect 7430 20186 7446 20220
rect 7614 20186 7630 20220
rect 7688 20186 7704 20220
rect 7872 20186 7888 20220
rect 6656 20078 6672 20112
rect 6840 20078 6856 20112
rect 6914 20078 6930 20112
rect 7098 20078 7114 20112
rect 7172 20078 7188 20112
rect 7356 20078 7372 20112
rect 7430 20078 7446 20112
rect 7614 20078 7630 20112
rect 7688 20078 7704 20112
rect 7872 20078 7888 20112
rect 6610 20028 6644 20044
rect 6610 19636 6644 19652
rect 6868 20028 6902 20044
rect 6868 19636 6902 19652
rect 7126 20028 7160 20044
rect 7126 19636 7160 19652
rect 7384 20028 7418 20044
rect 7384 19636 7418 19652
rect 7642 20028 7676 20044
rect 7642 19636 7676 19652
rect 7900 20028 7934 20044
rect 7900 19636 7934 19652
rect 6656 19568 6672 19602
rect 6840 19568 6856 19602
rect 6914 19568 6930 19602
rect 7098 19568 7114 19602
rect 7172 19568 7188 19602
rect 7356 19568 7372 19602
rect 7430 19568 7446 19602
rect 7614 19568 7630 19602
rect 7688 19568 7704 19602
rect 7872 19568 7888 19602
rect 6656 19460 6672 19494
rect 6840 19460 6856 19494
rect 6914 19460 6930 19494
rect 7098 19460 7114 19494
rect 7172 19460 7188 19494
rect 7356 19460 7372 19494
rect 7430 19460 7446 19494
rect 7614 19460 7630 19494
rect 7688 19460 7704 19494
rect 7872 19460 7888 19494
rect 6610 19410 6644 19426
rect 6610 19018 6644 19034
rect 6868 19410 6902 19426
rect 6868 19018 6902 19034
rect 7126 19410 7160 19426
rect 7126 19018 7160 19034
rect 7384 19410 7418 19426
rect 7384 19018 7418 19034
rect 7642 19410 7676 19426
rect 7642 19018 7676 19034
rect 7900 19410 7934 19426
rect 7900 19018 7934 19034
rect 6656 18950 6672 18984
rect 6840 18950 6856 18984
rect 6914 18950 6930 18984
rect 7098 18950 7114 18984
rect 7172 18950 7188 18984
rect 7356 18950 7372 18984
rect 7430 18950 7446 18984
rect 7614 18950 7630 18984
rect 7688 18950 7704 18984
rect 7872 18950 7888 18984
rect 6656 18842 6672 18876
rect 6840 18842 6856 18876
rect 6914 18842 6930 18876
rect 7098 18842 7114 18876
rect 7172 18842 7188 18876
rect 7356 18842 7372 18876
rect 7430 18842 7446 18876
rect 7614 18842 7630 18876
rect 7688 18842 7704 18876
rect 7872 18842 7888 18876
rect 6610 18792 6644 18808
rect 6610 18400 6644 18416
rect 6868 18792 6902 18808
rect 6868 18400 6902 18416
rect 7126 18792 7160 18808
rect 7126 18400 7160 18416
rect 7384 18792 7418 18808
rect 7384 18400 7418 18416
rect 7642 18792 7676 18808
rect 7642 18400 7676 18416
rect 7900 18792 7934 18808
rect 7900 18400 7934 18416
rect 6656 18332 6672 18366
rect 6840 18332 6856 18366
rect 6914 18332 6930 18366
rect 7098 18332 7114 18366
rect 7172 18332 7188 18366
rect 7356 18332 7372 18366
rect 7430 18332 7446 18366
rect 7614 18332 7630 18366
rect 7688 18332 7704 18366
rect 7872 18332 7888 18366
rect 6656 18224 6672 18258
rect 6840 18224 6856 18258
rect 6914 18224 6930 18258
rect 7098 18224 7114 18258
rect 7172 18224 7188 18258
rect 7356 18224 7372 18258
rect 7430 18224 7446 18258
rect 7614 18224 7630 18258
rect 7688 18224 7704 18258
rect 7872 18224 7888 18258
rect 6610 18174 6644 18190
rect 6610 17782 6644 17798
rect 6868 18174 6902 18190
rect 6868 17782 6902 17798
rect 7126 18174 7160 18190
rect 7126 17782 7160 17798
rect 7384 18174 7418 18190
rect 7384 17782 7418 17798
rect 7642 18174 7676 18190
rect 7642 17782 7676 17798
rect 7900 18174 7934 18190
rect 7900 17782 7934 17798
rect 8216 21416 8312 21450
rect 9672 21416 9768 21450
rect 8216 21354 8250 21416
rect 9734 21354 9768 21416
rect 8376 21314 8392 21348
rect 8560 21314 8576 21348
rect 8634 21314 8650 21348
rect 8818 21314 8834 21348
rect 8892 21314 8908 21348
rect 9076 21314 9092 21348
rect 9150 21314 9166 21348
rect 9334 21314 9350 21348
rect 9408 21314 9424 21348
rect 9592 21314 9608 21348
rect 8330 21264 8364 21280
rect 8330 20872 8364 20888
rect 8588 21264 8622 21280
rect 8588 20872 8622 20888
rect 8846 21264 8880 21280
rect 8846 20872 8880 20888
rect 9104 21264 9138 21280
rect 9104 20872 9138 20888
rect 9362 21264 9396 21280
rect 9362 20872 9396 20888
rect 9620 21264 9654 21280
rect 9620 20872 9654 20888
rect 8376 20804 8392 20838
rect 8560 20804 8576 20838
rect 8634 20804 8650 20838
rect 8818 20804 8834 20838
rect 8892 20804 8908 20838
rect 9076 20804 9092 20838
rect 9150 20804 9166 20838
rect 9334 20804 9350 20838
rect 9408 20804 9424 20838
rect 9592 20804 9608 20838
rect 8376 20696 8392 20730
rect 8560 20696 8576 20730
rect 8634 20696 8650 20730
rect 8818 20696 8834 20730
rect 8892 20696 8908 20730
rect 9076 20696 9092 20730
rect 9150 20696 9166 20730
rect 9334 20696 9350 20730
rect 9408 20696 9424 20730
rect 9592 20696 9608 20730
rect 8330 20646 8364 20662
rect 8330 20254 8364 20270
rect 8588 20646 8622 20662
rect 8588 20254 8622 20270
rect 8846 20646 8880 20662
rect 8846 20254 8880 20270
rect 9104 20646 9138 20662
rect 9104 20254 9138 20270
rect 9362 20646 9396 20662
rect 9362 20254 9396 20270
rect 9620 20646 9654 20662
rect 9620 20254 9654 20270
rect 8376 20186 8392 20220
rect 8560 20186 8576 20220
rect 8634 20186 8650 20220
rect 8818 20186 8834 20220
rect 8892 20186 8908 20220
rect 9076 20186 9092 20220
rect 9150 20186 9166 20220
rect 9334 20186 9350 20220
rect 9408 20186 9424 20220
rect 9592 20186 9608 20220
rect 8376 20078 8392 20112
rect 8560 20078 8576 20112
rect 8634 20078 8650 20112
rect 8818 20078 8834 20112
rect 8892 20078 8908 20112
rect 9076 20078 9092 20112
rect 9150 20078 9166 20112
rect 9334 20078 9350 20112
rect 9408 20078 9424 20112
rect 9592 20078 9608 20112
rect 8330 20028 8364 20044
rect 8330 19636 8364 19652
rect 8588 20028 8622 20044
rect 8588 19636 8622 19652
rect 8846 20028 8880 20044
rect 8846 19636 8880 19652
rect 9104 20028 9138 20044
rect 9104 19636 9138 19652
rect 9362 20028 9396 20044
rect 9362 19636 9396 19652
rect 9620 20028 9654 20044
rect 9620 19636 9654 19652
rect 8376 19568 8392 19602
rect 8560 19568 8576 19602
rect 8634 19568 8650 19602
rect 8818 19568 8834 19602
rect 8892 19568 8908 19602
rect 9076 19568 9092 19602
rect 9150 19568 9166 19602
rect 9334 19568 9350 19602
rect 9408 19568 9424 19602
rect 9592 19568 9608 19602
rect 8376 19460 8392 19494
rect 8560 19460 8576 19494
rect 8634 19460 8650 19494
rect 8818 19460 8834 19494
rect 8892 19460 8908 19494
rect 9076 19460 9092 19494
rect 9150 19460 9166 19494
rect 9334 19460 9350 19494
rect 9408 19460 9424 19494
rect 9592 19460 9608 19494
rect 8330 19410 8364 19426
rect 8330 19018 8364 19034
rect 8588 19410 8622 19426
rect 8588 19018 8622 19034
rect 8846 19410 8880 19426
rect 8846 19018 8880 19034
rect 9104 19410 9138 19426
rect 9104 19018 9138 19034
rect 9362 19410 9396 19426
rect 9362 19018 9396 19034
rect 9620 19410 9654 19426
rect 9620 19018 9654 19034
rect 8376 18950 8392 18984
rect 8560 18950 8576 18984
rect 8634 18950 8650 18984
rect 8818 18950 8834 18984
rect 8892 18950 8908 18984
rect 9076 18950 9092 18984
rect 9150 18950 9166 18984
rect 9334 18950 9350 18984
rect 9408 18950 9424 18984
rect 9592 18950 9608 18984
rect 8376 18842 8392 18876
rect 8560 18842 8576 18876
rect 8634 18842 8650 18876
rect 8818 18842 8834 18876
rect 8892 18842 8908 18876
rect 9076 18842 9092 18876
rect 9150 18842 9166 18876
rect 9334 18842 9350 18876
rect 9408 18842 9424 18876
rect 9592 18842 9608 18876
rect 8330 18792 8364 18808
rect 8330 18400 8364 18416
rect 8588 18792 8622 18808
rect 8588 18400 8622 18416
rect 8846 18792 8880 18808
rect 8846 18400 8880 18416
rect 9104 18792 9138 18808
rect 9104 18400 9138 18416
rect 9362 18792 9396 18808
rect 9362 18400 9396 18416
rect 9620 18792 9654 18808
rect 9620 18400 9654 18416
rect 8376 18332 8392 18366
rect 8560 18332 8576 18366
rect 8634 18332 8650 18366
rect 8818 18332 8834 18366
rect 8892 18332 8908 18366
rect 9076 18332 9092 18366
rect 9150 18332 9166 18366
rect 9334 18332 9350 18366
rect 9408 18332 9424 18366
rect 9592 18332 9608 18366
rect 8376 18224 8392 18258
rect 8560 18224 8576 18258
rect 8634 18224 8650 18258
rect 8818 18224 8834 18258
rect 8892 18224 8908 18258
rect 9076 18224 9092 18258
rect 9150 18224 9166 18258
rect 9334 18224 9350 18258
rect 9408 18224 9424 18258
rect 9592 18224 9608 18258
rect 8330 18174 8364 18190
rect 8330 17782 8364 17798
rect 8588 18174 8622 18190
rect 8588 17782 8622 17798
rect 8846 18174 8880 18190
rect 8846 17782 8880 17798
rect 9104 18174 9138 18190
rect 9104 17782 9138 17798
rect 9362 18174 9396 18190
rect 9362 17782 9396 17798
rect 9620 18174 9654 18190
rect 9620 17782 9654 17798
rect 6656 17714 6672 17748
rect 6840 17714 6856 17748
rect 6914 17714 6930 17748
rect 7098 17714 7114 17748
rect 7172 17714 7188 17748
rect 7356 17714 7372 17748
rect 7430 17714 7446 17748
rect 7614 17714 7630 17748
rect 7688 17714 7704 17748
rect 7872 17714 7888 17748
rect 6496 17646 6530 17708
rect 8376 17714 8392 17748
rect 8560 17714 8576 17748
rect 8634 17714 8650 17748
rect 8818 17714 8834 17748
rect 8892 17714 8908 17748
rect 9076 17714 9092 17748
rect 9150 17714 9166 17748
rect 9334 17714 9350 17748
rect 9408 17714 9424 17748
rect 9592 17714 9608 17748
rect 8014 17646 8040 17708
rect 6496 17612 6592 17646
rect 7952 17616 8040 17646
rect 8220 17646 8250 17708
rect 19384 22242 19418 22304
rect 18438 22202 18454 22236
rect 18488 22202 18504 22236
rect 18630 22202 18646 22236
rect 18680 22202 18696 22236
rect 18822 22202 18838 22236
rect 18872 22202 18888 22236
rect 19014 22202 19030 22236
rect 19064 22202 19080 22236
rect 19206 22202 19222 22236
rect 19256 22202 19272 22236
rect 18310 22152 18344 22168
rect 18310 21760 18344 21776
rect 18406 22152 18440 22168
rect 18406 21760 18440 21776
rect 18502 22152 18536 22168
rect 18502 21760 18536 21776
rect 18598 22152 18632 22168
rect 18598 21760 18632 21776
rect 18694 22152 18728 22168
rect 18694 21760 18728 21776
rect 18790 22152 18824 22168
rect 18790 21760 18824 21776
rect 18886 22152 18920 22168
rect 18886 21760 18920 21776
rect 18982 22152 19016 22168
rect 18982 21760 19016 21776
rect 19078 22152 19112 22168
rect 19078 21760 19112 21776
rect 19174 22152 19208 22168
rect 19174 21760 19208 21776
rect 19270 22152 19304 22168
rect 19270 21760 19304 21776
rect 18342 21692 18358 21726
rect 18392 21692 18408 21726
rect 18534 21692 18550 21726
rect 18584 21692 18600 21726
rect 18726 21692 18742 21726
rect 18776 21692 18792 21726
rect 18918 21692 18934 21726
rect 18968 21692 18984 21726
rect 19110 21692 19126 21726
rect 19160 21692 19176 21726
rect 18342 21584 18358 21618
rect 18392 21584 18408 21618
rect 18534 21584 18550 21618
rect 18584 21584 18600 21618
rect 18726 21584 18742 21618
rect 18776 21584 18792 21618
rect 18918 21584 18934 21618
rect 18968 21584 18984 21618
rect 19110 21584 19126 21618
rect 19160 21584 19176 21618
rect 18310 21534 18344 21550
rect 18310 21142 18344 21158
rect 18406 21534 18440 21550
rect 18406 21142 18440 21158
rect 18502 21534 18536 21550
rect 18502 21142 18536 21158
rect 18598 21534 18632 21550
rect 18598 21142 18632 21158
rect 18694 21534 18728 21550
rect 18694 21142 18728 21158
rect 18790 21534 18824 21550
rect 18790 21142 18824 21158
rect 18886 21534 18920 21550
rect 18886 21142 18920 21158
rect 18982 21534 19016 21550
rect 18982 21142 19016 21158
rect 19078 21534 19112 21550
rect 19078 21142 19112 21158
rect 19174 21534 19208 21550
rect 19174 21142 19208 21158
rect 19270 21534 19304 21550
rect 19270 21142 19304 21158
rect 18438 21074 18454 21108
rect 18488 21074 18504 21108
rect 18630 21074 18646 21108
rect 18680 21074 18696 21108
rect 18822 21074 18838 21108
rect 18872 21074 18888 21108
rect 19014 21074 19030 21108
rect 19064 21074 19080 21108
rect 19206 21074 19222 21108
rect 19256 21074 19272 21108
rect 18196 21006 18230 21068
rect 19384 21006 19418 21068
rect 18196 20972 18292 21006
rect 19322 20972 19418 21006
rect 18540 20854 18680 20972
rect 18196 20820 18292 20854
rect 19652 20820 19748 20854
rect 18196 20758 18230 20820
rect 10056 19866 10152 19900
rect 10894 19866 10990 19900
rect 10056 19804 10090 19866
rect 10956 19804 10990 19866
rect 10298 19764 10314 19798
rect 10348 19764 10364 19798
rect 10490 19764 10506 19798
rect 10540 19764 10556 19798
rect 10682 19764 10698 19798
rect 10732 19764 10748 19798
rect 10170 19714 10204 19730
rect 10170 19322 10204 19338
rect 10266 19714 10300 19730
rect 10266 19322 10300 19338
rect 10362 19714 10396 19730
rect 10362 19322 10396 19338
rect 10458 19714 10492 19730
rect 10458 19322 10492 19338
rect 10554 19714 10588 19730
rect 10554 19322 10588 19338
rect 10650 19714 10684 19730
rect 10650 19322 10684 19338
rect 10746 19714 10780 19730
rect 10746 19322 10780 19338
rect 10842 19714 10876 19730
rect 10842 19322 10876 19338
rect 10202 19254 10218 19288
rect 10252 19254 10268 19288
rect 10394 19254 10410 19288
rect 10444 19254 10460 19288
rect 10586 19254 10602 19288
rect 10636 19254 10652 19288
rect 10778 19254 10794 19288
rect 10828 19254 10844 19288
rect 10056 19186 10090 19248
rect 10956 19186 10990 19248
rect 10056 19152 10152 19186
rect 10894 19152 10990 19186
rect 10060 18978 10240 19152
rect 10056 18944 10152 18978
rect 11182 18944 11278 18978
rect 10056 18882 10090 18944
rect 9768 17708 10056 17776
rect 11244 18882 11278 18944
rect 10202 18842 10218 18876
rect 10252 18842 10268 18876
rect 10394 18842 10410 18876
rect 10444 18842 10460 18876
rect 10586 18842 10602 18876
rect 10636 18842 10652 18876
rect 10778 18842 10794 18876
rect 10828 18842 10844 18876
rect 10970 18842 10986 18876
rect 11020 18842 11036 18876
rect 10170 18792 10204 18808
rect 10170 18400 10204 18416
rect 10266 18792 10300 18808
rect 10266 18400 10300 18416
rect 10362 18792 10396 18808
rect 10362 18400 10396 18416
rect 10458 18792 10492 18808
rect 10458 18400 10492 18416
rect 10554 18792 10588 18808
rect 10554 18400 10588 18416
rect 10650 18792 10684 18808
rect 10650 18400 10684 18416
rect 10746 18792 10780 18808
rect 10746 18400 10780 18416
rect 10842 18792 10876 18808
rect 10842 18400 10876 18416
rect 10938 18792 10972 18808
rect 10938 18400 10972 18416
rect 11034 18792 11068 18808
rect 11034 18400 11068 18416
rect 11130 18792 11164 18808
rect 11130 18400 11164 18416
rect 10298 18332 10314 18366
rect 10348 18332 10364 18366
rect 10490 18332 10506 18366
rect 10540 18332 10556 18366
rect 10682 18332 10698 18366
rect 10732 18332 10748 18366
rect 10874 18332 10890 18366
rect 10924 18332 10940 18366
rect 11066 18332 11082 18366
rect 11116 18332 11132 18366
rect 10298 18224 10314 18258
rect 10348 18224 10364 18258
rect 10490 18224 10506 18258
rect 10540 18224 10556 18258
rect 10682 18224 10698 18258
rect 10732 18224 10748 18258
rect 10874 18224 10890 18258
rect 10924 18224 10940 18258
rect 11066 18224 11082 18258
rect 11116 18224 11132 18258
rect 10170 18174 10204 18190
rect 10170 17782 10204 17798
rect 10266 18174 10300 18190
rect 10266 17782 10300 17798
rect 10362 18174 10396 18190
rect 10362 17782 10396 17798
rect 10458 18174 10492 18190
rect 10458 17782 10492 17798
rect 10554 18174 10588 18190
rect 10554 17782 10588 17798
rect 10650 18174 10684 18190
rect 10650 17782 10684 17798
rect 10746 18174 10780 18190
rect 10746 17782 10780 17798
rect 10842 18174 10876 18190
rect 10842 17782 10876 17798
rect 10938 18174 10972 18190
rect 10938 17782 10972 17798
rect 11034 18174 11068 18190
rect 11034 17782 11068 17798
rect 11130 18174 11164 18190
rect 11130 17782 11164 17798
rect 10202 17714 10218 17748
rect 10252 17714 10268 17748
rect 10394 17714 10410 17748
rect 10444 17714 10460 17748
rect 10586 17714 10602 17748
rect 10636 17714 10652 17748
rect 10778 17714 10794 17748
rect 10828 17714 10844 17748
rect 10970 17714 10986 17748
rect 11020 17714 11036 17748
rect 9734 17646 10090 17708
rect 19714 20758 19748 20820
rect 18356 20718 18372 20752
rect 18540 20718 18556 20752
rect 18614 20718 18630 20752
rect 18798 20718 18814 20752
rect 18872 20718 18888 20752
rect 19056 20718 19072 20752
rect 19130 20718 19146 20752
rect 19314 20718 19330 20752
rect 19388 20718 19404 20752
rect 19572 20718 19588 20752
rect 18310 20668 18344 20684
rect 18310 20276 18344 20292
rect 18568 20668 18602 20684
rect 18568 20276 18602 20292
rect 18826 20668 18860 20684
rect 18826 20276 18860 20292
rect 19084 20668 19118 20684
rect 19084 20276 19118 20292
rect 19342 20668 19376 20684
rect 19342 20276 19376 20292
rect 19600 20668 19634 20684
rect 19600 20276 19634 20292
rect 18356 20208 18372 20242
rect 18540 20208 18556 20242
rect 18614 20208 18630 20242
rect 18798 20208 18814 20242
rect 18872 20208 18888 20242
rect 19056 20208 19072 20242
rect 19130 20208 19146 20242
rect 19314 20208 19330 20242
rect 19388 20208 19404 20242
rect 19572 20208 19588 20242
rect 18356 20100 18372 20134
rect 18540 20100 18556 20134
rect 18614 20100 18630 20134
rect 18798 20100 18814 20134
rect 18872 20100 18888 20134
rect 19056 20100 19072 20134
rect 19130 20100 19146 20134
rect 19314 20100 19330 20134
rect 19388 20100 19404 20134
rect 19572 20100 19588 20134
rect 18310 20050 18344 20066
rect 18310 19658 18344 19674
rect 18568 20050 18602 20066
rect 18568 19658 18602 19674
rect 18826 20050 18860 20066
rect 18826 19658 18860 19674
rect 19084 20050 19118 20066
rect 19084 19658 19118 19674
rect 19342 20050 19376 20066
rect 19342 19658 19376 19674
rect 19600 20050 19634 20066
rect 19600 19658 19634 19674
rect 18356 19590 18372 19624
rect 18540 19590 18556 19624
rect 18614 19590 18630 19624
rect 18798 19590 18814 19624
rect 18872 19590 18888 19624
rect 19056 19590 19072 19624
rect 19130 19590 19146 19624
rect 19314 19590 19330 19624
rect 19388 19590 19404 19624
rect 19572 19590 19588 19624
rect 18356 19482 18372 19516
rect 18540 19482 18556 19516
rect 18614 19482 18630 19516
rect 18798 19482 18814 19516
rect 18872 19482 18888 19516
rect 19056 19482 19072 19516
rect 19130 19482 19146 19516
rect 19314 19482 19330 19516
rect 19388 19482 19404 19516
rect 19572 19482 19588 19516
rect 18310 19432 18344 19448
rect 18310 19040 18344 19056
rect 18568 19432 18602 19448
rect 18568 19040 18602 19056
rect 18826 19432 18860 19448
rect 18826 19040 18860 19056
rect 19084 19432 19118 19448
rect 19084 19040 19118 19056
rect 19342 19432 19376 19448
rect 19342 19040 19376 19056
rect 19600 19432 19634 19448
rect 19600 19040 19634 19056
rect 18356 18972 18372 19006
rect 18540 18972 18556 19006
rect 18614 18972 18630 19006
rect 18798 18972 18814 19006
rect 18872 18972 18888 19006
rect 19056 18972 19072 19006
rect 19130 18972 19146 19006
rect 19314 18972 19330 19006
rect 19388 18972 19404 19006
rect 19572 18972 19588 19006
rect 18356 18864 18372 18898
rect 18540 18864 18556 18898
rect 18614 18864 18630 18898
rect 18798 18864 18814 18898
rect 18872 18864 18888 18898
rect 19056 18864 19072 18898
rect 19130 18864 19146 18898
rect 19314 18864 19330 18898
rect 19388 18864 19404 18898
rect 19572 18864 19588 18898
rect 18310 18814 18344 18830
rect 18310 18422 18344 18438
rect 18568 18814 18602 18830
rect 18568 18422 18602 18438
rect 18826 18814 18860 18830
rect 18826 18422 18860 18438
rect 19084 18814 19118 18830
rect 19084 18422 19118 18438
rect 19342 18814 19376 18830
rect 19342 18422 19376 18438
rect 19600 18814 19634 18830
rect 19600 18422 19634 18438
rect 18356 18354 18372 18388
rect 18540 18354 18556 18388
rect 18614 18354 18630 18388
rect 18798 18354 18814 18388
rect 18872 18354 18888 18388
rect 19056 18354 19072 18388
rect 19130 18354 19146 18388
rect 19314 18354 19330 18388
rect 19388 18354 19404 18388
rect 19572 18354 19588 18388
rect 18196 18286 18230 18348
rect 19714 18286 19748 18348
rect 18196 18252 18292 18286
rect 19652 18252 19748 18286
rect 18480 18156 18680 18252
rect 11244 17646 11278 17708
rect 8220 17616 8312 17646
rect 7952 17612 8048 17616
rect 8216 17612 8312 17616
rect 9672 17616 10152 17646
rect 9672 17612 9768 17616
rect 10056 17612 10152 17616
rect 11182 17612 11278 17646
rect 2472 11214 2568 11248
rect 4808 11214 4904 11248
rect 2472 11152 2506 11214
rect 1300 9183 1568 10532
rect 4870 11152 4904 11214
rect 2472 9358 2506 9420
rect 16872 11214 16968 11248
rect 19208 11214 19304 11248
rect 16872 11152 16906 11214
rect 6096 10466 6276 10608
rect 4870 9358 4904 9420
rect 2472 9324 2568 9358
rect 4808 9324 4904 9358
rect 5012 10432 5108 10466
rect 7098 10432 7194 10466
rect 5012 10370 5046 10432
rect 1297 9149 1357 9183
rect 3983 9149 4043 9183
rect 1297 9123 1331 9149
rect -10164 8374 -10068 8408
rect -9038 8374 -8942 8408
rect -10164 8312 -10130 8374
rect -8976 8312 -8942 8374
rect -9922 8272 -9906 8306
rect -9872 8272 -9856 8306
rect -9730 8272 -9714 8306
rect -9680 8272 -9664 8306
rect -9538 8272 -9522 8306
rect -9488 8272 -9472 8306
rect -9346 8272 -9330 8306
rect -9296 8272 -9280 8306
rect -9154 8272 -9138 8306
rect -9104 8272 -9088 8306
rect -10050 8222 -10016 8238
rect -10050 7830 -10016 7846
rect -9954 8222 -9920 8238
rect -9954 7830 -9920 7846
rect -9858 8222 -9824 8238
rect -9858 7830 -9824 7846
rect -9762 8222 -9728 8238
rect -9762 7830 -9728 7846
rect -9666 8222 -9632 8238
rect -9666 7830 -9632 7846
rect -9570 8222 -9536 8238
rect -9570 7830 -9536 7846
rect -9474 8222 -9440 8238
rect -9474 7830 -9440 7846
rect -9378 8222 -9344 8238
rect -9378 7830 -9344 7846
rect -9282 8222 -9248 8238
rect -9282 7830 -9248 7846
rect -9186 8222 -9152 8238
rect -9186 7830 -9152 7846
rect -9090 8222 -9056 8238
rect -9090 7830 -9056 7846
rect -10018 7762 -10002 7796
rect -9968 7762 -9952 7796
rect -9826 7762 -9810 7796
rect -9776 7762 -9760 7796
rect -9634 7762 -9618 7796
rect -9584 7762 -9568 7796
rect -9442 7762 -9426 7796
rect -9392 7762 -9376 7796
rect -9250 7762 -9234 7796
rect -9200 7762 -9184 7796
rect -10018 7654 -10002 7688
rect -9968 7654 -9952 7688
rect -9826 7654 -9810 7688
rect -9776 7654 -9760 7688
rect -9634 7654 -9618 7688
rect -9584 7654 -9568 7688
rect -9442 7654 -9426 7688
rect -9392 7654 -9376 7688
rect -9250 7654 -9234 7688
rect -9200 7654 -9184 7688
rect -10050 7604 -10016 7620
rect -10050 7212 -10016 7228
rect -9954 7604 -9920 7620
rect -9954 7212 -9920 7228
rect -9858 7604 -9824 7620
rect -9858 7212 -9824 7228
rect -9762 7604 -9728 7620
rect -9762 7212 -9728 7228
rect -9666 7604 -9632 7620
rect -9666 7212 -9632 7228
rect -9570 7604 -9536 7620
rect -9570 7212 -9536 7228
rect -9474 7604 -9440 7620
rect -9474 7212 -9440 7228
rect -9378 7604 -9344 7620
rect -9378 7212 -9344 7228
rect -9282 7604 -9248 7620
rect -9282 7212 -9248 7228
rect -9186 7604 -9152 7620
rect -9186 7212 -9152 7228
rect -9090 7604 -9056 7620
rect -9090 7212 -9056 7228
rect -9922 7144 -9906 7178
rect -9872 7144 -9856 7178
rect -9730 7144 -9714 7178
rect -9680 7144 -9664 7178
rect -9538 7144 -9522 7178
rect -9488 7144 -9472 7178
rect -9346 7144 -9330 7178
rect -9296 7144 -9280 7178
rect -9154 7144 -9138 7178
rect -9104 7144 -9088 7178
rect -9922 7036 -9906 7070
rect -9872 7036 -9856 7070
rect -9730 7036 -9714 7070
rect -9680 7036 -9664 7070
rect -9538 7036 -9522 7070
rect -9488 7036 -9472 7070
rect -9346 7036 -9330 7070
rect -9296 7036 -9280 7070
rect -9154 7036 -9138 7070
rect -9104 7036 -9088 7070
rect -10050 6986 -10016 7002
rect -10050 6594 -10016 6610
rect -9954 6986 -9920 7002
rect -9954 6594 -9920 6610
rect -9858 6986 -9824 7002
rect -9858 6594 -9824 6610
rect -9762 6986 -9728 7002
rect -9762 6594 -9728 6610
rect -9666 6986 -9632 7002
rect -9666 6594 -9632 6610
rect -9570 6986 -9536 7002
rect -9570 6594 -9536 6610
rect -9474 6986 -9440 7002
rect -9474 6594 -9440 6610
rect -9378 6986 -9344 7002
rect -9378 6594 -9344 6610
rect -9282 6986 -9248 7002
rect -9282 6594 -9248 6610
rect -9186 6986 -9152 7002
rect -9186 6594 -9152 6610
rect -9090 6986 -9056 7002
rect -9090 6594 -9056 6610
rect -10018 6526 -10002 6560
rect -9968 6526 -9952 6560
rect -9826 6526 -9810 6560
rect -9776 6526 -9760 6560
rect -9634 6526 -9618 6560
rect -9584 6526 -9568 6560
rect -9442 6526 -9426 6560
rect -9392 6526 -9376 6560
rect -9250 6526 -9234 6560
rect -9200 6526 -9184 6560
rect -10164 6458 -10130 6520
rect -8844 8310 -8748 8344
rect -8392 8310 -8296 8344
rect -8844 8248 -8810 8310
rect -8942 6520 -8844 6668
rect -8330 8248 -8296 8310
rect -8674 8196 -8658 8230
rect -8482 8196 -8466 8230
rect -8742 8168 -8708 8184
rect -8742 6584 -8708 6600
rect -8432 8168 -8398 8184
rect -8432 6584 -8398 6600
rect -8674 6538 -8658 6572
rect -8482 6538 -8466 6572
rect -8976 6458 -8810 6520
rect -8330 6458 -8296 6520
rect -10164 6424 -10068 6458
rect -9038 6448 -8748 6458
rect -9038 6424 -8942 6448
rect -8844 6424 -8748 6448
rect -8392 6424 -8296 6458
rect -10120 6328 -10020 6424
rect -10164 6294 -10068 6328
rect -9038 6294 -8942 6328
rect -10164 6232 -10130 6294
rect -8976 6232 -8942 6294
rect 4009 9123 4043 9149
rect 1528 8870 1672 8956
rect 1964 8904 2540 8956
rect 2832 8904 3476 8956
rect 3768 8904 3816 8956
rect 3662 8870 3816 8904
rect 1528 8808 1610 8870
rect 1528 8704 1576 8808
rect 3724 8808 3816 8870
rect 1818 8768 1834 8802
rect 1868 8768 1884 8802
rect 2010 8768 2026 8802
rect 2060 8768 2076 8802
rect 2202 8768 2218 8802
rect 2252 8768 2268 8802
rect 2394 8768 2410 8802
rect 2444 8768 2460 8802
rect 2586 8768 2602 8802
rect 2636 8768 2652 8802
rect 2778 8768 2794 8802
rect 2828 8768 2844 8802
rect 2970 8768 2986 8802
rect 3020 8768 3036 8802
rect 3162 8768 3178 8802
rect 3212 8768 3228 8802
rect 3354 8768 3370 8802
rect 3404 8768 3420 8802
rect 3546 8768 3562 8802
rect 3596 8768 3612 8802
rect 1528 8356 1540 8704
rect 1528 8252 1576 8356
rect 1690 8718 1724 8734
rect 1690 8326 1724 8342
rect 1786 8718 1820 8734
rect 1786 8326 1820 8342
rect 1882 8718 1916 8734
rect 1882 8326 1916 8342
rect 1978 8718 2012 8734
rect 1978 8326 2012 8342
rect 2074 8718 2108 8734
rect 2074 8326 2108 8342
rect 2170 8718 2204 8734
rect 2170 8326 2204 8342
rect 2266 8718 2300 8734
rect 2266 8326 2300 8342
rect 2362 8718 2396 8734
rect 2362 8326 2396 8342
rect 2458 8718 2492 8734
rect 2458 8326 2492 8342
rect 2554 8718 2588 8734
rect 2554 8326 2588 8342
rect 2650 8718 2684 8734
rect 2650 8326 2684 8342
rect 2746 8718 2780 8734
rect 2746 8326 2780 8342
rect 2842 8718 2876 8734
rect 2842 8326 2876 8342
rect 2938 8718 2972 8734
rect 2938 8326 2972 8342
rect 3034 8718 3068 8734
rect 3034 8326 3068 8342
rect 3130 8718 3164 8734
rect 3130 8326 3164 8342
rect 3226 8718 3260 8734
rect 3226 8326 3260 8342
rect 3322 8718 3356 8734
rect 3322 8326 3356 8342
rect 3418 8718 3452 8734
rect 3418 8326 3452 8342
rect 3514 8718 3548 8734
rect 3514 8326 3548 8342
rect 3610 8718 3644 8734
rect 3610 8326 3644 8342
rect 3758 8672 3816 8808
rect 3800 8416 3816 8672
rect 1722 8258 1738 8292
rect 1772 8258 1788 8292
rect 1914 8258 1930 8292
rect 1964 8258 1980 8292
rect 2106 8258 2122 8292
rect 2156 8258 2172 8292
rect 2298 8258 2314 8292
rect 2348 8258 2364 8292
rect 2490 8258 2506 8292
rect 2540 8258 2556 8292
rect 2682 8258 2698 8292
rect 2732 8258 2748 8292
rect 2874 8258 2890 8292
rect 2924 8258 2940 8292
rect 3066 8258 3082 8292
rect 3116 8258 3132 8292
rect 3258 8258 3274 8292
rect 3308 8258 3324 8292
rect 3450 8258 3466 8292
rect 3500 8258 3516 8292
rect 1528 8190 1610 8252
rect 3758 8252 3816 8416
rect 3724 8190 3816 8252
rect 1528 8156 1672 8190
rect 3662 8156 3816 8190
rect 1528 8152 3816 8156
rect 1528 8148 3476 8152
rect 1528 8088 1672 8148
rect 1964 8088 2540 8148
rect 2860 8092 3476 8148
rect 3768 8092 3816 8152
rect 2860 8088 3816 8092
rect 1528 8084 3816 8088
rect 1528 8050 1672 8084
rect 3662 8050 3816 8084
rect 1528 7988 1610 8050
rect 1528 7844 1576 7988
rect 3724 7988 3816 8050
rect 1818 7948 1834 7982
rect 1868 7948 1884 7982
rect 2010 7948 2026 7982
rect 2060 7948 2076 7982
rect 2202 7948 2218 7982
rect 2252 7948 2268 7982
rect 2394 7948 2410 7982
rect 2444 7948 2460 7982
rect 2586 7948 2602 7982
rect 2636 7948 2652 7982
rect 2778 7948 2794 7982
rect 2828 7948 2844 7982
rect 2970 7948 2986 7982
rect 3020 7948 3036 7982
rect 3162 7948 3178 7982
rect 3212 7948 3228 7982
rect 3354 7948 3370 7982
rect 3404 7948 3420 7982
rect 3546 7948 3562 7982
rect 3596 7948 3612 7982
rect 1528 7588 1540 7844
rect 1528 7432 1576 7588
rect 1690 7898 1724 7914
rect 1690 7506 1724 7522
rect 1786 7898 1820 7914
rect 1786 7506 1820 7522
rect 1882 7898 1916 7914
rect 1882 7506 1916 7522
rect 1978 7898 2012 7914
rect 1978 7506 2012 7522
rect 2074 7898 2108 7914
rect 2074 7506 2108 7522
rect 2170 7898 2204 7914
rect 2170 7506 2204 7522
rect 2266 7898 2300 7914
rect 2266 7506 2300 7522
rect 2362 7898 2396 7914
rect 2362 7506 2396 7522
rect 2458 7898 2492 7914
rect 2458 7506 2492 7522
rect 2554 7898 2588 7914
rect 2554 7506 2588 7522
rect 2650 7898 2684 7914
rect 2650 7506 2684 7522
rect 2746 7898 2780 7914
rect 2746 7506 2780 7522
rect 2842 7898 2876 7914
rect 2842 7506 2876 7522
rect 2938 7898 2972 7914
rect 2938 7506 2972 7522
rect 3034 7898 3068 7914
rect 3034 7506 3068 7522
rect 3130 7898 3164 7914
rect 3130 7506 3164 7522
rect 3226 7898 3260 7914
rect 3226 7506 3260 7522
rect 3322 7898 3356 7914
rect 3322 7506 3356 7522
rect 3418 7898 3452 7914
rect 3418 7506 3452 7522
rect 3514 7898 3548 7914
rect 3514 7506 3548 7522
rect 3610 7898 3644 7914
rect 3610 7506 3644 7522
rect 3758 7824 3816 7988
rect 3800 7568 3816 7824
rect 1722 7438 1738 7472
rect 1772 7438 1788 7472
rect 1914 7438 1930 7472
rect 1964 7438 1980 7472
rect 2106 7438 2122 7472
rect 2156 7438 2172 7472
rect 2298 7438 2314 7472
rect 2348 7438 2364 7472
rect 2490 7438 2506 7472
rect 2540 7438 2556 7472
rect 2682 7438 2698 7472
rect 2732 7438 2748 7472
rect 2874 7438 2890 7472
rect 2924 7438 2940 7472
rect 3066 7438 3082 7472
rect 3116 7438 3132 7472
rect 3258 7438 3274 7472
rect 3308 7438 3324 7472
rect 3450 7438 3466 7472
rect 3500 7438 3516 7472
rect 1528 7370 1610 7432
rect 3758 7432 3816 7568
rect 3724 7370 3816 7432
rect 1528 7336 1672 7370
rect 3662 7336 3816 7370
rect 1528 7328 3816 7336
rect 1528 7268 1672 7328
rect 1964 7268 2540 7328
rect 2832 7268 3476 7328
rect 3768 7268 3816 7328
rect 1528 7264 3816 7268
rect 1528 7230 1672 7264
rect 3662 7230 3816 7264
rect 1528 7168 1610 7230
rect 1528 7004 1576 7168
rect 3724 7168 3816 7230
rect 1818 7128 1834 7162
rect 1868 7128 1884 7162
rect 2010 7128 2026 7162
rect 2060 7128 2076 7162
rect 2202 7128 2218 7162
rect 2252 7128 2268 7162
rect 2394 7128 2410 7162
rect 2444 7128 2460 7162
rect 2586 7128 2602 7162
rect 2636 7128 2652 7162
rect 2778 7128 2794 7162
rect 2828 7128 2844 7162
rect 2970 7128 2986 7162
rect 3020 7128 3036 7162
rect 3162 7128 3178 7162
rect 3212 7128 3228 7162
rect 3354 7128 3370 7162
rect 3404 7128 3420 7162
rect 3546 7128 3562 7162
rect 3596 7128 3612 7162
rect 1528 6748 1536 7004
rect 1528 6612 1576 6748
rect 1690 7078 1724 7094
rect 1690 6686 1724 6702
rect 1786 7078 1820 7094
rect 1786 6686 1820 6702
rect 1882 7078 1916 7094
rect 1882 6686 1916 6702
rect 1978 7078 2012 7094
rect 1978 6686 2012 6702
rect 2074 7078 2108 7094
rect 2074 6686 2108 6702
rect 2170 7078 2204 7094
rect 2170 6686 2204 6702
rect 2266 7078 2300 7094
rect 2266 6686 2300 6702
rect 2362 7078 2396 7094
rect 2362 6686 2396 6702
rect 2458 7078 2492 7094
rect 2458 6686 2492 6702
rect 2554 7078 2588 7094
rect 2554 6686 2588 6702
rect 2650 7078 2684 7094
rect 2650 6686 2684 6702
rect 2746 7078 2780 7094
rect 2746 6686 2780 6702
rect 2842 7078 2876 7094
rect 2842 6686 2876 6702
rect 2938 7078 2972 7094
rect 2938 6686 2972 6702
rect 3034 7078 3068 7094
rect 3034 6686 3068 6702
rect 3130 7078 3164 7094
rect 3130 6686 3164 6702
rect 3226 7078 3260 7094
rect 3226 6686 3260 6702
rect 3322 7078 3356 7094
rect 3322 6686 3356 6702
rect 3418 7078 3452 7094
rect 3418 6686 3452 6702
rect 3514 7078 3548 7094
rect 3514 6686 3548 6702
rect 3610 7078 3644 7094
rect 3610 6686 3644 6702
rect 3758 7012 3816 7168
rect 3800 6756 3816 7012
rect 1722 6618 1738 6652
rect 1772 6618 1788 6652
rect 1914 6618 1930 6652
rect 1964 6618 1980 6652
rect 2106 6618 2122 6652
rect 2156 6618 2172 6652
rect 2298 6618 2314 6652
rect 2348 6618 2364 6652
rect 2490 6618 2506 6652
rect 2540 6618 2556 6652
rect 2682 6618 2698 6652
rect 2732 6618 2748 6652
rect 2874 6618 2890 6652
rect 2924 6618 2940 6652
rect 3066 6618 3082 6652
rect 3116 6618 3132 6652
rect 3258 6618 3274 6652
rect 3308 6618 3324 6652
rect 3450 6618 3466 6652
rect 3500 6618 3516 6652
rect 1528 6550 1610 6612
rect 3758 6612 3816 6756
rect 3724 6550 3816 6612
rect 1528 6468 1672 6550
rect 3662 6516 3816 6550
rect 1964 6468 2540 6516
rect 2832 6512 3816 6516
rect 2832 6468 3476 6512
rect 3768 6468 3816 6512
rect 1297 6271 1331 6297
rect 4492 8858 4724 9324
rect 7160 10370 7194 10432
rect 5158 10330 5174 10364
rect 5208 10330 5224 10364
rect 5350 10330 5366 10364
rect 5400 10330 5416 10364
rect 5542 10330 5558 10364
rect 5592 10330 5608 10364
rect 5734 10330 5750 10364
rect 5784 10330 5800 10364
rect 5926 10330 5942 10364
rect 5976 10330 5992 10364
rect 6118 10330 6134 10364
rect 6168 10330 6184 10364
rect 6310 10330 6326 10364
rect 6360 10330 6376 10364
rect 6502 10330 6518 10364
rect 6552 10330 6568 10364
rect 6694 10330 6710 10364
rect 6744 10330 6760 10364
rect 6886 10330 6902 10364
rect 6936 10330 6952 10364
rect 5126 10271 5160 10287
rect 5126 9879 5160 9895
rect 5222 10271 5256 10287
rect 5222 9879 5256 9895
rect 5318 10271 5352 10287
rect 5318 9879 5352 9895
rect 5414 10271 5448 10287
rect 5414 9879 5448 9895
rect 5510 10271 5544 10287
rect 5510 9879 5544 9895
rect 5606 10271 5640 10287
rect 5606 9879 5640 9895
rect 5702 10271 5736 10287
rect 5702 9879 5736 9895
rect 5798 10271 5832 10287
rect 5798 9879 5832 9895
rect 5894 10271 5928 10287
rect 5894 9879 5928 9895
rect 5990 10271 6024 10287
rect 5990 9879 6024 9895
rect 6086 10271 6120 10287
rect 6086 9879 6120 9895
rect 6182 10271 6216 10287
rect 6182 9879 6216 9895
rect 6278 10271 6312 10287
rect 6278 9879 6312 9895
rect 6374 10271 6408 10287
rect 6374 9879 6408 9895
rect 6470 10271 6504 10287
rect 6470 9879 6504 9895
rect 6566 10271 6600 10287
rect 6566 9879 6600 9895
rect 6662 10271 6696 10287
rect 6662 9879 6696 9895
rect 6758 10271 6792 10287
rect 6758 9879 6792 9895
rect 6854 10271 6888 10287
rect 6854 9879 6888 9895
rect 6950 10271 6984 10287
rect 6950 9879 6984 9895
rect 7046 10271 7080 10287
rect 7046 9879 7080 9895
rect 5254 9802 5270 9836
rect 5304 9802 5320 9836
rect 5446 9802 5462 9836
rect 5496 9802 5512 9836
rect 5638 9802 5654 9836
rect 5688 9802 5704 9836
rect 5830 9802 5846 9836
rect 5880 9802 5896 9836
rect 6022 9802 6038 9836
rect 6072 9802 6088 9836
rect 6214 9802 6230 9836
rect 6264 9802 6280 9836
rect 6406 9802 6422 9836
rect 6456 9802 6472 9836
rect 6598 9802 6614 9836
rect 6648 9802 6664 9836
rect 6790 9802 6806 9836
rect 6840 9802 6856 9836
rect 6982 9802 6998 9836
rect 7032 9802 7048 9836
rect 5254 9694 5270 9728
rect 5304 9694 5320 9728
rect 5446 9694 5462 9728
rect 5496 9694 5512 9728
rect 5638 9694 5654 9728
rect 5688 9694 5704 9728
rect 5830 9694 5846 9728
rect 5880 9694 5896 9728
rect 6022 9694 6038 9728
rect 6072 9694 6088 9728
rect 6214 9694 6230 9728
rect 6264 9694 6280 9728
rect 6406 9694 6422 9728
rect 6456 9694 6472 9728
rect 6598 9694 6614 9728
rect 6648 9694 6664 9728
rect 6790 9694 6806 9728
rect 6840 9694 6856 9728
rect 6982 9694 6998 9728
rect 7032 9694 7048 9728
rect 5126 9635 5160 9651
rect 5126 9243 5160 9259
rect 5222 9635 5256 9651
rect 5222 9243 5256 9259
rect 5318 9635 5352 9651
rect 5318 9243 5352 9259
rect 5414 9635 5448 9651
rect 5414 9243 5448 9259
rect 5510 9635 5544 9651
rect 5510 9243 5544 9259
rect 5606 9635 5640 9651
rect 5606 9243 5640 9259
rect 5702 9635 5736 9651
rect 5702 9243 5736 9259
rect 5798 9635 5832 9651
rect 5798 9243 5832 9259
rect 5894 9635 5928 9651
rect 5894 9243 5928 9259
rect 5990 9635 6024 9651
rect 5990 9243 6024 9259
rect 6086 9635 6120 9651
rect 6086 9243 6120 9259
rect 6182 9635 6216 9651
rect 6182 9243 6216 9259
rect 6278 9635 6312 9651
rect 6278 9243 6312 9259
rect 6374 9635 6408 9651
rect 6374 9243 6408 9259
rect 6470 9635 6504 9651
rect 6470 9243 6504 9259
rect 6566 9635 6600 9651
rect 6566 9243 6600 9259
rect 6662 9635 6696 9651
rect 6662 9243 6696 9259
rect 6758 9635 6792 9651
rect 6758 9243 6792 9259
rect 6854 9635 6888 9651
rect 6854 9243 6888 9259
rect 6950 9635 6984 9651
rect 6950 9243 6984 9259
rect 7046 9635 7080 9651
rect 7046 9243 7080 9259
rect 5158 9166 5174 9200
rect 5208 9166 5224 9200
rect 5350 9166 5366 9200
rect 5400 9166 5416 9200
rect 5542 9166 5558 9200
rect 5592 9166 5608 9200
rect 5734 9166 5750 9200
rect 5784 9166 5800 9200
rect 5926 9166 5942 9200
rect 5976 9166 5992 9200
rect 6118 9166 6134 9200
rect 6168 9166 6184 9200
rect 6310 9166 6326 9200
rect 6360 9166 6376 9200
rect 6502 9166 6518 9200
rect 6552 9166 6568 9200
rect 6694 9166 6710 9200
rect 6744 9166 6760 9200
rect 6886 9166 6902 9200
rect 6936 9166 6952 9200
rect 5012 9098 5046 9160
rect 7160 9098 7194 9160
rect 5012 9064 5108 9098
rect 7098 9064 7194 9098
rect 7512 10402 7608 10436
rect 9598 10402 9694 10436
rect 7512 10340 7546 10402
rect 5012 8858 5108 8870
rect 4492 8836 5108 8858
rect 7098 8836 7194 8870
rect 4492 8774 5046 8836
rect 4492 8750 5012 8774
rect 7160 8774 7194 8836
rect 5158 8734 5174 8768
rect 5208 8734 5224 8768
rect 5350 8734 5366 8768
rect 5400 8734 5416 8768
rect 5542 8734 5558 8768
rect 5592 8734 5608 8768
rect 5734 8734 5750 8768
rect 5784 8734 5800 8768
rect 5926 8734 5942 8768
rect 5976 8734 5992 8768
rect 6118 8734 6134 8768
rect 6168 8734 6184 8768
rect 6310 8734 6326 8768
rect 6360 8734 6376 8768
rect 6502 8734 6518 8768
rect 6552 8734 6568 8768
rect 6694 8734 6710 8768
rect 6744 8734 6760 8768
rect 6886 8734 6902 8768
rect 6936 8734 6952 8768
rect 5126 8684 5160 8700
rect 5126 8292 5160 8308
rect 5222 8684 5256 8700
rect 5222 8292 5256 8308
rect 5318 8684 5352 8700
rect 5318 8292 5352 8308
rect 5414 8684 5448 8700
rect 5414 8292 5448 8308
rect 5510 8684 5544 8700
rect 5510 8292 5544 8308
rect 5606 8684 5640 8700
rect 5606 8292 5640 8308
rect 5702 8684 5736 8700
rect 5702 8292 5736 8308
rect 5798 8684 5832 8700
rect 5798 8292 5832 8308
rect 5894 8684 5928 8700
rect 5894 8292 5928 8308
rect 5990 8684 6024 8700
rect 5990 8292 6024 8308
rect 6086 8684 6120 8700
rect 6086 8292 6120 8308
rect 6182 8684 6216 8700
rect 6182 8292 6216 8308
rect 6278 8684 6312 8700
rect 6278 8292 6312 8308
rect 6374 8684 6408 8700
rect 6374 8292 6408 8308
rect 6470 8684 6504 8700
rect 6470 8292 6504 8308
rect 6566 8684 6600 8700
rect 6566 8292 6600 8308
rect 6662 8684 6696 8700
rect 6662 8292 6696 8308
rect 6758 8684 6792 8700
rect 6758 8292 6792 8308
rect 6854 8684 6888 8700
rect 6854 8292 6888 8308
rect 6950 8684 6984 8700
rect 6950 8292 6984 8308
rect 7046 8684 7080 8700
rect 7046 8292 7080 8308
rect 5254 8224 5270 8258
rect 5304 8224 5320 8258
rect 5446 8224 5462 8258
rect 5496 8224 5512 8258
rect 5638 8224 5654 8258
rect 5688 8224 5704 8258
rect 5830 8224 5846 8258
rect 5880 8224 5896 8258
rect 6022 8224 6038 8258
rect 6072 8224 6088 8258
rect 6214 8224 6230 8258
rect 6264 8224 6280 8258
rect 6406 8224 6422 8258
rect 6456 8224 6472 8258
rect 6598 8224 6614 8258
rect 6648 8224 6664 8258
rect 6790 8224 6806 8258
rect 6840 8224 6856 8258
rect 6982 8224 6998 8258
rect 7032 8224 7048 8258
rect 5254 8116 5270 8150
rect 5304 8116 5320 8150
rect 5446 8116 5462 8150
rect 5496 8116 5512 8150
rect 5638 8116 5654 8150
rect 5688 8116 5704 8150
rect 5830 8116 5846 8150
rect 5880 8116 5896 8150
rect 6022 8116 6038 8150
rect 6072 8116 6088 8150
rect 6214 8116 6230 8150
rect 6264 8116 6280 8150
rect 6406 8116 6422 8150
rect 6456 8116 6472 8150
rect 6598 8116 6614 8150
rect 6648 8116 6664 8150
rect 6790 8116 6806 8150
rect 6840 8116 6856 8150
rect 6982 8116 6998 8150
rect 7032 8116 7048 8150
rect 5126 8066 5160 8082
rect 5126 7674 5160 7690
rect 5222 8066 5256 8082
rect 5222 7674 5256 7690
rect 5318 8066 5352 8082
rect 5318 7674 5352 7690
rect 5414 8066 5448 8082
rect 5414 7674 5448 7690
rect 5510 8066 5544 8082
rect 5510 7674 5544 7690
rect 5606 8066 5640 8082
rect 5606 7674 5640 7690
rect 5702 8066 5736 8082
rect 5702 7674 5736 7690
rect 5798 8066 5832 8082
rect 5798 7674 5832 7690
rect 5894 8066 5928 8082
rect 5894 7674 5928 7690
rect 5990 8066 6024 8082
rect 5990 7674 6024 7690
rect 6086 8066 6120 8082
rect 6086 7674 6120 7690
rect 6182 8066 6216 8082
rect 6182 7674 6216 7690
rect 6278 8066 6312 8082
rect 6278 7674 6312 7690
rect 6374 8066 6408 8082
rect 6374 7674 6408 7690
rect 6470 8066 6504 8082
rect 6470 7674 6504 7690
rect 6566 8066 6600 8082
rect 6566 7674 6600 7690
rect 6662 8066 6696 8082
rect 6662 7674 6696 7690
rect 6758 8066 6792 8082
rect 6758 7674 6792 7690
rect 6854 8066 6888 8082
rect 6854 7674 6888 7690
rect 6950 8066 6984 8082
rect 6950 7674 6984 7690
rect 7046 8066 7080 8082
rect 7046 7674 7080 7690
rect 5158 7606 5174 7640
rect 5208 7606 5224 7640
rect 5350 7606 5366 7640
rect 5400 7606 5416 7640
rect 5542 7606 5558 7640
rect 5592 7606 5608 7640
rect 5734 7606 5750 7640
rect 5784 7606 5800 7640
rect 5926 7606 5942 7640
rect 5976 7606 5992 7640
rect 6118 7606 6134 7640
rect 6168 7606 6184 7640
rect 6310 7606 6326 7640
rect 6360 7606 6376 7640
rect 6502 7606 6518 7640
rect 6552 7606 6568 7640
rect 6694 7606 6710 7640
rect 6744 7606 6760 7640
rect 6886 7606 6902 7640
rect 6936 7606 6952 7640
rect 5012 7538 5046 7600
rect 7160 7538 7194 7600
rect 5012 7528 5108 7538
rect 5008 7504 5108 7528
rect 7098 7504 7194 7538
rect 5008 7288 7188 7504
rect 4009 6271 4043 6297
rect 5248 6296 5540 7288
rect 1297 6237 1357 6271
rect 3983 6237 4043 6271
rect 4808 6248 5540 6296
rect -9922 6192 -9906 6226
rect -9872 6192 -9856 6226
rect -9730 6192 -9714 6226
rect -9680 6192 -9664 6226
rect -9538 6192 -9522 6226
rect -9488 6192 -9472 6226
rect -9346 6192 -9330 6226
rect -9296 6192 -9280 6226
rect -9154 6192 -9138 6226
rect -9104 6192 -9088 6226
rect -10050 6142 -10016 6158
rect -10050 5750 -10016 5766
rect -9954 6142 -9920 6158
rect -9954 5750 -9920 5766
rect -9858 6142 -9824 6158
rect -9858 5750 -9824 5766
rect -9762 6142 -9728 6158
rect -9762 5750 -9728 5766
rect -9666 6142 -9632 6158
rect -9666 5750 -9632 5766
rect -9570 6142 -9536 6158
rect -9570 5750 -9536 5766
rect -9474 6142 -9440 6158
rect -9474 5750 -9440 5766
rect -9378 6142 -9344 6158
rect -9378 5750 -9344 5766
rect -9282 6142 -9248 6158
rect -9282 5750 -9248 5766
rect -9186 6142 -9152 6158
rect -9186 5750 -9152 5766
rect -9090 6142 -9056 6158
rect -9090 5750 -9056 5766
rect -10018 5682 -10002 5716
rect -9968 5682 -9952 5716
rect -9826 5682 -9810 5716
rect -9776 5682 -9760 5716
rect -9634 5682 -9618 5716
rect -9584 5682 -9568 5716
rect -9442 5682 -9426 5716
rect -9392 5682 -9376 5716
rect -9250 5682 -9234 5716
rect -9200 5682 -9184 5716
rect -10018 5574 -10002 5608
rect -9968 5574 -9952 5608
rect -9826 5574 -9810 5608
rect -9776 5574 -9760 5608
rect -9634 5574 -9618 5608
rect -9584 5574 -9568 5608
rect -9442 5574 -9426 5608
rect -9392 5574 -9376 5608
rect -9250 5574 -9234 5608
rect -9200 5574 -9184 5608
rect -10050 5524 -10016 5540
rect -10050 5132 -10016 5148
rect -9954 5524 -9920 5540
rect -9954 5132 -9920 5148
rect -9858 5524 -9824 5540
rect -9858 5132 -9824 5148
rect -9762 5524 -9728 5540
rect -9762 5132 -9728 5148
rect -9666 5524 -9632 5540
rect -9666 5132 -9632 5148
rect -9570 5524 -9536 5540
rect -9570 5132 -9536 5148
rect -9474 5524 -9440 5540
rect -9474 5132 -9440 5148
rect -9378 5524 -9344 5540
rect -9378 5132 -9344 5148
rect -9282 5524 -9248 5540
rect -9282 5132 -9248 5148
rect -9186 5524 -9152 5540
rect -9186 5132 -9152 5148
rect -9090 5524 -9056 5540
rect -9090 5132 -9056 5148
rect -9922 5064 -9906 5098
rect -9872 5064 -9856 5098
rect -9730 5064 -9714 5098
rect -9680 5064 -9664 5098
rect -9538 5064 -9522 5098
rect -9488 5064 -9472 5098
rect -9346 5064 -9330 5098
rect -9296 5064 -9280 5098
rect -9154 5064 -9138 5098
rect -9104 5064 -9088 5098
rect -9922 4956 -9906 4990
rect -9872 4956 -9856 4990
rect -9730 4956 -9714 4990
rect -9680 4956 -9664 4990
rect -9538 4956 -9522 4990
rect -9488 4956 -9472 4990
rect -9346 4956 -9330 4990
rect -9296 4956 -9280 4990
rect -9154 4956 -9138 4990
rect -9104 4956 -9088 4990
rect -10050 4906 -10016 4922
rect -10050 4514 -10016 4530
rect -9954 4906 -9920 4922
rect -9954 4514 -9920 4530
rect -9858 4906 -9824 4922
rect -9858 4514 -9824 4530
rect -9762 4906 -9728 4922
rect -9762 4514 -9728 4530
rect -9666 4906 -9632 4922
rect -9666 4514 -9632 4530
rect -9570 4906 -9536 4922
rect -9570 4514 -9536 4530
rect -9474 4906 -9440 4922
rect -9474 4514 -9440 4530
rect -9378 4906 -9344 4922
rect -9378 4514 -9344 4530
rect -9282 4906 -9248 4922
rect -9282 4514 -9248 4530
rect -9186 4906 -9152 4922
rect -9186 4514 -9152 4530
rect -9090 4906 -9056 4922
rect -9090 4514 -9056 4530
rect -10018 4446 -10002 4480
rect -9968 4446 -9952 4480
rect -9826 4446 -9810 4480
rect -9776 4446 -9760 4480
rect -9634 4446 -9618 4480
rect -9584 4446 -9568 4480
rect -9442 4446 -9426 4480
rect -9392 4446 -9376 4480
rect -9250 4446 -9234 4480
rect -9200 4446 -9184 4480
rect -10164 4378 -10130 4440
rect 4330 6048 5540 6248
rect -8976 4378 -8942 4440
rect -10164 4344 -10068 4378
rect -9038 4344 -8942 4378
rect 112 6014 208 6048
rect 1238 6014 2008 6048
rect 3038 6014 3808 6048
rect 4838 6036 5608 6048
rect 4838 6014 4934 6036
rect 112 5952 146 6014
rect -10140 4182 -10040 4344
rect -10164 4148 -10068 4182
rect -8708 4148 -8612 4182
rect -10164 4086 -10130 4148
rect -8646 4086 -8612 4148
rect -10004 4046 -9988 4080
rect -9820 4046 -9804 4080
rect -9746 4046 -9730 4080
rect -9562 4046 -9546 4080
rect -9488 4046 -9472 4080
rect -9304 4046 -9288 4080
rect -9230 4046 -9214 4080
rect -9046 4046 -9030 4080
rect -8972 4046 -8956 4080
rect -8788 4046 -8772 4080
rect -10050 3996 -10016 4012
rect -10050 3604 -10016 3620
rect -9792 3996 -9758 4012
rect -9792 3604 -9758 3620
rect -9534 3996 -9500 4012
rect -9534 3604 -9500 3620
rect -9276 3996 -9242 4012
rect -9276 3604 -9242 3620
rect -9018 3996 -8984 4012
rect -9018 3604 -8984 3620
rect -8760 3996 -8726 4012
rect -8760 3604 -8726 3620
rect -10004 3536 -9988 3570
rect -9820 3536 -9804 3570
rect -9746 3536 -9730 3570
rect -9562 3536 -9546 3570
rect -9488 3536 -9472 3570
rect -9304 3536 -9288 3570
rect -9230 3536 -9214 3570
rect -9046 3536 -9030 3570
rect -8972 3536 -8956 3570
rect -8788 3536 -8772 3570
rect -10004 3428 -9988 3462
rect -9820 3428 -9804 3462
rect -9746 3428 -9730 3462
rect -9562 3428 -9546 3462
rect -9488 3428 -9472 3462
rect -9304 3428 -9288 3462
rect -9230 3428 -9214 3462
rect -9046 3428 -9030 3462
rect -8972 3428 -8956 3462
rect -8788 3428 -8772 3462
rect -10050 3378 -10016 3394
rect -10050 2986 -10016 3002
rect -9792 3378 -9758 3394
rect -9792 2986 -9758 3002
rect -9534 3378 -9500 3394
rect -9534 2986 -9500 3002
rect -9276 3378 -9242 3394
rect -9276 2986 -9242 3002
rect -9018 3378 -8984 3394
rect -9018 2986 -8984 3002
rect -8760 3378 -8726 3394
rect -8760 2986 -8726 3002
rect -10004 2918 -9988 2952
rect -9820 2918 -9804 2952
rect -9746 2918 -9730 2952
rect -9562 2918 -9546 2952
rect -9488 2918 -9472 2952
rect -9304 2918 -9288 2952
rect -9230 2918 -9214 2952
rect -9046 2918 -9030 2952
rect -8972 2918 -8956 2952
rect -8788 2918 -8772 2952
rect -10004 2810 -9988 2844
rect -9820 2810 -9804 2844
rect -9746 2810 -9730 2844
rect -9562 2810 -9546 2844
rect -9488 2810 -9472 2844
rect -9304 2810 -9288 2844
rect -9230 2810 -9214 2844
rect -9046 2810 -9030 2844
rect -8972 2810 -8956 2844
rect -8788 2810 -8772 2844
rect -10050 2760 -10016 2776
rect -10050 2368 -10016 2384
rect -9792 2760 -9758 2776
rect -9792 2368 -9758 2384
rect -9534 2760 -9500 2776
rect -9534 2368 -9500 2384
rect -9276 2760 -9242 2776
rect -9276 2368 -9242 2384
rect -9018 2760 -8984 2776
rect -9018 2368 -8984 2384
rect -8760 2760 -8726 2776
rect -8760 2368 -8726 2384
rect -10004 2300 -9988 2334
rect -9820 2300 -9804 2334
rect -9746 2300 -9730 2334
rect -9562 2300 -9546 2334
rect -9488 2300 -9472 2334
rect -9304 2300 -9288 2334
rect -9230 2300 -9214 2334
rect -9046 2300 -9030 2334
rect -8972 2300 -8956 2334
rect -8788 2300 -8772 2334
rect -10004 2192 -9988 2226
rect -9820 2192 -9804 2226
rect -9746 2192 -9730 2226
rect -9562 2192 -9546 2226
rect -9488 2192 -9472 2226
rect -9304 2192 -9288 2226
rect -9230 2192 -9214 2226
rect -9046 2192 -9030 2226
rect -8972 2192 -8956 2226
rect -8788 2192 -8772 2226
rect -10050 2142 -10016 2158
rect -10050 1750 -10016 1766
rect -9792 2142 -9758 2158
rect -9792 1750 -9758 1766
rect -9534 2142 -9500 2158
rect -9534 1750 -9500 1766
rect -9276 2142 -9242 2158
rect -9276 1750 -9242 1766
rect -9018 2142 -8984 2158
rect -9018 1750 -8984 1766
rect -8760 2142 -8726 2158
rect -8760 1750 -8726 1766
rect -10004 1682 -9988 1716
rect -9820 1682 -9804 1716
rect -9746 1682 -9730 1716
rect -9562 1682 -9546 1716
rect -9488 1682 -9472 1716
rect -9304 1682 -9288 1716
rect -9230 1682 -9214 1716
rect -9046 1682 -9030 1716
rect -8972 1682 -8956 1716
rect -8788 1682 -8772 1716
rect -10004 1574 -9988 1608
rect -9820 1574 -9804 1608
rect -9746 1574 -9730 1608
rect -9562 1574 -9546 1608
rect -9488 1574 -9472 1608
rect -9304 1574 -9288 1608
rect -9230 1574 -9214 1608
rect -9046 1574 -9030 1608
rect -8972 1574 -8956 1608
rect -8788 1574 -8772 1608
rect -10050 1524 -10016 1540
rect -10050 1132 -10016 1148
rect -9792 1524 -9758 1540
rect -9792 1132 -9758 1148
rect -9534 1524 -9500 1540
rect -9534 1132 -9500 1148
rect -9276 1524 -9242 1540
rect -9276 1132 -9242 1148
rect -9018 1524 -8984 1540
rect -9018 1132 -8984 1148
rect -8760 1524 -8726 1540
rect -8760 1132 -8726 1148
rect -10004 1064 -9988 1098
rect -9820 1064 -9804 1098
rect -9746 1064 -9730 1098
rect -9562 1064 -9546 1098
rect -9488 1064 -9472 1098
rect -9304 1064 -9288 1098
rect -9230 1064 -9214 1098
rect -9046 1064 -9030 1098
rect -8972 1064 -8956 1098
rect -8788 1064 -8772 1098
rect -10004 956 -9988 990
rect -9820 956 -9804 990
rect -9746 956 -9730 990
rect -9562 956 -9546 990
rect -9488 956 -9472 990
rect -9304 956 -9288 990
rect -9230 956 -9214 990
rect -9046 956 -9030 990
rect -8972 956 -8956 990
rect -8788 956 -8772 990
rect -10050 906 -10016 922
rect -10050 514 -10016 530
rect -9792 906 -9758 922
rect -9792 514 -9758 530
rect -9534 906 -9500 922
rect -9534 514 -9500 530
rect -9276 906 -9242 922
rect -9276 514 -9242 530
rect -9018 906 -8984 922
rect -9018 514 -8984 530
rect -8760 906 -8726 922
rect -8760 514 -8726 530
rect -10004 446 -9988 480
rect -9820 446 -9804 480
rect -9746 446 -9730 480
rect -9562 446 -9546 480
rect -9488 446 -9472 480
rect -9304 446 -9288 480
rect -9230 446 -9214 480
rect -9046 446 -9030 480
rect -8972 446 -8956 480
rect -8788 446 -8772 480
rect -10164 378 -10130 440
rect 1300 5952 1946 6014
rect 354 5912 370 5946
rect 404 5912 420 5946
rect 546 5912 562 5946
rect 596 5912 612 5946
rect 738 5912 754 5946
rect 788 5912 804 5946
rect 930 5912 946 5946
rect 980 5912 996 5946
rect 1122 5912 1138 5946
rect 1172 5912 1188 5946
rect 226 5862 260 5878
rect 226 5470 260 5486
rect 322 5862 356 5878
rect 322 5470 356 5486
rect 418 5862 452 5878
rect 418 5470 452 5486
rect 514 5862 548 5878
rect 514 5470 548 5486
rect 610 5862 644 5878
rect 610 5470 644 5486
rect 706 5862 740 5878
rect 706 5470 740 5486
rect 802 5862 836 5878
rect 802 5470 836 5486
rect 898 5862 932 5878
rect 898 5470 932 5486
rect 994 5862 1028 5878
rect 994 5470 1028 5486
rect 1090 5862 1124 5878
rect 1090 5470 1124 5486
rect 1186 5862 1220 5878
rect 1186 5470 1220 5486
rect 258 5402 274 5436
rect 308 5402 324 5436
rect 450 5402 466 5436
rect 500 5402 516 5436
rect 642 5402 658 5436
rect 692 5402 708 5436
rect 834 5402 850 5436
rect 884 5402 900 5436
rect 1026 5402 1042 5436
rect 1076 5402 1092 5436
rect 258 5294 274 5328
rect 308 5294 324 5328
rect 450 5294 466 5328
rect 500 5294 516 5328
rect 642 5294 658 5328
rect 692 5294 708 5328
rect 834 5294 850 5328
rect 884 5294 900 5328
rect 1026 5294 1042 5328
rect 1076 5294 1092 5328
rect 226 5244 260 5260
rect 226 4852 260 4868
rect 322 5244 356 5260
rect 322 4852 356 4868
rect 418 5244 452 5260
rect 418 4852 452 4868
rect 514 5244 548 5260
rect 514 4852 548 4868
rect 610 5244 644 5260
rect 610 4852 644 4868
rect 706 5244 740 5260
rect 706 4852 740 4868
rect 802 5244 836 5260
rect 802 4852 836 4868
rect 898 5244 932 5260
rect 898 4852 932 4868
rect 994 5244 1028 5260
rect 994 4852 1028 4868
rect 1090 5244 1124 5260
rect 1090 4852 1124 4868
rect 1186 5244 1220 5260
rect 1186 4852 1220 4868
rect 354 4784 370 4818
rect 404 4784 420 4818
rect 546 4784 562 4818
rect 596 4784 612 4818
rect 738 4784 754 4818
rect 788 4784 804 4818
rect 930 4784 946 4818
rect 980 4784 996 4818
rect 1122 4784 1138 4818
rect 1172 4784 1188 4818
rect 354 4676 370 4710
rect 404 4676 420 4710
rect 546 4676 562 4710
rect 596 4676 612 4710
rect 738 4676 754 4710
rect 788 4676 804 4710
rect 930 4676 946 4710
rect 980 4676 996 4710
rect 1122 4676 1138 4710
rect 1172 4676 1188 4710
rect 226 4626 260 4642
rect 226 4234 260 4250
rect 322 4626 356 4642
rect 322 4234 356 4250
rect 418 4626 452 4642
rect 418 4234 452 4250
rect 514 4626 548 4642
rect 514 4234 548 4250
rect 610 4626 644 4642
rect 610 4234 644 4250
rect 706 4626 740 4642
rect 706 4234 740 4250
rect 802 4626 836 4642
rect 802 4234 836 4250
rect 898 4626 932 4642
rect 898 4234 932 4250
rect 994 4626 1028 4642
rect 994 4234 1028 4250
rect 1090 4626 1124 4642
rect 1090 4234 1124 4250
rect 1186 4626 1220 4642
rect 1186 4234 1220 4250
rect 258 4166 274 4200
rect 308 4166 324 4200
rect 450 4166 466 4200
rect 500 4166 516 4200
rect 642 4166 658 4200
rect 692 4166 708 4200
rect 834 4166 850 4200
rect 884 4166 900 4200
rect 1026 4166 1042 4200
rect 1076 4166 1092 4200
rect 112 4098 146 4160
rect 1334 5808 1912 5952
rect 1300 4098 1334 4160
rect 112 4064 208 4098
rect 1238 4064 1334 4098
rect 1640 4160 1912 5808
rect 3100 5952 3746 6014
rect 2154 5912 2170 5946
rect 2204 5912 2220 5946
rect 2346 5912 2362 5946
rect 2396 5912 2412 5946
rect 2538 5912 2554 5946
rect 2588 5912 2604 5946
rect 2730 5912 2746 5946
rect 2780 5912 2796 5946
rect 2922 5912 2938 5946
rect 2972 5912 2988 5946
rect 2026 5862 2060 5878
rect 2026 5470 2060 5486
rect 2122 5862 2156 5878
rect 2122 5470 2156 5486
rect 2218 5862 2252 5878
rect 2218 5470 2252 5486
rect 2314 5862 2348 5878
rect 2314 5470 2348 5486
rect 2410 5862 2444 5878
rect 2410 5470 2444 5486
rect 2506 5862 2540 5878
rect 2506 5470 2540 5486
rect 2602 5862 2636 5878
rect 2602 5470 2636 5486
rect 2698 5862 2732 5878
rect 2698 5470 2732 5486
rect 2794 5862 2828 5878
rect 2794 5470 2828 5486
rect 2890 5862 2924 5878
rect 2890 5470 2924 5486
rect 2986 5862 3020 5878
rect 2986 5470 3020 5486
rect 2058 5402 2074 5436
rect 2108 5402 2124 5436
rect 2250 5402 2266 5436
rect 2300 5402 2316 5436
rect 2442 5402 2458 5436
rect 2492 5402 2508 5436
rect 2634 5402 2650 5436
rect 2684 5402 2700 5436
rect 2826 5402 2842 5436
rect 2876 5402 2892 5436
rect 2058 5294 2074 5328
rect 2108 5294 2124 5328
rect 2250 5294 2266 5328
rect 2300 5294 2316 5328
rect 2442 5294 2458 5328
rect 2492 5294 2508 5328
rect 2634 5294 2650 5328
rect 2684 5294 2700 5328
rect 2826 5294 2842 5328
rect 2876 5294 2892 5328
rect 2026 5244 2060 5260
rect 2026 4852 2060 4868
rect 2122 5244 2156 5260
rect 2122 4852 2156 4868
rect 2218 5244 2252 5260
rect 2218 4852 2252 4868
rect 2314 5244 2348 5260
rect 2314 4852 2348 4868
rect 2410 5244 2444 5260
rect 2410 4852 2444 4868
rect 2506 5244 2540 5260
rect 2506 4852 2540 4868
rect 2602 5244 2636 5260
rect 2602 4852 2636 4868
rect 2698 5244 2732 5260
rect 2698 4852 2732 4868
rect 2794 5244 2828 5260
rect 2794 4852 2828 4868
rect 2890 5244 2924 5260
rect 2890 4852 2924 4868
rect 2986 5244 3020 5260
rect 2986 4852 3020 4868
rect 2154 4784 2170 4818
rect 2204 4784 2220 4818
rect 2346 4784 2362 4818
rect 2396 4784 2412 4818
rect 2538 4784 2554 4818
rect 2588 4784 2604 4818
rect 2730 4784 2746 4818
rect 2780 4784 2796 4818
rect 2922 4784 2938 4818
rect 2972 4784 2988 4818
rect 2154 4676 2170 4710
rect 2204 4676 2220 4710
rect 2346 4676 2362 4710
rect 2396 4676 2412 4710
rect 2538 4676 2554 4710
rect 2588 4676 2604 4710
rect 2730 4676 2746 4710
rect 2780 4676 2796 4710
rect 2922 4676 2938 4710
rect 2972 4676 2988 4710
rect 2026 4626 2060 4642
rect 2026 4234 2060 4250
rect 2122 4626 2156 4642
rect 2122 4234 2156 4250
rect 2218 4626 2252 4642
rect 2218 4234 2252 4250
rect 2314 4626 2348 4642
rect 2314 4234 2348 4250
rect 2410 4626 2444 4642
rect 2410 4234 2444 4250
rect 2506 4626 2540 4642
rect 2506 4234 2540 4250
rect 2602 4626 2636 4642
rect 2602 4234 2636 4250
rect 2698 4626 2732 4642
rect 2698 4234 2732 4250
rect 2794 4626 2828 4642
rect 2794 4234 2828 4250
rect 2890 4626 2924 4642
rect 2890 4234 2924 4250
rect 2986 4626 3020 4642
rect 2986 4234 3020 4250
rect 2058 4166 2074 4200
rect 2108 4166 2124 4200
rect 2250 4166 2266 4200
rect 2300 4166 2316 4200
rect 2442 4166 2458 4200
rect 2492 4166 2508 4200
rect 2634 4166 2650 4200
rect 2684 4166 2700 4200
rect 2826 4166 2842 4200
rect 2876 4166 2892 4200
rect 1640 4098 1946 4160
rect 3134 5808 3712 5952
rect 3100 4098 3134 4160
rect 1640 4064 2008 4098
rect 3038 4064 3134 4098
rect 3440 4160 3712 5808
rect 4900 5952 4934 6014
rect 3954 5912 3970 5946
rect 4004 5912 4020 5946
rect 4146 5912 4162 5946
rect 4196 5912 4212 5946
rect 4338 5912 4354 5946
rect 4388 5912 4404 5946
rect 4530 5912 4546 5946
rect 4580 5912 4596 5946
rect 4722 5912 4738 5946
rect 4772 5912 4788 5946
rect 3826 5862 3860 5878
rect 3826 5470 3860 5486
rect 3922 5862 3956 5878
rect 3922 5470 3956 5486
rect 4018 5862 4052 5878
rect 4018 5470 4052 5486
rect 4114 5862 4148 5878
rect 4114 5470 4148 5486
rect 4210 5862 4244 5878
rect 4210 5470 4244 5486
rect 4306 5862 4340 5878
rect 4306 5470 4340 5486
rect 4402 5862 4436 5878
rect 4402 5470 4436 5486
rect 4498 5862 4532 5878
rect 4498 5470 4532 5486
rect 4594 5862 4628 5878
rect 4594 5470 4628 5486
rect 4690 5862 4724 5878
rect 4690 5470 4724 5486
rect 4786 5862 4820 5878
rect 4786 5470 4820 5486
rect 3858 5402 3874 5436
rect 3908 5402 3924 5436
rect 4050 5402 4066 5436
rect 4100 5402 4116 5436
rect 4242 5402 4258 5436
rect 4292 5402 4308 5436
rect 4434 5402 4450 5436
rect 4484 5402 4500 5436
rect 4626 5402 4642 5436
rect 4676 5402 4692 5436
rect 3858 5294 3874 5328
rect 3908 5294 3924 5328
rect 4050 5294 4066 5328
rect 4100 5294 4116 5328
rect 4242 5294 4258 5328
rect 4292 5294 4308 5328
rect 4434 5294 4450 5328
rect 4484 5294 4500 5328
rect 4626 5294 4642 5328
rect 4676 5294 4692 5328
rect 3826 5244 3860 5260
rect 3826 4852 3860 4868
rect 3922 5244 3956 5260
rect 3922 4852 3956 4868
rect 4018 5244 4052 5260
rect 4018 4852 4052 4868
rect 4114 5244 4148 5260
rect 4114 4852 4148 4868
rect 4210 5244 4244 5260
rect 4210 4852 4244 4868
rect 4306 5244 4340 5260
rect 4306 4852 4340 4868
rect 4402 5244 4436 5260
rect 4402 4852 4436 4868
rect 4498 5244 4532 5260
rect 4498 4852 4532 4868
rect 4594 5244 4628 5260
rect 4594 4852 4628 4868
rect 4690 5244 4724 5260
rect 4690 4852 4724 4868
rect 4786 5244 4820 5260
rect 4786 4852 4820 4868
rect 3954 4784 3970 4818
rect 4004 4784 4020 4818
rect 4146 4784 4162 4818
rect 4196 4784 4212 4818
rect 4338 4784 4354 4818
rect 4388 4784 4404 4818
rect 4530 4784 4546 4818
rect 4580 4784 4596 4818
rect 4722 4784 4738 4818
rect 4772 4784 4788 4818
rect 3954 4676 3970 4710
rect 4004 4676 4020 4710
rect 4146 4676 4162 4710
rect 4196 4676 4212 4710
rect 4338 4676 4354 4710
rect 4388 4676 4404 4710
rect 4530 4676 4546 4710
rect 4580 4676 4596 4710
rect 4722 4676 4738 4710
rect 4772 4676 4788 4710
rect 3826 4626 3860 4642
rect 3826 4234 3860 4250
rect 3922 4626 3956 4642
rect 3922 4234 3956 4250
rect 4018 4626 4052 4642
rect 4018 4234 4052 4250
rect 4114 4626 4148 4642
rect 4114 4234 4148 4250
rect 4210 4626 4244 4642
rect 4210 4234 4244 4250
rect 4306 4626 4340 4642
rect 4306 4234 4340 4250
rect 4402 4626 4436 4642
rect 4402 4234 4436 4250
rect 4498 4626 4532 4642
rect 4498 4234 4532 4250
rect 4594 4626 4628 4642
rect 4594 4234 4628 4250
rect 4690 4626 4724 4642
rect 4690 4234 4724 4250
rect 4786 4626 4820 4642
rect 4786 4234 4820 4250
rect 3858 4166 3874 4200
rect 3908 4166 3924 4200
rect 4050 4166 4066 4200
rect 4100 4166 4116 4200
rect 4242 4166 4258 4200
rect 4292 4166 4308 4200
rect 4434 4166 4450 4200
rect 4484 4166 4500 4200
rect 4626 4166 4642 4200
rect 4676 4166 4692 4200
rect 3440 4098 3746 4160
rect 4900 4098 4934 4160
rect 3440 4064 3808 4098
rect 4838 4064 4934 4098
rect 5248 6014 5608 6036
rect 6638 6014 6734 6048
rect 5248 5952 5546 6014
rect 5248 4160 5512 5952
rect 6700 5952 6734 6014
rect 5754 5912 5770 5946
rect 5804 5912 5820 5946
rect 5946 5912 5962 5946
rect 5996 5912 6012 5946
rect 6138 5912 6154 5946
rect 6188 5912 6204 5946
rect 6330 5912 6346 5946
rect 6380 5912 6396 5946
rect 6522 5912 6538 5946
rect 6572 5912 6588 5946
rect 5626 5862 5660 5878
rect 5626 5470 5660 5486
rect 5722 5862 5756 5878
rect 5722 5470 5756 5486
rect 5818 5862 5852 5878
rect 5818 5470 5852 5486
rect 5914 5862 5948 5878
rect 5914 5470 5948 5486
rect 6010 5862 6044 5878
rect 6010 5470 6044 5486
rect 6106 5862 6140 5878
rect 6106 5470 6140 5486
rect 6202 5862 6236 5878
rect 6202 5470 6236 5486
rect 6298 5862 6332 5878
rect 6298 5470 6332 5486
rect 6394 5862 6428 5878
rect 6394 5470 6428 5486
rect 6490 5862 6524 5878
rect 6490 5470 6524 5486
rect 6586 5862 6620 5878
rect 6586 5470 6620 5486
rect 5658 5402 5674 5436
rect 5708 5402 5724 5436
rect 5850 5402 5866 5436
rect 5900 5402 5916 5436
rect 6042 5402 6058 5436
rect 6092 5402 6108 5436
rect 6234 5402 6250 5436
rect 6284 5402 6300 5436
rect 6426 5402 6442 5436
rect 6476 5402 6492 5436
rect 5658 5294 5674 5328
rect 5708 5294 5724 5328
rect 5850 5294 5866 5328
rect 5900 5294 5916 5328
rect 6042 5294 6058 5328
rect 6092 5294 6108 5328
rect 6234 5294 6250 5328
rect 6284 5294 6300 5328
rect 6426 5294 6442 5328
rect 6476 5294 6492 5328
rect 5626 5244 5660 5260
rect 5626 4852 5660 4868
rect 5722 5244 5756 5260
rect 5722 4852 5756 4868
rect 5818 5244 5852 5260
rect 5818 4852 5852 4868
rect 5914 5244 5948 5260
rect 5914 4852 5948 4868
rect 6010 5244 6044 5260
rect 6010 4852 6044 4868
rect 6106 5244 6140 5260
rect 6106 4852 6140 4868
rect 6202 5244 6236 5260
rect 6202 4852 6236 4868
rect 6298 5244 6332 5260
rect 6298 4852 6332 4868
rect 6394 5244 6428 5260
rect 6394 4852 6428 4868
rect 6490 5244 6524 5260
rect 6490 4852 6524 4868
rect 6586 5244 6620 5260
rect 6586 4852 6620 4868
rect 5754 4784 5770 4818
rect 5804 4784 5820 4818
rect 5946 4784 5962 4818
rect 5996 4784 6012 4818
rect 6138 4784 6154 4818
rect 6188 4784 6204 4818
rect 6330 4784 6346 4818
rect 6380 4784 6396 4818
rect 6522 4784 6538 4818
rect 6572 4784 6588 4818
rect 5754 4676 5770 4710
rect 5804 4676 5820 4710
rect 5946 4676 5962 4710
rect 5996 4676 6012 4710
rect 6138 4676 6154 4710
rect 6188 4676 6204 4710
rect 6330 4676 6346 4710
rect 6380 4676 6396 4710
rect 6522 4676 6538 4710
rect 6572 4676 6588 4710
rect 5626 4626 5660 4642
rect 5626 4234 5660 4250
rect 5722 4626 5756 4642
rect 5722 4234 5756 4250
rect 5818 4626 5852 4642
rect 5818 4234 5852 4250
rect 5914 4626 5948 4642
rect 5914 4234 5948 4250
rect 6010 4626 6044 4642
rect 6010 4234 6044 4250
rect 6106 4626 6140 4642
rect 6106 4234 6140 4250
rect 6202 4626 6236 4642
rect 6202 4234 6236 4250
rect 6298 4626 6332 4642
rect 6298 4234 6332 4250
rect 6394 4626 6428 4642
rect 6394 4234 6428 4250
rect 6490 4626 6524 4642
rect 6490 4234 6524 4250
rect 6586 4626 6620 4642
rect 6586 4234 6620 4250
rect 5658 4166 5674 4200
rect 5708 4166 5724 4200
rect 5850 4166 5866 4200
rect 5900 4166 5916 4200
rect 6042 4166 6058 4200
rect 6092 4166 6108 4200
rect 6234 4166 6250 4200
rect 6284 4166 6300 4200
rect 6426 4166 6442 4200
rect 6476 4166 6492 4200
rect 5248 4098 5546 4160
rect 6734 4988 7512 5188
rect 9660 10340 9694 10402
rect 7754 10300 7770 10334
rect 7804 10300 7820 10334
rect 7946 10300 7962 10334
rect 7996 10300 8012 10334
rect 8138 10300 8154 10334
rect 8188 10300 8204 10334
rect 8330 10300 8346 10334
rect 8380 10300 8396 10334
rect 8522 10300 8538 10334
rect 8572 10300 8588 10334
rect 8714 10300 8730 10334
rect 8764 10300 8780 10334
rect 8906 10300 8922 10334
rect 8956 10300 8972 10334
rect 9098 10300 9114 10334
rect 9148 10300 9164 10334
rect 9290 10300 9306 10334
rect 9340 10300 9356 10334
rect 9482 10300 9498 10334
rect 9532 10300 9548 10334
rect 7626 10250 7660 10266
rect 7626 9858 7660 9874
rect 7722 10250 7756 10266
rect 7722 9858 7756 9874
rect 7818 10250 7852 10266
rect 7818 9858 7852 9874
rect 7914 10250 7948 10266
rect 7914 9858 7948 9874
rect 8010 10250 8044 10266
rect 8010 9858 8044 9874
rect 8106 10250 8140 10266
rect 8106 9858 8140 9874
rect 8202 10250 8236 10266
rect 8202 9858 8236 9874
rect 8298 10250 8332 10266
rect 8298 9858 8332 9874
rect 8394 10250 8428 10266
rect 8394 9858 8428 9874
rect 8490 10250 8524 10266
rect 8490 9858 8524 9874
rect 8586 10250 8620 10266
rect 8586 9858 8620 9874
rect 8682 10250 8716 10266
rect 8682 9858 8716 9874
rect 8778 10250 8812 10266
rect 8778 9858 8812 9874
rect 8874 10250 8908 10266
rect 8874 9858 8908 9874
rect 8970 10250 9004 10266
rect 8970 9858 9004 9874
rect 9066 10250 9100 10266
rect 9066 9858 9100 9874
rect 9162 10250 9196 10266
rect 9162 9858 9196 9874
rect 9258 10250 9292 10266
rect 9258 9858 9292 9874
rect 9354 10250 9388 10266
rect 9354 9858 9388 9874
rect 9450 10250 9484 10266
rect 9450 9858 9484 9874
rect 9546 10250 9580 10266
rect 9546 9858 9580 9874
rect 7658 9790 7674 9824
rect 7708 9790 7724 9824
rect 7850 9790 7866 9824
rect 7900 9790 7916 9824
rect 8042 9790 8058 9824
rect 8092 9790 8108 9824
rect 8234 9790 8250 9824
rect 8284 9790 8300 9824
rect 8426 9790 8442 9824
rect 8476 9790 8492 9824
rect 8618 9790 8634 9824
rect 8668 9790 8684 9824
rect 8810 9790 8826 9824
rect 8860 9790 8876 9824
rect 9002 9790 9018 9824
rect 9052 9790 9068 9824
rect 9194 9790 9210 9824
rect 9244 9790 9260 9824
rect 9386 9790 9402 9824
rect 9436 9790 9452 9824
rect 7658 9682 7674 9716
rect 7708 9682 7724 9716
rect 7850 9682 7866 9716
rect 7900 9682 7916 9716
rect 8042 9682 8058 9716
rect 8092 9682 8108 9716
rect 8234 9682 8250 9716
rect 8284 9682 8300 9716
rect 8426 9682 8442 9716
rect 8476 9682 8492 9716
rect 8618 9682 8634 9716
rect 8668 9682 8684 9716
rect 8810 9682 8826 9716
rect 8860 9682 8876 9716
rect 9002 9682 9018 9716
rect 9052 9682 9068 9716
rect 9194 9682 9210 9716
rect 9244 9682 9260 9716
rect 9386 9682 9402 9716
rect 9436 9682 9452 9716
rect 7626 9632 7660 9648
rect 7626 9240 7660 9256
rect 7722 9632 7756 9648
rect 7722 9240 7756 9256
rect 7818 9632 7852 9648
rect 7818 9240 7852 9256
rect 7914 9632 7948 9648
rect 7914 9240 7948 9256
rect 8010 9632 8044 9648
rect 8010 9240 8044 9256
rect 8106 9632 8140 9648
rect 8106 9240 8140 9256
rect 8202 9632 8236 9648
rect 8202 9240 8236 9256
rect 8298 9632 8332 9648
rect 8298 9240 8332 9256
rect 8394 9632 8428 9648
rect 8394 9240 8428 9256
rect 8490 9632 8524 9648
rect 8490 9240 8524 9256
rect 8586 9632 8620 9648
rect 8586 9240 8620 9256
rect 8682 9632 8716 9648
rect 8682 9240 8716 9256
rect 8778 9632 8812 9648
rect 8778 9240 8812 9256
rect 8874 9632 8908 9648
rect 8874 9240 8908 9256
rect 8970 9632 9004 9648
rect 8970 9240 9004 9256
rect 9066 9632 9100 9648
rect 9066 9240 9100 9256
rect 9162 9632 9196 9648
rect 9162 9240 9196 9256
rect 9258 9632 9292 9648
rect 9258 9240 9292 9256
rect 9354 9632 9388 9648
rect 9354 9240 9388 9256
rect 9450 9632 9484 9648
rect 9450 9240 9484 9256
rect 9546 9632 9580 9648
rect 9546 9240 9580 9256
rect 7754 9172 7770 9206
rect 7804 9172 7820 9206
rect 7946 9172 7962 9206
rect 7996 9172 8012 9206
rect 8138 9172 8154 9206
rect 8188 9172 8204 9206
rect 8330 9172 8346 9206
rect 8380 9172 8396 9206
rect 8522 9172 8538 9206
rect 8572 9172 8588 9206
rect 8714 9172 8730 9206
rect 8764 9172 8780 9206
rect 8906 9172 8922 9206
rect 8956 9172 8972 9206
rect 9098 9172 9114 9206
rect 9148 9172 9164 9206
rect 9290 9172 9306 9206
rect 9340 9172 9356 9206
rect 9482 9172 9498 9206
rect 9532 9172 9548 9206
rect 7754 9064 7770 9098
rect 7804 9064 7820 9098
rect 7946 9064 7962 9098
rect 7996 9064 8012 9098
rect 8138 9064 8154 9098
rect 8188 9064 8204 9098
rect 8330 9064 8346 9098
rect 8380 9064 8396 9098
rect 8522 9064 8538 9098
rect 8572 9064 8588 9098
rect 8714 9064 8730 9098
rect 8764 9064 8780 9098
rect 8906 9064 8922 9098
rect 8956 9064 8972 9098
rect 9098 9064 9114 9098
rect 9148 9064 9164 9098
rect 9290 9064 9306 9098
rect 9340 9064 9356 9098
rect 9482 9064 9498 9098
rect 9532 9064 9548 9098
rect 7626 9014 7660 9030
rect 7626 8622 7660 8638
rect 7722 9014 7756 9030
rect 7722 8622 7756 8638
rect 7818 9014 7852 9030
rect 7818 8622 7852 8638
rect 7914 9014 7948 9030
rect 7914 8622 7948 8638
rect 8010 9014 8044 9030
rect 8010 8622 8044 8638
rect 8106 9014 8140 9030
rect 8106 8622 8140 8638
rect 8202 9014 8236 9030
rect 8202 8622 8236 8638
rect 8298 9014 8332 9030
rect 8298 8622 8332 8638
rect 8394 9014 8428 9030
rect 8394 8622 8428 8638
rect 8490 9014 8524 9030
rect 8490 8622 8524 8638
rect 8586 9014 8620 9030
rect 8586 8622 8620 8638
rect 8682 9014 8716 9030
rect 8682 8622 8716 8638
rect 8778 9014 8812 9030
rect 8778 8622 8812 8638
rect 8874 9014 8908 9030
rect 8874 8622 8908 8638
rect 8970 9014 9004 9030
rect 8970 8622 9004 8638
rect 9066 9014 9100 9030
rect 9066 8622 9100 8638
rect 9162 9014 9196 9030
rect 9162 8622 9196 8638
rect 9258 9014 9292 9030
rect 9258 8622 9292 8638
rect 9354 9014 9388 9030
rect 9354 8622 9388 8638
rect 9450 9014 9484 9030
rect 9450 8622 9484 8638
rect 9546 9014 9580 9030
rect 9546 8622 9580 8638
rect 7658 8554 7674 8588
rect 7708 8554 7724 8588
rect 7850 8554 7866 8588
rect 7900 8554 7916 8588
rect 8042 8554 8058 8588
rect 8092 8554 8108 8588
rect 8234 8554 8250 8588
rect 8284 8554 8300 8588
rect 8426 8554 8442 8588
rect 8476 8554 8492 8588
rect 8618 8554 8634 8588
rect 8668 8554 8684 8588
rect 8810 8554 8826 8588
rect 8860 8554 8876 8588
rect 9002 8554 9018 8588
rect 9052 8554 9068 8588
rect 9194 8554 9210 8588
rect 9244 8554 9260 8588
rect 9386 8554 9402 8588
rect 9436 8554 9452 8588
rect 7658 8446 7674 8480
rect 7708 8446 7724 8480
rect 7850 8446 7866 8480
rect 7900 8446 7916 8480
rect 8042 8446 8058 8480
rect 8092 8446 8108 8480
rect 8234 8446 8250 8480
rect 8284 8446 8300 8480
rect 8426 8446 8442 8480
rect 8476 8446 8492 8480
rect 8618 8446 8634 8480
rect 8668 8446 8684 8480
rect 8810 8446 8826 8480
rect 8860 8446 8876 8480
rect 9002 8446 9018 8480
rect 9052 8446 9068 8480
rect 9194 8446 9210 8480
rect 9244 8446 9260 8480
rect 9386 8446 9402 8480
rect 9436 8446 9452 8480
rect 7626 8396 7660 8412
rect 7626 8004 7660 8020
rect 7722 8396 7756 8412
rect 7722 8004 7756 8020
rect 7818 8396 7852 8412
rect 7818 8004 7852 8020
rect 7914 8396 7948 8412
rect 7914 8004 7948 8020
rect 8010 8396 8044 8412
rect 8010 8004 8044 8020
rect 8106 8396 8140 8412
rect 8106 8004 8140 8020
rect 8202 8396 8236 8412
rect 8202 8004 8236 8020
rect 8298 8396 8332 8412
rect 8298 8004 8332 8020
rect 8394 8396 8428 8412
rect 8394 8004 8428 8020
rect 8490 8396 8524 8412
rect 8490 8004 8524 8020
rect 8586 8396 8620 8412
rect 8586 8004 8620 8020
rect 8682 8396 8716 8412
rect 8682 8004 8716 8020
rect 8778 8396 8812 8412
rect 8778 8004 8812 8020
rect 8874 8396 8908 8412
rect 8874 8004 8908 8020
rect 8970 8396 9004 8412
rect 8970 8004 9004 8020
rect 9066 8396 9100 8412
rect 9066 8004 9100 8020
rect 9162 8396 9196 8412
rect 9162 8004 9196 8020
rect 9258 8396 9292 8412
rect 9258 8004 9292 8020
rect 9354 8396 9388 8412
rect 9354 8004 9388 8020
rect 9450 8396 9484 8412
rect 9450 8004 9484 8020
rect 9546 8396 9580 8412
rect 9546 8004 9580 8020
rect 7754 7936 7770 7970
rect 7804 7936 7820 7970
rect 7946 7936 7962 7970
rect 7996 7936 8012 7970
rect 8138 7936 8154 7970
rect 8188 7936 8204 7970
rect 8330 7936 8346 7970
rect 8380 7936 8396 7970
rect 8522 7936 8538 7970
rect 8572 7936 8588 7970
rect 8714 7936 8730 7970
rect 8764 7936 8780 7970
rect 8906 7936 8922 7970
rect 8956 7936 8972 7970
rect 9098 7936 9114 7970
rect 9148 7936 9164 7970
rect 9290 7936 9306 7970
rect 9340 7936 9356 7970
rect 9482 7936 9498 7970
rect 9532 7936 9548 7970
rect 7754 7828 7770 7862
rect 7804 7828 7820 7862
rect 7946 7828 7962 7862
rect 7996 7828 8012 7862
rect 8138 7828 8154 7862
rect 8188 7828 8204 7862
rect 8330 7828 8346 7862
rect 8380 7828 8396 7862
rect 8522 7828 8538 7862
rect 8572 7828 8588 7862
rect 8714 7828 8730 7862
rect 8764 7828 8780 7862
rect 8906 7828 8922 7862
rect 8956 7828 8972 7862
rect 9098 7828 9114 7862
rect 9148 7828 9164 7862
rect 9290 7828 9306 7862
rect 9340 7828 9356 7862
rect 9482 7828 9498 7862
rect 9532 7828 9548 7862
rect 7626 7778 7660 7794
rect 7626 7386 7660 7402
rect 7722 7778 7756 7794
rect 7722 7386 7756 7402
rect 7818 7778 7852 7794
rect 7818 7386 7852 7402
rect 7914 7778 7948 7794
rect 7914 7386 7948 7402
rect 8010 7778 8044 7794
rect 8010 7386 8044 7402
rect 8106 7778 8140 7794
rect 8106 7386 8140 7402
rect 8202 7778 8236 7794
rect 8202 7386 8236 7402
rect 8298 7778 8332 7794
rect 8298 7386 8332 7402
rect 8394 7778 8428 7794
rect 8394 7386 8428 7402
rect 8490 7778 8524 7794
rect 8490 7386 8524 7402
rect 8586 7778 8620 7794
rect 8586 7386 8620 7402
rect 8682 7778 8716 7794
rect 8682 7386 8716 7402
rect 8778 7778 8812 7794
rect 8778 7386 8812 7402
rect 8874 7778 8908 7794
rect 8874 7386 8908 7402
rect 8970 7778 9004 7794
rect 8970 7386 9004 7402
rect 9066 7778 9100 7794
rect 9066 7386 9100 7402
rect 9162 7778 9196 7794
rect 9162 7386 9196 7402
rect 9258 7778 9292 7794
rect 9258 7386 9292 7402
rect 9354 7778 9388 7794
rect 9354 7386 9388 7402
rect 9450 7778 9484 7794
rect 9450 7386 9484 7402
rect 9546 7778 9580 7794
rect 9546 7386 9580 7402
rect 7658 7318 7674 7352
rect 7708 7318 7724 7352
rect 7850 7318 7866 7352
rect 7900 7318 7916 7352
rect 8042 7318 8058 7352
rect 8092 7318 8108 7352
rect 8234 7318 8250 7352
rect 8284 7318 8300 7352
rect 8426 7318 8442 7352
rect 8476 7318 8492 7352
rect 8618 7318 8634 7352
rect 8668 7318 8684 7352
rect 8810 7318 8826 7352
rect 8860 7318 8876 7352
rect 9002 7318 9018 7352
rect 9052 7318 9068 7352
rect 9194 7318 9210 7352
rect 9244 7318 9260 7352
rect 9386 7318 9402 7352
rect 9436 7318 9452 7352
rect 7658 7210 7674 7244
rect 7708 7210 7724 7244
rect 7850 7210 7866 7244
rect 7900 7210 7916 7244
rect 8042 7210 8058 7244
rect 8092 7210 8108 7244
rect 8234 7210 8250 7244
rect 8284 7210 8300 7244
rect 8426 7210 8442 7244
rect 8476 7210 8492 7244
rect 8618 7210 8634 7244
rect 8668 7210 8684 7244
rect 8810 7210 8826 7244
rect 8860 7210 8876 7244
rect 9002 7210 9018 7244
rect 9052 7210 9068 7244
rect 9194 7210 9210 7244
rect 9244 7210 9260 7244
rect 9386 7210 9402 7244
rect 9436 7210 9452 7244
rect 7626 7160 7660 7176
rect 7626 6768 7660 6784
rect 7722 7160 7756 7176
rect 7722 6768 7756 6784
rect 7818 7160 7852 7176
rect 7818 6768 7852 6784
rect 7914 7160 7948 7176
rect 7914 6768 7948 6784
rect 8010 7160 8044 7176
rect 8010 6768 8044 6784
rect 8106 7160 8140 7176
rect 8106 6768 8140 6784
rect 8202 7160 8236 7176
rect 8202 6768 8236 6784
rect 8298 7160 8332 7176
rect 8298 6768 8332 6784
rect 8394 7160 8428 7176
rect 8394 6768 8428 6784
rect 8490 7160 8524 7176
rect 8490 6768 8524 6784
rect 8586 7160 8620 7176
rect 8586 6768 8620 6784
rect 8682 7160 8716 7176
rect 8682 6768 8716 6784
rect 8778 7160 8812 7176
rect 8778 6768 8812 6784
rect 8874 7160 8908 7176
rect 8874 6768 8908 6784
rect 8970 7160 9004 7176
rect 8970 6768 9004 6784
rect 9066 7160 9100 7176
rect 9066 6768 9100 6784
rect 9162 7160 9196 7176
rect 9162 6768 9196 6784
rect 9258 7160 9292 7176
rect 9258 6768 9292 6784
rect 9354 7160 9388 7176
rect 9354 6768 9388 6784
rect 9450 7160 9484 7176
rect 9450 6768 9484 6784
rect 9546 7160 9580 7176
rect 9546 6768 9580 6784
rect 7754 6700 7770 6734
rect 7804 6700 7820 6734
rect 7946 6700 7962 6734
rect 7996 6700 8012 6734
rect 8138 6700 8154 6734
rect 8188 6700 8204 6734
rect 8330 6700 8346 6734
rect 8380 6700 8396 6734
rect 8522 6700 8538 6734
rect 8572 6700 8588 6734
rect 8714 6700 8730 6734
rect 8764 6700 8780 6734
rect 8906 6700 8922 6734
rect 8956 6700 8972 6734
rect 9098 6700 9114 6734
rect 9148 6700 9164 6734
rect 9290 6700 9306 6734
rect 9340 6700 9356 6734
rect 9482 6700 9498 6734
rect 9532 6700 9548 6734
rect 7754 6592 7770 6626
rect 7804 6592 7820 6626
rect 7946 6592 7962 6626
rect 7996 6592 8012 6626
rect 8138 6592 8154 6626
rect 8188 6592 8204 6626
rect 8330 6592 8346 6626
rect 8380 6592 8396 6626
rect 8522 6592 8538 6626
rect 8572 6592 8588 6626
rect 8714 6592 8730 6626
rect 8764 6592 8780 6626
rect 8906 6592 8922 6626
rect 8956 6592 8972 6626
rect 9098 6592 9114 6626
rect 9148 6592 9164 6626
rect 9290 6592 9306 6626
rect 9340 6592 9356 6626
rect 9482 6592 9498 6626
rect 9532 6592 9548 6626
rect 7626 6542 7660 6558
rect 7626 6150 7660 6166
rect 7722 6542 7756 6558
rect 7722 6150 7756 6166
rect 7818 6542 7852 6558
rect 7818 6150 7852 6166
rect 7914 6542 7948 6558
rect 7914 6150 7948 6166
rect 8010 6542 8044 6558
rect 8010 6150 8044 6166
rect 8106 6542 8140 6558
rect 8106 6150 8140 6166
rect 8202 6542 8236 6558
rect 8202 6150 8236 6166
rect 8298 6542 8332 6558
rect 8298 6150 8332 6166
rect 8394 6542 8428 6558
rect 8394 6150 8428 6166
rect 8490 6542 8524 6558
rect 8490 6150 8524 6166
rect 8586 6542 8620 6558
rect 8586 6150 8620 6166
rect 8682 6542 8716 6558
rect 8682 6150 8716 6166
rect 8778 6542 8812 6558
rect 8778 6150 8812 6166
rect 8874 6542 8908 6558
rect 8874 6150 8908 6166
rect 8970 6542 9004 6558
rect 8970 6150 9004 6166
rect 9066 6542 9100 6558
rect 9066 6150 9100 6166
rect 9162 6542 9196 6558
rect 9162 6150 9196 6166
rect 9258 6542 9292 6558
rect 9258 6150 9292 6166
rect 9354 6542 9388 6558
rect 9354 6150 9388 6166
rect 9450 6542 9484 6558
rect 9450 6150 9484 6166
rect 9546 6542 9580 6558
rect 9546 6150 9580 6166
rect 7658 6082 7674 6116
rect 7708 6082 7724 6116
rect 7850 6082 7866 6116
rect 7900 6082 7916 6116
rect 8042 6082 8058 6116
rect 8092 6082 8108 6116
rect 8234 6082 8250 6116
rect 8284 6082 8300 6116
rect 8426 6082 8442 6116
rect 8476 6082 8492 6116
rect 8618 6082 8634 6116
rect 8668 6082 8684 6116
rect 8810 6082 8826 6116
rect 8860 6082 8876 6116
rect 9002 6082 9018 6116
rect 9052 6082 9068 6116
rect 9194 6082 9210 6116
rect 9244 6082 9260 6116
rect 9386 6082 9402 6116
rect 9436 6082 9452 6116
rect 7658 5974 7674 6008
rect 7708 5974 7724 6008
rect 7850 5974 7866 6008
rect 7900 5974 7916 6008
rect 8042 5974 8058 6008
rect 8092 5974 8108 6008
rect 8234 5974 8250 6008
rect 8284 5974 8300 6008
rect 8426 5974 8442 6008
rect 8476 5974 8492 6008
rect 8618 5974 8634 6008
rect 8668 5974 8684 6008
rect 8810 5974 8826 6008
rect 8860 5974 8876 6008
rect 9002 5974 9018 6008
rect 9052 5974 9068 6008
rect 9194 5974 9210 6008
rect 9244 5974 9260 6008
rect 9386 5974 9402 6008
rect 9436 5974 9452 6008
rect 7626 5924 7660 5940
rect 7626 5532 7660 5548
rect 7722 5924 7756 5940
rect 7722 5532 7756 5548
rect 7818 5924 7852 5940
rect 7818 5532 7852 5548
rect 7914 5924 7948 5940
rect 7914 5532 7948 5548
rect 8010 5924 8044 5940
rect 8010 5532 8044 5548
rect 8106 5924 8140 5940
rect 8106 5532 8140 5548
rect 8202 5924 8236 5940
rect 8202 5532 8236 5548
rect 8298 5924 8332 5940
rect 8298 5532 8332 5548
rect 8394 5924 8428 5940
rect 8394 5532 8428 5548
rect 8490 5924 8524 5940
rect 8490 5532 8524 5548
rect 8586 5924 8620 5940
rect 8586 5532 8620 5548
rect 8682 5924 8716 5940
rect 8682 5532 8716 5548
rect 8778 5924 8812 5940
rect 8778 5532 8812 5548
rect 8874 5924 8908 5940
rect 8874 5532 8908 5548
rect 8970 5924 9004 5940
rect 8970 5532 9004 5548
rect 9066 5924 9100 5940
rect 9066 5532 9100 5548
rect 9162 5924 9196 5940
rect 9162 5532 9196 5548
rect 9258 5924 9292 5940
rect 9258 5532 9292 5548
rect 9354 5924 9388 5940
rect 9354 5532 9388 5548
rect 9450 5924 9484 5940
rect 9450 5532 9484 5548
rect 9546 5924 9580 5940
rect 9546 5532 9580 5548
rect 7754 5464 7770 5498
rect 7804 5464 7820 5498
rect 7946 5464 7962 5498
rect 7996 5464 8012 5498
rect 8138 5464 8154 5498
rect 8188 5464 8204 5498
rect 8330 5464 8346 5498
rect 8380 5464 8396 5498
rect 8522 5464 8538 5498
rect 8572 5464 8588 5498
rect 8714 5464 8730 5498
rect 8764 5464 8780 5498
rect 8906 5464 8922 5498
rect 8956 5464 8972 5498
rect 9098 5464 9114 5498
rect 9148 5464 9164 5498
rect 9290 5464 9306 5498
rect 9340 5464 9356 5498
rect 9482 5464 9498 5498
rect 9532 5464 9548 5498
rect 7754 5356 7770 5390
rect 7804 5356 7820 5390
rect 7946 5356 7962 5390
rect 7996 5356 8012 5390
rect 8138 5356 8154 5390
rect 8188 5356 8204 5390
rect 8330 5356 8346 5390
rect 8380 5356 8396 5390
rect 8522 5356 8538 5390
rect 8572 5356 8588 5390
rect 8714 5356 8730 5390
rect 8764 5356 8780 5390
rect 8906 5356 8922 5390
rect 8956 5356 8972 5390
rect 9098 5356 9114 5390
rect 9148 5356 9164 5390
rect 9290 5356 9306 5390
rect 9340 5356 9356 5390
rect 9482 5356 9498 5390
rect 9532 5356 9548 5390
rect 7626 5306 7660 5322
rect 7626 4914 7660 4930
rect 7722 5306 7756 5322
rect 7722 4914 7756 4930
rect 7818 5306 7852 5322
rect 7818 4914 7852 4930
rect 7914 5306 7948 5322
rect 7914 4914 7948 4930
rect 8010 5306 8044 5322
rect 8010 4914 8044 4930
rect 8106 5306 8140 5322
rect 8106 4914 8140 4930
rect 8202 5306 8236 5322
rect 8202 4914 8236 4930
rect 8298 5306 8332 5322
rect 8298 4914 8332 4930
rect 8394 5306 8428 5322
rect 8394 4914 8428 4930
rect 8490 5306 8524 5322
rect 8490 4914 8524 4930
rect 8586 5306 8620 5322
rect 8586 4914 8620 4930
rect 8682 5306 8716 5322
rect 8682 4914 8716 4930
rect 8778 5306 8812 5322
rect 8778 4914 8812 4930
rect 8874 5306 8908 5322
rect 8874 4914 8908 4930
rect 8970 5306 9004 5322
rect 8970 4914 9004 4930
rect 9066 5306 9100 5322
rect 9066 4914 9100 4930
rect 9162 5306 9196 5322
rect 9162 4914 9196 4930
rect 9258 5306 9292 5322
rect 9258 4914 9292 4930
rect 9354 5306 9388 5322
rect 9354 4914 9388 4930
rect 9450 5306 9484 5322
rect 9450 4914 9484 4930
rect 9546 5306 9580 5322
rect 9546 4914 9580 4930
rect 7658 4846 7674 4880
rect 7708 4846 7724 4880
rect 7850 4846 7866 4880
rect 7900 4846 7916 4880
rect 8042 4846 8058 4880
rect 8092 4846 8108 4880
rect 8234 4846 8250 4880
rect 8284 4846 8300 4880
rect 8426 4846 8442 4880
rect 8476 4846 8492 4880
rect 8618 4846 8634 4880
rect 8668 4846 8684 4880
rect 8810 4846 8826 4880
rect 8860 4846 8876 4880
rect 9002 4846 9018 4880
rect 9052 4846 9068 4880
rect 9194 4846 9210 4880
rect 9244 4846 9260 4880
rect 9386 4846 9402 4880
rect 9436 4846 9452 4880
rect 7512 4778 7546 4840
rect 15700 9183 15968 10532
rect 19270 11152 19304 11214
rect 16872 9358 16906 9420
rect 20496 10466 20676 10608
rect 19270 9358 19304 9420
rect 16872 9324 16968 9358
rect 19208 9324 19304 9358
rect 19412 10432 19508 10466
rect 21498 10432 21594 10466
rect 19412 10370 19446 10432
rect 15697 9149 15757 9183
rect 18383 9149 18443 9183
rect 15697 9123 15731 9149
rect 18409 9123 18443 9149
rect 15928 8870 16072 8956
rect 16364 8904 16940 8956
rect 17232 8904 17876 8956
rect 18168 8904 18216 8956
rect 18062 8870 18216 8904
rect 15928 8808 16010 8870
rect 15928 8704 15976 8808
rect 18124 8808 18216 8870
rect 16218 8768 16234 8802
rect 16268 8768 16284 8802
rect 16410 8768 16426 8802
rect 16460 8768 16476 8802
rect 16602 8768 16618 8802
rect 16652 8768 16668 8802
rect 16794 8768 16810 8802
rect 16844 8768 16860 8802
rect 16986 8768 17002 8802
rect 17036 8768 17052 8802
rect 17178 8768 17194 8802
rect 17228 8768 17244 8802
rect 17370 8768 17386 8802
rect 17420 8768 17436 8802
rect 17562 8768 17578 8802
rect 17612 8768 17628 8802
rect 17754 8768 17770 8802
rect 17804 8768 17820 8802
rect 17946 8768 17962 8802
rect 17996 8768 18012 8802
rect 15928 8356 15940 8704
rect 15928 8252 15976 8356
rect 16090 8718 16124 8734
rect 16090 8326 16124 8342
rect 16186 8718 16220 8734
rect 16186 8326 16220 8342
rect 16282 8718 16316 8734
rect 16282 8326 16316 8342
rect 16378 8718 16412 8734
rect 16378 8326 16412 8342
rect 16474 8718 16508 8734
rect 16474 8326 16508 8342
rect 16570 8718 16604 8734
rect 16570 8326 16604 8342
rect 16666 8718 16700 8734
rect 16666 8326 16700 8342
rect 16762 8718 16796 8734
rect 16762 8326 16796 8342
rect 16858 8718 16892 8734
rect 16858 8326 16892 8342
rect 16954 8718 16988 8734
rect 16954 8326 16988 8342
rect 17050 8718 17084 8734
rect 17050 8326 17084 8342
rect 17146 8718 17180 8734
rect 17146 8326 17180 8342
rect 17242 8718 17276 8734
rect 17242 8326 17276 8342
rect 17338 8718 17372 8734
rect 17338 8326 17372 8342
rect 17434 8718 17468 8734
rect 17434 8326 17468 8342
rect 17530 8718 17564 8734
rect 17530 8326 17564 8342
rect 17626 8718 17660 8734
rect 17626 8326 17660 8342
rect 17722 8718 17756 8734
rect 17722 8326 17756 8342
rect 17818 8718 17852 8734
rect 17818 8326 17852 8342
rect 17914 8718 17948 8734
rect 17914 8326 17948 8342
rect 18010 8718 18044 8734
rect 18010 8326 18044 8342
rect 18158 8672 18216 8808
rect 18200 8416 18216 8672
rect 16122 8258 16138 8292
rect 16172 8258 16188 8292
rect 16314 8258 16330 8292
rect 16364 8258 16380 8292
rect 16506 8258 16522 8292
rect 16556 8258 16572 8292
rect 16698 8258 16714 8292
rect 16748 8258 16764 8292
rect 16890 8258 16906 8292
rect 16940 8258 16956 8292
rect 17082 8258 17098 8292
rect 17132 8258 17148 8292
rect 17274 8258 17290 8292
rect 17324 8258 17340 8292
rect 17466 8258 17482 8292
rect 17516 8258 17532 8292
rect 17658 8258 17674 8292
rect 17708 8258 17724 8292
rect 17850 8258 17866 8292
rect 17900 8258 17916 8292
rect 15928 8190 16010 8252
rect 18158 8252 18216 8416
rect 18124 8190 18216 8252
rect 15928 8156 16072 8190
rect 18062 8156 18216 8190
rect 15928 8152 18216 8156
rect 15928 8148 17876 8152
rect 15928 8088 16072 8148
rect 16364 8088 16940 8148
rect 17260 8092 17876 8148
rect 18168 8092 18216 8152
rect 17260 8088 18216 8092
rect 15928 8084 18216 8088
rect 15928 8050 16072 8084
rect 18062 8050 18216 8084
rect 15928 7988 16010 8050
rect 15928 7844 15976 7988
rect 18124 7988 18216 8050
rect 16218 7948 16234 7982
rect 16268 7948 16284 7982
rect 16410 7948 16426 7982
rect 16460 7948 16476 7982
rect 16602 7948 16618 7982
rect 16652 7948 16668 7982
rect 16794 7948 16810 7982
rect 16844 7948 16860 7982
rect 16986 7948 17002 7982
rect 17036 7948 17052 7982
rect 17178 7948 17194 7982
rect 17228 7948 17244 7982
rect 17370 7948 17386 7982
rect 17420 7948 17436 7982
rect 17562 7948 17578 7982
rect 17612 7948 17628 7982
rect 17754 7948 17770 7982
rect 17804 7948 17820 7982
rect 17946 7948 17962 7982
rect 17996 7948 18012 7982
rect 15928 7588 15940 7844
rect 15928 7432 15976 7588
rect 16090 7898 16124 7914
rect 16090 7506 16124 7522
rect 16186 7898 16220 7914
rect 16186 7506 16220 7522
rect 16282 7898 16316 7914
rect 16282 7506 16316 7522
rect 16378 7898 16412 7914
rect 16378 7506 16412 7522
rect 16474 7898 16508 7914
rect 16474 7506 16508 7522
rect 16570 7898 16604 7914
rect 16570 7506 16604 7522
rect 16666 7898 16700 7914
rect 16666 7506 16700 7522
rect 16762 7898 16796 7914
rect 16762 7506 16796 7522
rect 16858 7898 16892 7914
rect 16858 7506 16892 7522
rect 16954 7898 16988 7914
rect 16954 7506 16988 7522
rect 17050 7898 17084 7914
rect 17050 7506 17084 7522
rect 17146 7898 17180 7914
rect 17146 7506 17180 7522
rect 17242 7898 17276 7914
rect 17242 7506 17276 7522
rect 17338 7898 17372 7914
rect 17338 7506 17372 7522
rect 17434 7898 17468 7914
rect 17434 7506 17468 7522
rect 17530 7898 17564 7914
rect 17530 7506 17564 7522
rect 17626 7898 17660 7914
rect 17626 7506 17660 7522
rect 17722 7898 17756 7914
rect 17722 7506 17756 7522
rect 17818 7898 17852 7914
rect 17818 7506 17852 7522
rect 17914 7898 17948 7914
rect 17914 7506 17948 7522
rect 18010 7898 18044 7914
rect 18010 7506 18044 7522
rect 18158 7824 18216 7988
rect 18200 7568 18216 7824
rect 16122 7438 16138 7472
rect 16172 7438 16188 7472
rect 16314 7438 16330 7472
rect 16364 7438 16380 7472
rect 16506 7438 16522 7472
rect 16556 7438 16572 7472
rect 16698 7438 16714 7472
rect 16748 7438 16764 7472
rect 16890 7438 16906 7472
rect 16940 7438 16956 7472
rect 17082 7438 17098 7472
rect 17132 7438 17148 7472
rect 17274 7438 17290 7472
rect 17324 7438 17340 7472
rect 17466 7438 17482 7472
rect 17516 7438 17532 7472
rect 17658 7438 17674 7472
rect 17708 7438 17724 7472
rect 17850 7438 17866 7472
rect 17900 7438 17916 7472
rect 15928 7370 16010 7432
rect 18158 7432 18216 7568
rect 18124 7370 18216 7432
rect 15928 7336 16072 7370
rect 18062 7336 18216 7370
rect 15928 7328 18216 7336
rect 15928 7268 16072 7328
rect 16364 7268 16940 7328
rect 17232 7268 17876 7328
rect 18168 7268 18216 7328
rect 15928 7264 18216 7268
rect 15928 7230 16072 7264
rect 18062 7230 18216 7264
rect 15928 7168 16010 7230
rect 15928 7004 15976 7168
rect 18124 7168 18216 7230
rect 16218 7128 16234 7162
rect 16268 7128 16284 7162
rect 16410 7128 16426 7162
rect 16460 7128 16476 7162
rect 16602 7128 16618 7162
rect 16652 7128 16668 7162
rect 16794 7128 16810 7162
rect 16844 7128 16860 7162
rect 16986 7128 17002 7162
rect 17036 7128 17052 7162
rect 17178 7128 17194 7162
rect 17228 7128 17244 7162
rect 17370 7128 17386 7162
rect 17420 7128 17436 7162
rect 17562 7128 17578 7162
rect 17612 7128 17628 7162
rect 17754 7128 17770 7162
rect 17804 7128 17820 7162
rect 17946 7128 17962 7162
rect 17996 7128 18012 7162
rect 15928 6748 15936 7004
rect 15928 6612 15976 6748
rect 16090 7078 16124 7094
rect 16090 6686 16124 6702
rect 16186 7078 16220 7094
rect 16186 6686 16220 6702
rect 16282 7078 16316 7094
rect 16282 6686 16316 6702
rect 16378 7078 16412 7094
rect 16378 6686 16412 6702
rect 16474 7078 16508 7094
rect 16474 6686 16508 6702
rect 16570 7078 16604 7094
rect 16570 6686 16604 6702
rect 16666 7078 16700 7094
rect 16666 6686 16700 6702
rect 16762 7078 16796 7094
rect 16762 6686 16796 6702
rect 16858 7078 16892 7094
rect 16858 6686 16892 6702
rect 16954 7078 16988 7094
rect 16954 6686 16988 6702
rect 17050 7078 17084 7094
rect 17050 6686 17084 6702
rect 17146 7078 17180 7094
rect 17146 6686 17180 6702
rect 17242 7078 17276 7094
rect 17242 6686 17276 6702
rect 17338 7078 17372 7094
rect 17338 6686 17372 6702
rect 17434 7078 17468 7094
rect 17434 6686 17468 6702
rect 17530 7078 17564 7094
rect 17530 6686 17564 6702
rect 17626 7078 17660 7094
rect 17626 6686 17660 6702
rect 17722 7078 17756 7094
rect 17722 6686 17756 6702
rect 17818 7078 17852 7094
rect 17818 6686 17852 6702
rect 17914 7078 17948 7094
rect 17914 6686 17948 6702
rect 18010 7078 18044 7094
rect 18010 6686 18044 6702
rect 18158 7012 18216 7168
rect 18200 6756 18216 7012
rect 16122 6618 16138 6652
rect 16172 6618 16188 6652
rect 16314 6618 16330 6652
rect 16364 6618 16380 6652
rect 16506 6618 16522 6652
rect 16556 6618 16572 6652
rect 16698 6618 16714 6652
rect 16748 6618 16764 6652
rect 16890 6618 16906 6652
rect 16940 6618 16956 6652
rect 17082 6618 17098 6652
rect 17132 6618 17148 6652
rect 17274 6618 17290 6652
rect 17324 6618 17340 6652
rect 17466 6618 17482 6652
rect 17516 6618 17532 6652
rect 17658 6618 17674 6652
rect 17708 6618 17724 6652
rect 17850 6618 17866 6652
rect 17900 6618 17916 6652
rect 15928 6550 16010 6612
rect 18158 6612 18216 6756
rect 18124 6550 18216 6612
rect 15928 6468 16072 6550
rect 18062 6516 18216 6550
rect 16364 6468 16940 6516
rect 17232 6512 18216 6516
rect 17232 6468 17876 6512
rect 18168 6468 18216 6512
rect 15697 6271 15731 6297
rect 18892 8858 19124 9324
rect 21560 10370 21594 10432
rect 19558 10330 19574 10364
rect 19608 10330 19624 10364
rect 19750 10330 19766 10364
rect 19800 10330 19816 10364
rect 19942 10330 19958 10364
rect 19992 10330 20008 10364
rect 20134 10330 20150 10364
rect 20184 10330 20200 10364
rect 20326 10330 20342 10364
rect 20376 10330 20392 10364
rect 20518 10330 20534 10364
rect 20568 10330 20584 10364
rect 20710 10330 20726 10364
rect 20760 10330 20776 10364
rect 20902 10330 20918 10364
rect 20952 10330 20968 10364
rect 21094 10330 21110 10364
rect 21144 10330 21160 10364
rect 21286 10330 21302 10364
rect 21336 10330 21352 10364
rect 19526 10271 19560 10287
rect 19526 9879 19560 9895
rect 19622 10271 19656 10287
rect 19622 9879 19656 9895
rect 19718 10271 19752 10287
rect 19718 9879 19752 9895
rect 19814 10271 19848 10287
rect 19814 9879 19848 9895
rect 19910 10271 19944 10287
rect 19910 9879 19944 9895
rect 20006 10271 20040 10287
rect 20006 9879 20040 9895
rect 20102 10271 20136 10287
rect 20102 9879 20136 9895
rect 20198 10271 20232 10287
rect 20198 9879 20232 9895
rect 20294 10271 20328 10287
rect 20294 9879 20328 9895
rect 20390 10271 20424 10287
rect 20390 9879 20424 9895
rect 20486 10271 20520 10287
rect 20486 9879 20520 9895
rect 20582 10271 20616 10287
rect 20582 9879 20616 9895
rect 20678 10271 20712 10287
rect 20678 9879 20712 9895
rect 20774 10271 20808 10287
rect 20774 9879 20808 9895
rect 20870 10271 20904 10287
rect 20870 9879 20904 9895
rect 20966 10271 21000 10287
rect 20966 9879 21000 9895
rect 21062 10271 21096 10287
rect 21062 9879 21096 9895
rect 21158 10271 21192 10287
rect 21158 9879 21192 9895
rect 21254 10271 21288 10287
rect 21254 9879 21288 9895
rect 21350 10271 21384 10287
rect 21350 9879 21384 9895
rect 21446 10271 21480 10287
rect 21446 9879 21480 9895
rect 19654 9802 19670 9836
rect 19704 9802 19720 9836
rect 19846 9802 19862 9836
rect 19896 9802 19912 9836
rect 20038 9802 20054 9836
rect 20088 9802 20104 9836
rect 20230 9802 20246 9836
rect 20280 9802 20296 9836
rect 20422 9802 20438 9836
rect 20472 9802 20488 9836
rect 20614 9802 20630 9836
rect 20664 9802 20680 9836
rect 20806 9802 20822 9836
rect 20856 9802 20872 9836
rect 20998 9802 21014 9836
rect 21048 9802 21064 9836
rect 21190 9802 21206 9836
rect 21240 9802 21256 9836
rect 21382 9802 21398 9836
rect 21432 9802 21448 9836
rect 19654 9694 19670 9728
rect 19704 9694 19720 9728
rect 19846 9694 19862 9728
rect 19896 9694 19912 9728
rect 20038 9694 20054 9728
rect 20088 9694 20104 9728
rect 20230 9694 20246 9728
rect 20280 9694 20296 9728
rect 20422 9694 20438 9728
rect 20472 9694 20488 9728
rect 20614 9694 20630 9728
rect 20664 9694 20680 9728
rect 20806 9694 20822 9728
rect 20856 9694 20872 9728
rect 20998 9694 21014 9728
rect 21048 9694 21064 9728
rect 21190 9694 21206 9728
rect 21240 9694 21256 9728
rect 21382 9694 21398 9728
rect 21432 9694 21448 9728
rect 19526 9635 19560 9651
rect 19526 9243 19560 9259
rect 19622 9635 19656 9651
rect 19622 9243 19656 9259
rect 19718 9635 19752 9651
rect 19718 9243 19752 9259
rect 19814 9635 19848 9651
rect 19814 9243 19848 9259
rect 19910 9635 19944 9651
rect 19910 9243 19944 9259
rect 20006 9635 20040 9651
rect 20006 9243 20040 9259
rect 20102 9635 20136 9651
rect 20102 9243 20136 9259
rect 20198 9635 20232 9651
rect 20198 9243 20232 9259
rect 20294 9635 20328 9651
rect 20294 9243 20328 9259
rect 20390 9635 20424 9651
rect 20390 9243 20424 9259
rect 20486 9635 20520 9651
rect 20486 9243 20520 9259
rect 20582 9635 20616 9651
rect 20582 9243 20616 9259
rect 20678 9635 20712 9651
rect 20678 9243 20712 9259
rect 20774 9635 20808 9651
rect 20774 9243 20808 9259
rect 20870 9635 20904 9651
rect 20870 9243 20904 9259
rect 20966 9635 21000 9651
rect 20966 9243 21000 9259
rect 21062 9635 21096 9651
rect 21062 9243 21096 9259
rect 21158 9635 21192 9651
rect 21158 9243 21192 9259
rect 21254 9635 21288 9651
rect 21254 9243 21288 9259
rect 21350 9635 21384 9651
rect 21350 9243 21384 9259
rect 21446 9635 21480 9651
rect 21446 9243 21480 9259
rect 19558 9166 19574 9200
rect 19608 9166 19624 9200
rect 19750 9166 19766 9200
rect 19800 9166 19816 9200
rect 19942 9166 19958 9200
rect 19992 9166 20008 9200
rect 20134 9166 20150 9200
rect 20184 9166 20200 9200
rect 20326 9166 20342 9200
rect 20376 9166 20392 9200
rect 20518 9166 20534 9200
rect 20568 9166 20584 9200
rect 20710 9166 20726 9200
rect 20760 9166 20776 9200
rect 20902 9166 20918 9200
rect 20952 9166 20968 9200
rect 21094 9166 21110 9200
rect 21144 9166 21160 9200
rect 21286 9166 21302 9200
rect 21336 9166 21352 9200
rect 19412 9098 19446 9160
rect 21560 9098 21594 9160
rect 19412 9064 19508 9098
rect 21498 9064 21594 9098
rect 21912 10402 22008 10436
rect 23998 10402 24094 10436
rect 21912 10340 21946 10402
rect 19412 8858 19508 8870
rect 18892 8836 19508 8858
rect 21498 8836 21594 8870
rect 18892 8774 19446 8836
rect 18892 8750 19412 8774
rect 21560 8774 21594 8836
rect 19558 8734 19574 8768
rect 19608 8734 19624 8768
rect 19750 8734 19766 8768
rect 19800 8734 19816 8768
rect 19942 8734 19958 8768
rect 19992 8734 20008 8768
rect 20134 8734 20150 8768
rect 20184 8734 20200 8768
rect 20326 8734 20342 8768
rect 20376 8734 20392 8768
rect 20518 8734 20534 8768
rect 20568 8734 20584 8768
rect 20710 8734 20726 8768
rect 20760 8734 20776 8768
rect 20902 8734 20918 8768
rect 20952 8734 20968 8768
rect 21094 8734 21110 8768
rect 21144 8734 21160 8768
rect 21286 8734 21302 8768
rect 21336 8734 21352 8768
rect 19526 8684 19560 8700
rect 19526 8292 19560 8308
rect 19622 8684 19656 8700
rect 19622 8292 19656 8308
rect 19718 8684 19752 8700
rect 19718 8292 19752 8308
rect 19814 8684 19848 8700
rect 19814 8292 19848 8308
rect 19910 8684 19944 8700
rect 19910 8292 19944 8308
rect 20006 8684 20040 8700
rect 20006 8292 20040 8308
rect 20102 8684 20136 8700
rect 20102 8292 20136 8308
rect 20198 8684 20232 8700
rect 20198 8292 20232 8308
rect 20294 8684 20328 8700
rect 20294 8292 20328 8308
rect 20390 8684 20424 8700
rect 20390 8292 20424 8308
rect 20486 8684 20520 8700
rect 20486 8292 20520 8308
rect 20582 8684 20616 8700
rect 20582 8292 20616 8308
rect 20678 8684 20712 8700
rect 20678 8292 20712 8308
rect 20774 8684 20808 8700
rect 20774 8292 20808 8308
rect 20870 8684 20904 8700
rect 20870 8292 20904 8308
rect 20966 8684 21000 8700
rect 20966 8292 21000 8308
rect 21062 8684 21096 8700
rect 21062 8292 21096 8308
rect 21158 8684 21192 8700
rect 21158 8292 21192 8308
rect 21254 8684 21288 8700
rect 21254 8292 21288 8308
rect 21350 8684 21384 8700
rect 21350 8292 21384 8308
rect 21446 8684 21480 8700
rect 21446 8292 21480 8308
rect 19654 8224 19670 8258
rect 19704 8224 19720 8258
rect 19846 8224 19862 8258
rect 19896 8224 19912 8258
rect 20038 8224 20054 8258
rect 20088 8224 20104 8258
rect 20230 8224 20246 8258
rect 20280 8224 20296 8258
rect 20422 8224 20438 8258
rect 20472 8224 20488 8258
rect 20614 8224 20630 8258
rect 20664 8224 20680 8258
rect 20806 8224 20822 8258
rect 20856 8224 20872 8258
rect 20998 8224 21014 8258
rect 21048 8224 21064 8258
rect 21190 8224 21206 8258
rect 21240 8224 21256 8258
rect 21382 8224 21398 8258
rect 21432 8224 21448 8258
rect 19654 8116 19670 8150
rect 19704 8116 19720 8150
rect 19846 8116 19862 8150
rect 19896 8116 19912 8150
rect 20038 8116 20054 8150
rect 20088 8116 20104 8150
rect 20230 8116 20246 8150
rect 20280 8116 20296 8150
rect 20422 8116 20438 8150
rect 20472 8116 20488 8150
rect 20614 8116 20630 8150
rect 20664 8116 20680 8150
rect 20806 8116 20822 8150
rect 20856 8116 20872 8150
rect 20998 8116 21014 8150
rect 21048 8116 21064 8150
rect 21190 8116 21206 8150
rect 21240 8116 21256 8150
rect 21382 8116 21398 8150
rect 21432 8116 21448 8150
rect 19526 8066 19560 8082
rect 19526 7674 19560 7690
rect 19622 8066 19656 8082
rect 19622 7674 19656 7690
rect 19718 8066 19752 8082
rect 19718 7674 19752 7690
rect 19814 8066 19848 8082
rect 19814 7674 19848 7690
rect 19910 8066 19944 8082
rect 19910 7674 19944 7690
rect 20006 8066 20040 8082
rect 20006 7674 20040 7690
rect 20102 8066 20136 8082
rect 20102 7674 20136 7690
rect 20198 8066 20232 8082
rect 20198 7674 20232 7690
rect 20294 8066 20328 8082
rect 20294 7674 20328 7690
rect 20390 8066 20424 8082
rect 20390 7674 20424 7690
rect 20486 8066 20520 8082
rect 20486 7674 20520 7690
rect 20582 8066 20616 8082
rect 20582 7674 20616 7690
rect 20678 8066 20712 8082
rect 20678 7674 20712 7690
rect 20774 8066 20808 8082
rect 20774 7674 20808 7690
rect 20870 8066 20904 8082
rect 20870 7674 20904 7690
rect 20966 8066 21000 8082
rect 20966 7674 21000 7690
rect 21062 8066 21096 8082
rect 21062 7674 21096 7690
rect 21158 8066 21192 8082
rect 21158 7674 21192 7690
rect 21254 8066 21288 8082
rect 21254 7674 21288 7690
rect 21350 8066 21384 8082
rect 21350 7674 21384 7690
rect 21446 8066 21480 8082
rect 21446 7674 21480 7690
rect 19558 7606 19574 7640
rect 19608 7606 19624 7640
rect 19750 7606 19766 7640
rect 19800 7606 19816 7640
rect 19942 7606 19958 7640
rect 19992 7606 20008 7640
rect 20134 7606 20150 7640
rect 20184 7606 20200 7640
rect 20326 7606 20342 7640
rect 20376 7606 20392 7640
rect 20518 7606 20534 7640
rect 20568 7606 20584 7640
rect 20710 7606 20726 7640
rect 20760 7606 20776 7640
rect 20902 7606 20918 7640
rect 20952 7606 20968 7640
rect 21094 7606 21110 7640
rect 21144 7606 21160 7640
rect 21286 7606 21302 7640
rect 21336 7606 21352 7640
rect 19412 7538 19446 7600
rect 21560 7538 21594 7600
rect 19412 7528 19508 7538
rect 19408 7504 19508 7528
rect 21498 7504 21594 7538
rect 19408 7288 21588 7504
rect 18409 6271 18443 6297
rect 19648 6296 19940 7288
rect 15697 6237 15757 6271
rect 18383 6237 18443 6271
rect 19208 6248 19940 6296
rect 18730 6048 19940 6248
rect 9660 4778 9694 4840
rect 7512 4744 7608 4778
rect 9598 4744 9694 4778
rect 14512 6014 14608 6048
rect 15638 6014 16408 6048
rect 17438 6014 18208 6048
rect 19238 6036 20008 6048
rect 19238 6014 19334 6036
rect 14512 5952 14546 6014
rect 6700 4098 6734 4160
rect 5248 4064 5608 4098
rect 6638 4064 6734 4098
rect 15700 5952 16346 6014
rect 14754 5912 14770 5946
rect 14804 5912 14820 5946
rect 14946 5912 14962 5946
rect 14996 5912 15012 5946
rect 15138 5912 15154 5946
rect 15188 5912 15204 5946
rect 15330 5912 15346 5946
rect 15380 5912 15396 5946
rect 15522 5912 15538 5946
rect 15572 5912 15588 5946
rect 14626 5862 14660 5878
rect 14626 5470 14660 5486
rect 14722 5862 14756 5878
rect 14722 5470 14756 5486
rect 14818 5862 14852 5878
rect 14818 5470 14852 5486
rect 14914 5862 14948 5878
rect 14914 5470 14948 5486
rect 15010 5862 15044 5878
rect 15010 5470 15044 5486
rect 15106 5862 15140 5878
rect 15106 5470 15140 5486
rect 15202 5862 15236 5878
rect 15202 5470 15236 5486
rect 15298 5862 15332 5878
rect 15298 5470 15332 5486
rect 15394 5862 15428 5878
rect 15394 5470 15428 5486
rect 15490 5862 15524 5878
rect 15490 5470 15524 5486
rect 15586 5862 15620 5878
rect 15586 5470 15620 5486
rect 14658 5402 14674 5436
rect 14708 5402 14724 5436
rect 14850 5402 14866 5436
rect 14900 5402 14916 5436
rect 15042 5402 15058 5436
rect 15092 5402 15108 5436
rect 15234 5402 15250 5436
rect 15284 5402 15300 5436
rect 15426 5402 15442 5436
rect 15476 5402 15492 5436
rect 14658 5294 14674 5328
rect 14708 5294 14724 5328
rect 14850 5294 14866 5328
rect 14900 5294 14916 5328
rect 15042 5294 15058 5328
rect 15092 5294 15108 5328
rect 15234 5294 15250 5328
rect 15284 5294 15300 5328
rect 15426 5294 15442 5328
rect 15476 5294 15492 5328
rect 14626 5244 14660 5260
rect 14626 4852 14660 4868
rect 14722 5244 14756 5260
rect 14722 4852 14756 4868
rect 14818 5244 14852 5260
rect 14818 4852 14852 4868
rect 14914 5244 14948 5260
rect 14914 4852 14948 4868
rect 15010 5244 15044 5260
rect 15010 4852 15044 4868
rect 15106 5244 15140 5260
rect 15106 4852 15140 4868
rect 15202 5244 15236 5260
rect 15202 4852 15236 4868
rect 15298 5244 15332 5260
rect 15298 4852 15332 4868
rect 15394 5244 15428 5260
rect 15394 4852 15428 4868
rect 15490 5244 15524 5260
rect 15490 4852 15524 4868
rect 15586 5244 15620 5260
rect 15586 4852 15620 4868
rect 14754 4784 14770 4818
rect 14804 4784 14820 4818
rect 14946 4784 14962 4818
rect 14996 4784 15012 4818
rect 15138 4784 15154 4818
rect 15188 4784 15204 4818
rect 15330 4784 15346 4818
rect 15380 4784 15396 4818
rect 15522 4784 15538 4818
rect 15572 4784 15588 4818
rect 14754 4676 14770 4710
rect 14804 4676 14820 4710
rect 14946 4676 14962 4710
rect 14996 4676 15012 4710
rect 15138 4676 15154 4710
rect 15188 4676 15204 4710
rect 15330 4676 15346 4710
rect 15380 4676 15396 4710
rect 15522 4676 15538 4710
rect 15572 4676 15588 4710
rect 14626 4626 14660 4642
rect 14626 4234 14660 4250
rect 14722 4626 14756 4642
rect 14722 4234 14756 4250
rect 14818 4626 14852 4642
rect 14818 4234 14852 4250
rect 14914 4626 14948 4642
rect 14914 4234 14948 4250
rect 15010 4626 15044 4642
rect 15010 4234 15044 4250
rect 15106 4626 15140 4642
rect 15106 4234 15140 4250
rect 15202 4626 15236 4642
rect 15202 4234 15236 4250
rect 15298 4626 15332 4642
rect 15298 4234 15332 4250
rect 15394 4626 15428 4642
rect 15394 4234 15428 4250
rect 15490 4626 15524 4642
rect 15490 4234 15524 4250
rect 15586 4626 15620 4642
rect 15586 4234 15620 4250
rect 14658 4166 14674 4200
rect 14708 4166 14724 4200
rect 14850 4166 14866 4200
rect 14900 4166 14916 4200
rect 15042 4166 15058 4200
rect 15092 4166 15108 4200
rect 15234 4166 15250 4200
rect 15284 4166 15300 4200
rect 15426 4166 15442 4200
rect 15476 4166 15492 4200
rect 14512 4098 14546 4160
rect 15734 5808 16312 5952
rect 15700 4098 15734 4160
rect 14512 4064 14608 4098
rect 15638 4064 15734 4098
rect 16040 4160 16312 5808
rect 17500 5952 18146 6014
rect 16554 5912 16570 5946
rect 16604 5912 16620 5946
rect 16746 5912 16762 5946
rect 16796 5912 16812 5946
rect 16938 5912 16954 5946
rect 16988 5912 17004 5946
rect 17130 5912 17146 5946
rect 17180 5912 17196 5946
rect 17322 5912 17338 5946
rect 17372 5912 17388 5946
rect 16426 5862 16460 5878
rect 16426 5470 16460 5486
rect 16522 5862 16556 5878
rect 16522 5470 16556 5486
rect 16618 5862 16652 5878
rect 16618 5470 16652 5486
rect 16714 5862 16748 5878
rect 16714 5470 16748 5486
rect 16810 5862 16844 5878
rect 16810 5470 16844 5486
rect 16906 5862 16940 5878
rect 16906 5470 16940 5486
rect 17002 5862 17036 5878
rect 17002 5470 17036 5486
rect 17098 5862 17132 5878
rect 17098 5470 17132 5486
rect 17194 5862 17228 5878
rect 17194 5470 17228 5486
rect 17290 5862 17324 5878
rect 17290 5470 17324 5486
rect 17386 5862 17420 5878
rect 17386 5470 17420 5486
rect 16458 5402 16474 5436
rect 16508 5402 16524 5436
rect 16650 5402 16666 5436
rect 16700 5402 16716 5436
rect 16842 5402 16858 5436
rect 16892 5402 16908 5436
rect 17034 5402 17050 5436
rect 17084 5402 17100 5436
rect 17226 5402 17242 5436
rect 17276 5402 17292 5436
rect 16458 5294 16474 5328
rect 16508 5294 16524 5328
rect 16650 5294 16666 5328
rect 16700 5294 16716 5328
rect 16842 5294 16858 5328
rect 16892 5294 16908 5328
rect 17034 5294 17050 5328
rect 17084 5294 17100 5328
rect 17226 5294 17242 5328
rect 17276 5294 17292 5328
rect 16426 5244 16460 5260
rect 16426 4852 16460 4868
rect 16522 5244 16556 5260
rect 16522 4852 16556 4868
rect 16618 5244 16652 5260
rect 16618 4852 16652 4868
rect 16714 5244 16748 5260
rect 16714 4852 16748 4868
rect 16810 5244 16844 5260
rect 16810 4852 16844 4868
rect 16906 5244 16940 5260
rect 16906 4852 16940 4868
rect 17002 5244 17036 5260
rect 17002 4852 17036 4868
rect 17098 5244 17132 5260
rect 17098 4852 17132 4868
rect 17194 5244 17228 5260
rect 17194 4852 17228 4868
rect 17290 5244 17324 5260
rect 17290 4852 17324 4868
rect 17386 5244 17420 5260
rect 17386 4852 17420 4868
rect 16554 4784 16570 4818
rect 16604 4784 16620 4818
rect 16746 4784 16762 4818
rect 16796 4784 16812 4818
rect 16938 4784 16954 4818
rect 16988 4784 17004 4818
rect 17130 4784 17146 4818
rect 17180 4784 17196 4818
rect 17322 4784 17338 4818
rect 17372 4784 17388 4818
rect 16554 4676 16570 4710
rect 16604 4676 16620 4710
rect 16746 4676 16762 4710
rect 16796 4676 16812 4710
rect 16938 4676 16954 4710
rect 16988 4676 17004 4710
rect 17130 4676 17146 4710
rect 17180 4676 17196 4710
rect 17322 4676 17338 4710
rect 17372 4676 17388 4710
rect 16426 4626 16460 4642
rect 16426 4234 16460 4250
rect 16522 4626 16556 4642
rect 16522 4234 16556 4250
rect 16618 4626 16652 4642
rect 16618 4234 16652 4250
rect 16714 4626 16748 4642
rect 16714 4234 16748 4250
rect 16810 4626 16844 4642
rect 16810 4234 16844 4250
rect 16906 4626 16940 4642
rect 16906 4234 16940 4250
rect 17002 4626 17036 4642
rect 17002 4234 17036 4250
rect 17098 4626 17132 4642
rect 17098 4234 17132 4250
rect 17194 4626 17228 4642
rect 17194 4234 17228 4250
rect 17290 4626 17324 4642
rect 17290 4234 17324 4250
rect 17386 4626 17420 4642
rect 17386 4234 17420 4250
rect 16458 4166 16474 4200
rect 16508 4166 16524 4200
rect 16650 4166 16666 4200
rect 16700 4166 16716 4200
rect 16842 4166 16858 4200
rect 16892 4166 16908 4200
rect 17034 4166 17050 4200
rect 17084 4166 17100 4200
rect 17226 4166 17242 4200
rect 17276 4166 17292 4200
rect 16040 4098 16346 4160
rect 17534 5808 18112 5952
rect 17500 4098 17534 4160
rect 16040 4064 16408 4098
rect 17438 4064 17534 4098
rect 17840 4160 18112 5808
rect 19300 5952 19334 6014
rect 18354 5912 18370 5946
rect 18404 5912 18420 5946
rect 18546 5912 18562 5946
rect 18596 5912 18612 5946
rect 18738 5912 18754 5946
rect 18788 5912 18804 5946
rect 18930 5912 18946 5946
rect 18980 5912 18996 5946
rect 19122 5912 19138 5946
rect 19172 5912 19188 5946
rect 18226 5862 18260 5878
rect 18226 5470 18260 5486
rect 18322 5862 18356 5878
rect 18322 5470 18356 5486
rect 18418 5862 18452 5878
rect 18418 5470 18452 5486
rect 18514 5862 18548 5878
rect 18514 5470 18548 5486
rect 18610 5862 18644 5878
rect 18610 5470 18644 5486
rect 18706 5862 18740 5878
rect 18706 5470 18740 5486
rect 18802 5862 18836 5878
rect 18802 5470 18836 5486
rect 18898 5862 18932 5878
rect 18898 5470 18932 5486
rect 18994 5862 19028 5878
rect 18994 5470 19028 5486
rect 19090 5862 19124 5878
rect 19090 5470 19124 5486
rect 19186 5862 19220 5878
rect 19186 5470 19220 5486
rect 18258 5402 18274 5436
rect 18308 5402 18324 5436
rect 18450 5402 18466 5436
rect 18500 5402 18516 5436
rect 18642 5402 18658 5436
rect 18692 5402 18708 5436
rect 18834 5402 18850 5436
rect 18884 5402 18900 5436
rect 19026 5402 19042 5436
rect 19076 5402 19092 5436
rect 18258 5294 18274 5328
rect 18308 5294 18324 5328
rect 18450 5294 18466 5328
rect 18500 5294 18516 5328
rect 18642 5294 18658 5328
rect 18692 5294 18708 5328
rect 18834 5294 18850 5328
rect 18884 5294 18900 5328
rect 19026 5294 19042 5328
rect 19076 5294 19092 5328
rect 18226 5244 18260 5260
rect 18226 4852 18260 4868
rect 18322 5244 18356 5260
rect 18322 4852 18356 4868
rect 18418 5244 18452 5260
rect 18418 4852 18452 4868
rect 18514 5244 18548 5260
rect 18514 4852 18548 4868
rect 18610 5244 18644 5260
rect 18610 4852 18644 4868
rect 18706 5244 18740 5260
rect 18706 4852 18740 4868
rect 18802 5244 18836 5260
rect 18802 4852 18836 4868
rect 18898 5244 18932 5260
rect 18898 4852 18932 4868
rect 18994 5244 19028 5260
rect 18994 4852 19028 4868
rect 19090 5244 19124 5260
rect 19090 4852 19124 4868
rect 19186 5244 19220 5260
rect 19186 4852 19220 4868
rect 18354 4784 18370 4818
rect 18404 4784 18420 4818
rect 18546 4784 18562 4818
rect 18596 4784 18612 4818
rect 18738 4784 18754 4818
rect 18788 4784 18804 4818
rect 18930 4784 18946 4818
rect 18980 4784 18996 4818
rect 19122 4784 19138 4818
rect 19172 4784 19188 4818
rect 18354 4676 18370 4710
rect 18404 4676 18420 4710
rect 18546 4676 18562 4710
rect 18596 4676 18612 4710
rect 18738 4676 18754 4710
rect 18788 4676 18804 4710
rect 18930 4676 18946 4710
rect 18980 4676 18996 4710
rect 19122 4676 19138 4710
rect 19172 4676 19188 4710
rect 18226 4626 18260 4642
rect 18226 4234 18260 4250
rect 18322 4626 18356 4642
rect 18322 4234 18356 4250
rect 18418 4626 18452 4642
rect 18418 4234 18452 4250
rect 18514 4626 18548 4642
rect 18514 4234 18548 4250
rect 18610 4626 18644 4642
rect 18610 4234 18644 4250
rect 18706 4626 18740 4642
rect 18706 4234 18740 4250
rect 18802 4626 18836 4642
rect 18802 4234 18836 4250
rect 18898 4626 18932 4642
rect 18898 4234 18932 4250
rect 18994 4626 19028 4642
rect 18994 4234 19028 4250
rect 19090 4626 19124 4642
rect 19090 4234 19124 4250
rect 19186 4626 19220 4642
rect 19186 4234 19220 4250
rect 18258 4166 18274 4200
rect 18308 4166 18324 4200
rect 18450 4166 18466 4200
rect 18500 4166 18516 4200
rect 18642 4166 18658 4200
rect 18692 4166 18708 4200
rect 18834 4166 18850 4200
rect 18884 4166 18900 4200
rect 19026 4166 19042 4200
rect 19076 4166 19092 4200
rect 17840 4098 18146 4160
rect 19300 4098 19334 4160
rect 17840 4064 18208 4098
rect 19238 4064 19334 4098
rect 19648 6014 20008 6036
rect 21038 6014 21134 6048
rect 19648 5952 19946 6014
rect 19648 4160 19912 5952
rect 21100 5952 21134 6014
rect 20154 5912 20170 5946
rect 20204 5912 20220 5946
rect 20346 5912 20362 5946
rect 20396 5912 20412 5946
rect 20538 5912 20554 5946
rect 20588 5912 20604 5946
rect 20730 5912 20746 5946
rect 20780 5912 20796 5946
rect 20922 5912 20938 5946
rect 20972 5912 20988 5946
rect 20026 5862 20060 5878
rect 20026 5470 20060 5486
rect 20122 5862 20156 5878
rect 20122 5470 20156 5486
rect 20218 5862 20252 5878
rect 20218 5470 20252 5486
rect 20314 5862 20348 5878
rect 20314 5470 20348 5486
rect 20410 5862 20444 5878
rect 20410 5470 20444 5486
rect 20506 5862 20540 5878
rect 20506 5470 20540 5486
rect 20602 5862 20636 5878
rect 20602 5470 20636 5486
rect 20698 5862 20732 5878
rect 20698 5470 20732 5486
rect 20794 5862 20828 5878
rect 20794 5470 20828 5486
rect 20890 5862 20924 5878
rect 20890 5470 20924 5486
rect 20986 5862 21020 5878
rect 20986 5470 21020 5486
rect 20058 5402 20074 5436
rect 20108 5402 20124 5436
rect 20250 5402 20266 5436
rect 20300 5402 20316 5436
rect 20442 5402 20458 5436
rect 20492 5402 20508 5436
rect 20634 5402 20650 5436
rect 20684 5402 20700 5436
rect 20826 5402 20842 5436
rect 20876 5402 20892 5436
rect 20058 5294 20074 5328
rect 20108 5294 20124 5328
rect 20250 5294 20266 5328
rect 20300 5294 20316 5328
rect 20442 5294 20458 5328
rect 20492 5294 20508 5328
rect 20634 5294 20650 5328
rect 20684 5294 20700 5328
rect 20826 5294 20842 5328
rect 20876 5294 20892 5328
rect 20026 5244 20060 5260
rect 20026 4852 20060 4868
rect 20122 5244 20156 5260
rect 20122 4852 20156 4868
rect 20218 5244 20252 5260
rect 20218 4852 20252 4868
rect 20314 5244 20348 5260
rect 20314 4852 20348 4868
rect 20410 5244 20444 5260
rect 20410 4852 20444 4868
rect 20506 5244 20540 5260
rect 20506 4852 20540 4868
rect 20602 5244 20636 5260
rect 20602 4852 20636 4868
rect 20698 5244 20732 5260
rect 20698 4852 20732 4868
rect 20794 5244 20828 5260
rect 20794 4852 20828 4868
rect 20890 5244 20924 5260
rect 20890 4852 20924 4868
rect 20986 5244 21020 5260
rect 20986 4852 21020 4868
rect 20154 4784 20170 4818
rect 20204 4784 20220 4818
rect 20346 4784 20362 4818
rect 20396 4784 20412 4818
rect 20538 4784 20554 4818
rect 20588 4784 20604 4818
rect 20730 4784 20746 4818
rect 20780 4784 20796 4818
rect 20922 4784 20938 4818
rect 20972 4784 20988 4818
rect 20154 4676 20170 4710
rect 20204 4676 20220 4710
rect 20346 4676 20362 4710
rect 20396 4676 20412 4710
rect 20538 4676 20554 4710
rect 20588 4676 20604 4710
rect 20730 4676 20746 4710
rect 20780 4676 20796 4710
rect 20922 4676 20938 4710
rect 20972 4676 20988 4710
rect 20026 4626 20060 4642
rect 20026 4234 20060 4250
rect 20122 4626 20156 4642
rect 20122 4234 20156 4250
rect 20218 4626 20252 4642
rect 20218 4234 20252 4250
rect 20314 4626 20348 4642
rect 20314 4234 20348 4250
rect 20410 4626 20444 4642
rect 20410 4234 20444 4250
rect 20506 4626 20540 4642
rect 20506 4234 20540 4250
rect 20602 4626 20636 4642
rect 20602 4234 20636 4250
rect 20698 4626 20732 4642
rect 20698 4234 20732 4250
rect 20794 4626 20828 4642
rect 20794 4234 20828 4250
rect 20890 4626 20924 4642
rect 20890 4234 20924 4250
rect 20986 4626 21020 4642
rect 20986 4234 21020 4250
rect 20058 4166 20074 4200
rect 20108 4166 20124 4200
rect 20250 4166 20266 4200
rect 20300 4166 20316 4200
rect 20442 4166 20458 4200
rect 20492 4166 20508 4200
rect 20634 4166 20650 4200
rect 20684 4166 20700 4200
rect 20826 4166 20842 4200
rect 20876 4166 20892 4200
rect 19648 4098 19946 4160
rect 21134 4988 21912 5188
rect 24060 10340 24094 10402
rect 22154 10300 22170 10334
rect 22204 10300 22220 10334
rect 22346 10300 22362 10334
rect 22396 10300 22412 10334
rect 22538 10300 22554 10334
rect 22588 10300 22604 10334
rect 22730 10300 22746 10334
rect 22780 10300 22796 10334
rect 22922 10300 22938 10334
rect 22972 10300 22988 10334
rect 23114 10300 23130 10334
rect 23164 10300 23180 10334
rect 23306 10300 23322 10334
rect 23356 10300 23372 10334
rect 23498 10300 23514 10334
rect 23548 10300 23564 10334
rect 23690 10300 23706 10334
rect 23740 10300 23756 10334
rect 23882 10300 23898 10334
rect 23932 10300 23948 10334
rect 22026 10250 22060 10266
rect 22026 9858 22060 9874
rect 22122 10250 22156 10266
rect 22122 9858 22156 9874
rect 22218 10250 22252 10266
rect 22218 9858 22252 9874
rect 22314 10250 22348 10266
rect 22314 9858 22348 9874
rect 22410 10250 22444 10266
rect 22410 9858 22444 9874
rect 22506 10250 22540 10266
rect 22506 9858 22540 9874
rect 22602 10250 22636 10266
rect 22602 9858 22636 9874
rect 22698 10250 22732 10266
rect 22698 9858 22732 9874
rect 22794 10250 22828 10266
rect 22794 9858 22828 9874
rect 22890 10250 22924 10266
rect 22890 9858 22924 9874
rect 22986 10250 23020 10266
rect 22986 9858 23020 9874
rect 23082 10250 23116 10266
rect 23082 9858 23116 9874
rect 23178 10250 23212 10266
rect 23178 9858 23212 9874
rect 23274 10250 23308 10266
rect 23274 9858 23308 9874
rect 23370 10250 23404 10266
rect 23370 9858 23404 9874
rect 23466 10250 23500 10266
rect 23466 9858 23500 9874
rect 23562 10250 23596 10266
rect 23562 9858 23596 9874
rect 23658 10250 23692 10266
rect 23658 9858 23692 9874
rect 23754 10250 23788 10266
rect 23754 9858 23788 9874
rect 23850 10250 23884 10266
rect 23850 9858 23884 9874
rect 23946 10250 23980 10266
rect 23946 9858 23980 9874
rect 22058 9790 22074 9824
rect 22108 9790 22124 9824
rect 22250 9790 22266 9824
rect 22300 9790 22316 9824
rect 22442 9790 22458 9824
rect 22492 9790 22508 9824
rect 22634 9790 22650 9824
rect 22684 9790 22700 9824
rect 22826 9790 22842 9824
rect 22876 9790 22892 9824
rect 23018 9790 23034 9824
rect 23068 9790 23084 9824
rect 23210 9790 23226 9824
rect 23260 9790 23276 9824
rect 23402 9790 23418 9824
rect 23452 9790 23468 9824
rect 23594 9790 23610 9824
rect 23644 9790 23660 9824
rect 23786 9790 23802 9824
rect 23836 9790 23852 9824
rect 22058 9682 22074 9716
rect 22108 9682 22124 9716
rect 22250 9682 22266 9716
rect 22300 9682 22316 9716
rect 22442 9682 22458 9716
rect 22492 9682 22508 9716
rect 22634 9682 22650 9716
rect 22684 9682 22700 9716
rect 22826 9682 22842 9716
rect 22876 9682 22892 9716
rect 23018 9682 23034 9716
rect 23068 9682 23084 9716
rect 23210 9682 23226 9716
rect 23260 9682 23276 9716
rect 23402 9682 23418 9716
rect 23452 9682 23468 9716
rect 23594 9682 23610 9716
rect 23644 9682 23660 9716
rect 23786 9682 23802 9716
rect 23836 9682 23852 9716
rect 22026 9632 22060 9648
rect 22026 9240 22060 9256
rect 22122 9632 22156 9648
rect 22122 9240 22156 9256
rect 22218 9632 22252 9648
rect 22218 9240 22252 9256
rect 22314 9632 22348 9648
rect 22314 9240 22348 9256
rect 22410 9632 22444 9648
rect 22410 9240 22444 9256
rect 22506 9632 22540 9648
rect 22506 9240 22540 9256
rect 22602 9632 22636 9648
rect 22602 9240 22636 9256
rect 22698 9632 22732 9648
rect 22698 9240 22732 9256
rect 22794 9632 22828 9648
rect 22794 9240 22828 9256
rect 22890 9632 22924 9648
rect 22890 9240 22924 9256
rect 22986 9632 23020 9648
rect 22986 9240 23020 9256
rect 23082 9632 23116 9648
rect 23082 9240 23116 9256
rect 23178 9632 23212 9648
rect 23178 9240 23212 9256
rect 23274 9632 23308 9648
rect 23274 9240 23308 9256
rect 23370 9632 23404 9648
rect 23370 9240 23404 9256
rect 23466 9632 23500 9648
rect 23466 9240 23500 9256
rect 23562 9632 23596 9648
rect 23562 9240 23596 9256
rect 23658 9632 23692 9648
rect 23658 9240 23692 9256
rect 23754 9632 23788 9648
rect 23754 9240 23788 9256
rect 23850 9632 23884 9648
rect 23850 9240 23884 9256
rect 23946 9632 23980 9648
rect 23946 9240 23980 9256
rect 22154 9172 22170 9206
rect 22204 9172 22220 9206
rect 22346 9172 22362 9206
rect 22396 9172 22412 9206
rect 22538 9172 22554 9206
rect 22588 9172 22604 9206
rect 22730 9172 22746 9206
rect 22780 9172 22796 9206
rect 22922 9172 22938 9206
rect 22972 9172 22988 9206
rect 23114 9172 23130 9206
rect 23164 9172 23180 9206
rect 23306 9172 23322 9206
rect 23356 9172 23372 9206
rect 23498 9172 23514 9206
rect 23548 9172 23564 9206
rect 23690 9172 23706 9206
rect 23740 9172 23756 9206
rect 23882 9172 23898 9206
rect 23932 9172 23948 9206
rect 22154 9064 22170 9098
rect 22204 9064 22220 9098
rect 22346 9064 22362 9098
rect 22396 9064 22412 9098
rect 22538 9064 22554 9098
rect 22588 9064 22604 9098
rect 22730 9064 22746 9098
rect 22780 9064 22796 9098
rect 22922 9064 22938 9098
rect 22972 9064 22988 9098
rect 23114 9064 23130 9098
rect 23164 9064 23180 9098
rect 23306 9064 23322 9098
rect 23356 9064 23372 9098
rect 23498 9064 23514 9098
rect 23548 9064 23564 9098
rect 23690 9064 23706 9098
rect 23740 9064 23756 9098
rect 23882 9064 23898 9098
rect 23932 9064 23948 9098
rect 22026 9014 22060 9030
rect 22026 8622 22060 8638
rect 22122 9014 22156 9030
rect 22122 8622 22156 8638
rect 22218 9014 22252 9030
rect 22218 8622 22252 8638
rect 22314 9014 22348 9030
rect 22314 8622 22348 8638
rect 22410 9014 22444 9030
rect 22410 8622 22444 8638
rect 22506 9014 22540 9030
rect 22506 8622 22540 8638
rect 22602 9014 22636 9030
rect 22602 8622 22636 8638
rect 22698 9014 22732 9030
rect 22698 8622 22732 8638
rect 22794 9014 22828 9030
rect 22794 8622 22828 8638
rect 22890 9014 22924 9030
rect 22890 8622 22924 8638
rect 22986 9014 23020 9030
rect 22986 8622 23020 8638
rect 23082 9014 23116 9030
rect 23082 8622 23116 8638
rect 23178 9014 23212 9030
rect 23178 8622 23212 8638
rect 23274 9014 23308 9030
rect 23274 8622 23308 8638
rect 23370 9014 23404 9030
rect 23370 8622 23404 8638
rect 23466 9014 23500 9030
rect 23466 8622 23500 8638
rect 23562 9014 23596 9030
rect 23562 8622 23596 8638
rect 23658 9014 23692 9030
rect 23658 8622 23692 8638
rect 23754 9014 23788 9030
rect 23754 8622 23788 8638
rect 23850 9014 23884 9030
rect 23850 8622 23884 8638
rect 23946 9014 23980 9030
rect 23946 8622 23980 8638
rect 22058 8554 22074 8588
rect 22108 8554 22124 8588
rect 22250 8554 22266 8588
rect 22300 8554 22316 8588
rect 22442 8554 22458 8588
rect 22492 8554 22508 8588
rect 22634 8554 22650 8588
rect 22684 8554 22700 8588
rect 22826 8554 22842 8588
rect 22876 8554 22892 8588
rect 23018 8554 23034 8588
rect 23068 8554 23084 8588
rect 23210 8554 23226 8588
rect 23260 8554 23276 8588
rect 23402 8554 23418 8588
rect 23452 8554 23468 8588
rect 23594 8554 23610 8588
rect 23644 8554 23660 8588
rect 23786 8554 23802 8588
rect 23836 8554 23852 8588
rect 22058 8446 22074 8480
rect 22108 8446 22124 8480
rect 22250 8446 22266 8480
rect 22300 8446 22316 8480
rect 22442 8446 22458 8480
rect 22492 8446 22508 8480
rect 22634 8446 22650 8480
rect 22684 8446 22700 8480
rect 22826 8446 22842 8480
rect 22876 8446 22892 8480
rect 23018 8446 23034 8480
rect 23068 8446 23084 8480
rect 23210 8446 23226 8480
rect 23260 8446 23276 8480
rect 23402 8446 23418 8480
rect 23452 8446 23468 8480
rect 23594 8446 23610 8480
rect 23644 8446 23660 8480
rect 23786 8446 23802 8480
rect 23836 8446 23852 8480
rect 22026 8396 22060 8412
rect 22026 8004 22060 8020
rect 22122 8396 22156 8412
rect 22122 8004 22156 8020
rect 22218 8396 22252 8412
rect 22218 8004 22252 8020
rect 22314 8396 22348 8412
rect 22314 8004 22348 8020
rect 22410 8396 22444 8412
rect 22410 8004 22444 8020
rect 22506 8396 22540 8412
rect 22506 8004 22540 8020
rect 22602 8396 22636 8412
rect 22602 8004 22636 8020
rect 22698 8396 22732 8412
rect 22698 8004 22732 8020
rect 22794 8396 22828 8412
rect 22794 8004 22828 8020
rect 22890 8396 22924 8412
rect 22890 8004 22924 8020
rect 22986 8396 23020 8412
rect 22986 8004 23020 8020
rect 23082 8396 23116 8412
rect 23082 8004 23116 8020
rect 23178 8396 23212 8412
rect 23178 8004 23212 8020
rect 23274 8396 23308 8412
rect 23274 8004 23308 8020
rect 23370 8396 23404 8412
rect 23370 8004 23404 8020
rect 23466 8396 23500 8412
rect 23466 8004 23500 8020
rect 23562 8396 23596 8412
rect 23562 8004 23596 8020
rect 23658 8396 23692 8412
rect 23658 8004 23692 8020
rect 23754 8396 23788 8412
rect 23754 8004 23788 8020
rect 23850 8396 23884 8412
rect 23850 8004 23884 8020
rect 23946 8396 23980 8412
rect 23946 8004 23980 8020
rect 22154 7936 22170 7970
rect 22204 7936 22220 7970
rect 22346 7936 22362 7970
rect 22396 7936 22412 7970
rect 22538 7936 22554 7970
rect 22588 7936 22604 7970
rect 22730 7936 22746 7970
rect 22780 7936 22796 7970
rect 22922 7936 22938 7970
rect 22972 7936 22988 7970
rect 23114 7936 23130 7970
rect 23164 7936 23180 7970
rect 23306 7936 23322 7970
rect 23356 7936 23372 7970
rect 23498 7936 23514 7970
rect 23548 7936 23564 7970
rect 23690 7936 23706 7970
rect 23740 7936 23756 7970
rect 23882 7936 23898 7970
rect 23932 7936 23948 7970
rect 22154 7828 22170 7862
rect 22204 7828 22220 7862
rect 22346 7828 22362 7862
rect 22396 7828 22412 7862
rect 22538 7828 22554 7862
rect 22588 7828 22604 7862
rect 22730 7828 22746 7862
rect 22780 7828 22796 7862
rect 22922 7828 22938 7862
rect 22972 7828 22988 7862
rect 23114 7828 23130 7862
rect 23164 7828 23180 7862
rect 23306 7828 23322 7862
rect 23356 7828 23372 7862
rect 23498 7828 23514 7862
rect 23548 7828 23564 7862
rect 23690 7828 23706 7862
rect 23740 7828 23756 7862
rect 23882 7828 23898 7862
rect 23932 7828 23948 7862
rect 22026 7778 22060 7794
rect 22026 7386 22060 7402
rect 22122 7778 22156 7794
rect 22122 7386 22156 7402
rect 22218 7778 22252 7794
rect 22218 7386 22252 7402
rect 22314 7778 22348 7794
rect 22314 7386 22348 7402
rect 22410 7778 22444 7794
rect 22410 7386 22444 7402
rect 22506 7778 22540 7794
rect 22506 7386 22540 7402
rect 22602 7778 22636 7794
rect 22602 7386 22636 7402
rect 22698 7778 22732 7794
rect 22698 7386 22732 7402
rect 22794 7778 22828 7794
rect 22794 7386 22828 7402
rect 22890 7778 22924 7794
rect 22890 7386 22924 7402
rect 22986 7778 23020 7794
rect 22986 7386 23020 7402
rect 23082 7778 23116 7794
rect 23082 7386 23116 7402
rect 23178 7778 23212 7794
rect 23178 7386 23212 7402
rect 23274 7778 23308 7794
rect 23274 7386 23308 7402
rect 23370 7778 23404 7794
rect 23370 7386 23404 7402
rect 23466 7778 23500 7794
rect 23466 7386 23500 7402
rect 23562 7778 23596 7794
rect 23562 7386 23596 7402
rect 23658 7778 23692 7794
rect 23658 7386 23692 7402
rect 23754 7778 23788 7794
rect 23754 7386 23788 7402
rect 23850 7778 23884 7794
rect 23850 7386 23884 7402
rect 23946 7778 23980 7794
rect 23946 7386 23980 7402
rect 22058 7318 22074 7352
rect 22108 7318 22124 7352
rect 22250 7318 22266 7352
rect 22300 7318 22316 7352
rect 22442 7318 22458 7352
rect 22492 7318 22508 7352
rect 22634 7318 22650 7352
rect 22684 7318 22700 7352
rect 22826 7318 22842 7352
rect 22876 7318 22892 7352
rect 23018 7318 23034 7352
rect 23068 7318 23084 7352
rect 23210 7318 23226 7352
rect 23260 7318 23276 7352
rect 23402 7318 23418 7352
rect 23452 7318 23468 7352
rect 23594 7318 23610 7352
rect 23644 7318 23660 7352
rect 23786 7318 23802 7352
rect 23836 7318 23852 7352
rect 22058 7210 22074 7244
rect 22108 7210 22124 7244
rect 22250 7210 22266 7244
rect 22300 7210 22316 7244
rect 22442 7210 22458 7244
rect 22492 7210 22508 7244
rect 22634 7210 22650 7244
rect 22684 7210 22700 7244
rect 22826 7210 22842 7244
rect 22876 7210 22892 7244
rect 23018 7210 23034 7244
rect 23068 7210 23084 7244
rect 23210 7210 23226 7244
rect 23260 7210 23276 7244
rect 23402 7210 23418 7244
rect 23452 7210 23468 7244
rect 23594 7210 23610 7244
rect 23644 7210 23660 7244
rect 23786 7210 23802 7244
rect 23836 7210 23852 7244
rect 22026 7160 22060 7176
rect 22026 6768 22060 6784
rect 22122 7160 22156 7176
rect 22122 6768 22156 6784
rect 22218 7160 22252 7176
rect 22218 6768 22252 6784
rect 22314 7160 22348 7176
rect 22314 6768 22348 6784
rect 22410 7160 22444 7176
rect 22410 6768 22444 6784
rect 22506 7160 22540 7176
rect 22506 6768 22540 6784
rect 22602 7160 22636 7176
rect 22602 6768 22636 6784
rect 22698 7160 22732 7176
rect 22698 6768 22732 6784
rect 22794 7160 22828 7176
rect 22794 6768 22828 6784
rect 22890 7160 22924 7176
rect 22890 6768 22924 6784
rect 22986 7160 23020 7176
rect 22986 6768 23020 6784
rect 23082 7160 23116 7176
rect 23082 6768 23116 6784
rect 23178 7160 23212 7176
rect 23178 6768 23212 6784
rect 23274 7160 23308 7176
rect 23274 6768 23308 6784
rect 23370 7160 23404 7176
rect 23370 6768 23404 6784
rect 23466 7160 23500 7176
rect 23466 6768 23500 6784
rect 23562 7160 23596 7176
rect 23562 6768 23596 6784
rect 23658 7160 23692 7176
rect 23658 6768 23692 6784
rect 23754 7160 23788 7176
rect 23754 6768 23788 6784
rect 23850 7160 23884 7176
rect 23850 6768 23884 6784
rect 23946 7160 23980 7176
rect 23946 6768 23980 6784
rect 22154 6700 22170 6734
rect 22204 6700 22220 6734
rect 22346 6700 22362 6734
rect 22396 6700 22412 6734
rect 22538 6700 22554 6734
rect 22588 6700 22604 6734
rect 22730 6700 22746 6734
rect 22780 6700 22796 6734
rect 22922 6700 22938 6734
rect 22972 6700 22988 6734
rect 23114 6700 23130 6734
rect 23164 6700 23180 6734
rect 23306 6700 23322 6734
rect 23356 6700 23372 6734
rect 23498 6700 23514 6734
rect 23548 6700 23564 6734
rect 23690 6700 23706 6734
rect 23740 6700 23756 6734
rect 23882 6700 23898 6734
rect 23932 6700 23948 6734
rect 22154 6592 22170 6626
rect 22204 6592 22220 6626
rect 22346 6592 22362 6626
rect 22396 6592 22412 6626
rect 22538 6592 22554 6626
rect 22588 6592 22604 6626
rect 22730 6592 22746 6626
rect 22780 6592 22796 6626
rect 22922 6592 22938 6626
rect 22972 6592 22988 6626
rect 23114 6592 23130 6626
rect 23164 6592 23180 6626
rect 23306 6592 23322 6626
rect 23356 6592 23372 6626
rect 23498 6592 23514 6626
rect 23548 6592 23564 6626
rect 23690 6592 23706 6626
rect 23740 6592 23756 6626
rect 23882 6592 23898 6626
rect 23932 6592 23948 6626
rect 22026 6542 22060 6558
rect 22026 6150 22060 6166
rect 22122 6542 22156 6558
rect 22122 6150 22156 6166
rect 22218 6542 22252 6558
rect 22218 6150 22252 6166
rect 22314 6542 22348 6558
rect 22314 6150 22348 6166
rect 22410 6542 22444 6558
rect 22410 6150 22444 6166
rect 22506 6542 22540 6558
rect 22506 6150 22540 6166
rect 22602 6542 22636 6558
rect 22602 6150 22636 6166
rect 22698 6542 22732 6558
rect 22698 6150 22732 6166
rect 22794 6542 22828 6558
rect 22794 6150 22828 6166
rect 22890 6542 22924 6558
rect 22890 6150 22924 6166
rect 22986 6542 23020 6558
rect 22986 6150 23020 6166
rect 23082 6542 23116 6558
rect 23082 6150 23116 6166
rect 23178 6542 23212 6558
rect 23178 6150 23212 6166
rect 23274 6542 23308 6558
rect 23274 6150 23308 6166
rect 23370 6542 23404 6558
rect 23370 6150 23404 6166
rect 23466 6542 23500 6558
rect 23466 6150 23500 6166
rect 23562 6542 23596 6558
rect 23562 6150 23596 6166
rect 23658 6542 23692 6558
rect 23658 6150 23692 6166
rect 23754 6542 23788 6558
rect 23754 6150 23788 6166
rect 23850 6542 23884 6558
rect 23850 6150 23884 6166
rect 23946 6542 23980 6558
rect 23946 6150 23980 6166
rect 22058 6082 22074 6116
rect 22108 6082 22124 6116
rect 22250 6082 22266 6116
rect 22300 6082 22316 6116
rect 22442 6082 22458 6116
rect 22492 6082 22508 6116
rect 22634 6082 22650 6116
rect 22684 6082 22700 6116
rect 22826 6082 22842 6116
rect 22876 6082 22892 6116
rect 23018 6082 23034 6116
rect 23068 6082 23084 6116
rect 23210 6082 23226 6116
rect 23260 6082 23276 6116
rect 23402 6082 23418 6116
rect 23452 6082 23468 6116
rect 23594 6082 23610 6116
rect 23644 6082 23660 6116
rect 23786 6082 23802 6116
rect 23836 6082 23852 6116
rect 22058 5974 22074 6008
rect 22108 5974 22124 6008
rect 22250 5974 22266 6008
rect 22300 5974 22316 6008
rect 22442 5974 22458 6008
rect 22492 5974 22508 6008
rect 22634 5974 22650 6008
rect 22684 5974 22700 6008
rect 22826 5974 22842 6008
rect 22876 5974 22892 6008
rect 23018 5974 23034 6008
rect 23068 5974 23084 6008
rect 23210 5974 23226 6008
rect 23260 5974 23276 6008
rect 23402 5974 23418 6008
rect 23452 5974 23468 6008
rect 23594 5974 23610 6008
rect 23644 5974 23660 6008
rect 23786 5974 23802 6008
rect 23836 5974 23852 6008
rect 22026 5924 22060 5940
rect 22026 5532 22060 5548
rect 22122 5924 22156 5940
rect 22122 5532 22156 5548
rect 22218 5924 22252 5940
rect 22218 5532 22252 5548
rect 22314 5924 22348 5940
rect 22314 5532 22348 5548
rect 22410 5924 22444 5940
rect 22410 5532 22444 5548
rect 22506 5924 22540 5940
rect 22506 5532 22540 5548
rect 22602 5924 22636 5940
rect 22602 5532 22636 5548
rect 22698 5924 22732 5940
rect 22698 5532 22732 5548
rect 22794 5924 22828 5940
rect 22794 5532 22828 5548
rect 22890 5924 22924 5940
rect 22890 5532 22924 5548
rect 22986 5924 23020 5940
rect 22986 5532 23020 5548
rect 23082 5924 23116 5940
rect 23082 5532 23116 5548
rect 23178 5924 23212 5940
rect 23178 5532 23212 5548
rect 23274 5924 23308 5940
rect 23274 5532 23308 5548
rect 23370 5924 23404 5940
rect 23370 5532 23404 5548
rect 23466 5924 23500 5940
rect 23466 5532 23500 5548
rect 23562 5924 23596 5940
rect 23562 5532 23596 5548
rect 23658 5924 23692 5940
rect 23658 5532 23692 5548
rect 23754 5924 23788 5940
rect 23754 5532 23788 5548
rect 23850 5924 23884 5940
rect 23850 5532 23884 5548
rect 23946 5924 23980 5940
rect 23946 5532 23980 5548
rect 22154 5464 22170 5498
rect 22204 5464 22220 5498
rect 22346 5464 22362 5498
rect 22396 5464 22412 5498
rect 22538 5464 22554 5498
rect 22588 5464 22604 5498
rect 22730 5464 22746 5498
rect 22780 5464 22796 5498
rect 22922 5464 22938 5498
rect 22972 5464 22988 5498
rect 23114 5464 23130 5498
rect 23164 5464 23180 5498
rect 23306 5464 23322 5498
rect 23356 5464 23372 5498
rect 23498 5464 23514 5498
rect 23548 5464 23564 5498
rect 23690 5464 23706 5498
rect 23740 5464 23756 5498
rect 23882 5464 23898 5498
rect 23932 5464 23948 5498
rect 22154 5356 22170 5390
rect 22204 5356 22220 5390
rect 22346 5356 22362 5390
rect 22396 5356 22412 5390
rect 22538 5356 22554 5390
rect 22588 5356 22604 5390
rect 22730 5356 22746 5390
rect 22780 5356 22796 5390
rect 22922 5356 22938 5390
rect 22972 5356 22988 5390
rect 23114 5356 23130 5390
rect 23164 5356 23180 5390
rect 23306 5356 23322 5390
rect 23356 5356 23372 5390
rect 23498 5356 23514 5390
rect 23548 5356 23564 5390
rect 23690 5356 23706 5390
rect 23740 5356 23756 5390
rect 23882 5356 23898 5390
rect 23932 5356 23948 5390
rect 22026 5306 22060 5322
rect 22026 4914 22060 4930
rect 22122 5306 22156 5322
rect 22122 4914 22156 4930
rect 22218 5306 22252 5322
rect 22218 4914 22252 4930
rect 22314 5306 22348 5322
rect 22314 4914 22348 4930
rect 22410 5306 22444 5322
rect 22410 4914 22444 4930
rect 22506 5306 22540 5322
rect 22506 4914 22540 4930
rect 22602 5306 22636 5322
rect 22602 4914 22636 4930
rect 22698 5306 22732 5322
rect 22698 4914 22732 4930
rect 22794 5306 22828 5322
rect 22794 4914 22828 4930
rect 22890 5306 22924 5322
rect 22890 4914 22924 4930
rect 22986 5306 23020 5322
rect 22986 4914 23020 4930
rect 23082 5306 23116 5322
rect 23082 4914 23116 4930
rect 23178 5306 23212 5322
rect 23178 4914 23212 4930
rect 23274 5306 23308 5322
rect 23274 4914 23308 4930
rect 23370 5306 23404 5322
rect 23370 4914 23404 4930
rect 23466 5306 23500 5322
rect 23466 4914 23500 4930
rect 23562 5306 23596 5322
rect 23562 4914 23596 4930
rect 23658 5306 23692 5322
rect 23658 4914 23692 4930
rect 23754 5306 23788 5322
rect 23754 4914 23788 4930
rect 23850 5306 23884 5322
rect 23850 4914 23884 4930
rect 23946 5306 23980 5322
rect 23946 4914 23980 4930
rect 22058 4846 22074 4880
rect 22108 4846 22124 4880
rect 22250 4846 22266 4880
rect 22300 4846 22316 4880
rect 22442 4846 22458 4880
rect 22492 4846 22508 4880
rect 22634 4846 22650 4880
rect 22684 4846 22700 4880
rect 22826 4846 22842 4880
rect 22876 4846 22892 4880
rect 23018 4846 23034 4880
rect 23068 4846 23084 4880
rect 23210 4846 23226 4880
rect 23260 4846 23276 4880
rect 23402 4846 23418 4880
rect 23452 4846 23468 4880
rect 23594 4846 23610 4880
rect 23644 4846 23660 4880
rect 23786 4846 23802 4880
rect 23836 4846 23852 4880
rect 21912 4778 21946 4840
rect 24060 4778 24094 4840
rect 21912 4744 22008 4778
rect 23998 4744 24094 4778
rect 21100 4098 21134 4160
rect 19648 4064 20008 4098
rect 21038 4064 21134 4098
rect 116 3902 416 4064
rect 1640 3902 2216 4064
rect 3440 3902 4016 4064
rect 5248 3902 5816 4064
rect 14516 3902 14816 4064
rect 16040 3902 16616 4064
rect 17840 3902 18416 4064
rect 19648 3902 20216 4064
rect 112 3868 208 3902
rect 1568 3868 2008 3902
rect 3368 3868 3808 3902
rect 5168 3868 5608 3902
rect 6968 3868 7064 3902
rect 112 3806 146 3868
rect -8500 958 -8290 974
rect -8290 708 -8250 818
rect -8500 692 -8250 708
rect -8440 508 -8250 692
rect -8612 440 -8500 508
rect -8646 378 -8500 440
rect -10164 344 -10068 378
rect -8708 348 -8500 378
rect -8360 398 -8250 508
rect -8708 344 -8612 348
rect 1630 3806 1946 3868
rect 272 3766 288 3800
rect 456 3766 472 3800
rect 530 3766 546 3800
rect 714 3766 730 3800
rect 788 3766 804 3800
rect 972 3766 988 3800
rect 1046 3766 1062 3800
rect 1230 3766 1246 3800
rect 1304 3766 1320 3800
rect 1488 3766 1504 3800
rect 226 3716 260 3732
rect 226 3324 260 3340
rect 484 3716 518 3732
rect 484 3324 518 3340
rect 742 3716 776 3732
rect 742 3324 776 3340
rect 1000 3716 1034 3732
rect 1000 3324 1034 3340
rect 1258 3716 1292 3732
rect 1258 3324 1292 3340
rect 1516 3716 1550 3732
rect 1516 3324 1550 3340
rect 272 3256 288 3290
rect 456 3256 472 3290
rect 530 3256 546 3290
rect 714 3256 730 3290
rect 788 3256 804 3290
rect 972 3256 988 3290
rect 1046 3256 1062 3290
rect 1230 3256 1246 3290
rect 1304 3256 1320 3290
rect 1488 3256 1504 3290
rect 272 3148 288 3182
rect 456 3148 472 3182
rect 530 3148 546 3182
rect 714 3148 730 3182
rect 788 3148 804 3182
rect 972 3148 988 3182
rect 1046 3148 1062 3182
rect 1230 3148 1246 3182
rect 1304 3148 1320 3182
rect 1488 3148 1504 3182
rect 226 3098 260 3114
rect 226 2706 260 2722
rect 484 3098 518 3114
rect 484 2706 518 2722
rect 742 3098 776 3114
rect 742 2706 776 2722
rect 1000 3098 1034 3114
rect 1000 2706 1034 2722
rect 1258 3098 1292 3114
rect 1258 2706 1292 2722
rect 1516 3098 1550 3114
rect 1516 2706 1550 2722
rect 272 2638 288 2672
rect 456 2638 472 2672
rect 530 2638 546 2672
rect 714 2638 730 2672
rect 788 2638 804 2672
rect 972 2638 988 2672
rect 1046 2638 1062 2672
rect 1230 2638 1246 2672
rect 1304 2638 1320 2672
rect 1488 2638 1504 2672
rect 272 2530 288 2564
rect 456 2530 472 2564
rect 530 2530 546 2564
rect 714 2530 730 2564
rect 788 2530 804 2564
rect 972 2530 988 2564
rect 1046 2530 1062 2564
rect 1230 2530 1246 2564
rect 1304 2530 1320 2564
rect 1488 2530 1504 2564
rect 226 2480 260 2496
rect 226 2088 260 2104
rect 484 2480 518 2496
rect 484 2088 518 2104
rect 742 2480 776 2496
rect 742 2088 776 2104
rect 1000 2480 1034 2496
rect 1000 2088 1034 2104
rect 1258 2480 1292 2496
rect 1258 2088 1292 2104
rect 1516 2480 1550 2496
rect 1516 2088 1550 2104
rect 272 2020 288 2054
rect 456 2020 472 2054
rect 530 2020 546 2054
rect 714 2020 730 2054
rect 788 2020 804 2054
rect 972 2020 988 2054
rect 1046 2020 1062 2054
rect 1230 2020 1246 2054
rect 1304 2020 1320 2054
rect 1488 2020 1504 2054
rect 272 1912 288 1946
rect 456 1912 472 1946
rect 530 1912 546 1946
rect 714 1912 730 1946
rect 788 1912 804 1946
rect 972 1912 988 1946
rect 1046 1912 1062 1946
rect 1230 1912 1246 1946
rect 1304 1912 1320 1946
rect 1488 1912 1504 1946
rect 226 1862 260 1878
rect 226 1470 260 1486
rect 484 1862 518 1878
rect 484 1470 518 1486
rect 742 1862 776 1878
rect 742 1470 776 1486
rect 1000 1862 1034 1878
rect 1000 1470 1034 1486
rect 1258 1862 1292 1878
rect 1258 1470 1292 1486
rect 1516 1862 1550 1878
rect 1516 1470 1550 1486
rect 272 1402 288 1436
rect 456 1402 472 1436
rect 530 1402 546 1436
rect 714 1402 730 1436
rect 788 1402 804 1436
rect 972 1402 988 1436
rect 1046 1402 1062 1436
rect 1230 1402 1246 1436
rect 1304 1402 1320 1436
rect 1488 1402 1504 1436
rect 272 1294 288 1328
rect 456 1294 472 1328
rect 530 1294 546 1328
rect 714 1294 730 1328
rect 788 1294 804 1328
rect 972 1294 988 1328
rect 1046 1294 1062 1328
rect 1230 1294 1246 1328
rect 1304 1294 1320 1328
rect 1488 1294 1504 1328
rect 226 1244 260 1260
rect 226 852 260 868
rect 484 1244 518 1260
rect 484 852 518 868
rect 742 1244 776 1260
rect 742 852 776 868
rect 1000 1244 1034 1260
rect 1000 852 1034 868
rect 1258 1244 1292 1260
rect 1258 852 1292 868
rect 1516 1244 1550 1260
rect 1516 852 1550 868
rect 272 784 288 818
rect 456 784 472 818
rect 530 784 546 818
rect 714 784 730 818
rect 788 784 804 818
rect 972 784 988 818
rect 1046 784 1062 818
rect 1230 784 1246 818
rect 1304 784 1320 818
rect 1488 784 1504 818
rect 272 676 288 710
rect 456 676 472 710
rect 530 676 546 710
rect 714 676 730 710
rect 788 676 804 710
rect 972 676 988 710
rect 1046 676 1062 710
rect 1230 676 1246 710
rect 1304 676 1320 710
rect 1488 676 1504 710
rect 226 626 260 642
rect 226 234 260 250
rect 484 626 518 642
rect 484 234 518 250
rect 742 626 776 642
rect 742 234 776 250
rect 1000 626 1034 642
rect 1000 234 1034 250
rect 1258 626 1292 642
rect 1258 234 1292 250
rect 1516 626 1550 642
rect 1516 234 1550 250
rect 272 166 288 200
rect 456 166 472 200
rect 530 166 546 200
rect 714 166 730 200
rect 788 166 804 200
rect 972 166 988 200
rect 1046 166 1062 200
rect 1230 166 1246 200
rect 1304 166 1320 200
rect 1488 166 1504 200
rect 112 98 146 160
rect 1664 268 1912 3806
rect 1664 160 1696 268
rect 1630 98 1696 160
rect 112 64 208 98
rect 1568 68 1696 98
rect 1876 160 1912 268
rect 3430 3806 3746 3868
rect 2072 3766 2088 3800
rect 2256 3766 2272 3800
rect 2330 3766 2346 3800
rect 2514 3766 2530 3800
rect 2588 3766 2604 3800
rect 2772 3766 2788 3800
rect 2846 3766 2862 3800
rect 3030 3766 3046 3800
rect 3104 3766 3120 3800
rect 3288 3766 3304 3800
rect 2026 3716 2060 3732
rect 2026 3324 2060 3340
rect 2284 3716 2318 3732
rect 2284 3324 2318 3340
rect 2542 3716 2576 3732
rect 2542 3324 2576 3340
rect 2800 3716 2834 3732
rect 2800 3324 2834 3340
rect 3058 3716 3092 3732
rect 3058 3324 3092 3340
rect 3316 3716 3350 3732
rect 3316 3324 3350 3340
rect 2072 3256 2088 3290
rect 2256 3256 2272 3290
rect 2330 3256 2346 3290
rect 2514 3256 2530 3290
rect 2588 3256 2604 3290
rect 2772 3256 2788 3290
rect 2846 3256 2862 3290
rect 3030 3256 3046 3290
rect 3104 3256 3120 3290
rect 3288 3256 3304 3290
rect 2072 3148 2088 3182
rect 2256 3148 2272 3182
rect 2330 3148 2346 3182
rect 2514 3148 2530 3182
rect 2588 3148 2604 3182
rect 2772 3148 2788 3182
rect 2846 3148 2862 3182
rect 3030 3148 3046 3182
rect 3104 3148 3120 3182
rect 3288 3148 3304 3182
rect 2026 3098 2060 3114
rect 2026 2706 2060 2722
rect 2284 3098 2318 3114
rect 2284 2706 2318 2722
rect 2542 3098 2576 3114
rect 2542 2706 2576 2722
rect 2800 3098 2834 3114
rect 2800 2706 2834 2722
rect 3058 3098 3092 3114
rect 3058 2706 3092 2722
rect 3316 3098 3350 3114
rect 3316 2706 3350 2722
rect 2072 2638 2088 2672
rect 2256 2638 2272 2672
rect 2330 2638 2346 2672
rect 2514 2638 2530 2672
rect 2588 2638 2604 2672
rect 2772 2638 2788 2672
rect 2846 2638 2862 2672
rect 3030 2638 3046 2672
rect 3104 2638 3120 2672
rect 3288 2638 3304 2672
rect 2072 2530 2088 2564
rect 2256 2530 2272 2564
rect 2330 2530 2346 2564
rect 2514 2530 2530 2564
rect 2588 2530 2604 2564
rect 2772 2530 2788 2564
rect 2846 2530 2862 2564
rect 3030 2530 3046 2564
rect 3104 2530 3120 2564
rect 3288 2530 3304 2564
rect 2026 2480 2060 2496
rect 2026 2088 2060 2104
rect 2284 2480 2318 2496
rect 2284 2088 2318 2104
rect 2542 2480 2576 2496
rect 2542 2088 2576 2104
rect 2800 2480 2834 2496
rect 2800 2088 2834 2104
rect 3058 2480 3092 2496
rect 3058 2088 3092 2104
rect 3316 2480 3350 2496
rect 3316 2088 3350 2104
rect 2072 2020 2088 2054
rect 2256 2020 2272 2054
rect 2330 2020 2346 2054
rect 2514 2020 2530 2054
rect 2588 2020 2604 2054
rect 2772 2020 2788 2054
rect 2846 2020 2862 2054
rect 3030 2020 3046 2054
rect 3104 2020 3120 2054
rect 3288 2020 3304 2054
rect 2072 1912 2088 1946
rect 2256 1912 2272 1946
rect 2330 1912 2346 1946
rect 2514 1912 2530 1946
rect 2588 1912 2604 1946
rect 2772 1912 2788 1946
rect 2846 1912 2862 1946
rect 3030 1912 3046 1946
rect 3104 1912 3120 1946
rect 3288 1912 3304 1946
rect 2026 1862 2060 1878
rect 2026 1470 2060 1486
rect 2284 1862 2318 1878
rect 2284 1470 2318 1486
rect 2542 1862 2576 1878
rect 2542 1470 2576 1486
rect 2800 1862 2834 1878
rect 2800 1470 2834 1486
rect 3058 1862 3092 1878
rect 3058 1470 3092 1486
rect 3316 1862 3350 1878
rect 3316 1470 3350 1486
rect 2072 1402 2088 1436
rect 2256 1402 2272 1436
rect 2330 1402 2346 1436
rect 2514 1402 2530 1436
rect 2588 1402 2604 1436
rect 2772 1402 2788 1436
rect 2846 1402 2862 1436
rect 3030 1402 3046 1436
rect 3104 1402 3120 1436
rect 3288 1402 3304 1436
rect 2072 1294 2088 1328
rect 2256 1294 2272 1328
rect 2330 1294 2346 1328
rect 2514 1294 2530 1328
rect 2588 1294 2604 1328
rect 2772 1294 2788 1328
rect 2846 1294 2862 1328
rect 3030 1294 3046 1328
rect 3104 1294 3120 1328
rect 3288 1294 3304 1328
rect 2026 1244 2060 1260
rect 2026 852 2060 868
rect 2284 1244 2318 1260
rect 2284 852 2318 868
rect 2542 1244 2576 1260
rect 2542 852 2576 868
rect 2800 1244 2834 1260
rect 2800 852 2834 868
rect 3058 1244 3092 1260
rect 3058 852 3092 868
rect 3316 1244 3350 1260
rect 3316 852 3350 868
rect 2072 784 2088 818
rect 2256 784 2272 818
rect 2330 784 2346 818
rect 2514 784 2530 818
rect 2588 784 2604 818
rect 2772 784 2788 818
rect 2846 784 2862 818
rect 3030 784 3046 818
rect 3104 784 3120 818
rect 3288 784 3304 818
rect 2072 676 2088 710
rect 2256 676 2272 710
rect 2330 676 2346 710
rect 2514 676 2530 710
rect 2588 676 2604 710
rect 2772 676 2788 710
rect 2846 676 2862 710
rect 3030 676 3046 710
rect 3104 676 3120 710
rect 3288 676 3304 710
rect 2026 626 2060 642
rect 2026 234 2060 250
rect 2284 626 2318 642
rect 2284 234 2318 250
rect 2542 626 2576 642
rect 2542 234 2576 250
rect 2800 626 2834 642
rect 2800 234 2834 250
rect 3058 626 3092 642
rect 3058 234 3092 250
rect 3316 626 3350 642
rect 3316 234 3350 250
rect 2072 166 2088 200
rect 2256 166 2272 200
rect 2330 166 2346 200
rect 2514 166 2530 200
rect 2588 166 2604 200
rect 2772 166 2788 200
rect 2846 166 2862 200
rect 3030 166 3046 200
rect 3104 166 3120 200
rect 3288 166 3304 200
rect 1876 98 1946 160
rect 3464 276 3712 3806
rect 3464 160 3512 276
rect 3430 98 3512 160
rect 1876 68 2008 98
rect 1568 64 1664 68
rect 1912 64 2008 68
rect 3368 64 3512 98
rect 3692 160 3712 276
rect 5230 3806 5546 3868
rect 3872 3766 3888 3800
rect 4056 3766 4072 3800
rect 4130 3766 4146 3800
rect 4314 3766 4330 3800
rect 4388 3766 4404 3800
rect 4572 3766 4588 3800
rect 4646 3766 4662 3800
rect 4830 3766 4846 3800
rect 4904 3766 4920 3800
rect 5088 3766 5104 3800
rect 3826 3716 3860 3732
rect 3826 3324 3860 3340
rect 4084 3716 4118 3732
rect 4084 3324 4118 3340
rect 4342 3716 4376 3732
rect 4342 3324 4376 3340
rect 4600 3716 4634 3732
rect 4600 3324 4634 3340
rect 4858 3716 4892 3732
rect 4858 3324 4892 3340
rect 5116 3716 5150 3732
rect 5116 3324 5150 3340
rect 3872 3256 3888 3290
rect 4056 3256 4072 3290
rect 4130 3256 4146 3290
rect 4314 3256 4330 3290
rect 4388 3256 4404 3290
rect 4572 3256 4588 3290
rect 4646 3256 4662 3290
rect 4830 3256 4846 3290
rect 4904 3256 4920 3290
rect 5088 3256 5104 3290
rect 3872 3148 3888 3182
rect 4056 3148 4072 3182
rect 4130 3148 4146 3182
rect 4314 3148 4330 3182
rect 4388 3148 4404 3182
rect 4572 3148 4588 3182
rect 4646 3148 4662 3182
rect 4830 3148 4846 3182
rect 4904 3148 4920 3182
rect 5088 3148 5104 3182
rect 3826 3098 3860 3114
rect 3826 2706 3860 2722
rect 4084 3098 4118 3114
rect 4084 2706 4118 2722
rect 4342 3098 4376 3114
rect 4342 2706 4376 2722
rect 4600 3098 4634 3114
rect 4600 2706 4634 2722
rect 4858 3098 4892 3114
rect 4858 2706 4892 2722
rect 5116 3098 5150 3114
rect 5116 2706 5150 2722
rect 3872 2638 3888 2672
rect 4056 2638 4072 2672
rect 4130 2638 4146 2672
rect 4314 2638 4330 2672
rect 4388 2638 4404 2672
rect 4572 2638 4588 2672
rect 4646 2638 4662 2672
rect 4830 2638 4846 2672
rect 4904 2638 4920 2672
rect 5088 2638 5104 2672
rect 3872 2530 3888 2564
rect 4056 2530 4072 2564
rect 4130 2530 4146 2564
rect 4314 2530 4330 2564
rect 4388 2530 4404 2564
rect 4572 2530 4588 2564
rect 4646 2530 4662 2564
rect 4830 2530 4846 2564
rect 4904 2530 4920 2564
rect 5088 2530 5104 2564
rect 3826 2480 3860 2496
rect 3826 2088 3860 2104
rect 4084 2480 4118 2496
rect 4084 2088 4118 2104
rect 4342 2480 4376 2496
rect 4342 2088 4376 2104
rect 4600 2480 4634 2496
rect 4600 2088 4634 2104
rect 4858 2480 4892 2496
rect 4858 2088 4892 2104
rect 5116 2480 5150 2496
rect 5116 2088 5150 2104
rect 3872 2020 3888 2054
rect 4056 2020 4072 2054
rect 4130 2020 4146 2054
rect 4314 2020 4330 2054
rect 4388 2020 4404 2054
rect 4572 2020 4588 2054
rect 4646 2020 4662 2054
rect 4830 2020 4846 2054
rect 4904 2020 4920 2054
rect 5088 2020 5104 2054
rect 3872 1912 3888 1946
rect 4056 1912 4072 1946
rect 4130 1912 4146 1946
rect 4314 1912 4330 1946
rect 4388 1912 4404 1946
rect 4572 1912 4588 1946
rect 4646 1912 4662 1946
rect 4830 1912 4846 1946
rect 4904 1912 4920 1946
rect 5088 1912 5104 1946
rect 3826 1862 3860 1878
rect 3826 1470 3860 1486
rect 4084 1862 4118 1878
rect 4084 1470 4118 1486
rect 4342 1862 4376 1878
rect 4342 1470 4376 1486
rect 4600 1862 4634 1878
rect 4600 1470 4634 1486
rect 4858 1862 4892 1878
rect 4858 1470 4892 1486
rect 5116 1862 5150 1878
rect 5116 1470 5150 1486
rect 3872 1402 3888 1436
rect 4056 1402 4072 1436
rect 4130 1402 4146 1436
rect 4314 1402 4330 1436
rect 4388 1402 4404 1436
rect 4572 1402 4588 1436
rect 4646 1402 4662 1436
rect 4830 1402 4846 1436
rect 4904 1402 4920 1436
rect 5088 1402 5104 1436
rect 3872 1294 3888 1328
rect 4056 1294 4072 1328
rect 4130 1294 4146 1328
rect 4314 1294 4330 1328
rect 4388 1294 4404 1328
rect 4572 1294 4588 1328
rect 4646 1294 4662 1328
rect 4830 1294 4846 1328
rect 4904 1294 4920 1328
rect 5088 1294 5104 1328
rect 3826 1244 3860 1260
rect 3826 852 3860 868
rect 4084 1244 4118 1260
rect 4084 852 4118 868
rect 4342 1244 4376 1260
rect 4342 852 4376 868
rect 4600 1244 4634 1260
rect 4600 852 4634 868
rect 4858 1244 4892 1260
rect 4858 852 4892 868
rect 5116 1244 5150 1260
rect 5116 852 5150 868
rect 3872 784 3888 818
rect 4056 784 4072 818
rect 4130 784 4146 818
rect 4314 784 4330 818
rect 4388 784 4404 818
rect 4572 784 4588 818
rect 4646 784 4662 818
rect 4830 784 4846 818
rect 4904 784 4920 818
rect 5088 784 5104 818
rect 3872 676 3888 710
rect 4056 676 4072 710
rect 4130 676 4146 710
rect 4314 676 4330 710
rect 4388 676 4404 710
rect 4572 676 4588 710
rect 4646 676 4662 710
rect 4830 676 4846 710
rect 4904 676 4920 710
rect 5088 676 5104 710
rect 3826 626 3860 642
rect 3826 234 3860 250
rect 4084 626 4118 642
rect 4084 234 4118 250
rect 4342 626 4376 642
rect 4342 234 4376 250
rect 4600 626 4634 642
rect 4600 234 4634 250
rect 4858 626 4892 642
rect 4858 234 4892 250
rect 5116 626 5150 642
rect 5116 234 5150 250
rect 3872 166 3888 200
rect 4056 166 4072 200
rect 4130 166 4146 200
rect 4314 166 4330 200
rect 4388 166 4404 200
rect 4572 166 4588 200
rect 4646 166 4662 200
rect 4830 166 4846 200
rect 4904 166 4920 200
rect 5088 166 5104 200
rect 3692 98 3746 160
rect 5264 276 5512 3806
rect 5264 160 5288 276
rect 5230 98 5288 160
rect 3692 64 3808 98
rect 5168 64 5288 98
rect 5468 160 5512 276
rect 7030 3806 7064 3868
rect 5672 3766 5688 3800
rect 5856 3766 5872 3800
rect 5930 3766 5946 3800
rect 6114 3766 6130 3800
rect 6188 3766 6204 3800
rect 6372 3766 6388 3800
rect 6446 3766 6462 3800
rect 6630 3766 6646 3800
rect 6704 3766 6720 3800
rect 6888 3766 6904 3800
rect 5626 3716 5660 3732
rect 5626 3324 5660 3340
rect 5884 3716 5918 3732
rect 5884 3324 5918 3340
rect 6142 3716 6176 3732
rect 6142 3324 6176 3340
rect 6400 3716 6434 3732
rect 6400 3324 6434 3340
rect 6658 3716 6692 3732
rect 6658 3324 6692 3340
rect 6916 3716 6950 3732
rect 6916 3324 6950 3340
rect 5672 3256 5688 3290
rect 5856 3256 5872 3290
rect 5930 3256 5946 3290
rect 6114 3256 6130 3290
rect 6188 3256 6204 3290
rect 6372 3256 6388 3290
rect 6446 3256 6462 3290
rect 6630 3256 6646 3290
rect 6704 3256 6720 3290
rect 6888 3256 6904 3290
rect 5672 3148 5688 3182
rect 5856 3148 5872 3182
rect 5930 3148 5946 3182
rect 6114 3148 6130 3182
rect 6188 3148 6204 3182
rect 6372 3148 6388 3182
rect 6446 3148 6462 3182
rect 6630 3148 6646 3182
rect 6704 3148 6720 3182
rect 6888 3148 6904 3182
rect 5626 3098 5660 3114
rect 5626 2706 5660 2722
rect 5884 3098 5918 3114
rect 5884 2706 5918 2722
rect 6142 3098 6176 3114
rect 6142 2706 6176 2722
rect 6400 3098 6434 3114
rect 6400 2706 6434 2722
rect 6658 3098 6692 3114
rect 6658 2706 6692 2722
rect 6916 3098 6950 3114
rect 6916 2706 6950 2722
rect 5672 2638 5688 2672
rect 5856 2638 5872 2672
rect 5930 2638 5946 2672
rect 6114 2638 6130 2672
rect 6188 2638 6204 2672
rect 6372 2638 6388 2672
rect 6446 2638 6462 2672
rect 6630 2638 6646 2672
rect 6704 2638 6720 2672
rect 6888 2638 6904 2672
rect 5672 2530 5688 2564
rect 5856 2530 5872 2564
rect 5930 2530 5946 2564
rect 6114 2530 6130 2564
rect 6188 2530 6204 2564
rect 6372 2530 6388 2564
rect 6446 2530 6462 2564
rect 6630 2530 6646 2564
rect 6704 2530 6720 2564
rect 6888 2530 6904 2564
rect 5626 2480 5660 2496
rect 5626 2088 5660 2104
rect 5884 2480 5918 2496
rect 5884 2088 5918 2104
rect 6142 2480 6176 2496
rect 6142 2088 6176 2104
rect 6400 2480 6434 2496
rect 6400 2088 6434 2104
rect 6658 2480 6692 2496
rect 6658 2088 6692 2104
rect 6916 2480 6950 2496
rect 6916 2088 6950 2104
rect 5672 2020 5688 2054
rect 5856 2020 5872 2054
rect 5930 2020 5946 2054
rect 6114 2020 6130 2054
rect 6188 2020 6204 2054
rect 6372 2020 6388 2054
rect 6446 2020 6462 2054
rect 6630 2020 6646 2054
rect 6704 2020 6720 2054
rect 6888 2020 6904 2054
rect 5672 1912 5688 1946
rect 5856 1912 5872 1946
rect 5930 1912 5946 1946
rect 6114 1912 6130 1946
rect 6188 1912 6204 1946
rect 6372 1912 6388 1946
rect 6446 1912 6462 1946
rect 6630 1912 6646 1946
rect 6704 1912 6720 1946
rect 6888 1912 6904 1946
rect 5626 1862 5660 1878
rect 5626 1470 5660 1486
rect 5884 1862 5918 1878
rect 5884 1470 5918 1486
rect 6142 1862 6176 1878
rect 6142 1470 6176 1486
rect 6400 1862 6434 1878
rect 6400 1470 6434 1486
rect 6658 1862 6692 1878
rect 6658 1470 6692 1486
rect 6916 1862 6950 1878
rect 6916 1470 6950 1486
rect 5672 1402 5688 1436
rect 5856 1402 5872 1436
rect 5930 1402 5946 1436
rect 6114 1402 6130 1436
rect 6188 1402 6204 1436
rect 6372 1402 6388 1436
rect 6446 1402 6462 1436
rect 6630 1402 6646 1436
rect 6704 1402 6720 1436
rect 6888 1402 6904 1436
rect 5672 1294 5688 1328
rect 5856 1294 5872 1328
rect 5930 1294 5946 1328
rect 6114 1294 6130 1328
rect 6188 1294 6204 1328
rect 6372 1294 6388 1328
rect 6446 1294 6462 1328
rect 6630 1294 6646 1328
rect 6704 1294 6720 1328
rect 6888 1294 6904 1328
rect 5626 1244 5660 1260
rect 5626 852 5660 868
rect 5884 1244 5918 1260
rect 5884 852 5918 868
rect 6142 1244 6176 1260
rect 6142 852 6176 868
rect 6400 1244 6434 1260
rect 6400 852 6434 868
rect 6658 1244 6692 1260
rect 6658 852 6692 868
rect 6916 1244 6950 1260
rect 6916 852 6950 868
rect 5672 784 5688 818
rect 5856 784 5872 818
rect 5930 784 5946 818
rect 6114 784 6130 818
rect 6188 784 6204 818
rect 6372 784 6388 818
rect 6446 784 6462 818
rect 6630 784 6646 818
rect 6704 784 6720 818
rect 6888 784 6904 818
rect 5672 676 5688 710
rect 5856 676 5872 710
rect 5930 676 5946 710
rect 6114 676 6130 710
rect 6188 676 6204 710
rect 6372 676 6388 710
rect 6446 676 6462 710
rect 6630 676 6646 710
rect 6704 676 6720 710
rect 6888 676 6904 710
rect 5626 626 5660 642
rect 5626 234 5660 250
rect 5884 626 5918 642
rect 5884 234 5918 250
rect 6142 626 6176 642
rect 6142 234 6176 250
rect 6400 626 6434 642
rect 6400 234 6434 250
rect 6658 626 6692 642
rect 6658 234 6692 250
rect 6916 626 6950 642
rect 6916 234 6950 250
rect 5672 166 5688 200
rect 5856 166 5872 200
rect 5930 166 5946 200
rect 6114 166 6130 200
rect 6188 166 6204 200
rect 6372 166 6388 200
rect 6446 166 6462 200
rect 6630 166 6646 200
rect 6704 166 6720 200
rect 6888 166 6904 200
rect 5468 98 5546 160
rect 7030 98 7064 160
rect 5468 64 5608 98
rect 6968 64 7064 98
rect 14512 3868 14608 3902
rect 15968 3868 16408 3902
rect 17768 3868 18208 3902
rect 19568 3868 20008 3902
rect 21368 3868 21464 3902
rect 14512 3806 14546 3868
rect 16030 3806 16346 3868
rect 14672 3766 14688 3800
rect 14856 3766 14872 3800
rect 14930 3766 14946 3800
rect 15114 3766 15130 3800
rect 15188 3766 15204 3800
rect 15372 3766 15388 3800
rect 15446 3766 15462 3800
rect 15630 3766 15646 3800
rect 15704 3766 15720 3800
rect 15888 3766 15904 3800
rect 14626 3716 14660 3732
rect 14626 3324 14660 3340
rect 14884 3716 14918 3732
rect 14884 3324 14918 3340
rect 15142 3716 15176 3732
rect 15142 3324 15176 3340
rect 15400 3716 15434 3732
rect 15400 3324 15434 3340
rect 15658 3716 15692 3732
rect 15658 3324 15692 3340
rect 15916 3716 15950 3732
rect 15916 3324 15950 3340
rect 14672 3256 14688 3290
rect 14856 3256 14872 3290
rect 14930 3256 14946 3290
rect 15114 3256 15130 3290
rect 15188 3256 15204 3290
rect 15372 3256 15388 3290
rect 15446 3256 15462 3290
rect 15630 3256 15646 3290
rect 15704 3256 15720 3290
rect 15888 3256 15904 3290
rect 14672 3148 14688 3182
rect 14856 3148 14872 3182
rect 14930 3148 14946 3182
rect 15114 3148 15130 3182
rect 15188 3148 15204 3182
rect 15372 3148 15388 3182
rect 15446 3148 15462 3182
rect 15630 3148 15646 3182
rect 15704 3148 15720 3182
rect 15888 3148 15904 3182
rect 14626 3098 14660 3114
rect 14626 2706 14660 2722
rect 14884 3098 14918 3114
rect 14884 2706 14918 2722
rect 15142 3098 15176 3114
rect 15142 2706 15176 2722
rect 15400 3098 15434 3114
rect 15400 2706 15434 2722
rect 15658 3098 15692 3114
rect 15658 2706 15692 2722
rect 15916 3098 15950 3114
rect 15916 2706 15950 2722
rect 14672 2638 14688 2672
rect 14856 2638 14872 2672
rect 14930 2638 14946 2672
rect 15114 2638 15130 2672
rect 15188 2638 15204 2672
rect 15372 2638 15388 2672
rect 15446 2638 15462 2672
rect 15630 2638 15646 2672
rect 15704 2638 15720 2672
rect 15888 2638 15904 2672
rect 14672 2530 14688 2564
rect 14856 2530 14872 2564
rect 14930 2530 14946 2564
rect 15114 2530 15130 2564
rect 15188 2530 15204 2564
rect 15372 2530 15388 2564
rect 15446 2530 15462 2564
rect 15630 2530 15646 2564
rect 15704 2530 15720 2564
rect 15888 2530 15904 2564
rect 14626 2480 14660 2496
rect 14626 2088 14660 2104
rect 14884 2480 14918 2496
rect 14884 2088 14918 2104
rect 15142 2480 15176 2496
rect 15142 2088 15176 2104
rect 15400 2480 15434 2496
rect 15400 2088 15434 2104
rect 15658 2480 15692 2496
rect 15658 2088 15692 2104
rect 15916 2480 15950 2496
rect 15916 2088 15950 2104
rect 14672 2020 14688 2054
rect 14856 2020 14872 2054
rect 14930 2020 14946 2054
rect 15114 2020 15130 2054
rect 15188 2020 15204 2054
rect 15372 2020 15388 2054
rect 15446 2020 15462 2054
rect 15630 2020 15646 2054
rect 15704 2020 15720 2054
rect 15888 2020 15904 2054
rect 14672 1912 14688 1946
rect 14856 1912 14872 1946
rect 14930 1912 14946 1946
rect 15114 1912 15130 1946
rect 15188 1912 15204 1946
rect 15372 1912 15388 1946
rect 15446 1912 15462 1946
rect 15630 1912 15646 1946
rect 15704 1912 15720 1946
rect 15888 1912 15904 1946
rect 14626 1862 14660 1878
rect 14626 1470 14660 1486
rect 14884 1862 14918 1878
rect 14884 1470 14918 1486
rect 15142 1862 15176 1878
rect 15142 1470 15176 1486
rect 15400 1862 15434 1878
rect 15400 1470 15434 1486
rect 15658 1862 15692 1878
rect 15658 1470 15692 1486
rect 15916 1862 15950 1878
rect 15916 1470 15950 1486
rect 14672 1402 14688 1436
rect 14856 1402 14872 1436
rect 14930 1402 14946 1436
rect 15114 1402 15130 1436
rect 15188 1402 15204 1436
rect 15372 1402 15388 1436
rect 15446 1402 15462 1436
rect 15630 1402 15646 1436
rect 15704 1402 15720 1436
rect 15888 1402 15904 1436
rect 14672 1294 14688 1328
rect 14856 1294 14872 1328
rect 14930 1294 14946 1328
rect 15114 1294 15130 1328
rect 15188 1294 15204 1328
rect 15372 1294 15388 1328
rect 15446 1294 15462 1328
rect 15630 1294 15646 1328
rect 15704 1294 15720 1328
rect 15888 1294 15904 1328
rect 14626 1244 14660 1260
rect 14626 852 14660 868
rect 14884 1244 14918 1260
rect 14884 852 14918 868
rect 15142 1244 15176 1260
rect 15142 852 15176 868
rect 15400 1244 15434 1260
rect 15400 852 15434 868
rect 15658 1244 15692 1260
rect 15658 852 15692 868
rect 15916 1244 15950 1260
rect 15916 852 15950 868
rect 14672 784 14688 818
rect 14856 784 14872 818
rect 14930 784 14946 818
rect 15114 784 15130 818
rect 15188 784 15204 818
rect 15372 784 15388 818
rect 15446 784 15462 818
rect 15630 784 15646 818
rect 15704 784 15720 818
rect 15888 784 15904 818
rect 14672 676 14688 710
rect 14856 676 14872 710
rect 14930 676 14946 710
rect 15114 676 15130 710
rect 15188 676 15204 710
rect 15372 676 15388 710
rect 15446 676 15462 710
rect 15630 676 15646 710
rect 15704 676 15720 710
rect 15888 676 15904 710
rect 14626 626 14660 642
rect 14626 234 14660 250
rect 14884 626 14918 642
rect 14884 234 14918 250
rect 15142 626 15176 642
rect 15142 234 15176 250
rect 15400 626 15434 642
rect 15400 234 15434 250
rect 15658 626 15692 642
rect 15658 234 15692 250
rect 15916 626 15950 642
rect 15916 234 15950 250
rect 14672 166 14688 200
rect 14856 166 14872 200
rect 14930 166 14946 200
rect 15114 166 15130 200
rect 15188 166 15204 200
rect 15372 166 15388 200
rect 15446 166 15462 200
rect 15630 166 15646 200
rect 15704 166 15720 200
rect 15888 166 15904 200
rect 14512 98 14546 160
rect 16064 268 16312 3806
rect 16064 160 16096 268
rect 16030 98 16096 160
rect 14512 64 14608 98
rect 15968 68 16096 98
rect 16276 160 16312 268
rect 17830 3806 18146 3868
rect 16472 3766 16488 3800
rect 16656 3766 16672 3800
rect 16730 3766 16746 3800
rect 16914 3766 16930 3800
rect 16988 3766 17004 3800
rect 17172 3766 17188 3800
rect 17246 3766 17262 3800
rect 17430 3766 17446 3800
rect 17504 3766 17520 3800
rect 17688 3766 17704 3800
rect 16426 3716 16460 3732
rect 16426 3324 16460 3340
rect 16684 3716 16718 3732
rect 16684 3324 16718 3340
rect 16942 3716 16976 3732
rect 16942 3324 16976 3340
rect 17200 3716 17234 3732
rect 17200 3324 17234 3340
rect 17458 3716 17492 3732
rect 17458 3324 17492 3340
rect 17716 3716 17750 3732
rect 17716 3324 17750 3340
rect 16472 3256 16488 3290
rect 16656 3256 16672 3290
rect 16730 3256 16746 3290
rect 16914 3256 16930 3290
rect 16988 3256 17004 3290
rect 17172 3256 17188 3290
rect 17246 3256 17262 3290
rect 17430 3256 17446 3290
rect 17504 3256 17520 3290
rect 17688 3256 17704 3290
rect 16472 3148 16488 3182
rect 16656 3148 16672 3182
rect 16730 3148 16746 3182
rect 16914 3148 16930 3182
rect 16988 3148 17004 3182
rect 17172 3148 17188 3182
rect 17246 3148 17262 3182
rect 17430 3148 17446 3182
rect 17504 3148 17520 3182
rect 17688 3148 17704 3182
rect 16426 3098 16460 3114
rect 16426 2706 16460 2722
rect 16684 3098 16718 3114
rect 16684 2706 16718 2722
rect 16942 3098 16976 3114
rect 16942 2706 16976 2722
rect 17200 3098 17234 3114
rect 17200 2706 17234 2722
rect 17458 3098 17492 3114
rect 17458 2706 17492 2722
rect 17716 3098 17750 3114
rect 17716 2706 17750 2722
rect 16472 2638 16488 2672
rect 16656 2638 16672 2672
rect 16730 2638 16746 2672
rect 16914 2638 16930 2672
rect 16988 2638 17004 2672
rect 17172 2638 17188 2672
rect 17246 2638 17262 2672
rect 17430 2638 17446 2672
rect 17504 2638 17520 2672
rect 17688 2638 17704 2672
rect 16472 2530 16488 2564
rect 16656 2530 16672 2564
rect 16730 2530 16746 2564
rect 16914 2530 16930 2564
rect 16988 2530 17004 2564
rect 17172 2530 17188 2564
rect 17246 2530 17262 2564
rect 17430 2530 17446 2564
rect 17504 2530 17520 2564
rect 17688 2530 17704 2564
rect 16426 2480 16460 2496
rect 16426 2088 16460 2104
rect 16684 2480 16718 2496
rect 16684 2088 16718 2104
rect 16942 2480 16976 2496
rect 16942 2088 16976 2104
rect 17200 2480 17234 2496
rect 17200 2088 17234 2104
rect 17458 2480 17492 2496
rect 17458 2088 17492 2104
rect 17716 2480 17750 2496
rect 17716 2088 17750 2104
rect 16472 2020 16488 2054
rect 16656 2020 16672 2054
rect 16730 2020 16746 2054
rect 16914 2020 16930 2054
rect 16988 2020 17004 2054
rect 17172 2020 17188 2054
rect 17246 2020 17262 2054
rect 17430 2020 17446 2054
rect 17504 2020 17520 2054
rect 17688 2020 17704 2054
rect 16472 1912 16488 1946
rect 16656 1912 16672 1946
rect 16730 1912 16746 1946
rect 16914 1912 16930 1946
rect 16988 1912 17004 1946
rect 17172 1912 17188 1946
rect 17246 1912 17262 1946
rect 17430 1912 17446 1946
rect 17504 1912 17520 1946
rect 17688 1912 17704 1946
rect 16426 1862 16460 1878
rect 16426 1470 16460 1486
rect 16684 1862 16718 1878
rect 16684 1470 16718 1486
rect 16942 1862 16976 1878
rect 16942 1470 16976 1486
rect 17200 1862 17234 1878
rect 17200 1470 17234 1486
rect 17458 1862 17492 1878
rect 17458 1470 17492 1486
rect 17716 1862 17750 1878
rect 17716 1470 17750 1486
rect 16472 1402 16488 1436
rect 16656 1402 16672 1436
rect 16730 1402 16746 1436
rect 16914 1402 16930 1436
rect 16988 1402 17004 1436
rect 17172 1402 17188 1436
rect 17246 1402 17262 1436
rect 17430 1402 17446 1436
rect 17504 1402 17520 1436
rect 17688 1402 17704 1436
rect 16472 1294 16488 1328
rect 16656 1294 16672 1328
rect 16730 1294 16746 1328
rect 16914 1294 16930 1328
rect 16988 1294 17004 1328
rect 17172 1294 17188 1328
rect 17246 1294 17262 1328
rect 17430 1294 17446 1328
rect 17504 1294 17520 1328
rect 17688 1294 17704 1328
rect 16426 1244 16460 1260
rect 16426 852 16460 868
rect 16684 1244 16718 1260
rect 16684 852 16718 868
rect 16942 1244 16976 1260
rect 16942 852 16976 868
rect 17200 1244 17234 1260
rect 17200 852 17234 868
rect 17458 1244 17492 1260
rect 17458 852 17492 868
rect 17716 1244 17750 1260
rect 17716 852 17750 868
rect 16472 784 16488 818
rect 16656 784 16672 818
rect 16730 784 16746 818
rect 16914 784 16930 818
rect 16988 784 17004 818
rect 17172 784 17188 818
rect 17246 784 17262 818
rect 17430 784 17446 818
rect 17504 784 17520 818
rect 17688 784 17704 818
rect 16472 676 16488 710
rect 16656 676 16672 710
rect 16730 676 16746 710
rect 16914 676 16930 710
rect 16988 676 17004 710
rect 17172 676 17188 710
rect 17246 676 17262 710
rect 17430 676 17446 710
rect 17504 676 17520 710
rect 17688 676 17704 710
rect 16426 626 16460 642
rect 16426 234 16460 250
rect 16684 626 16718 642
rect 16684 234 16718 250
rect 16942 626 16976 642
rect 16942 234 16976 250
rect 17200 626 17234 642
rect 17200 234 17234 250
rect 17458 626 17492 642
rect 17458 234 17492 250
rect 17716 626 17750 642
rect 17716 234 17750 250
rect 16472 166 16488 200
rect 16656 166 16672 200
rect 16730 166 16746 200
rect 16914 166 16930 200
rect 16988 166 17004 200
rect 17172 166 17188 200
rect 17246 166 17262 200
rect 17430 166 17446 200
rect 17504 166 17520 200
rect 17688 166 17704 200
rect 16276 98 16346 160
rect 17864 276 18112 3806
rect 17864 160 17912 276
rect 17830 98 17912 160
rect 16276 68 16408 98
rect 15968 64 16064 68
rect 16312 64 16408 68
rect 17768 64 17912 98
rect 18092 160 18112 276
rect 19630 3806 19946 3868
rect 18272 3766 18288 3800
rect 18456 3766 18472 3800
rect 18530 3766 18546 3800
rect 18714 3766 18730 3800
rect 18788 3766 18804 3800
rect 18972 3766 18988 3800
rect 19046 3766 19062 3800
rect 19230 3766 19246 3800
rect 19304 3766 19320 3800
rect 19488 3766 19504 3800
rect 18226 3716 18260 3732
rect 18226 3324 18260 3340
rect 18484 3716 18518 3732
rect 18484 3324 18518 3340
rect 18742 3716 18776 3732
rect 18742 3324 18776 3340
rect 19000 3716 19034 3732
rect 19000 3324 19034 3340
rect 19258 3716 19292 3732
rect 19258 3324 19292 3340
rect 19516 3716 19550 3732
rect 19516 3324 19550 3340
rect 18272 3256 18288 3290
rect 18456 3256 18472 3290
rect 18530 3256 18546 3290
rect 18714 3256 18730 3290
rect 18788 3256 18804 3290
rect 18972 3256 18988 3290
rect 19046 3256 19062 3290
rect 19230 3256 19246 3290
rect 19304 3256 19320 3290
rect 19488 3256 19504 3290
rect 18272 3148 18288 3182
rect 18456 3148 18472 3182
rect 18530 3148 18546 3182
rect 18714 3148 18730 3182
rect 18788 3148 18804 3182
rect 18972 3148 18988 3182
rect 19046 3148 19062 3182
rect 19230 3148 19246 3182
rect 19304 3148 19320 3182
rect 19488 3148 19504 3182
rect 18226 3098 18260 3114
rect 18226 2706 18260 2722
rect 18484 3098 18518 3114
rect 18484 2706 18518 2722
rect 18742 3098 18776 3114
rect 18742 2706 18776 2722
rect 19000 3098 19034 3114
rect 19000 2706 19034 2722
rect 19258 3098 19292 3114
rect 19258 2706 19292 2722
rect 19516 3098 19550 3114
rect 19516 2706 19550 2722
rect 18272 2638 18288 2672
rect 18456 2638 18472 2672
rect 18530 2638 18546 2672
rect 18714 2638 18730 2672
rect 18788 2638 18804 2672
rect 18972 2638 18988 2672
rect 19046 2638 19062 2672
rect 19230 2638 19246 2672
rect 19304 2638 19320 2672
rect 19488 2638 19504 2672
rect 18272 2530 18288 2564
rect 18456 2530 18472 2564
rect 18530 2530 18546 2564
rect 18714 2530 18730 2564
rect 18788 2530 18804 2564
rect 18972 2530 18988 2564
rect 19046 2530 19062 2564
rect 19230 2530 19246 2564
rect 19304 2530 19320 2564
rect 19488 2530 19504 2564
rect 18226 2480 18260 2496
rect 18226 2088 18260 2104
rect 18484 2480 18518 2496
rect 18484 2088 18518 2104
rect 18742 2480 18776 2496
rect 18742 2088 18776 2104
rect 19000 2480 19034 2496
rect 19000 2088 19034 2104
rect 19258 2480 19292 2496
rect 19258 2088 19292 2104
rect 19516 2480 19550 2496
rect 19516 2088 19550 2104
rect 18272 2020 18288 2054
rect 18456 2020 18472 2054
rect 18530 2020 18546 2054
rect 18714 2020 18730 2054
rect 18788 2020 18804 2054
rect 18972 2020 18988 2054
rect 19046 2020 19062 2054
rect 19230 2020 19246 2054
rect 19304 2020 19320 2054
rect 19488 2020 19504 2054
rect 18272 1912 18288 1946
rect 18456 1912 18472 1946
rect 18530 1912 18546 1946
rect 18714 1912 18730 1946
rect 18788 1912 18804 1946
rect 18972 1912 18988 1946
rect 19046 1912 19062 1946
rect 19230 1912 19246 1946
rect 19304 1912 19320 1946
rect 19488 1912 19504 1946
rect 18226 1862 18260 1878
rect 18226 1470 18260 1486
rect 18484 1862 18518 1878
rect 18484 1470 18518 1486
rect 18742 1862 18776 1878
rect 18742 1470 18776 1486
rect 19000 1862 19034 1878
rect 19000 1470 19034 1486
rect 19258 1862 19292 1878
rect 19258 1470 19292 1486
rect 19516 1862 19550 1878
rect 19516 1470 19550 1486
rect 18272 1402 18288 1436
rect 18456 1402 18472 1436
rect 18530 1402 18546 1436
rect 18714 1402 18730 1436
rect 18788 1402 18804 1436
rect 18972 1402 18988 1436
rect 19046 1402 19062 1436
rect 19230 1402 19246 1436
rect 19304 1402 19320 1436
rect 19488 1402 19504 1436
rect 18272 1294 18288 1328
rect 18456 1294 18472 1328
rect 18530 1294 18546 1328
rect 18714 1294 18730 1328
rect 18788 1294 18804 1328
rect 18972 1294 18988 1328
rect 19046 1294 19062 1328
rect 19230 1294 19246 1328
rect 19304 1294 19320 1328
rect 19488 1294 19504 1328
rect 18226 1244 18260 1260
rect 18226 852 18260 868
rect 18484 1244 18518 1260
rect 18484 852 18518 868
rect 18742 1244 18776 1260
rect 18742 852 18776 868
rect 19000 1244 19034 1260
rect 19000 852 19034 868
rect 19258 1244 19292 1260
rect 19258 852 19292 868
rect 19516 1244 19550 1260
rect 19516 852 19550 868
rect 18272 784 18288 818
rect 18456 784 18472 818
rect 18530 784 18546 818
rect 18714 784 18730 818
rect 18788 784 18804 818
rect 18972 784 18988 818
rect 19046 784 19062 818
rect 19230 784 19246 818
rect 19304 784 19320 818
rect 19488 784 19504 818
rect 18272 676 18288 710
rect 18456 676 18472 710
rect 18530 676 18546 710
rect 18714 676 18730 710
rect 18788 676 18804 710
rect 18972 676 18988 710
rect 19046 676 19062 710
rect 19230 676 19246 710
rect 19304 676 19320 710
rect 19488 676 19504 710
rect 18226 626 18260 642
rect 18226 234 18260 250
rect 18484 626 18518 642
rect 18484 234 18518 250
rect 18742 626 18776 642
rect 18742 234 18776 250
rect 19000 626 19034 642
rect 19000 234 19034 250
rect 19258 626 19292 642
rect 19258 234 19292 250
rect 19516 626 19550 642
rect 19516 234 19550 250
rect 18272 166 18288 200
rect 18456 166 18472 200
rect 18530 166 18546 200
rect 18714 166 18730 200
rect 18788 166 18804 200
rect 18972 166 18988 200
rect 19046 166 19062 200
rect 19230 166 19246 200
rect 19304 166 19320 200
rect 19488 166 19504 200
rect 18092 98 18146 160
rect 19664 276 19912 3806
rect 19664 160 19688 276
rect 19630 98 19688 160
rect 18092 64 18208 98
rect 19568 64 19688 98
rect 19868 160 19912 276
rect 21430 3806 21464 3868
rect 20072 3766 20088 3800
rect 20256 3766 20272 3800
rect 20330 3766 20346 3800
rect 20514 3766 20530 3800
rect 20588 3766 20604 3800
rect 20772 3766 20788 3800
rect 20846 3766 20862 3800
rect 21030 3766 21046 3800
rect 21104 3766 21120 3800
rect 21288 3766 21304 3800
rect 20026 3716 20060 3732
rect 20026 3324 20060 3340
rect 20284 3716 20318 3732
rect 20284 3324 20318 3340
rect 20542 3716 20576 3732
rect 20542 3324 20576 3340
rect 20800 3716 20834 3732
rect 20800 3324 20834 3340
rect 21058 3716 21092 3732
rect 21058 3324 21092 3340
rect 21316 3716 21350 3732
rect 21316 3324 21350 3340
rect 20072 3256 20088 3290
rect 20256 3256 20272 3290
rect 20330 3256 20346 3290
rect 20514 3256 20530 3290
rect 20588 3256 20604 3290
rect 20772 3256 20788 3290
rect 20846 3256 20862 3290
rect 21030 3256 21046 3290
rect 21104 3256 21120 3290
rect 21288 3256 21304 3290
rect 20072 3148 20088 3182
rect 20256 3148 20272 3182
rect 20330 3148 20346 3182
rect 20514 3148 20530 3182
rect 20588 3148 20604 3182
rect 20772 3148 20788 3182
rect 20846 3148 20862 3182
rect 21030 3148 21046 3182
rect 21104 3148 21120 3182
rect 21288 3148 21304 3182
rect 20026 3098 20060 3114
rect 20026 2706 20060 2722
rect 20284 3098 20318 3114
rect 20284 2706 20318 2722
rect 20542 3098 20576 3114
rect 20542 2706 20576 2722
rect 20800 3098 20834 3114
rect 20800 2706 20834 2722
rect 21058 3098 21092 3114
rect 21058 2706 21092 2722
rect 21316 3098 21350 3114
rect 21316 2706 21350 2722
rect 20072 2638 20088 2672
rect 20256 2638 20272 2672
rect 20330 2638 20346 2672
rect 20514 2638 20530 2672
rect 20588 2638 20604 2672
rect 20772 2638 20788 2672
rect 20846 2638 20862 2672
rect 21030 2638 21046 2672
rect 21104 2638 21120 2672
rect 21288 2638 21304 2672
rect 20072 2530 20088 2564
rect 20256 2530 20272 2564
rect 20330 2530 20346 2564
rect 20514 2530 20530 2564
rect 20588 2530 20604 2564
rect 20772 2530 20788 2564
rect 20846 2530 20862 2564
rect 21030 2530 21046 2564
rect 21104 2530 21120 2564
rect 21288 2530 21304 2564
rect 20026 2480 20060 2496
rect 20026 2088 20060 2104
rect 20284 2480 20318 2496
rect 20284 2088 20318 2104
rect 20542 2480 20576 2496
rect 20542 2088 20576 2104
rect 20800 2480 20834 2496
rect 20800 2088 20834 2104
rect 21058 2480 21092 2496
rect 21058 2088 21092 2104
rect 21316 2480 21350 2496
rect 21316 2088 21350 2104
rect 20072 2020 20088 2054
rect 20256 2020 20272 2054
rect 20330 2020 20346 2054
rect 20514 2020 20530 2054
rect 20588 2020 20604 2054
rect 20772 2020 20788 2054
rect 20846 2020 20862 2054
rect 21030 2020 21046 2054
rect 21104 2020 21120 2054
rect 21288 2020 21304 2054
rect 20072 1912 20088 1946
rect 20256 1912 20272 1946
rect 20330 1912 20346 1946
rect 20514 1912 20530 1946
rect 20588 1912 20604 1946
rect 20772 1912 20788 1946
rect 20846 1912 20862 1946
rect 21030 1912 21046 1946
rect 21104 1912 21120 1946
rect 21288 1912 21304 1946
rect 20026 1862 20060 1878
rect 20026 1470 20060 1486
rect 20284 1862 20318 1878
rect 20284 1470 20318 1486
rect 20542 1862 20576 1878
rect 20542 1470 20576 1486
rect 20800 1862 20834 1878
rect 20800 1470 20834 1486
rect 21058 1862 21092 1878
rect 21058 1470 21092 1486
rect 21316 1862 21350 1878
rect 21316 1470 21350 1486
rect 20072 1402 20088 1436
rect 20256 1402 20272 1436
rect 20330 1402 20346 1436
rect 20514 1402 20530 1436
rect 20588 1402 20604 1436
rect 20772 1402 20788 1436
rect 20846 1402 20862 1436
rect 21030 1402 21046 1436
rect 21104 1402 21120 1436
rect 21288 1402 21304 1436
rect 20072 1294 20088 1328
rect 20256 1294 20272 1328
rect 20330 1294 20346 1328
rect 20514 1294 20530 1328
rect 20588 1294 20604 1328
rect 20772 1294 20788 1328
rect 20846 1294 20862 1328
rect 21030 1294 21046 1328
rect 21104 1294 21120 1328
rect 21288 1294 21304 1328
rect 20026 1244 20060 1260
rect 20026 852 20060 868
rect 20284 1244 20318 1260
rect 20284 852 20318 868
rect 20542 1244 20576 1260
rect 20542 852 20576 868
rect 20800 1244 20834 1260
rect 20800 852 20834 868
rect 21058 1244 21092 1260
rect 21058 852 21092 868
rect 21316 1244 21350 1260
rect 21316 852 21350 868
rect 20072 784 20088 818
rect 20256 784 20272 818
rect 20330 784 20346 818
rect 20514 784 20530 818
rect 20588 784 20604 818
rect 20772 784 20788 818
rect 20846 784 20862 818
rect 21030 784 21046 818
rect 21104 784 21120 818
rect 21288 784 21304 818
rect 20072 676 20088 710
rect 20256 676 20272 710
rect 20330 676 20346 710
rect 20514 676 20530 710
rect 20588 676 20604 710
rect 20772 676 20788 710
rect 20846 676 20862 710
rect 21030 676 21046 710
rect 21104 676 21120 710
rect 21288 676 21304 710
rect 20026 626 20060 642
rect 20026 234 20060 250
rect 20284 626 20318 642
rect 20284 234 20318 250
rect 20542 626 20576 642
rect 20542 234 20576 250
rect 20800 626 20834 642
rect 20800 234 20834 250
rect 21058 626 21092 642
rect 21058 234 21092 250
rect 21316 626 21350 642
rect 21316 234 21350 250
rect 20072 166 20088 200
rect 20256 166 20272 200
rect 20330 166 20346 200
rect 20514 166 20530 200
rect 20588 166 20604 200
rect 20772 166 20788 200
rect 20846 166 20862 200
rect 21030 166 21046 200
rect 21104 166 21120 200
rect 21288 166 21304 200
rect 19868 98 19946 160
rect 21430 98 21464 160
rect 19868 64 20008 98
rect 21368 64 21464 98
rect 3456 48 3736 64
rect 5252 40 5528 64
rect 17856 48 18136 64
rect 19652 40 19928 64
rect -2784 -1188 -2768 -382
rect -1960 -1188 -1944 -382
rect 11616 -1188 11632 -382
rect 12440 -1188 12456 -382
<< viali >>
rect 7440 27336 7540 27436
rect 6552 27134 6620 27168
rect 6710 27134 6778 27168
rect 6868 27134 6936 27168
rect 7026 27134 7094 27168
rect 7184 27134 7252 27168
rect 7342 27134 7410 27168
rect 7500 27134 7568 27168
rect 7658 27134 7726 27168
rect 7816 27134 7884 27168
rect 7974 27134 8042 27168
rect 6490 26699 6524 27075
rect 6648 26699 6682 27075
rect 6806 26699 6840 27075
rect 6964 26699 6998 27075
rect 7122 26699 7156 27075
rect 7280 26699 7314 27075
rect 7438 26699 7472 27075
rect 7596 26699 7630 27075
rect 7754 26699 7788 27075
rect 7912 26699 7946 27075
rect 8070 26699 8104 27075
rect 6552 26606 6620 26640
rect 6710 26606 6778 26640
rect 6868 26606 6936 26640
rect 7026 26606 7094 26640
rect 7184 26606 7252 26640
rect 7342 26606 7410 26640
rect 7500 26606 7568 26640
rect 7658 26606 7726 26640
rect 7816 26606 7884 26640
rect 7974 26606 8042 26640
rect 6552 26498 6620 26532
rect 6710 26498 6778 26532
rect 6868 26498 6936 26532
rect 7026 26498 7094 26532
rect 7184 26498 7252 26532
rect 7342 26498 7410 26532
rect 7500 26498 7568 26532
rect 7658 26498 7726 26532
rect 7816 26498 7884 26532
rect 7974 26498 8042 26532
rect 6490 26063 6524 26439
rect 6648 26063 6682 26439
rect 6806 26063 6840 26439
rect 6964 26063 6998 26439
rect 7122 26063 7156 26439
rect 7280 26063 7314 26439
rect 7438 26063 7472 26439
rect 7596 26063 7630 26439
rect 7754 26063 7788 26439
rect 7912 26063 7946 26439
rect 8070 26063 8104 26439
rect 6552 25970 6620 26004
rect 6710 25970 6778 26004
rect 6868 25970 6936 26004
rect 7026 25970 7094 26004
rect 7184 25970 7252 26004
rect 7342 25970 7410 26004
rect 7500 25970 7568 26004
rect 7658 25970 7726 26004
rect 7816 25970 7884 26004
rect 7974 25970 8042 26004
rect 6552 25862 6620 25896
rect 6710 25862 6778 25896
rect 6868 25862 6936 25896
rect 7026 25862 7094 25896
rect 7184 25862 7252 25896
rect 7342 25862 7410 25896
rect 7500 25862 7568 25896
rect 7658 25862 7726 25896
rect 7816 25862 7884 25896
rect 7974 25862 8042 25896
rect 6490 25427 6524 25803
rect 6648 25427 6682 25803
rect 6806 25427 6840 25803
rect 6964 25427 6998 25803
rect 7122 25427 7156 25803
rect 7280 25427 7314 25803
rect 7438 25427 7472 25803
rect 7596 25427 7630 25803
rect 7754 25427 7788 25803
rect 7912 25427 7946 25803
rect 8070 25427 8104 25803
rect 6552 25334 6620 25368
rect 6710 25334 6778 25368
rect 6868 25334 6936 25368
rect 7026 25334 7094 25368
rect 7184 25334 7252 25368
rect 7342 25334 7410 25368
rect 7500 25334 7568 25368
rect 7658 25334 7726 25368
rect 7816 25334 7884 25368
rect 7974 25334 8042 25368
rect 8772 27134 8840 27168
rect 8930 27134 8998 27168
rect 9088 27134 9156 27168
rect 9246 27134 9314 27168
rect 9404 27134 9472 27168
rect 9562 27134 9630 27168
rect 9720 27134 9788 27168
rect 9878 27134 9946 27168
rect 10036 27134 10104 27168
rect 10194 27134 10262 27168
rect 8710 26699 8744 27075
rect 8868 26699 8902 27075
rect 9026 26699 9060 27075
rect 9184 26699 9218 27075
rect 9342 26699 9376 27075
rect 9500 26699 9534 27075
rect 9658 26699 9692 27075
rect 9816 26699 9850 27075
rect 9974 26699 10008 27075
rect 10132 26699 10166 27075
rect 10290 26699 10324 27075
rect 8772 26606 8840 26640
rect 8930 26606 8998 26640
rect 9088 26606 9156 26640
rect 9246 26606 9314 26640
rect 9404 26606 9472 26640
rect 9562 26606 9630 26640
rect 9720 26606 9788 26640
rect 9878 26606 9946 26640
rect 10036 26606 10104 26640
rect 10194 26606 10262 26640
rect 8772 26498 8840 26532
rect 8930 26498 8998 26532
rect 9088 26498 9156 26532
rect 9246 26498 9314 26532
rect 9404 26498 9472 26532
rect 9562 26498 9630 26532
rect 9720 26498 9788 26532
rect 9878 26498 9946 26532
rect 10036 26498 10104 26532
rect 10194 26498 10262 26532
rect 8710 26063 8744 26439
rect 8868 26063 8902 26439
rect 9026 26063 9060 26439
rect 9184 26063 9218 26439
rect 9342 26063 9376 26439
rect 9500 26063 9534 26439
rect 9658 26063 9692 26439
rect 9816 26063 9850 26439
rect 9974 26063 10008 26439
rect 10132 26063 10166 26439
rect 10290 26063 10324 26439
rect 8772 25970 8840 26004
rect 8930 25970 8998 26004
rect 9088 25970 9156 26004
rect 9246 25970 9314 26004
rect 9404 25970 9472 26004
rect 9562 25970 9630 26004
rect 9720 25970 9788 26004
rect 9878 25970 9946 26004
rect 10036 25970 10104 26004
rect 10194 25970 10262 26004
rect 8772 25862 8840 25896
rect 8930 25862 8998 25896
rect 9088 25862 9156 25896
rect 9246 25862 9314 25896
rect 9404 25862 9472 25896
rect 9562 25862 9630 25896
rect 9720 25862 9788 25896
rect 9878 25862 9946 25896
rect 10036 25862 10104 25896
rect 10194 25862 10262 25896
rect 8710 25427 8744 25803
rect 8868 25427 8902 25803
rect 9026 25427 9060 25803
rect 9184 25427 9218 25803
rect 9342 25427 9376 25803
rect 9500 25427 9534 25803
rect 9658 25427 9692 25803
rect 9816 25427 9850 25803
rect 9974 25427 10008 25803
rect 10132 25427 10166 25803
rect 10290 25427 10324 25803
rect 8772 25334 8840 25368
rect 8930 25334 8998 25368
rect 9088 25334 9156 25368
rect 9246 25334 9314 25368
rect 9404 25334 9472 25368
rect 9562 25334 9630 25368
rect 9720 25334 9788 25368
rect 9878 25334 9946 25368
rect 10036 25334 10104 25368
rect 10194 25334 10262 25368
rect 10952 27134 11020 27168
rect 11110 27134 11178 27168
rect 11268 27134 11336 27168
rect 11426 27134 11494 27168
rect 11584 27134 11652 27168
rect 11742 27134 11810 27168
rect 11900 27134 11968 27168
rect 12058 27134 12126 27168
rect 12216 27134 12284 27168
rect 12374 27134 12442 27168
rect 10890 26699 10924 27075
rect 11048 26699 11082 27075
rect 11206 26699 11240 27075
rect 11364 26699 11398 27075
rect 11522 26699 11556 27075
rect 11680 26699 11714 27075
rect 11838 26699 11872 27075
rect 11996 26699 12030 27075
rect 12154 26699 12188 27075
rect 12312 26699 12346 27075
rect 12470 26699 12504 27075
rect 10952 26606 11020 26640
rect 11110 26606 11178 26640
rect 11268 26606 11336 26640
rect 11426 26606 11494 26640
rect 11584 26606 11652 26640
rect 11742 26606 11810 26640
rect 11900 26606 11968 26640
rect 12058 26606 12126 26640
rect 12216 26606 12284 26640
rect 12374 26606 12442 26640
rect 10952 26498 11020 26532
rect 11110 26498 11178 26532
rect 11268 26498 11336 26532
rect 11426 26498 11494 26532
rect 11584 26498 11652 26532
rect 11742 26498 11810 26532
rect 11900 26498 11968 26532
rect 12058 26498 12126 26532
rect 12216 26498 12284 26532
rect 12374 26498 12442 26532
rect 10890 26063 10924 26439
rect 11048 26063 11082 26439
rect 11206 26063 11240 26439
rect 11364 26063 11398 26439
rect 11522 26063 11556 26439
rect 11680 26063 11714 26439
rect 11838 26063 11872 26439
rect 11996 26063 12030 26439
rect 12154 26063 12188 26439
rect 12312 26063 12346 26439
rect 12470 26063 12504 26439
rect 10952 25970 11020 26004
rect 11110 25970 11178 26004
rect 11268 25970 11336 26004
rect 11426 25970 11494 26004
rect 11584 25970 11652 26004
rect 11742 25970 11810 26004
rect 11900 25970 11968 26004
rect 12058 25970 12126 26004
rect 12216 25970 12284 26004
rect 12374 25970 12442 26004
rect 10952 25862 11020 25896
rect 11110 25862 11178 25896
rect 11268 25862 11336 25896
rect 11426 25862 11494 25896
rect 11584 25862 11652 25896
rect 11742 25862 11810 25896
rect 11900 25862 11968 25896
rect 12058 25862 12126 25896
rect 12216 25862 12284 25896
rect 12374 25862 12442 25896
rect 10890 25427 10924 25803
rect 11048 25427 11082 25803
rect 11206 25427 11240 25803
rect 11364 25427 11398 25803
rect 11522 25427 11556 25803
rect 11680 25427 11714 25803
rect 11838 25427 11872 25803
rect 11996 25427 12030 25803
rect 12154 25427 12188 25803
rect 12312 25427 12346 25803
rect 12470 25427 12504 25803
rect 10952 25334 11020 25368
rect 11110 25334 11178 25368
rect 11268 25334 11336 25368
rect 11426 25334 11494 25368
rect 11584 25334 11652 25368
rect 11742 25334 11810 25368
rect 11900 25334 11968 25368
rect 12058 25334 12126 25368
rect 12216 25334 12284 25368
rect 12374 25334 12442 25368
rect 13132 27134 13200 27168
rect 13290 27134 13358 27168
rect 13448 27134 13516 27168
rect 13606 27134 13674 27168
rect 13764 27134 13832 27168
rect 13922 27134 13990 27168
rect 14080 27134 14148 27168
rect 14238 27134 14306 27168
rect 14396 27134 14464 27168
rect 14554 27134 14622 27168
rect 13070 26699 13104 27075
rect 13228 26699 13262 27075
rect 13386 26699 13420 27075
rect 13544 26699 13578 27075
rect 13702 26699 13736 27075
rect 13860 26699 13894 27075
rect 14018 26699 14052 27075
rect 14176 26699 14210 27075
rect 14334 26699 14368 27075
rect 14492 26699 14526 27075
rect 14650 26699 14684 27075
rect 13132 26606 13200 26640
rect 13290 26606 13358 26640
rect 13448 26606 13516 26640
rect 13606 26606 13674 26640
rect 13764 26606 13832 26640
rect 13922 26606 13990 26640
rect 14080 26606 14148 26640
rect 14238 26606 14306 26640
rect 14396 26606 14464 26640
rect 14554 26606 14622 26640
rect 13132 26498 13200 26532
rect 13290 26498 13358 26532
rect 13448 26498 13516 26532
rect 13606 26498 13674 26532
rect 13764 26498 13832 26532
rect 13922 26498 13990 26532
rect 14080 26498 14148 26532
rect 14238 26498 14306 26532
rect 14396 26498 14464 26532
rect 14554 26498 14622 26532
rect 13070 26063 13104 26439
rect 13228 26063 13262 26439
rect 13386 26063 13420 26439
rect 13544 26063 13578 26439
rect 13702 26063 13736 26439
rect 13860 26063 13894 26439
rect 14018 26063 14052 26439
rect 14176 26063 14210 26439
rect 14334 26063 14368 26439
rect 14492 26063 14526 26439
rect 14650 26063 14684 26439
rect 13132 25970 13200 26004
rect 13290 25970 13358 26004
rect 13448 25970 13516 26004
rect 13606 25970 13674 26004
rect 13764 25970 13832 26004
rect 13922 25970 13990 26004
rect 14080 25970 14148 26004
rect 14238 25970 14306 26004
rect 14396 25970 14464 26004
rect 14554 25970 14622 26004
rect 13132 25862 13200 25896
rect 13290 25862 13358 25896
rect 13448 25862 13516 25896
rect 13606 25862 13674 25896
rect 13764 25862 13832 25896
rect 13922 25862 13990 25896
rect 14080 25862 14148 25896
rect 14238 25862 14306 25896
rect 14396 25862 14464 25896
rect 14554 25862 14622 25896
rect 13070 25427 13104 25803
rect 13228 25427 13262 25803
rect 13386 25427 13420 25803
rect 13544 25427 13578 25803
rect 13702 25427 13736 25803
rect 13860 25427 13894 25803
rect 14018 25427 14052 25803
rect 14176 25427 14210 25803
rect 14334 25427 14368 25803
rect 14492 25427 14526 25803
rect 14650 25427 14684 25803
rect 13132 25334 13200 25368
rect 13290 25334 13358 25368
rect 13448 25334 13516 25368
rect 13606 25334 13674 25368
rect 13764 25334 13832 25368
rect 13922 25334 13990 25368
rect 14080 25334 14148 25368
rect 14238 25334 14306 25368
rect 14396 25334 14464 25368
rect 14554 25334 14622 25368
rect 15332 27134 15400 27168
rect 15490 27134 15558 27168
rect 15648 27134 15716 27168
rect 15806 27134 15874 27168
rect 15964 27134 16032 27168
rect 16122 27134 16190 27168
rect 16280 27134 16348 27168
rect 16438 27134 16506 27168
rect 16596 27134 16664 27168
rect 16754 27134 16822 27168
rect 15270 26699 15304 27075
rect 15428 26699 15462 27075
rect 15586 26699 15620 27075
rect 15744 26699 15778 27075
rect 15902 26699 15936 27075
rect 16060 26699 16094 27075
rect 16218 26699 16252 27075
rect 16376 26699 16410 27075
rect 16534 26699 16568 27075
rect 16692 26699 16726 27075
rect 16850 26699 16884 27075
rect 15332 26606 15400 26640
rect 15490 26606 15558 26640
rect 15648 26606 15716 26640
rect 15806 26606 15874 26640
rect 15964 26606 16032 26640
rect 16122 26606 16190 26640
rect 16280 26606 16348 26640
rect 16438 26606 16506 26640
rect 16596 26606 16664 26640
rect 16754 26606 16822 26640
rect 15332 26498 15400 26532
rect 15490 26498 15558 26532
rect 15648 26498 15716 26532
rect 15806 26498 15874 26532
rect 15964 26498 16032 26532
rect 16122 26498 16190 26532
rect 16280 26498 16348 26532
rect 16438 26498 16506 26532
rect 16596 26498 16664 26532
rect 16754 26498 16822 26532
rect 15270 26063 15304 26439
rect 15428 26063 15462 26439
rect 15586 26063 15620 26439
rect 15744 26063 15778 26439
rect 15902 26063 15936 26439
rect 16060 26063 16094 26439
rect 16218 26063 16252 26439
rect 16376 26063 16410 26439
rect 16534 26063 16568 26439
rect 16692 26063 16726 26439
rect 16850 26063 16884 26439
rect 15332 25970 15400 26004
rect 15490 25970 15558 26004
rect 15648 25970 15716 26004
rect 15806 25970 15874 26004
rect 15964 25970 16032 26004
rect 16122 25970 16190 26004
rect 16280 25970 16348 26004
rect 16438 25970 16506 26004
rect 16596 25970 16664 26004
rect 16754 25970 16822 26004
rect 15332 25862 15400 25896
rect 15490 25862 15558 25896
rect 15648 25862 15716 25896
rect 15806 25862 15874 25896
rect 15964 25862 16032 25896
rect 16122 25862 16190 25896
rect 16280 25862 16348 25896
rect 16438 25862 16506 25896
rect 16596 25862 16664 25896
rect 16754 25862 16822 25896
rect 15270 25427 15304 25803
rect 15428 25427 15462 25803
rect 15586 25427 15620 25803
rect 15744 25427 15778 25803
rect 15902 25427 15936 25803
rect 16060 25427 16094 25803
rect 16218 25427 16252 25803
rect 16376 25427 16410 25803
rect 16534 25427 16568 25803
rect 16692 25427 16726 25803
rect 16850 25427 16884 25803
rect 15332 25334 15400 25368
rect 15490 25334 15558 25368
rect 15648 25334 15716 25368
rect 15806 25334 15874 25368
rect 15964 25334 16032 25368
rect 16122 25334 16190 25368
rect 16280 25334 16348 25368
rect 16438 25334 16506 25368
rect 16596 25334 16664 25368
rect 16754 25334 16822 25368
rect 19060 25296 19220 25436
rect 6538 25038 6572 25072
rect 6730 25038 6764 25072
rect 6922 25038 6956 25072
rect 7114 25038 7148 25072
rect 7306 25038 7340 25072
rect 7498 25038 7532 25072
rect 7690 25038 7724 25072
rect 7882 25038 7916 25072
rect 6490 24603 6524 24979
rect 6586 24603 6620 24979
rect 6682 24603 6716 24979
rect 6778 24603 6812 24979
rect 6874 24603 6908 24979
rect 6970 24603 7004 24979
rect 7066 24603 7100 24979
rect 7162 24603 7196 24979
rect 7258 24603 7292 24979
rect 7354 24603 7388 24979
rect 7450 24603 7484 24979
rect 7546 24603 7580 24979
rect 7642 24603 7676 24979
rect 7738 24603 7772 24979
rect 7834 24603 7868 24979
rect 7930 24603 7964 24979
rect 6634 24510 6668 24544
rect 6826 24510 6860 24544
rect 7018 24510 7052 24544
rect 7210 24510 7244 24544
rect 7402 24510 7436 24544
rect 7594 24510 7628 24544
rect 7786 24510 7820 24544
rect 6634 24402 6668 24436
rect 6826 24402 6860 24436
rect 7018 24402 7052 24436
rect 7210 24402 7244 24436
rect 7402 24402 7436 24436
rect 7594 24402 7628 24436
rect 7786 24402 7820 24436
rect 6490 23967 6524 24343
rect 6586 23967 6620 24343
rect 6682 23967 6716 24343
rect 6778 23967 6812 24343
rect 6874 23967 6908 24343
rect 6970 23967 7004 24343
rect 7066 23967 7100 24343
rect 7162 23967 7196 24343
rect 7258 23967 7292 24343
rect 7354 23967 7388 24343
rect 7450 23967 7484 24343
rect 7546 23967 7580 24343
rect 7642 23967 7676 24343
rect 7738 23967 7772 24343
rect 7834 23967 7868 24343
rect 7930 23967 7964 24343
rect 6538 23874 6572 23908
rect 6730 23874 6764 23908
rect 6922 23874 6956 23908
rect 7114 23874 7148 23908
rect 7306 23874 7340 23908
rect 7498 23874 7532 23908
rect 7690 23874 7724 23908
rect 7882 23874 7916 23908
rect 8758 25038 8792 25072
rect 8950 25038 8984 25072
rect 9142 25038 9176 25072
rect 9334 25038 9368 25072
rect 9526 25038 9560 25072
rect 9718 25038 9752 25072
rect 9910 25038 9944 25072
rect 10102 25038 10136 25072
rect 8710 24603 8744 24979
rect 8806 24603 8840 24979
rect 8902 24603 8936 24979
rect 8998 24603 9032 24979
rect 9094 24603 9128 24979
rect 9190 24603 9224 24979
rect 9286 24603 9320 24979
rect 9382 24603 9416 24979
rect 9478 24603 9512 24979
rect 9574 24603 9608 24979
rect 9670 24603 9704 24979
rect 9766 24603 9800 24979
rect 9862 24603 9896 24979
rect 9958 24603 9992 24979
rect 10054 24603 10088 24979
rect 10150 24603 10184 24979
rect 8854 24510 8888 24544
rect 9046 24510 9080 24544
rect 9238 24510 9272 24544
rect 9430 24510 9464 24544
rect 9622 24510 9656 24544
rect 9814 24510 9848 24544
rect 10006 24510 10040 24544
rect 8854 24402 8888 24436
rect 9046 24402 9080 24436
rect 9238 24402 9272 24436
rect 9430 24402 9464 24436
rect 9622 24402 9656 24436
rect 9814 24402 9848 24436
rect 10006 24402 10040 24436
rect 8710 23967 8744 24343
rect 8806 23967 8840 24343
rect 8902 23967 8936 24343
rect 8998 23967 9032 24343
rect 9094 23967 9128 24343
rect 9190 23967 9224 24343
rect 9286 23967 9320 24343
rect 9382 23967 9416 24343
rect 9478 23967 9512 24343
rect 9574 23967 9608 24343
rect 9670 23967 9704 24343
rect 9766 23967 9800 24343
rect 9862 23967 9896 24343
rect 9958 23967 9992 24343
rect 10054 23967 10088 24343
rect 10150 23967 10184 24343
rect 8758 23874 8792 23908
rect 8950 23874 8984 23908
rect 9142 23874 9176 23908
rect 9334 23874 9368 23908
rect 9526 23874 9560 23908
rect 9718 23874 9752 23908
rect 9910 23874 9944 23908
rect 10102 23874 10136 23908
rect 10938 25038 10972 25072
rect 11130 25038 11164 25072
rect 11322 25038 11356 25072
rect 11514 25038 11548 25072
rect 11706 25038 11740 25072
rect 11898 25038 11932 25072
rect 12090 25038 12124 25072
rect 12282 25038 12316 25072
rect 10890 24603 10924 24979
rect 10986 24603 11020 24979
rect 11082 24603 11116 24979
rect 11178 24603 11212 24979
rect 11274 24603 11308 24979
rect 11370 24603 11404 24979
rect 11466 24603 11500 24979
rect 11562 24603 11596 24979
rect 11658 24603 11692 24979
rect 11754 24603 11788 24979
rect 11850 24603 11884 24979
rect 11946 24603 11980 24979
rect 12042 24603 12076 24979
rect 12138 24603 12172 24979
rect 12234 24603 12268 24979
rect 12330 24603 12364 24979
rect 11034 24510 11068 24544
rect 11226 24510 11260 24544
rect 11418 24510 11452 24544
rect 11610 24510 11644 24544
rect 11802 24510 11836 24544
rect 11994 24510 12028 24544
rect 12186 24510 12220 24544
rect 11034 24402 11068 24436
rect 11226 24402 11260 24436
rect 11418 24402 11452 24436
rect 11610 24402 11644 24436
rect 11802 24402 11836 24436
rect 11994 24402 12028 24436
rect 12186 24402 12220 24436
rect 10890 23967 10924 24343
rect 10986 23967 11020 24343
rect 11082 23967 11116 24343
rect 11178 23967 11212 24343
rect 11274 23967 11308 24343
rect 11370 23967 11404 24343
rect 11466 23967 11500 24343
rect 11562 23967 11596 24343
rect 11658 23967 11692 24343
rect 11754 23967 11788 24343
rect 11850 23967 11884 24343
rect 11946 23967 11980 24343
rect 12042 23967 12076 24343
rect 12138 23967 12172 24343
rect 12234 23967 12268 24343
rect 12330 23967 12364 24343
rect 10938 23874 10972 23908
rect 11130 23874 11164 23908
rect 11322 23874 11356 23908
rect 11514 23874 11548 23908
rect 11706 23874 11740 23908
rect 11898 23874 11932 23908
rect 12090 23874 12124 23908
rect 12282 23874 12316 23908
rect 13118 25038 13152 25072
rect 13310 25038 13344 25072
rect 13502 25038 13536 25072
rect 13694 25038 13728 25072
rect 13886 25038 13920 25072
rect 14078 25038 14112 25072
rect 14270 25038 14304 25072
rect 14462 25038 14496 25072
rect 13070 24603 13104 24979
rect 13166 24603 13200 24979
rect 13262 24603 13296 24979
rect 13358 24603 13392 24979
rect 13454 24603 13488 24979
rect 13550 24603 13584 24979
rect 13646 24603 13680 24979
rect 13742 24603 13776 24979
rect 13838 24603 13872 24979
rect 13934 24603 13968 24979
rect 14030 24603 14064 24979
rect 14126 24603 14160 24979
rect 14222 24603 14256 24979
rect 14318 24603 14352 24979
rect 14414 24603 14448 24979
rect 14510 24603 14544 24979
rect 13214 24510 13248 24544
rect 13406 24510 13440 24544
rect 13598 24510 13632 24544
rect 13790 24510 13824 24544
rect 13982 24510 14016 24544
rect 14174 24510 14208 24544
rect 14366 24510 14400 24544
rect 13214 24402 13248 24436
rect 13406 24402 13440 24436
rect 13598 24402 13632 24436
rect 13790 24402 13824 24436
rect 13982 24402 14016 24436
rect 14174 24402 14208 24436
rect 14366 24402 14400 24436
rect 13070 23967 13104 24343
rect 13166 23967 13200 24343
rect 13262 23967 13296 24343
rect 13358 23967 13392 24343
rect 13454 23967 13488 24343
rect 13550 23967 13584 24343
rect 13646 23967 13680 24343
rect 13742 23967 13776 24343
rect 13838 23967 13872 24343
rect 13934 23967 13968 24343
rect 14030 23967 14064 24343
rect 14126 23967 14160 24343
rect 14222 23967 14256 24343
rect 14318 23967 14352 24343
rect 14414 23967 14448 24343
rect 14510 23967 14544 24343
rect 13118 23874 13152 23908
rect 13310 23874 13344 23908
rect 13502 23874 13536 23908
rect 13694 23874 13728 23908
rect 13886 23874 13920 23908
rect 14078 23874 14112 23908
rect 14270 23874 14304 23908
rect 14462 23874 14496 23908
rect 15318 25038 15352 25072
rect 15510 25038 15544 25072
rect 15702 25038 15736 25072
rect 15894 25038 15928 25072
rect 16086 25038 16120 25072
rect 16278 25038 16312 25072
rect 16470 25038 16504 25072
rect 16662 25038 16696 25072
rect 15270 24603 15304 24979
rect 15366 24603 15400 24979
rect 15462 24603 15496 24979
rect 15558 24603 15592 24979
rect 15654 24603 15688 24979
rect 15750 24603 15784 24979
rect 15846 24603 15880 24979
rect 15942 24603 15976 24979
rect 16038 24603 16072 24979
rect 16134 24603 16168 24979
rect 16230 24603 16264 24979
rect 16326 24603 16360 24979
rect 16422 24603 16456 24979
rect 16518 24603 16552 24979
rect 16614 24603 16648 24979
rect 16710 24603 16744 24979
rect 15414 24510 15448 24544
rect 15606 24510 15640 24544
rect 15798 24510 15832 24544
rect 15990 24510 16024 24544
rect 16182 24510 16216 24544
rect 16374 24510 16408 24544
rect 16566 24510 16600 24544
rect 15414 24402 15448 24436
rect 15606 24402 15640 24436
rect 15798 24402 15832 24436
rect 15990 24402 16024 24436
rect 16182 24402 16216 24436
rect 16374 24402 16408 24436
rect 16566 24402 16600 24436
rect 15270 23967 15304 24343
rect 15366 23967 15400 24343
rect 15462 23967 15496 24343
rect 15558 23967 15592 24343
rect 15654 23967 15688 24343
rect 15750 23967 15784 24343
rect 15846 23967 15880 24343
rect 15942 23967 15976 24343
rect 16038 23967 16072 24343
rect 16134 23967 16168 24343
rect 16230 23967 16264 24343
rect 16326 23967 16360 24343
rect 16422 23967 16456 24343
rect 16518 23967 16552 24343
rect 16614 23967 16648 24343
rect 16710 23967 16744 24343
rect 15318 23874 15352 23908
rect 15510 23874 15544 23908
rect 15702 23874 15736 23908
rect 15894 23874 15928 23908
rect 16086 23874 16120 23908
rect 16278 23874 16312 23908
rect 16470 23874 16504 23908
rect 16662 23874 16696 23908
rect 6754 23460 6788 23494
rect 6946 23460 6980 23494
rect 7138 23460 7172 23494
rect 7330 23460 7364 23494
rect 7522 23460 7556 23494
rect 6610 23034 6644 23410
rect 6706 23034 6740 23410
rect 6802 23034 6836 23410
rect 6898 23034 6932 23410
rect 6994 23034 7028 23410
rect 7090 23034 7124 23410
rect 7186 23034 7220 23410
rect 7282 23034 7316 23410
rect 7378 23034 7412 23410
rect 7474 23034 7508 23410
rect 7570 23034 7604 23410
rect 6658 22950 6692 22984
rect 6850 22950 6884 22984
rect 7042 22950 7076 22984
rect 7234 22950 7268 22984
rect 7426 22950 7460 22984
rect 6658 22842 6692 22876
rect 6850 22842 6884 22876
rect 7042 22842 7076 22876
rect 7234 22842 7268 22876
rect 7426 22842 7460 22876
rect 6610 22416 6644 22792
rect 6706 22416 6740 22792
rect 6802 22416 6836 22792
rect 6898 22416 6932 22792
rect 6994 22416 7028 22792
rect 7090 22416 7124 22792
rect 7186 22416 7220 22792
rect 7282 22416 7316 22792
rect 7378 22416 7412 22792
rect 7474 22416 7508 22792
rect 7570 22416 7604 22792
rect 6754 22332 6788 22366
rect 6946 22332 6980 22366
rect 7138 22332 7172 22366
rect 7330 22332 7364 22366
rect 7522 22332 7556 22366
rect 6754 22224 6788 22258
rect 6946 22224 6980 22258
rect 7138 22224 7172 22258
rect 7330 22224 7364 22258
rect 7522 22224 7556 22258
rect 6610 21798 6644 22174
rect 6706 21798 6740 22174
rect 6802 21798 6836 22174
rect 6898 21798 6932 22174
rect 6994 21798 7028 22174
rect 7090 21798 7124 22174
rect 7186 21798 7220 22174
rect 7282 21798 7316 22174
rect 7378 21798 7412 22174
rect 7474 21798 7508 22174
rect 7570 21798 7604 22174
rect 6658 21714 6692 21748
rect 6850 21714 6884 21748
rect 7042 21714 7076 21748
rect 7234 21714 7268 21748
rect 7426 21714 7460 21748
rect 8474 23460 8508 23494
rect 8666 23460 8700 23494
rect 8858 23460 8892 23494
rect 9050 23460 9084 23494
rect 9242 23460 9276 23494
rect 8330 23034 8364 23410
rect 8426 23034 8460 23410
rect 8522 23034 8556 23410
rect 8618 23034 8652 23410
rect 8714 23034 8748 23410
rect 8810 23034 8844 23410
rect 8906 23034 8940 23410
rect 9002 23034 9036 23410
rect 9098 23034 9132 23410
rect 9194 23034 9228 23410
rect 9290 23034 9324 23410
rect 8378 22950 8412 22984
rect 8570 22950 8604 22984
rect 8762 22950 8796 22984
rect 8954 22950 8988 22984
rect 9146 22950 9180 22984
rect 8378 22842 8412 22876
rect 8570 22842 8604 22876
rect 8762 22842 8796 22876
rect 8954 22842 8988 22876
rect 9146 22842 9180 22876
rect 8330 22416 8364 22792
rect 8426 22416 8460 22792
rect 8522 22416 8556 22792
rect 8618 22416 8652 22792
rect 8714 22416 8748 22792
rect 8810 22416 8844 22792
rect 8906 22416 8940 22792
rect 9002 22416 9036 22792
rect 9098 22416 9132 22792
rect 9194 22416 9228 22792
rect 9290 22416 9324 22792
rect 8474 22332 8508 22366
rect 8666 22332 8700 22366
rect 8858 22332 8892 22366
rect 9050 22332 9084 22366
rect 9242 22332 9276 22366
rect 8474 22224 8508 22258
rect 8666 22224 8700 22258
rect 8858 22224 8892 22258
rect 9050 22224 9084 22258
rect 9242 22224 9276 22258
rect 8330 21798 8364 22174
rect 8426 21798 8460 22174
rect 8522 21798 8556 22174
rect 8618 21798 8652 22174
rect 8714 21798 8748 22174
rect 8810 21798 8844 22174
rect 8906 21798 8940 22174
rect 9002 21798 9036 22174
rect 9098 21798 9132 22174
rect 9194 21798 9228 22174
rect 9290 21798 9324 22174
rect 8378 21714 8412 21748
rect 8570 21714 8604 21748
rect 8762 21714 8796 21748
rect 8954 21714 8988 21748
rect 9146 21714 9180 21748
rect 18342 24671 18592 25068
rect 18342 23440 18592 23837
rect 19051 25048 19227 25082
rect 18958 23452 18992 25020
rect 19286 23452 19320 25020
rect 19051 23390 19227 23424
rect 18454 23070 18488 23104
rect 18646 23070 18680 23104
rect 18838 23070 18872 23104
rect 19030 23070 19064 23104
rect 19222 23070 19256 23104
rect 18310 22635 18344 23011
rect 18406 22635 18440 23011
rect 18502 22635 18536 23011
rect 18598 22635 18632 23011
rect 18694 22635 18728 23011
rect 18790 22635 18824 23011
rect 18886 22635 18920 23011
rect 18982 22635 19016 23011
rect 19078 22635 19112 23011
rect 19174 22635 19208 23011
rect 19270 22635 19304 23011
rect 18358 22542 18392 22576
rect 18550 22542 18584 22576
rect 18742 22542 18776 22576
rect 18934 22542 18968 22576
rect 19126 22542 19160 22576
rect 6672 21314 6840 21348
rect 6930 21314 7098 21348
rect 7188 21314 7356 21348
rect 7446 21314 7614 21348
rect 7704 21314 7872 21348
rect 6610 20888 6644 21264
rect 6868 20888 6902 21264
rect 7126 20888 7160 21264
rect 7384 20888 7418 21264
rect 7642 20888 7676 21264
rect 7900 20888 7934 21264
rect 6672 20804 6840 20838
rect 6930 20804 7098 20838
rect 7188 20804 7356 20838
rect 7446 20804 7614 20838
rect 7704 20804 7872 20838
rect 6672 20696 6840 20730
rect 6930 20696 7098 20730
rect 7188 20696 7356 20730
rect 7446 20696 7614 20730
rect 7704 20696 7872 20730
rect 6610 20270 6644 20646
rect 6868 20270 6902 20646
rect 7126 20270 7160 20646
rect 7384 20270 7418 20646
rect 7642 20270 7676 20646
rect 7900 20270 7934 20646
rect 6672 20186 6840 20220
rect 6930 20186 7098 20220
rect 7188 20186 7356 20220
rect 7446 20186 7614 20220
rect 7704 20186 7872 20220
rect 6672 20078 6840 20112
rect 6930 20078 7098 20112
rect 7188 20078 7356 20112
rect 7446 20078 7614 20112
rect 7704 20078 7872 20112
rect 6610 19652 6644 20028
rect 6868 19652 6902 20028
rect 7126 19652 7160 20028
rect 7384 19652 7418 20028
rect 7642 19652 7676 20028
rect 7900 19652 7934 20028
rect 6672 19568 6840 19602
rect 6930 19568 7098 19602
rect 7188 19568 7356 19602
rect 7446 19568 7614 19602
rect 7704 19568 7872 19602
rect 6672 19460 6840 19494
rect 6930 19460 7098 19494
rect 7188 19460 7356 19494
rect 7446 19460 7614 19494
rect 7704 19460 7872 19494
rect 6610 19034 6644 19410
rect 6868 19034 6902 19410
rect 7126 19034 7160 19410
rect 7384 19034 7418 19410
rect 7642 19034 7676 19410
rect 7900 19034 7934 19410
rect 6672 18950 6840 18984
rect 6930 18950 7098 18984
rect 7188 18950 7356 18984
rect 7446 18950 7614 18984
rect 7704 18950 7872 18984
rect 6672 18842 6840 18876
rect 6930 18842 7098 18876
rect 7188 18842 7356 18876
rect 7446 18842 7614 18876
rect 7704 18842 7872 18876
rect 6610 18416 6644 18792
rect 6868 18416 6902 18792
rect 7126 18416 7160 18792
rect 7384 18416 7418 18792
rect 7642 18416 7676 18792
rect 7900 18416 7934 18792
rect 6672 18332 6840 18366
rect 6930 18332 7098 18366
rect 7188 18332 7356 18366
rect 7446 18332 7614 18366
rect 7704 18332 7872 18366
rect 6672 18224 6840 18258
rect 6930 18224 7098 18258
rect 7188 18224 7356 18258
rect 7446 18224 7614 18258
rect 7704 18224 7872 18258
rect 6610 17798 6644 18174
rect 6868 17798 6902 18174
rect 7126 17798 7160 18174
rect 7384 17798 7418 18174
rect 7642 17798 7676 18174
rect 7900 17798 7934 18174
rect 8392 21314 8560 21348
rect 8650 21314 8818 21348
rect 8908 21314 9076 21348
rect 9166 21314 9334 21348
rect 9424 21314 9592 21348
rect 8330 20888 8364 21264
rect 8588 20888 8622 21264
rect 8846 20888 8880 21264
rect 9104 20888 9138 21264
rect 9362 20888 9396 21264
rect 9620 20888 9654 21264
rect 8392 20804 8560 20838
rect 8650 20804 8818 20838
rect 8908 20804 9076 20838
rect 9166 20804 9334 20838
rect 9424 20804 9592 20838
rect 8392 20696 8560 20730
rect 8650 20696 8818 20730
rect 8908 20696 9076 20730
rect 9166 20696 9334 20730
rect 9424 20696 9592 20730
rect 8330 20270 8364 20646
rect 8588 20270 8622 20646
rect 8846 20270 8880 20646
rect 9104 20270 9138 20646
rect 9362 20270 9396 20646
rect 9620 20270 9654 20646
rect 8392 20186 8560 20220
rect 8650 20186 8818 20220
rect 8908 20186 9076 20220
rect 9166 20186 9334 20220
rect 9424 20186 9592 20220
rect 8392 20078 8560 20112
rect 8650 20078 8818 20112
rect 8908 20078 9076 20112
rect 9166 20078 9334 20112
rect 9424 20078 9592 20112
rect 8330 19652 8364 20028
rect 8588 19652 8622 20028
rect 8846 19652 8880 20028
rect 9104 19652 9138 20028
rect 9362 19652 9396 20028
rect 9620 19652 9654 20028
rect 8392 19568 8560 19602
rect 8650 19568 8818 19602
rect 8908 19568 9076 19602
rect 9166 19568 9334 19602
rect 9424 19568 9592 19602
rect 8392 19460 8560 19494
rect 8650 19460 8818 19494
rect 8908 19460 9076 19494
rect 9166 19460 9334 19494
rect 9424 19460 9592 19494
rect 8330 19034 8364 19410
rect 8588 19034 8622 19410
rect 8846 19034 8880 19410
rect 9104 19034 9138 19410
rect 9362 19034 9396 19410
rect 9620 19034 9654 19410
rect 8392 18950 8560 18984
rect 8650 18950 8818 18984
rect 8908 18950 9076 18984
rect 9166 18950 9334 18984
rect 9424 18950 9592 18984
rect 8392 18842 8560 18876
rect 8650 18842 8818 18876
rect 8908 18842 9076 18876
rect 9166 18842 9334 18876
rect 9424 18842 9592 18876
rect 8330 18416 8364 18792
rect 8588 18416 8622 18792
rect 8846 18416 8880 18792
rect 9104 18416 9138 18792
rect 9362 18416 9396 18792
rect 9620 18416 9654 18792
rect 8392 18332 8560 18366
rect 8650 18332 8818 18366
rect 8908 18332 9076 18366
rect 9166 18332 9334 18366
rect 9424 18332 9592 18366
rect 8392 18224 8560 18258
rect 8650 18224 8818 18258
rect 8908 18224 9076 18258
rect 9166 18224 9334 18258
rect 9424 18224 9592 18258
rect 8330 17798 8364 18174
rect 8588 17798 8622 18174
rect 8846 17798 8880 18174
rect 9104 17798 9138 18174
rect 9362 17798 9396 18174
rect 9620 17798 9654 18174
rect 6672 17714 6840 17748
rect 6930 17714 7098 17748
rect 7188 17714 7356 17748
rect 7446 17714 7614 17748
rect 7704 17714 7872 17748
rect 8040 17708 8048 17776
rect 8048 17708 8216 17776
rect 8216 17708 8220 17776
rect 8392 17714 8560 17748
rect 8650 17714 8818 17748
rect 8908 17714 9076 17748
rect 9166 17714 9334 17748
rect 9424 17714 9592 17748
rect 8040 17616 8220 17708
rect 18454 22202 18488 22236
rect 18646 22202 18680 22236
rect 18838 22202 18872 22236
rect 19030 22202 19064 22236
rect 19222 22202 19256 22236
rect 18310 21776 18344 22152
rect 18406 21776 18440 22152
rect 18502 21776 18536 22152
rect 18598 21776 18632 22152
rect 18694 21776 18728 22152
rect 18790 21776 18824 22152
rect 18886 21776 18920 22152
rect 18982 21776 19016 22152
rect 19078 21776 19112 22152
rect 19174 21776 19208 22152
rect 19270 21776 19304 22152
rect 18358 21692 18392 21726
rect 18550 21692 18584 21726
rect 18742 21692 18776 21726
rect 18934 21692 18968 21726
rect 19126 21692 19160 21726
rect 18358 21584 18392 21618
rect 18550 21584 18584 21618
rect 18742 21584 18776 21618
rect 18934 21584 18968 21618
rect 19126 21584 19160 21618
rect 18310 21158 18344 21534
rect 18406 21158 18440 21534
rect 18502 21158 18536 21534
rect 18598 21158 18632 21534
rect 18694 21158 18728 21534
rect 18790 21158 18824 21534
rect 18886 21158 18920 21534
rect 18982 21158 19016 21534
rect 19078 21158 19112 21534
rect 19174 21158 19208 21534
rect 19270 21158 19304 21534
rect 18454 21074 18488 21108
rect 18646 21074 18680 21108
rect 18838 21074 18872 21108
rect 19030 21074 19064 21108
rect 19222 21074 19256 21108
rect 10314 19764 10348 19798
rect 10506 19764 10540 19798
rect 10698 19764 10732 19798
rect 10170 19338 10204 19714
rect 10266 19338 10300 19714
rect 10362 19338 10396 19714
rect 10458 19338 10492 19714
rect 10554 19338 10588 19714
rect 10650 19338 10684 19714
rect 10746 19338 10780 19714
rect 10842 19338 10876 19714
rect 10218 19254 10252 19288
rect 10410 19254 10444 19288
rect 10602 19254 10636 19288
rect 10794 19254 10828 19288
rect 10218 18842 10252 18876
rect 10410 18842 10444 18876
rect 10602 18842 10636 18876
rect 10794 18842 10828 18876
rect 10986 18842 11020 18876
rect 10170 18416 10204 18792
rect 10266 18416 10300 18792
rect 10362 18416 10396 18792
rect 10458 18416 10492 18792
rect 10554 18416 10588 18792
rect 10650 18416 10684 18792
rect 10746 18416 10780 18792
rect 10842 18416 10876 18792
rect 10938 18416 10972 18792
rect 11034 18416 11068 18792
rect 11130 18416 11164 18792
rect 10314 18332 10348 18366
rect 10506 18332 10540 18366
rect 10698 18332 10732 18366
rect 10890 18332 10924 18366
rect 11082 18332 11116 18366
rect 10314 18224 10348 18258
rect 10506 18224 10540 18258
rect 10698 18224 10732 18258
rect 10890 18224 10924 18258
rect 11082 18224 11116 18258
rect 10170 17798 10204 18174
rect 10266 17798 10300 18174
rect 10362 17798 10396 18174
rect 10458 17798 10492 18174
rect 10554 17798 10588 18174
rect 10650 17798 10684 18174
rect 10746 17798 10780 18174
rect 10842 17798 10876 18174
rect 10938 17798 10972 18174
rect 11034 17798 11068 18174
rect 11130 17798 11164 18174
rect 10218 17714 10252 17748
rect 10410 17714 10444 17748
rect 10602 17714 10636 17748
rect 10794 17714 10828 17748
rect 10986 17714 11020 17748
rect 18372 20718 18540 20752
rect 18630 20718 18798 20752
rect 18888 20718 19056 20752
rect 19146 20718 19314 20752
rect 19404 20718 19572 20752
rect 18310 20292 18344 20668
rect 18568 20292 18602 20668
rect 18826 20292 18860 20668
rect 19084 20292 19118 20668
rect 19342 20292 19376 20668
rect 19600 20292 19634 20668
rect 18372 20208 18540 20242
rect 18630 20208 18798 20242
rect 18888 20208 19056 20242
rect 19146 20208 19314 20242
rect 19404 20208 19572 20242
rect 18372 20100 18540 20134
rect 18630 20100 18798 20134
rect 18888 20100 19056 20134
rect 19146 20100 19314 20134
rect 19404 20100 19572 20134
rect 18310 19674 18344 20050
rect 18568 19674 18602 20050
rect 18826 19674 18860 20050
rect 19084 19674 19118 20050
rect 19342 19674 19376 20050
rect 19600 19674 19634 20050
rect 18372 19590 18540 19624
rect 18630 19590 18798 19624
rect 18888 19590 19056 19624
rect 19146 19590 19314 19624
rect 19404 19590 19572 19624
rect 18372 19482 18540 19516
rect 18630 19482 18798 19516
rect 18888 19482 19056 19516
rect 19146 19482 19314 19516
rect 19404 19482 19572 19516
rect 18310 19056 18344 19432
rect 18568 19056 18602 19432
rect 18826 19056 18860 19432
rect 19084 19056 19118 19432
rect 19342 19056 19376 19432
rect 19600 19056 19634 19432
rect 18372 18972 18540 19006
rect 18630 18972 18798 19006
rect 18888 18972 19056 19006
rect 19146 18972 19314 19006
rect 19404 18972 19572 19006
rect 18372 18864 18540 18898
rect 18630 18864 18798 18898
rect 18888 18864 19056 18898
rect 19146 18864 19314 18898
rect 19404 18864 19572 18898
rect 18310 18438 18344 18814
rect 18568 18438 18602 18814
rect 18826 18438 18860 18814
rect 19084 18438 19118 18814
rect 19342 18438 19376 18814
rect 19600 18438 19634 18814
rect 18372 18354 18540 18388
rect 18630 18354 18798 18388
rect 18888 18354 19056 18388
rect 19146 18354 19314 18388
rect 19404 18354 19572 18388
rect 18480 18056 18680 18156
rect 1300 10532 1568 10768
rect 2618 10703 2868 11100
rect 2996 10703 3246 11100
rect 3374 10703 3624 11100
rect 3752 10703 4002 11100
rect 4130 10703 4380 11100
rect 4508 10703 4758 11100
rect 2618 9472 2868 9869
rect 2996 9472 3246 9869
rect 3374 9472 3624 9869
rect 3752 9472 4002 9869
rect 4130 9472 4380 9869
rect 4508 9472 4758 9869
rect 6096 10608 6276 10808
rect 15700 10532 15968 10768
rect -9906 8272 -9872 8306
rect -9714 8272 -9680 8306
rect -9522 8272 -9488 8306
rect -9330 8272 -9296 8306
rect -9138 8272 -9104 8306
rect -10050 7846 -10016 8222
rect -9954 7846 -9920 8222
rect -9858 7846 -9824 8222
rect -9762 7846 -9728 8222
rect -9666 7846 -9632 8222
rect -9570 7846 -9536 8222
rect -9474 7846 -9440 8222
rect -9378 7846 -9344 8222
rect -9282 7846 -9248 8222
rect -9186 7846 -9152 8222
rect -9090 7846 -9056 8222
rect -10002 7762 -9968 7796
rect -9810 7762 -9776 7796
rect -9618 7762 -9584 7796
rect -9426 7762 -9392 7796
rect -9234 7762 -9200 7796
rect -10002 7654 -9968 7688
rect -9810 7654 -9776 7688
rect -9618 7654 -9584 7688
rect -9426 7654 -9392 7688
rect -9234 7654 -9200 7688
rect -10050 7228 -10016 7604
rect -9954 7228 -9920 7604
rect -9858 7228 -9824 7604
rect -9762 7228 -9728 7604
rect -9666 7228 -9632 7604
rect -9570 7228 -9536 7604
rect -9474 7228 -9440 7604
rect -9378 7228 -9344 7604
rect -9282 7228 -9248 7604
rect -9186 7228 -9152 7604
rect -9090 7228 -9056 7604
rect -9906 7144 -9872 7178
rect -9714 7144 -9680 7178
rect -9522 7144 -9488 7178
rect -9330 7144 -9296 7178
rect -9138 7144 -9104 7178
rect -9906 7036 -9872 7070
rect -9714 7036 -9680 7070
rect -9522 7036 -9488 7070
rect -9330 7036 -9296 7070
rect -9138 7036 -9104 7070
rect -10050 6610 -10016 6986
rect -9954 6610 -9920 6986
rect -9858 6610 -9824 6986
rect -9762 6610 -9728 6986
rect -9666 6610 -9632 6986
rect -9570 6610 -9536 6986
rect -9474 6610 -9440 6986
rect -9378 6610 -9344 6986
rect -9282 6610 -9248 6986
rect -9186 6610 -9152 6986
rect -9090 6610 -9056 6986
rect -10002 6526 -9968 6560
rect -9810 6526 -9776 6560
rect -9618 6526 -9584 6560
rect -9426 6526 -9392 6560
rect -9234 6526 -9200 6560
rect -8658 8196 -8482 8230
rect -8742 6600 -8708 8168
rect -8432 6600 -8398 8168
rect -8658 6538 -8482 6572
rect 1672 8904 1964 8964
rect 2540 8904 2832 8964
rect 3476 8904 3768 8964
rect 1834 8768 1868 8802
rect 2026 8768 2060 8802
rect 2218 8768 2252 8802
rect 2410 8768 2444 8802
rect 2602 8768 2636 8802
rect 2794 8768 2828 8802
rect 2986 8768 3020 8802
rect 3178 8768 3212 8802
rect 3370 8768 3404 8802
rect 3562 8768 3596 8802
rect 1540 8356 1576 8704
rect 1576 8356 1596 8704
rect 1690 8342 1724 8718
rect 1786 8342 1820 8718
rect 1882 8342 1916 8718
rect 1978 8342 2012 8718
rect 2074 8342 2108 8718
rect 2170 8342 2204 8718
rect 2266 8342 2300 8718
rect 2362 8342 2396 8718
rect 2458 8342 2492 8718
rect 2554 8342 2588 8718
rect 2650 8342 2684 8718
rect 2746 8342 2780 8718
rect 2842 8342 2876 8718
rect 2938 8342 2972 8718
rect 3034 8342 3068 8718
rect 3130 8342 3164 8718
rect 3226 8342 3260 8718
rect 3322 8342 3356 8718
rect 3418 8342 3452 8718
rect 3514 8342 3548 8718
rect 3610 8342 3644 8718
rect 3740 8416 3758 8672
rect 3758 8416 3800 8672
rect 1738 8258 1772 8292
rect 1930 8258 1964 8292
rect 2122 8258 2156 8292
rect 2314 8258 2348 8292
rect 2506 8258 2540 8292
rect 2698 8258 2732 8292
rect 2890 8258 2924 8292
rect 3082 8258 3116 8292
rect 3274 8258 3308 8292
rect 3466 8258 3500 8292
rect 1672 8088 1964 8148
rect 2540 8088 2860 8148
rect 3476 8092 3768 8152
rect 1834 7948 1868 7982
rect 2026 7948 2060 7982
rect 2218 7948 2252 7982
rect 2410 7948 2444 7982
rect 2602 7948 2636 7982
rect 2794 7948 2828 7982
rect 2986 7948 3020 7982
rect 3178 7948 3212 7982
rect 3370 7948 3404 7982
rect 3562 7948 3596 7982
rect 1540 7588 1576 7844
rect 1576 7588 1600 7844
rect 1690 7522 1724 7898
rect 1786 7522 1820 7898
rect 1882 7522 1916 7898
rect 1978 7522 2012 7898
rect 2074 7522 2108 7898
rect 2170 7522 2204 7898
rect 2266 7522 2300 7898
rect 2362 7522 2396 7898
rect 2458 7522 2492 7898
rect 2554 7522 2588 7898
rect 2650 7522 2684 7898
rect 2746 7522 2780 7898
rect 2842 7522 2876 7898
rect 2938 7522 2972 7898
rect 3034 7522 3068 7898
rect 3130 7522 3164 7898
rect 3226 7522 3260 7898
rect 3322 7522 3356 7898
rect 3418 7522 3452 7898
rect 3514 7522 3548 7898
rect 3610 7522 3644 7898
rect 3740 7568 3758 7824
rect 3758 7568 3800 7824
rect 1738 7438 1772 7472
rect 1930 7438 1964 7472
rect 2122 7438 2156 7472
rect 2314 7438 2348 7472
rect 2506 7438 2540 7472
rect 2698 7438 2732 7472
rect 2890 7438 2924 7472
rect 3082 7438 3116 7472
rect 3274 7438 3308 7472
rect 3466 7438 3500 7472
rect 1672 7268 1964 7328
rect 2540 7268 2832 7328
rect 3476 7268 3768 7328
rect 1834 7128 1868 7162
rect 2026 7128 2060 7162
rect 2218 7128 2252 7162
rect 2410 7128 2444 7162
rect 2602 7128 2636 7162
rect 2794 7128 2828 7162
rect 2986 7128 3020 7162
rect 3178 7128 3212 7162
rect 3370 7128 3404 7162
rect 3562 7128 3596 7162
rect 1536 6748 1576 7004
rect 1576 6748 1596 7004
rect 1690 6702 1724 7078
rect 1786 6702 1820 7078
rect 1882 6702 1916 7078
rect 1978 6702 2012 7078
rect 2074 6702 2108 7078
rect 2170 6702 2204 7078
rect 2266 6702 2300 7078
rect 2362 6702 2396 7078
rect 2458 6702 2492 7078
rect 2554 6702 2588 7078
rect 2650 6702 2684 7078
rect 2746 6702 2780 7078
rect 2842 6702 2876 7078
rect 2938 6702 2972 7078
rect 3034 6702 3068 7078
rect 3130 6702 3164 7078
rect 3226 6702 3260 7078
rect 3322 6702 3356 7078
rect 3418 6702 3452 7078
rect 3514 6702 3548 7078
rect 3610 6702 3644 7078
rect 3740 6756 3758 7012
rect 3758 6756 3800 7012
rect 1738 6618 1772 6652
rect 1930 6618 1964 6652
rect 2122 6618 2156 6652
rect 2314 6618 2348 6652
rect 2506 6618 2540 6652
rect 2698 6618 2732 6652
rect 2890 6618 2924 6652
rect 3082 6618 3116 6652
rect 3274 6618 3308 6652
rect 3466 6618 3500 6652
rect 1672 6456 1964 6516
rect 2540 6456 2832 6516
rect 3476 6452 3768 6512
rect 5174 10330 5208 10364
rect 5366 10330 5400 10364
rect 5558 10330 5592 10364
rect 5750 10330 5784 10364
rect 5942 10330 5976 10364
rect 6134 10330 6168 10364
rect 6326 10330 6360 10364
rect 6518 10330 6552 10364
rect 6710 10330 6744 10364
rect 6902 10330 6936 10364
rect 5126 9895 5160 10271
rect 5222 9895 5256 10271
rect 5318 9895 5352 10271
rect 5414 9895 5448 10271
rect 5510 9895 5544 10271
rect 5606 9895 5640 10271
rect 5702 9895 5736 10271
rect 5798 9895 5832 10271
rect 5894 9895 5928 10271
rect 5990 9895 6024 10271
rect 6086 9895 6120 10271
rect 6182 9895 6216 10271
rect 6278 9895 6312 10271
rect 6374 9895 6408 10271
rect 6470 9895 6504 10271
rect 6566 9895 6600 10271
rect 6662 9895 6696 10271
rect 6758 9895 6792 10271
rect 6854 9895 6888 10271
rect 6950 9895 6984 10271
rect 7046 9895 7080 10271
rect 5270 9802 5304 9836
rect 5462 9802 5496 9836
rect 5654 9802 5688 9836
rect 5846 9802 5880 9836
rect 6038 9802 6072 9836
rect 6230 9802 6264 9836
rect 6422 9802 6456 9836
rect 6614 9802 6648 9836
rect 6806 9802 6840 9836
rect 6998 9802 7032 9836
rect 5270 9694 5304 9728
rect 5462 9694 5496 9728
rect 5654 9694 5688 9728
rect 5846 9694 5880 9728
rect 6038 9694 6072 9728
rect 6230 9694 6264 9728
rect 6422 9694 6456 9728
rect 6614 9694 6648 9728
rect 6806 9694 6840 9728
rect 6998 9694 7032 9728
rect 5126 9259 5160 9635
rect 5222 9259 5256 9635
rect 5318 9259 5352 9635
rect 5414 9259 5448 9635
rect 5510 9259 5544 9635
rect 5606 9259 5640 9635
rect 5702 9259 5736 9635
rect 5798 9259 5832 9635
rect 5894 9259 5928 9635
rect 5990 9259 6024 9635
rect 6086 9259 6120 9635
rect 6182 9259 6216 9635
rect 6278 9259 6312 9635
rect 6374 9259 6408 9635
rect 6470 9259 6504 9635
rect 6566 9259 6600 9635
rect 6662 9259 6696 9635
rect 6758 9259 6792 9635
rect 6854 9259 6888 9635
rect 6950 9259 6984 9635
rect 7046 9259 7080 9635
rect 5174 9166 5208 9200
rect 5366 9166 5400 9200
rect 5558 9166 5592 9200
rect 5750 9166 5784 9200
rect 5942 9166 5976 9200
rect 6134 9166 6168 9200
rect 6326 9166 6360 9200
rect 6518 9166 6552 9200
rect 6710 9166 6744 9200
rect 6902 9166 6936 9200
rect 5174 8734 5208 8768
rect 5366 8734 5400 8768
rect 5558 8734 5592 8768
rect 5750 8734 5784 8768
rect 5942 8734 5976 8768
rect 6134 8734 6168 8768
rect 6326 8734 6360 8768
rect 6518 8734 6552 8768
rect 6710 8734 6744 8768
rect 6902 8734 6936 8768
rect 5126 8308 5160 8684
rect 5222 8308 5256 8684
rect 5318 8308 5352 8684
rect 5414 8308 5448 8684
rect 5510 8308 5544 8684
rect 5606 8308 5640 8684
rect 5702 8308 5736 8684
rect 5798 8308 5832 8684
rect 5894 8308 5928 8684
rect 5990 8308 6024 8684
rect 6086 8308 6120 8684
rect 6182 8308 6216 8684
rect 6278 8308 6312 8684
rect 6374 8308 6408 8684
rect 6470 8308 6504 8684
rect 6566 8308 6600 8684
rect 6662 8308 6696 8684
rect 6758 8308 6792 8684
rect 6854 8308 6888 8684
rect 6950 8308 6984 8684
rect 7046 8308 7080 8684
rect 5270 8224 5304 8258
rect 5462 8224 5496 8258
rect 5654 8224 5688 8258
rect 5846 8224 5880 8258
rect 6038 8224 6072 8258
rect 6230 8224 6264 8258
rect 6422 8224 6456 8258
rect 6614 8224 6648 8258
rect 6806 8224 6840 8258
rect 6998 8224 7032 8258
rect 5270 8116 5304 8150
rect 5462 8116 5496 8150
rect 5654 8116 5688 8150
rect 5846 8116 5880 8150
rect 6038 8116 6072 8150
rect 6230 8116 6264 8150
rect 6422 8116 6456 8150
rect 6614 8116 6648 8150
rect 6806 8116 6840 8150
rect 6998 8116 7032 8150
rect 5126 7690 5160 8066
rect 5222 7690 5256 8066
rect 5318 7690 5352 8066
rect 5414 7690 5448 8066
rect 5510 7690 5544 8066
rect 5606 7690 5640 8066
rect 5702 7690 5736 8066
rect 5798 7690 5832 8066
rect 5894 7690 5928 8066
rect 5990 7690 6024 8066
rect 6086 7690 6120 8066
rect 6182 7690 6216 8066
rect 6278 7690 6312 8066
rect 6374 7690 6408 8066
rect 6470 7690 6504 8066
rect 6566 7690 6600 8066
rect 6662 7690 6696 8066
rect 6758 7690 6792 8066
rect 6854 7690 6888 8066
rect 6950 7690 6984 8066
rect 7046 7690 7080 8066
rect 5174 7606 5208 7640
rect 5366 7606 5400 7640
rect 5558 7606 5592 7640
rect 5750 7606 5784 7640
rect 5942 7606 5976 7640
rect 6134 7606 6168 7640
rect 6326 7606 6360 7640
rect 6518 7606 6552 7640
rect 6710 7606 6744 7640
rect 6902 7606 6936 7640
rect -9906 6192 -9872 6226
rect -9714 6192 -9680 6226
rect -9522 6192 -9488 6226
rect -9330 6192 -9296 6226
rect -9138 6192 -9104 6226
rect -10050 5766 -10016 6142
rect -9954 5766 -9920 6142
rect -9858 5766 -9824 6142
rect -9762 5766 -9728 6142
rect -9666 5766 -9632 6142
rect -9570 5766 -9536 6142
rect -9474 5766 -9440 6142
rect -9378 5766 -9344 6142
rect -9282 5766 -9248 6142
rect -9186 5766 -9152 6142
rect -9090 5766 -9056 6142
rect -10002 5682 -9968 5716
rect -9810 5682 -9776 5716
rect -9618 5682 -9584 5716
rect -9426 5682 -9392 5716
rect -9234 5682 -9200 5716
rect -10002 5574 -9968 5608
rect -9810 5574 -9776 5608
rect -9618 5574 -9584 5608
rect -9426 5574 -9392 5608
rect -9234 5574 -9200 5608
rect -10050 5148 -10016 5524
rect -9954 5148 -9920 5524
rect -9858 5148 -9824 5524
rect -9762 5148 -9728 5524
rect -9666 5148 -9632 5524
rect -9570 5148 -9536 5524
rect -9474 5148 -9440 5524
rect -9378 5148 -9344 5524
rect -9282 5148 -9248 5524
rect -9186 5148 -9152 5524
rect -9090 5148 -9056 5524
rect -9906 5064 -9872 5098
rect -9714 5064 -9680 5098
rect -9522 5064 -9488 5098
rect -9330 5064 -9296 5098
rect -9138 5064 -9104 5098
rect -9906 4956 -9872 4990
rect -9714 4956 -9680 4990
rect -9522 4956 -9488 4990
rect -9330 4956 -9296 4990
rect -9138 4956 -9104 4990
rect -10050 4530 -10016 4906
rect -9954 4530 -9920 4906
rect -9858 4530 -9824 4906
rect -9762 4530 -9728 4906
rect -9666 4530 -9632 4906
rect -9570 4530 -9536 4906
rect -9474 4530 -9440 4906
rect -9378 4530 -9344 4906
rect -9282 4530 -9248 4906
rect -9186 4530 -9152 4906
rect -9090 4530 -9056 4906
rect -10002 4446 -9968 4480
rect -9810 4446 -9776 4480
rect -9618 4446 -9584 4480
rect -9426 4446 -9392 4480
rect -9234 4446 -9200 4480
rect -9988 4046 -9820 4080
rect -9730 4046 -9562 4080
rect -9472 4046 -9304 4080
rect -9214 4046 -9046 4080
rect -8956 4046 -8788 4080
rect -10050 3620 -10016 3996
rect -9792 3620 -9758 3996
rect -9534 3620 -9500 3996
rect -9276 3620 -9242 3996
rect -9018 3620 -8984 3996
rect -8760 3620 -8726 3996
rect -9988 3536 -9820 3570
rect -9730 3536 -9562 3570
rect -9472 3536 -9304 3570
rect -9214 3536 -9046 3570
rect -8956 3536 -8788 3570
rect -9988 3428 -9820 3462
rect -9730 3428 -9562 3462
rect -9472 3428 -9304 3462
rect -9214 3428 -9046 3462
rect -8956 3428 -8788 3462
rect -10050 3002 -10016 3378
rect -9792 3002 -9758 3378
rect -9534 3002 -9500 3378
rect -9276 3002 -9242 3378
rect -9018 3002 -8984 3378
rect -8760 3002 -8726 3378
rect -9988 2918 -9820 2952
rect -9730 2918 -9562 2952
rect -9472 2918 -9304 2952
rect -9214 2918 -9046 2952
rect -8956 2918 -8788 2952
rect -9988 2810 -9820 2844
rect -9730 2810 -9562 2844
rect -9472 2810 -9304 2844
rect -9214 2810 -9046 2844
rect -8956 2810 -8788 2844
rect -10050 2384 -10016 2760
rect -9792 2384 -9758 2760
rect -9534 2384 -9500 2760
rect -9276 2384 -9242 2760
rect -9018 2384 -8984 2760
rect -8760 2384 -8726 2760
rect -9988 2300 -9820 2334
rect -9730 2300 -9562 2334
rect -9472 2300 -9304 2334
rect -9214 2300 -9046 2334
rect -8956 2300 -8788 2334
rect -9988 2192 -9820 2226
rect -9730 2192 -9562 2226
rect -9472 2192 -9304 2226
rect -9214 2192 -9046 2226
rect -8956 2192 -8788 2226
rect -10050 1766 -10016 2142
rect -9792 1766 -9758 2142
rect -9534 1766 -9500 2142
rect -9276 1766 -9242 2142
rect -9018 1766 -8984 2142
rect -8760 1766 -8726 2142
rect -9988 1682 -9820 1716
rect -9730 1682 -9562 1716
rect -9472 1682 -9304 1716
rect -9214 1682 -9046 1716
rect -8956 1682 -8788 1716
rect -9988 1574 -9820 1608
rect -9730 1574 -9562 1608
rect -9472 1574 -9304 1608
rect -9214 1574 -9046 1608
rect -8956 1574 -8788 1608
rect -10050 1148 -10016 1524
rect -9792 1148 -9758 1524
rect -9534 1148 -9500 1524
rect -9276 1148 -9242 1524
rect -9018 1148 -8984 1524
rect -8760 1148 -8726 1524
rect -9988 1064 -9820 1098
rect -9730 1064 -9562 1098
rect -9472 1064 -9304 1098
rect -9214 1064 -9046 1098
rect -8956 1064 -8788 1098
rect -9988 956 -9820 990
rect -9730 956 -9562 990
rect -9472 956 -9304 990
rect -9214 956 -9046 990
rect -8956 956 -8788 990
rect -10050 530 -10016 906
rect -9792 530 -9758 906
rect -9534 530 -9500 906
rect -9276 530 -9242 906
rect -9018 530 -8984 906
rect -8760 530 -8726 906
rect -9988 446 -9820 480
rect -9730 446 -9562 480
rect -9472 446 -9304 480
rect -9214 446 -9046 480
rect -8956 446 -8788 480
rect 370 5912 404 5946
rect 562 5912 596 5946
rect 754 5912 788 5946
rect 946 5912 980 5946
rect 1138 5912 1172 5946
rect 226 5486 260 5862
rect 322 5486 356 5862
rect 418 5486 452 5862
rect 514 5486 548 5862
rect 610 5486 644 5862
rect 706 5486 740 5862
rect 802 5486 836 5862
rect 898 5486 932 5862
rect 994 5486 1028 5862
rect 1090 5486 1124 5862
rect 1186 5486 1220 5862
rect 274 5402 308 5436
rect 466 5402 500 5436
rect 658 5402 692 5436
rect 850 5402 884 5436
rect 1042 5402 1076 5436
rect 274 5294 308 5328
rect 466 5294 500 5328
rect 658 5294 692 5328
rect 850 5294 884 5328
rect 1042 5294 1076 5328
rect 226 4868 260 5244
rect 322 4868 356 5244
rect 418 4868 452 5244
rect 514 4868 548 5244
rect 610 4868 644 5244
rect 706 4868 740 5244
rect 802 4868 836 5244
rect 898 4868 932 5244
rect 994 4868 1028 5244
rect 1090 4868 1124 5244
rect 1186 4868 1220 5244
rect 370 4784 404 4818
rect 562 4784 596 4818
rect 754 4784 788 4818
rect 946 4784 980 4818
rect 1138 4784 1172 4818
rect 370 4676 404 4710
rect 562 4676 596 4710
rect 754 4676 788 4710
rect 946 4676 980 4710
rect 1138 4676 1172 4710
rect 226 4250 260 4626
rect 322 4250 356 4626
rect 418 4250 452 4626
rect 514 4250 548 4626
rect 610 4250 644 4626
rect 706 4250 740 4626
rect 802 4250 836 4626
rect 898 4250 932 4626
rect 994 4250 1028 4626
rect 1090 4250 1124 4626
rect 1186 4250 1220 4626
rect 274 4166 308 4200
rect 466 4166 500 4200
rect 658 4166 692 4200
rect 850 4166 884 4200
rect 1042 4166 1076 4200
rect 2170 5912 2204 5946
rect 2362 5912 2396 5946
rect 2554 5912 2588 5946
rect 2746 5912 2780 5946
rect 2938 5912 2972 5946
rect 2026 5486 2060 5862
rect 2122 5486 2156 5862
rect 2218 5486 2252 5862
rect 2314 5486 2348 5862
rect 2410 5486 2444 5862
rect 2506 5486 2540 5862
rect 2602 5486 2636 5862
rect 2698 5486 2732 5862
rect 2794 5486 2828 5862
rect 2890 5486 2924 5862
rect 2986 5486 3020 5862
rect 2074 5402 2108 5436
rect 2266 5402 2300 5436
rect 2458 5402 2492 5436
rect 2650 5402 2684 5436
rect 2842 5402 2876 5436
rect 2074 5294 2108 5328
rect 2266 5294 2300 5328
rect 2458 5294 2492 5328
rect 2650 5294 2684 5328
rect 2842 5294 2876 5328
rect 2026 4868 2060 5244
rect 2122 4868 2156 5244
rect 2218 4868 2252 5244
rect 2314 4868 2348 5244
rect 2410 4868 2444 5244
rect 2506 4868 2540 5244
rect 2602 4868 2636 5244
rect 2698 4868 2732 5244
rect 2794 4868 2828 5244
rect 2890 4868 2924 5244
rect 2986 4868 3020 5244
rect 2170 4784 2204 4818
rect 2362 4784 2396 4818
rect 2554 4784 2588 4818
rect 2746 4784 2780 4818
rect 2938 4784 2972 4818
rect 2170 4676 2204 4710
rect 2362 4676 2396 4710
rect 2554 4676 2588 4710
rect 2746 4676 2780 4710
rect 2938 4676 2972 4710
rect 2026 4250 2060 4626
rect 2122 4250 2156 4626
rect 2218 4250 2252 4626
rect 2314 4250 2348 4626
rect 2410 4250 2444 4626
rect 2506 4250 2540 4626
rect 2602 4250 2636 4626
rect 2698 4250 2732 4626
rect 2794 4250 2828 4626
rect 2890 4250 2924 4626
rect 2986 4250 3020 4626
rect 2074 4166 2108 4200
rect 2266 4166 2300 4200
rect 2458 4166 2492 4200
rect 2650 4166 2684 4200
rect 2842 4166 2876 4200
rect 3970 5912 4004 5946
rect 4162 5912 4196 5946
rect 4354 5912 4388 5946
rect 4546 5912 4580 5946
rect 4738 5912 4772 5946
rect 3826 5486 3860 5862
rect 3922 5486 3956 5862
rect 4018 5486 4052 5862
rect 4114 5486 4148 5862
rect 4210 5486 4244 5862
rect 4306 5486 4340 5862
rect 4402 5486 4436 5862
rect 4498 5486 4532 5862
rect 4594 5486 4628 5862
rect 4690 5486 4724 5862
rect 4786 5486 4820 5862
rect 3874 5402 3908 5436
rect 4066 5402 4100 5436
rect 4258 5402 4292 5436
rect 4450 5402 4484 5436
rect 4642 5402 4676 5436
rect 3874 5294 3908 5328
rect 4066 5294 4100 5328
rect 4258 5294 4292 5328
rect 4450 5294 4484 5328
rect 4642 5294 4676 5328
rect 3826 4868 3860 5244
rect 3922 4868 3956 5244
rect 4018 4868 4052 5244
rect 4114 4868 4148 5244
rect 4210 4868 4244 5244
rect 4306 4868 4340 5244
rect 4402 4868 4436 5244
rect 4498 4868 4532 5244
rect 4594 4868 4628 5244
rect 4690 4868 4724 5244
rect 4786 4868 4820 5244
rect 3970 4784 4004 4818
rect 4162 4784 4196 4818
rect 4354 4784 4388 4818
rect 4546 4784 4580 4818
rect 4738 4784 4772 4818
rect 3970 4676 4004 4710
rect 4162 4676 4196 4710
rect 4354 4676 4388 4710
rect 4546 4676 4580 4710
rect 4738 4676 4772 4710
rect 3826 4250 3860 4626
rect 3922 4250 3956 4626
rect 4018 4250 4052 4626
rect 4114 4250 4148 4626
rect 4210 4250 4244 4626
rect 4306 4250 4340 4626
rect 4402 4250 4436 4626
rect 4498 4250 4532 4626
rect 4594 4250 4628 4626
rect 4690 4250 4724 4626
rect 4786 4250 4820 4626
rect 3874 4166 3908 4200
rect 4066 4166 4100 4200
rect 4258 4166 4292 4200
rect 4450 4166 4484 4200
rect 4642 4166 4676 4200
rect 5770 5912 5804 5946
rect 5962 5912 5996 5946
rect 6154 5912 6188 5946
rect 6346 5912 6380 5946
rect 6538 5912 6572 5946
rect 5626 5486 5660 5862
rect 5722 5486 5756 5862
rect 5818 5486 5852 5862
rect 5914 5486 5948 5862
rect 6010 5486 6044 5862
rect 6106 5486 6140 5862
rect 6202 5486 6236 5862
rect 6298 5486 6332 5862
rect 6394 5486 6428 5862
rect 6490 5486 6524 5862
rect 6586 5486 6620 5862
rect 5674 5402 5708 5436
rect 5866 5402 5900 5436
rect 6058 5402 6092 5436
rect 6250 5402 6284 5436
rect 6442 5402 6476 5436
rect 5674 5294 5708 5328
rect 5866 5294 5900 5328
rect 6058 5294 6092 5328
rect 6250 5294 6284 5328
rect 6442 5294 6476 5328
rect 5626 4868 5660 5244
rect 5722 4868 5756 5244
rect 5818 4868 5852 5244
rect 5914 4868 5948 5244
rect 6010 4868 6044 5244
rect 6106 4868 6140 5244
rect 6202 4868 6236 5244
rect 6298 4868 6332 5244
rect 6394 4868 6428 5244
rect 6490 4868 6524 5244
rect 6586 4868 6620 5244
rect 5770 4784 5804 4818
rect 5962 4784 5996 4818
rect 6154 4784 6188 4818
rect 6346 4784 6380 4818
rect 6538 4784 6572 4818
rect 5770 4676 5804 4710
rect 5962 4676 5996 4710
rect 6154 4676 6188 4710
rect 6346 4676 6380 4710
rect 6538 4676 6572 4710
rect 5626 4250 5660 4626
rect 5722 4250 5756 4626
rect 5818 4250 5852 4626
rect 5914 4250 5948 4626
rect 6010 4250 6044 4626
rect 6106 4250 6140 4626
rect 6202 4250 6236 4626
rect 6298 4250 6332 4626
rect 6394 4250 6428 4626
rect 6490 4250 6524 4626
rect 6586 4250 6620 4626
rect 5674 4166 5708 4200
rect 5866 4166 5900 4200
rect 6058 4166 6092 4200
rect 6250 4166 6284 4200
rect 6442 4166 6476 4200
rect 7770 10300 7804 10334
rect 7962 10300 7996 10334
rect 8154 10300 8188 10334
rect 8346 10300 8380 10334
rect 8538 10300 8572 10334
rect 8730 10300 8764 10334
rect 8922 10300 8956 10334
rect 9114 10300 9148 10334
rect 9306 10300 9340 10334
rect 9498 10300 9532 10334
rect 7626 9874 7660 10250
rect 7722 9874 7756 10250
rect 7818 9874 7852 10250
rect 7914 9874 7948 10250
rect 8010 9874 8044 10250
rect 8106 9874 8140 10250
rect 8202 9874 8236 10250
rect 8298 9874 8332 10250
rect 8394 9874 8428 10250
rect 8490 9874 8524 10250
rect 8586 9874 8620 10250
rect 8682 9874 8716 10250
rect 8778 9874 8812 10250
rect 8874 9874 8908 10250
rect 8970 9874 9004 10250
rect 9066 9874 9100 10250
rect 9162 9874 9196 10250
rect 9258 9874 9292 10250
rect 9354 9874 9388 10250
rect 9450 9874 9484 10250
rect 9546 9874 9580 10250
rect 7674 9790 7708 9824
rect 7866 9790 7900 9824
rect 8058 9790 8092 9824
rect 8250 9790 8284 9824
rect 8442 9790 8476 9824
rect 8634 9790 8668 9824
rect 8826 9790 8860 9824
rect 9018 9790 9052 9824
rect 9210 9790 9244 9824
rect 9402 9790 9436 9824
rect 7674 9682 7708 9716
rect 7866 9682 7900 9716
rect 8058 9682 8092 9716
rect 8250 9682 8284 9716
rect 8442 9682 8476 9716
rect 8634 9682 8668 9716
rect 8826 9682 8860 9716
rect 9018 9682 9052 9716
rect 9210 9682 9244 9716
rect 9402 9682 9436 9716
rect 7626 9256 7660 9632
rect 7722 9256 7756 9632
rect 7818 9256 7852 9632
rect 7914 9256 7948 9632
rect 8010 9256 8044 9632
rect 8106 9256 8140 9632
rect 8202 9256 8236 9632
rect 8298 9256 8332 9632
rect 8394 9256 8428 9632
rect 8490 9256 8524 9632
rect 8586 9256 8620 9632
rect 8682 9256 8716 9632
rect 8778 9256 8812 9632
rect 8874 9256 8908 9632
rect 8970 9256 9004 9632
rect 9066 9256 9100 9632
rect 9162 9256 9196 9632
rect 9258 9256 9292 9632
rect 9354 9256 9388 9632
rect 9450 9256 9484 9632
rect 9546 9256 9580 9632
rect 7770 9172 7804 9206
rect 7962 9172 7996 9206
rect 8154 9172 8188 9206
rect 8346 9172 8380 9206
rect 8538 9172 8572 9206
rect 8730 9172 8764 9206
rect 8922 9172 8956 9206
rect 9114 9172 9148 9206
rect 9306 9172 9340 9206
rect 9498 9172 9532 9206
rect 7770 9064 7804 9098
rect 7962 9064 7996 9098
rect 8154 9064 8188 9098
rect 8346 9064 8380 9098
rect 8538 9064 8572 9098
rect 8730 9064 8764 9098
rect 8922 9064 8956 9098
rect 9114 9064 9148 9098
rect 9306 9064 9340 9098
rect 9498 9064 9532 9098
rect 7626 8638 7660 9014
rect 7722 8638 7756 9014
rect 7818 8638 7852 9014
rect 7914 8638 7948 9014
rect 8010 8638 8044 9014
rect 8106 8638 8140 9014
rect 8202 8638 8236 9014
rect 8298 8638 8332 9014
rect 8394 8638 8428 9014
rect 8490 8638 8524 9014
rect 8586 8638 8620 9014
rect 8682 8638 8716 9014
rect 8778 8638 8812 9014
rect 8874 8638 8908 9014
rect 8970 8638 9004 9014
rect 9066 8638 9100 9014
rect 9162 8638 9196 9014
rect 9258 8638 9292 9014
rect 9354 8638 9388 9014
rect 9450 8638 9484 9014
rect 9546 8638 9580 9014
rect 7674 8554 7708 8588
rect 7866 8554 7900 8588
rect 8058 8554 8092 8588
rect 8250 8554 8284 8588
rect 8442 8554 8476 8588
rect 8634 8554 8668 8588
rect 8826 8554 8860 8588
rect 9018 8554 9052 8588
rect 9210 8554 9244 8588
rect 9402 8554 9436 8588
rect 7674 8446 7708 8480
rect 7866 8446 7900 8480
rect 8058 8446 8092 8480
rect 8250 8446 8284 8480
rect 8442 8446 8476 8480
rect 8634 8446 8668 8480
rect 8826 8446 8860 8480
rect 9018 8446 9052 8480
rect 9210 8446 9244 8480
rect 9402 8446 9436 8480
rect 7626 8020 7660 8396
rect 7722 8020 7756 8396
rect 7818 8020 7852 8396
rect 7914 8020 7948 8396
rect 8010 8020 8044 8396
rect 8106 8020 8140 8396
rect 8202 8020 8236 8396
rect 8298 8020 8332 8396
rect 8394 8020 8428 8396
rect 8490 8020 8524 8396
rect 8586 8020 8620 8396
rect 8682 8020 8716 8396
rect 8778 8020 8812 8396
rect 8874 8020 8908 8396
rect 8970 8020 9004 8396
rect 9066 8020 9100 8396
rect 9162 8020 9196 8396
rect 9258 8020 9292 8396
rect 9354 8020 9388 8396
rect 9450 8020 9484 8396
rect 9546 8020 9580 8396
rect 7770 7936 7804 7970
rect 7962 7936 7996 7970
rect 8154 7936 8188 7970
rect 8346 7936 8380 7970
rect 8538 7936 8572 7970
rect 8730 7936 8764 7970
rect 8922 7936 8956 7970
rect 9114 7936 9148 7970
rect 9306 7936 9340 7970
rect 9498 7936 9532 7970
rect 7770 7828 7804 7862
rect 7962 7828 7996 7862
rect 8154 7828 8188 7862
rect 8346 7828 8380 7862
rect 8538 7828 8572 7862
rect 8730 7828 8764 7862
rect 8922 7828 8956 7862
rect 9114 7828 9148 7862
rect 9306 7828 9340 7862
rect 9498 7828 9532 7862
rect 7626 7402 7660 7778
rect 7722 7402 7756 7778
rect 7818 7402 7852 7778
rect 7914 7402 7948 7778
rect 8010 7402 8044 7778
rect 8106 7402 8140 7778
rect 8202 7402 8236 7778
rect 8298 7402 8332 7778
rect 8394 7402 8428 7778
rect 8490 7402 8524 7778
rect 8586 7402 8620 7778
rect 8682 7402 8716 7778
rect 8778 7402 8812 7778
rect 8874 7402 8908 7778
rect 8970 7402 9004 7778
rect 9066 7402 9100 7778
rect 9162 7402 9196 7778
rect 9258 7402 9292 7778
rect 9354 7402 9388 7778
rect 9450 7402 9484 7778
rect 9546 7402 9580 7778
rect 7674 7318 7708 7352
rect 7866 7318 7900 7352
rect 8058 7318 8092 7352
rect 8250 7318 8284 7352
rect 8442 7318 8476 7352
rect 8634 7318 8668 7352
rect 8826 7318 8860 7352
rect 9018 7318 9052 7352
rect 9210 7318 9244 7352
rect 9402 7318 9436 7352
rect 7674 7210 7708 7244
rect 7866 7210 7900 7244
rect 8058 7210 8092 7244
rect 8250 7210 8284 7244
rect 8442 7210 8476 7244
rect 8634 7210 8668 7244
rect 8826 7210 8860 7244
rect 9018 7210 9052 7244
rect 9210 7210 9244 7244
rect 9402 7210 9436 7244
rect 7626 6784 7660 7160
rect 7722 6784 7756 7160
rect 7818 6784 7852 7160
rect 7914 6784 7948 7160
rect 8010 6784 8044 7160
rect 8106 6784 8140 7160
rect 8202 6784 8236 7160
rect 8298 6784 8332 7160
rect 8394 6784 8428 7160
rect 8490 6784 8524 7160
rect 8586 6784 8620 7160
rect 8682 6784 8716 7160
rect 8778 6784 8812 7160
rect 8874 6784 8908 7160
rect 8970 6784 9004 7160
rect 9066 6784 9100 7160
rect 9162 6784 9196 7160
rect 9258 6784 9292 7160
rect 9354 6784 9388 7160
rect 9450 6784 9484 7160
rect 9546 6784 9580 7160
rect 7770 6700 7804 6734
rect 7962 6700 7996 6734
rect 8154 6700 8188 6734
rect 8346 6700 8380 6734
rect 8538 6700 8572 6734
rect 8730 6700 8764 6734
rect 8922 6700 8956 6734
rect 9114 6700 9148 6734
rect 9306 6700 9340 6734
rect 9498 6700 9532 6734
rect 7770 6592 7804 6626
rect 7962 6592 7996 6626
rect 8154 6592 8188 6626
rect 8346 6592 8380 6626
rect 8538 6592 8572 6626
rect 8730 6592 8764 6626
rect 8922 6592 8956 6626
rect 9114 6592 9148 6626
rect 9306 6592 9340 6626
rect 9498 6592 9532 6626
rect 7626 6166 7660 6542
rect 7722 6166 7756 6542
rect 7818 6166 7852 6542
rect 7914 6166 7948 6542
rect 8010 6166 8044 6542
rect 8106 6166 8140 6542
rect 8202 6166 8236 6542
rect 8298 6166 8332 6542
rect 8394 6166 8428 6542
rect 8490 6166 8524 6542
rect 8586 6166 8620 6542
rect 8682 6166 8716 6542
rect 8778 6166 8812 6542
rect 8874 6166 8908 6542
rect 8970 6166 9004 6542
rect 9066 6166 9100 6542
rect 9162 6166 9196 6542
rect 9258 6166 9292 6542
rect 9354 6166 9388 6542
rect 9450 6166 9484 6542
rect 9546 6166 9580 6542
rect 7674 6082 7708 6116
rect 7866 6082 7900 6116
rect 8058 6082 8092 6116
rect 8250 6082 8284 6116
rect 8442 6082 8476 6116
rect 8634 6082 8668 6116
rect 8826 6082 8860 6116
rect 9018 6082 9052 6116
rect 9210 6082 9244 6116
rect 9402 6082 9436 6116
rect 7674 5974 7708 6008
rect 7866 5974 7900 6008
rect 8058 5974 8092 6008
rect 8250 5974 8284 6008
rect 8442 5974 8476 6008
rect 8634 5974 8668 6008
rect 8826 5974 8860 6008
rect 9018 5974 9052 6008
rect 9210 5974 9244 6008
rect 9402 5974 9436 6008
rect 7626 5548 7660 5924
rect 7722 5548 7756 5924
rect 7818 5548 7852 5924
rect 7914 5548 7948 5924
rect 8010 5548 8044 5924
rect 8106 5548 8140 5924
rect 8202 5548 8236 5924
rect 8298 5548 8332 5924
rect 8394 5548 8428 5924
rect 8490 5548 8524 5924
rect 8586 5548 8620 5924
rect 8682 5548 8716 5924
rect 8778 5548 8812 5924
rect 8874 5548 8908 5924
rect 8970 5548 9004 5924
rect 9066 5548 9100 5924
rect 9162 5548 9196 5924
rect 9258 5548 9292 5924
rect 9354 5548 9388 5924
rect 9450 5548 9484 5924
rect 9546 5548 9580 5924
rect 7770 5464 7804 5498
rect 7962 5464 7996 5498
rect 8154 5464 8188 5498
rect 8346 5464 8380 5498
rect 8538 5464 8572 5498
rect 8730 5464 8764 5498
rect 8922 5464 8956 5498
rect 9114 5464 9148 5498
rect 9306 5464 9340 5498
rect 9498 5464 9532 5498
rect 7770 5356 7804 5390
rect 7962 5356 7996 5390
rect 8154 5356 8188 5390
rect 8346 5356 8380 5390
rect 8538 5356 8572 5390
rect 8730 5356 8764 5390
rect 8922 5356 8956 5390
rect 9114 5356 9148 5390
rect 9306 5356 9340 5390
rect 9498 5356 9532 5390
rect 7626 4930 7660 5306
rect 7722 4930 7756 5306
rect 7818 4930 7852 5306
rect 7914 4930 7948 5306
rect 8010 4930 8044 5306
rect 8106 4930 8140 5306
rect 8202 4930 8236 5306
rect 8298 4930 8332 5306
rect 8394 4930 8428 5306
rect 8490 4930 8524 5306
rect 8586 4930 8620 5306
rect 8682 4930 8716 5306
rect 8778 4930 8812 5306
rect 8874 4930 8908 5306
rect 8970 4930 9004 5306
rect 9066 4930 9100 5306
rect 9162 4930 9196 5306
rect 9258 4930 9292 5306
rect 9354 4930 9388 5306
rect 9450 4930 9484 5306
rect 9546 4930 9580 5306
rect 7674 4846 7708 4880
rect 7866 4846 7900 4880
rect 8058 4846 8092 4880
rect 8250 4846 8284 4880
rect 8442 4846 8476 4880
rect 8634 4846 8668 4880
rect 8826 4846 8860 4880
rect 9018 4846 9052 4880
rect 9210 4846 9244 4880
rect 9402 4846 9436 4880
rect 17018 10703 17268 11100
rect 17396 10703 17646 11100
rect 17774 10703 18024 11100
rect 18152 10703 18402 11100
rect 18530 10703 18780 11100
rect 18908 10703 19158 11100
rect 17018 9472 17268 9869
rect 17396 9472 17646 9869
rect 17774 9472 18024 9869
rect 18152 9472 18402 9869
rect 18530 9472 18780 9869
rect 18908 9472 19158 9869
rect 20496 10608 20676 10808
rect 16072 8904 16364 8964
rect 16940 8904 17232 8964
rect 17876 8904 18168 8964
rect 16234 8768 16268 8802
rect 16426 8768 16460 8802
rect 16618 8768 16652 8802
rect 16810 8768 16844 8802
rect 17002 8768 17036 8802
rect 17194 8768 17228 8802
rect 17386 8768 17420 8802
rect 17578 8768 17612 8802
rect 17770 8768 17804 8802
rect 17962 8768 17996 8802
rect 15940 8356 15976 8704
rect 15976 8356 15996 8704
rect 16090 8342 16124 8718
rect 16186 8342 16220 8718
rect 16282 8342 16316 8718
rect 16378 8342 16412 8718
rect 16474 8342 16508 8718
rect 16570 8342 16604 8718
rect 16666 8342 16700 8718
rect 16762 8342 16796 8718
rect 16858 8342 16892 8718
rect 16954 8342 16988 8718
rect 17050 8342 17084 8718
rect 17146 8342 17180 8718
rect 17242 8342 17276 8718
rect 17338 8342 17372 8718
rect 17434 8342 17468 8718
rect 17530 8342 17564 8718
rect 17626 8342 17660 8718
rect 17722 8342 17756 8718
rect 17818 8342 17852 8718
rect 17914 8342 17948 8718
rect 18010 8342 18044 8718
rect 18140 8416 18158 8672
rect 18158 8416 18200 8672
rect 16138 8258 16172 8292
rect 16330 8258 16364 8292
rect 16522 8258 16556 8292
rect 16714 8258 16748 8292
rect 16906 8258 16940 8292
rect 17098 8258 17132 8292
rect 17290 8258 17324 8292
rect 17482 8258 17516 8292
rect 17674 8258 17708 8292
rect 17866 8258 17900 8292
rect 16072 8088 16364 8148
rect 16940 8088 17260 8148
rect 17876 8092 18168 8152
rect 16234 7948 16268 7982
rect 16426 7948 16460 7982
rect 16618 7948 16652 7982
rect 16810 7948 16844 7982
rect 17002 7948 17036 7982
rect 17194 7948 17228 7982
rect 17386 7948 17420 7982
rect 17578 7948 17612 7982
rect 17770 7948 17804 7982
rect 17962 7948 17996 7982
rect 15940 7588 15976 7844
rect 15976 7588 16000 7844
rect 16090 7522 16124 7898
rect 16186 7522 16220 7898
rect 16282 7522 16316 7898
rect 16378 7522 16412 7898
rect 16474 7522 16508 7898
rect 16570 7522 16604 7898
rect 16666 7522 16700 7898
rect 16762 7522 16796 7898
rect 16858 7522 16892 7898
rect 16954 7522 16988 7898
rect 17050 7522 17084 7898
rect 17146 7522 17180 7898
rect 17242 7522 17276 7898
rect 17338 7522 17372 7898
rect 17434 7522 17468 7898
rect 17530 7522 17564 7898
rect 17626 7522 17660 7898
rect 17722 7522 17756 7898
rect 17818 7522 17852 7898
rect 17914 7522 17948 7898
rect 18010 7522 18044 7898
rect 18140 7568 18158 7824
rect 18158 7568 18200 7824
rect 16138 7438 16172 7472
rect 16330 7438 16364 7472
rect 16522 7438 16556 7472
rect 16714 7438 16748 7472
rect 16906 7438 16940 7472
rect 17098 7438 17132 7472
rect 17290 7438 17324 7472
rect 17482 7438 17516 7472
rect 17674 7438 17708 7472
rect 17866 7438 17900 7472
rect 16072 7268 16364 7328
rect 16940 7268 17232 7328
rect 17876 7268 18168 7328
rect 16234 7128 16268 7162
rect 16426 7128 16460 7162
rect 16618 7128 16652 7162
rect 16810 7128 16844 7162
rect 17002 7128 17036 7162
rect 17194 7128 17228 7162
rect 17386 7128 17420 7162
rect 17578 7128 17612 7162
rect 17770 7128 17804 7162
rect 17962 7128 17996 7162
rect 15936 6748 15976 7004
rect 15976 6748 15996 7004
rect 16090 6702 16124 7078
rect 16186 6702 16220 7078
rect 16282 6702 16316 7078
rect 16378 6702 16412 7078
rect 16474 6702 16508 7078
rect 16570 6702 16604 7078
rect 16666 6702 16700 7078
rect 16762 6702 16796 7078
rect 16858 6702 16892 7078
rect 16954 6702 16988 7078
rect 17050 6702 17084 7078
rect 17146 6702 17180 7078
rect 17242 6702 17276 7078
rect 17338 6702 17372 7078
rect 17434 6702 17468 7078
rect 17530 6702 17564 7078
rect 17626 6702 17660 7078
rect 17722 6702 17756 7078
rect 17818 6702 17852 7078
rect 17914 6702 17948 7078
rect 18010 6702 18044 7078
rect 18140 6756 18158 7012
rect 18158 6756 18200 7012
rect 16138 6618 16172 6652
rect 16330 6618 16364 6652
rect 16522 6618 16556 6652
rect 16714 6618 16748 6652
rect 16906 6618 16940 6652
rect 17098 6618 17132 6652
rect 17290 6618 17324 6652
rect 17482 6618 17516 6652
rect 17674 6618 17708 6652
rect 17866 6618 17900 6652
rect 16072 6456 16364 6516
rect 16940 6456 17232 6516
rect 17876 6452 18168 6512
rect 19574 10330 19608 10364
rect 19766 10330 19800 10364
rect 19958 10330 19992 10364
rect 20150 10330 20184 10364
rect 20342 10330 20376 10364
rect 20534 10330 20568 10364
rect 20726 10330 20760 10364
rect 20918 10330 20952 10364
rect 21110 10330 21144 10364
rect 21302 10330 21336 10364
rect 19526 9895 19560 10271
rect 19622 9895 19656 10271
rect 19718 9895 19752 10271
rect 19814 9895 19848 10271
rect 19910 9895 19944 10271
rect 20006 9895 20040 10271
rect 20102 9895 20136 10271
rect 20198 9895 20232 10271
rect 20294 9895 20328 10271
rect 20390 9895 20424 10271
rect 20486 9895 20520 10271
rect 20582 9895 20616 10271
rect 20678 9895 20712 10271
rect 20774 9895 20808 10271
rect 20870 9895 20904 10271
rect 20966 9895 21000 10271
rect 21062 9895 21096 10271
rect 21158 9895 21192 10271
rect 21254 9895 21288 10271
rect 21350 9895 21384 10271
rect 21446 9895 21480 10271
rect 19670 9802 19704 9836
rect 19862 9802 19896 9836
rect 20054 9802 20088 9836
rect 20246 9802 20280 9836
rect 20438 9802 20472 9836
rect 20630 9802 20664 9836
rect 20822 9802 20856 9836
rect 21014 9802 21048 9836
rect 21206 9802 21240 9836
rect 21398 9802 21432 9836
rect 19670 9694 19704 9728
rect 19862 9694 19896 9728
rect 20054 9694 20088 9728
rect 20246 9694 20280 9728
rect 20438 9694 20472 9728
rect 20630 9694 20664 9728
rect 20822 9694 20856 9728
rect 21014 9694 21048 9728
rect 21206 9694 21240 9728
rect 21398 9694 21432 9728
rect 19526 9259 19560 9635
rect 19622 9259 19656 9635
rect 19718 9259 19752 9635
rect 19814 9259 19848 9635
rect 19910 9259 19944 9635
rect 20006 9259 20040 9635
rect 20102 9259 20136 9635
rect 20198 9259 20232 9635
rect 20294 9259 20328 9635
rect 20390 9259 20424 9635
rect 20486 9259 20520 9635
rect 20582 9259 20616 9635
rect 20678 9259 20712 9635
rect 20774 9259 20808 9635
rect 20870 9259 20904 9635
rect 20966 9259 21000 9635
rect 21062 9259 21096 9635
rect 21158 9259 21192 9635
rect 21254 9259 21288 9635
rect 21350 9259 21384 9635
rect 21446 9259 21480 9635
rect 19574 9166 19608 9200
rect 19766 9166 19800 9200
rect 19958 9166 19992 9200
rect 20150 9166 20184 9200
rect 20342 9166 20376 9200
rect 20534 9166 20568 9200
rect 20726 9166 20760 9200
rect 20918 9166 20952 9200
rect 21110 9166 21144 9200
rect 21302 9166 21336 9200
rect 19574 8734 19608 8768
rect 19766 8734 19800 8768
rect 19958 8734 19992 8768
rect 20150 8734 20184 8768
rect 20342 8734 20376 8768
rect 20534 8734 20568 8768
rect 20726 8734 20760 8768
rect 20918 8734 20952 8768
rect 21110 8734 21144 8768
rect 21302 8734 21336 8768
rect 19526 8308 19560 8684
rect 19622 8308 19656 8684
rect 19718 8308 19752 8684
rect 19814 8308 19848 8684
rect 19910 8308 19944 8684
rect 20006 8308 20040 8684
rect 20102 8308 20136 8684
rect 20198 8308 20232 8684
rect 20294 8308 20328 8684
rect 20390 8308 20424 8684
rect 20486 8308 20520 8684
rect 20582 8308 20616 8684
rect 20678 8308 20712 8684
rect 20774 8308 20808 8684
rect 20870 8308 20904 8684
rect 20966 8308 21000 8684
rect 21062 8308 21096 8684
rect 21158 8308 21192 8684
rect 21254 8308 21288 8684
rect 21350 8308 21384 8684
rect 21446 8308 21480 8684
rect 19670 8224 19704 8258
rect 19862 8224 19896 8258
rect 20054 8224 20088 8258
rect 20246 8224 20280 8258
rect 20438 8224 20472 8258
rect 20630 8224 20664 8258
rect 20822 8224 20856 8258
rect 21014 8224 21048 8258
rect 21206 8224 21240 8258
rect 21398 8224 21432 8258
rect 19670 8116 19704 8150
rect 19862 8116 19896 8150
rect 20054 8116 20088 8150
rect 20246 8116 20280 8150
rect 20438 8116 20472 8150
rect 20630 8116 20664 8150
rect 20822 8116 20856 8150
rect 21014 8116 21048 8150
rect 21206 8116 21240 8150
rect 21398 8116 21432 8150
rect 19526 7690 19560 8066
rect 19622 7690 19656 8066
rect 19718 7690 19752 8066
rect 19814 7690 19848 8066
rect 19910 7690 19944 8066
rect 20006 7690 20040 8066
rect 20102 7690 20136 8066
rect 20198 7690 20232 8066
rect 20294 7690 20328 8066
rect 20390 7690 20424 8066
rect 20486 7690 20520 8066
rect 20582 7690 20616 8066
rect 20678 7690 20712 8066
rect 20774 7690 20808 8066
rect 20870 7690 20904 8066
rect 20966 7690 21000 8066
rect 21062 7690 21096 8066
rect 21158 7690 21192 8066
rect 21254 7690 21288 8066
rect 21350 7690 21384 8066
rect 21446 7690 21480 8066
rect 19574 7606 19608 7640
rect 19766 7606 19800 7640
rect 19958 7606 19992 7640
rect 20150 7606 20184 7640
rect 20342 7606 20376 7640
rect 20534 7606 20568 7640
rect 20726 7606 20760 7640
rect 20918 7606 20952 7640
rect 21110 7606 21144 7640
rect 21302 7606 21336 7640
rect 14770 5912 14804 5946
rect 14962 5912 14996 5946
rect 15154 5912 15188 5946
rect 15346 5912 15380 5946
rect 15538 5912 15572 5946
rect 14626 5486 14660 5862
rect 14722 5486 14756 5862
rect 14818 5486 14852 5862
rect 14914 5486 14948 5862
rect 15010 5486 15044 5862
rect 15106 5486 15140 5862
rect 15202 5486 15236 5862
rect 15298 5486 15332 5862
rect 15394 5486 15428 5862
rect 15490 5486 15524 5862
rect 15586 5486 15620 5862
rect 14674 5402 14708 5436
rect 14866 5402 14900 5436
rect 15058 5402 15092 5436
rect 15250 5402 15284 5436
rect 15442 5402 15476 5436
rect 14674 5294 14708 5328
rect 14866 5294 14900 5328
rect 15058 5294 15092 5328
rect 15250 5294 15284 5328
rect 15442 5294 15476 5328
rect 14626 4868 14660 5244
rect 14722 4868 14756 5244
rect 14818 4868 14852 5244
rect 14914 4868 14948 5244
rect 15010 4868 15044 5244
rect 15106 4868 15140 5244
rect 15202 4868 15236 5244
rect 15298 4868 15332 5244
rect 15394 4868 15428 5244
rect 15490 4868 15524 5244
rect 15586 4868 15620 5244
rect 14770 4784 14804 4818
rect 14962 4784 14996 4818
rect 15154 4784 15188 4818
rect 15346 4784 15380 4818
rect 15538 4784 15572 4818
rect 14770 4676 14804 4710
rect 14962 4676 14996 4710
rect 15154 4676 15188 4710
rect 15346 4676 15380 4710
rect 15538 4676 15572 4710
rect 14626 4250 14660 4626
rect 14722 4250 14756 4626
rect 14818 4250 14852 4626
rect 14914 4250 14948 4626
rect 15010 4250 15044 4626
rect 15106 4250 15140 4626
rect 15202 4250 15236 4626
rect 15298 4250 15332 4626
rect 15394 4250 15428 4626
rect 15490 4250 15524 4626
rect 15586 4250 15620 4626
rect 14674 4166 14708 4200
rect 14866 4166 14900 4200
rect 15058 4166 15092 4200
rect 15250 4166 15284 4200
rect 15442 4166 15476 4200
rect 16570 5912 16604 5946
rect 16762 5912 16796 5946
rect 16954 5912 16988 5946
rect 17146 5912 17180 5946
rect 17338 5912 17372 5946
rect 16426 5486 16460 5862
rect 16522 5486 16556 5862
rect 16618 5486 16652 5862
rect 16714 5486 16748 5862
rect 16810 5486 16844 5862
rect 16906 5486 16940 5862
rect 17002 5486 17036 5862
rect 17098 5486 17132 5862
rect 17194 5486 17228 5862
rect 17290 5486 17324 5862
rect 17386 5486 17420 5862
rect 16474 5402 16508 5436
rect 16666 5402 16700 5436
rect 16858 5402 16892 5436
rect 17050 5402 17084 5436
rect 17242 5402 17276 5436
rect 16474 5294 16508 5328
rect 16666 5294 16700 5328
rect 16858 5294 16892 5328
rect 17050 5294 17084 5328
rect 17242 5294 17276 5328
rect 16426 4868 16460 5244
rect 16522 4868 16556 5244
rect 16618 4868 16652 5244
rect 16714 4868 16748 5244
rect 16810 4868 16844 5244
rect 16906 4868 16940 5244
rect 17002 4868 17036 5244
rect 17098 4868 17132 5244
rect 17194 4868 17228 5244
rect 17290 4868 17324 5244
rect 17386 4868 17420 5244
rect 16570 4784 16604 4818
rect 16762 4784 16796 4818
rect 16954 4784 16988 4818
rect 17146 4784 17180 4818
rect 17338 4784 17372 4818
rect 16570 4676 16604 4710
rect 16762 4676 16796 4710
rect 16954 4676 16988 4710
rect 17146 4676 17180 4710
rect 17338 4676 17372 4710
rect 16426 4250 16460 4626
rect 16522 4250 16556 4626
rect 16618 4250 16652 4626
rect 16714 4250 16748 4626
rect 16810 4250 16844 4626
rect 16906 4250 16940 4626
rect 17002 4250 17036 4626
rect 17098 4250 17132 4626
rect 17194 4250 17228 4626
rect 17290 4250 17324 4626
rect 17386 4250 17420 4626
rect 16474 4166 16508 4200
rect 16666 4166 16700 4200
rect 16858 4166 16892 4200
rect 17050 4166 17084 4200
rect 17242 4166 17276 4200
rect 18370 5912 18404 5946
rect 18562 5912 18596 5946
rect 18754 5912 18788 5946
rect 18946 5912 18980 5946
rect 19138 5912 19172 5946
rect 18226 5486 18260 5862
rect 18322 5486 18356 5862
rect 18418 5486 18452 5862
rect 18514 5486 18548 5862
rect 18610 5486 18644 5862
rect 18706 5486 18740 5862
rect 18802 5486 18836 5862
rect 18898 5486 18932 5862
rect 18994 5486 19028 5862
rect 19090 5486 19124 5862
rect 19186 5486 19220 5862
rect 18274 5402 18308 5436
rect 18466 5402 18500 5436
rect 18658 5402 18692 5436
rect 18850 5402 18884 5436
rect 19042 5402 19076 5436
rect 18274 5294 18308 5328
rect 18466 5294 18500 5328
rect 18658 5294 18692 5328
rect 18850 5294 18884 5328
rect 19042 5294 19076 5328
rect 18226 4868 18260 5244
rect 18322 4868 18356 5244
rect 18418 4868 18452 5244
rect 18514 4868 18548 5244
rect 18610 4868 18644 5244
rect 18706 4868 18740 5244
rect 18802 4868 18836 5244
rect 18898 4868 18932 5244
rect 18994 4868 19028 5244
rect 19090 4868 19124 5244
rect 19186 4868 19220 5244
rect 18370 4784 18404 4818
rect 18562 4784 18596 4818
rect 18754 4784 18788 4818
rect 18946 4784 18980 4818
rect 19138 4784 19172 4818
rect 18370 4676 18404 4710
rect 18562 4676 18596 4710
rect 18754 4676 18788 4710
rect 18946 4676 18980 4710
rect 19138 4676 19172 4710
rect 18226 4250 18260 4626
rect 18322 4250 18356 4626
rect 18418 4250 18452 4626
rect 18514 4250 18548 4626
rect 18610 4250 18644 4626
rect 18706 4250 18740 4626
rect 18802 4250 18836 4626
rect 18898 4250 18932 4626
rect 18994 4250 19028 4626
rect 19090 4250 19124 4626
rect 19186 4250 19220 4626
rect 18274 4166 18308 4200
rect 18466 4166 18500 4200
rect 18658 4166 18692 4200
rect 18850 4166 18884 4200
rect 19042 4166 19076 4200
rect 20170 5912 20204 5946
rect 20362 5912 20396 5946
rect 20554 5912 20588 5946
rect 20746 5912 20780 5946
rect 20938 5912 20972 5946
rect 20026 5486 20060 5862
rect 20122 5486 20156 5862
rect 20218 5486 20252 5862
rect 20314 5486 20348 5862
rect 20410 5486 20444 5862
rect 20506 5486 20540 5862
rect 20602 5486 20636 5862
rect 20698 5486 20732 5862
rect 20794 5486 20828 5862
rect 20890 5486 20924 5862
rect 20986 5486 21020 5862
rect 20074 5402 20108 5436
rect 20266 5402 20300 5436
rect 20458 5402 20492 5436
rect 20650 5402 20684 5436
rect 20842 5402 20876 5436
rect 20074 5294 20108 5328
rect 20266 5294 20300 5328
rect 20458 5294 20492 5328
rect 20650 5294 20684 5328
rect 20842 5294 20876 5328
rect 20026 4868 20060 5244
rect 20122 4868 20156 5244
rect 20218 4868 20252 5244
rect 20314 4868 20348 5244
rect 20410 4868 20444 5244
rect 20506 4868 20540 5244
rect 20602 4868 20636 5244
rect 20698 4868 20732 5244
rect 20794 4868 20828 5244
rect 20890 4868 20924 5244
rect 20986 4868 21020 5244
rect 20170 4784 20204 4818
rect 20362 4784 20396 4818
rect 20554 4784 20588 4818
rect 20746 4784 20780 4818
rect 20938 4784 20972 4818
rect 20170 4676 20204 4710
rect 20362 4676 20396 4710
rect 20554 4676 20588 4710
rect 20746 4676 20780 4710
rect 20938 4676 20972 4710
rect 20026 4250 20060 4626
rect 20122 4250 20156 4626
rect 20218 4250 20252 4626
rect 20314 4250 20348 4626
rect 20410 4250 20444 4626
rect 20506 4250 20540 4626
rect 20602 4250 20636 4626
rect 20698 4250 20732 4626
rect 20794 4250 20828 4626
rect 20890 4250 20924 4626
rect 20986 4250 21020 4626
rect 20074 4166 20108 4200
rect 20266 4166 20300 4200
rect 20458 4166 20492 4200
rect 20650 4166 20684 4200
rect 20842 4166 20876 4200
rect 22170 10300 22204 10334
rect 22362 10300 22396 10334
rect 22554 10300 22588 10334
rect 22746 10300 22780 10334
rect 22938 10300 22972 10334
rect 23130 10300 23164 10334
rect 23322 10300 23356 10334
rect 23514 10300 23548 10334
rect 23706 10300 23740 10334
rect 23898 10300 23932 10334
rect 22026 9874 22060 10250
rect 22122 9874 22156 10250
rect 22218 9874 22252 10250
rect 22314 9874 22348 10250
rect 22410 9874 22444 10250
rect 22506 9874 22540 10250
rect 22602 9874 22636 10250
rect 22698 9874 22732 10250
rect 22794 9874 22828 10250
rect 22890 9874 22924 10250
rect 22986 9874 23020 10250
rect 23082 9874 23116 10250
rect 23178 9874 23212 10250
rect 23274 9874 23308 10250
rect 23370 9874 23404 10250
rect 23466 9874 23500 10250
rect 23562 9874 23596 10250
rect 23658 9874 23692 10250
rect 23754 9874 23788 10250
rect 23850 9874 23884 10250
rect 23946 9874 23980 10250
rect 22074 9790 22108 9824
rect 22266 9790 22300 9824
rect 22458 9790 22492 9824
rect 22650 9790 22684 9824
rect 22842 9790 22876 9824
rect 23034 9790 23068 9824
rect 23226 9790 23260 9824
rect 23418 9790 23452 9824
rect 23610 9790 23644 9824
rect 23802 9790 23836 9824
rect 22074 9682 22108 9716
rect 22266 9682 22300 9716
rect 22458 9682 22492 9716
rect 22650 9682 22684 9716
rect 22842 9682 22876 9716
rect 23034 9682 23068 9716
rect 23226 9682 23260 9716
rect 23418 9682 23452 9716
rect 23610 9682 23644 9716
rect 23802 9682 23836 9716
rect 22026 9256 22060 9632
rect 22122 9256 22156 9632
rect 22218 9256 22252 9632
rect 22314 9256 22348 9632
rect 22410 9256 22444 9632
rect 22506 9256 22540 9632
rect 22602 9256 22636 9632
rect 22698 9256 22732 9632
rect 22794 9256 22828 9632
rect 22890 9256 22924 9632
rect 22986 9256 23020 9632
rect 23082 9256 23116 9632
rect 23178 9256 23212 9632
rect 23274 9256 23308 9632
rect 23370 9256 23404 9632
rect 23466 9256 23500 9632
rect 23562 9256 23596 9632
rect 23658 9256 23692 9632
rect 23754 9256 23788 9632
rect 23850 9256 23884 9632
rect 23946 9256 23980 9632
rect 22170 9172 22204 9206
rect 22362 9172 22396 9206
rect 22554 9172 22588 9206
rect 22746 9172 22780 9206
rect 22938 9172 22972 9206
rect 23130 9172 23164 9206
rect 23322 9172 23356 9206
rect 23514 9172 23548 9206
rect 23706 9172 23740 9206
rect 23898 9172 23932 9206
rect 22170 9064 22204 9098
rect 22362 9064 22396 9098
rect 22554 9064 22588 9098
rect 22746 9064 22780 9098
rect 22938 9064 22972 9098
rect 23130 9064 23164 9098
rect 23322 9064 23356 9098
rect 23514 9064 23548 9098
rect 23706 9064 23740 9098
rect 23898 9064 23932 9098
rect 22026 8638 22060 9014
rect 22122 8638 22156 9014
rect 22218 8638 22252 9014
rect 22314 8638 22348 9014
rect 22410 8638 22444 9014
rect 22506 8638 22540 9014
rect 22602 8638 22636 9014
rect 22698 8638 22732 9014
rect 22794 8638 22828 9014
rect 22890 8638 22924 9014
rect 22986 8638 23020 9014
rect 23082 8638 23116 9014
rect 23178 8638 23212 9014
rect 23274 8638 23308 9014
rect 23370 8638 23404 9014
rect 23466 8638 23500 9014
rect 23562 8638 23596 9014
rect 23658 8638 23692 9014
rect 23754 8638 23788 9014
rect 23850 8638 23884 9014
rect 23946 8638 23980 9014
rect 22074 8554 22108 8588
rect 22266 8554 22300 8588
rect 22458 8554 22492 8588
rect 22650 8554 22684 8588
rect 22842 8554 22876 8588
rect 23034 8554 23068 8588
rect 23226 8554 23260 8588
rect 23418 8554 23452 8588
rect 23610 8554 23644 8588
rect 23802 8554 23836 8588
rect 22074 8446 22108 8480
rect 22266 8446 22300 8480
rect 22458 8446 22492 8480
rect 22650 8446 22684 8480
rect 22842 8446 22876 8480
rect 23034 8446 23068 8480
rect 23226 8446 23260 8480
rect 23418 8446 23452 8480
rect 23610 8446 23644 8480
rect 23802 8446 23836 8480
rect 22026 8020 22060 8396
rect 22122 8020 22156 8396
rect 22218 8020 22252 8396
rect 22314 8020 22348 8396
rect 22410 8020 22444 8396
rect 22506 8020 22540 8396
rect 22602 8020 22636 8396
rect 22698 8020 22732 8396
rect 22794 8020 22828 8396
rect 22890 8020 22924 8396
rect 22986 8020 23020 8396
rect 23082 8020 23116 8396
rect 23178 8020 23212 8396
rect 23274 8020 23308 8396
rect 23370 8020 23404 8396
rect 23466 8020 23500 8396
rect 23562 8020 23596 8396
rect 23658 8020 23692 8396
rect 23754 8020 23788 8396
rect 23850 8020 23884 8396
rect 23946 8020 23980 8396
rect 22170 7936 22204 7970
rect 22362 7936 22396 7970
rect 22554 7936 22588 7970
rect 22746 7936 22780 7970
rect 22938 7936 22972 7970
rect 23130 7936 23164 7970
rect 23322 7936 23356 7970
rect 23514 7936 23548 7970
rect 23706 7936 23740 7970
rect 23898 7936 23932 7970
rect 22170 7828 22204 7862
rect 22362 7828 22396 7862
rect 22554 7828 22588 7862
rect 22746 7828 22780 7862
rect 22938 7828 22972 7862
rect 23130 7828 23164 7862
rect 23322 7828 23356 7862
rect 23514 7828 23548 7862
rect 23706 7828 23740 7862
rect 23898 7828 23932 7862
rect 22026 7402 22060 7778
rect 22122 7402 22156 7778
rect 22218 7402 22252 7778
rect 22314 7402 22348 7778
rect 22410 7402 22444 7778
rect 22506 7402 22540 7778
rect 22602 7402 22636 7778
rect 22698 7402 22732 7778
rect 22794 7402 22828 7778
rect 22890 7402 22924 7778
rect 22986 7402 23020 7778
rect 23082 7402 23116 7778
rect 23178 7402 23212 7778
rect 23274 7402 23308 7778
rect 23370 7402 23404 7778
rect 23466 7402 23500 7778
rect 23562 7402 23596 7778
rect 23658 7402 23692 7778
rect 23754 7402 23788 7778
rect 23850 7402 23884 7778
rect 23946 7402 23980 7778
rect 22074 7318 22108 7352
rect 22266 7318 22300 7352
rect 22458 7318 22492 7352
rect 22650 7318 22684 7352
rect 22842 7318 22876 7352
rect 23034 7318 23068 7352
rect 23226 7318 23260 7352
rect 23418 7318 23452 7352
rect 23610 7318 23644 7352
rect 23802 7318 23836 7352
rect 22074 7210 22108 7244
rect 22266 7210 22300 7244
rect 22458 7210 22492 7244
rect 22650 7210 22684 7244
rect 22842 7210 22876 7244
rect 23034 7210 23068 7244
rect 23226 7210 23260 7244
rect 23418 7210 23452 7244
rect 23610 7210 23644 7244
rect 23802 7210 23836 7244
rect 22026 6784 22060 7160
rect 22122 6784 22156 7160
rect 22218 6784 22252 7160
rect 22314 6784 22348 7160
rect 22410 6784 22444 7160
rect 22506 6784 22540 7160
rect 22602 6784 22636 7160
rect 22698 6784 22732 7160
rect 22794 6784 22828 7160
rect 22890 6784 22924 7160
rect 22986 6784 23020 7160
rect 23082 6784 23116 7160
rect 23178 6784 23212 7160
rect 23274 6784 23308 7160
rect 23370 6784 23404 7160
rect 23466 6784 23500 7160
rect 23562 6784 23596 7160
rect 23658 6784 23692 7160
rect 23754 6784 23788 7160
rect 23850 6784 23884 7160
rect 23946 6784 23980 7160
rect 22170 6700 22204 6734
rect 22362 6700 22396 6734
rect 22554 6700 22588 6734
rect 22746 6700 22780 6734
rect 22938 6700 22972 6734
rect 23130 6700 23164 6734
rect 23322 6700 23356 6734
rect 23514 6700 23548 6734
rect 23706 6700 23740 6734
rect 23898 6700 23932 6734
rect 22170 6592 22204 6626
rect 22362 6592 22396 6626
rect 22554 6592 22588 6626
rect 22746 6592 22780 6626
rect 22938 6592 22972 6626
rect 23130 6592 23164 6626
rect 23322 6592 23356 6626
rect 23514 6592 23548 6626
rect 23706 6592 23740 6626
rect 23898 6592 23932 6626
rect 22026 6166 22060 6542
rect 22122 6166 22156 6542
rect 22218 6166 22252 6542
rect 22314 6166 22348 6542
rect 22410 6166 22444 6542
rect 22506 6166 22540 6542
rect 22602 6166 22636 6542
rect 22698 6166 22732 6542
rect 22794 6166 22828 6542
rect 22890 6166 22924 6542
rect 22986 6166 23020 6542
rect 23082 6166 23116 6542
rect 23178 6166 23212 6542
rect 23274 6166 23308 6542
rect 23370 6166 23404 6542
rect 23466 6166 23500 6542
rect 23562 6166 23596 6542
rect 23658 6166 23692 6542
rect 23754 6166 23788 6542
rect 23850 6166 23884 6542
rect 23946 6166 23980 6542
rect 22074 6082 22108 6116
rect 22266 6082 22300 6116
rect 22458 6082 22492 6116
rect 22650 6082 22684 6116
rect 22842 6082 22876 6116
rect 23034 6082 23068 6116
rect 23226 6082 23260 6116
rect 23418 6082 23452 6116
rect 23610 6082 23644 6116
rect 23802 6082 23836 6116
rect 22074 5974 22108 6008
rect 22266 5974 22300 6008
rect 22458 5974 22492 6008
rect 22650 5974 22684 6008
rect 22842 5974 22876 6008
rect 23034 5974 23068 6008
rect 23226 5974 23260 6008
rect 23418 5974 23452 6008
rect 23610 5974 23644 6008
rect 23802 5974 23836 6008
rect 22026 5548 22060 5924
rect 22122 5548 22156 5924
rect 22218 5548 22252 5924
rect 22314 5548 22348 5924
rect 22410 5548 22444 5924
rect 22506 5548 22540 5924
rect 22602 5548 22636 5924
rect 22698 5548 22732 5924
rect 22794 5548 22828 5924
rect 22890 5548 22924 5924
rect 22986 5548 23020 5924
rect 23082 5548 23116 5924
rect 23178 5548 23212 5924
rect 23274 5548 23308 5924
rect 23370 5548 23404 5924
rect 23466 5548 23500 5924
rect 23562 5548 23596 5924
rect 23658 5548 23692 5924
rect 23754 5548 23788 5924
rect 23850 5548 23884 5924
rect 23946 5548 23980 5924
rect 22170 5464 22204 5498
rect 22362 5464 22396 5498
rect 22554 5464 22588 5498
rect 22746 5464 22780 5498
rect 22938 5464 22972 5498
rect 23130 5464 23164 5498
rect 23322 5464 23356 5498
rect 23514 5464 23548 5498
rect 23706 5464 23740 5498
rect 23898 5464 23932 5498
rect 22170 5356 22204 5390
rect 22362 5356 22396 5390
rect 22554 5356 22588 5390
rect 22746 5356 22780 5390
rect 22938 5356 22972 5390
rect 23130 5356 23164 5390
rect 23322 5356 23356 5390
rect 23514 5356 23548 5390
rect 23706 5356 23740 5390
rect 23898 5356 23932 5390
rect 22026 4930 22060 5306
rect 22122 4930 22156 5306
rect 22218 4930 22252 5306
rect 22314 4930 22348 5306
rect 22410 4930 22444 5306
rect 22506 4930 22540 5306
rect 22602 4930 22636 5306
rect 22698 4930 22732 5306
rect 22794 4930 22828 5306
rect 22890 4930 22924 5306
rect 22986 4930 23020 5306
rect 23082 4930 23116 5306
rect 23178 4930 23212 5306
rect 23274 4930 23308 5306
rect 23370 4930 23404 5306
rect 23466 4930 23500 5306
rect 23562 4930 23596 5306
rect 23658 4930 23692 5306
rect 23754 4930 23788 5306
rect 23850 4930 23884 5306
rect 23946 4930 23980 5306
rect 22074 4846 22108 4880
rect 22266 4846 22300 4880
rect 22458 4846 22492 4880
rect 22650 4846 22684 4880
rect 22842 4846 22876 4880
rect 23034 4846 23068 4880
rect 23226 4846 23260 4880
rect 23418 4846 23452 4880
rect 23610 4846 23644 4880
rect 23802 4846 23836 4880
rect -8500 348 -8360 508
rect 288 3766 456 3800
rect 546 3766 714 3800
rect 804 3766 972 3800
rect 1062 3766 1230 3800
rect 1320 3766 1488 3800
rect 226 3340 260 3716
rect 484 3340 518 3716
rect 742 3340 776 3716
rect 1000 3340 1034 3716
rect 1258 3340 1292 3716
rect 1516 3340 1550 3716
rect 288 3256 456 3290
rect 546 3256 714 3290
rect 804 3256 972 3290
rect 1062 3256 1230 3290
rect 1320 3256 1488 3290
rect 288 3148 456 3182
rect 546 3148 714 3182
rect 804 3148 972 3182
rect 1062 3148 1230 3182
rect 1320 3148 1488 3182
rect 226 2722 260 3098
rect 484 2722 518 3098
rect 742 2722 776 3098
rect 1000 2722 1034 3098
rect 1258 2722 1292 3098
rect 1516 2722 1550 3098
rect 288 2638 456 2672
rect 546 2638 714 2672
rect 804 2638 972 2672
rect 1062 2638 1230 2672
rect 1320 2638 1488 2672
rect 288 2530 456 2564
rect 546 2530 714 2564
rect 804 2530 972 2564
rect 1062 2530 1230 2564
rect 1320 2530 1488 2564
rect 226 2104 260 2480
rect 484 2104 518 2480
rect 742 2104 776 2480
rect 1000 2104 1034 2480
rect 1258 2104 1292 2480
rect 1516 2104 1550 2480
rect 288 2020 456 2054
rect 546 2020 714 2054
rect 804 2020 972 2054
rect 1062 2020 1230 2054
rect 1320 2020 1488 2054
rect 288 1912 456 1946
rect 546 1912 714 1946
rect 804 1912 972 1946
rect 1062 1912 1230 1946
rect 1320 1912 1488 1946
rect 226 1486 260 1862
rect 484 1486 518 1862
rect 742 1486 776 1862
rect 1000 1486 1034 1862
rect 1258 1486 1292 1862
rect 1516 1486 1550 1862
rect 288 1402 456 1436
rect 546 1402 714 1436
rect 804 1402 972 1436
rect 1062 1402 1230 1436
rect 1320 1402 1488 1436
rect 288 1294 456 1328
rect 546 1294 714 1328
rect 804 1294 972 1328
rect 1062 1294 1230 1328
rect 1320 1294 1488 1328
rect 226 868 260 1244
rect 484 868 518 1244
rect 742 868 776 1244
rect 1000 868 1034 1244
rect 1258 868 1292 1244
rect 1516 868 1550 1244
rect 288 784 456 818
rect 546 784 714 818
rect 804 784 972 818
rect 1062 784 1230 818
rect 1320 784 1488 818
rect 288 676 456 710
rect 546 676 714 710
rect 804 676 972 710
rect 1062 676 1230 710
rect 1320 676 1488 710
rect 226 250 260 626
rect 484 250 518 626
rect 742 250 776 626
rect 1000 250 1034 626
rect 1258 250 1292 626
rect 1516 250 1550 626
rect 288 166 456 200
rect 546 166 714 200
rect 804 166 972 200
rect 1062 166 1230 200
rect 1320 166 1488 200
rect 1696 68 1876 268
rect 2088 3766 2256 3800
rect 2346 3766 2514 3800
rect 2604 3766 2772 3800
rect 2862 3766 3030 3800
rect 3120 3766 3288 3800
rect 2026 3340 2060 3716
rect 2284 3340 2318 3716
rect 2542 3340 2576 3716
rect 2800 3340 2834 3716
rect 3058 3340 3092 3716
rect 3316 3340 3350 3716
rect 2088 3256 2256 3290
rect 2346 3256 2514 3290
rect 2604 3256 2772 3290
rect 2862 3256 3030 3290
rect 3120 3256 3288 3290
rect 2088 3148 2256 3182
rect 2346 3148 2514 3182
rect 2604 3148 2772 3182
rect 2862 3148 3030 3182
rect 3120 3148 3288 3182
rect 2026 2722 2060 3098
rect 2284 2722 2318 3098
rect 2542 2722 2576 3098
rect 2800 2722 2834 3098
rect 3058 2722 3092 3098
rect 3316 2722 3350 3098
rect 2088 2638 2256 2672
rect 2346 2638 2514 2672
rect 2604 2638 2772 2672
rect 2862 2638 3030 2672
rect 3120 2638 3288 2672
rect 2088 2530 2256 2564
rect 2346 2530 2514 2564
rect 2604 2530 2772 2564
rect 2862 2530 3030 2564
rect 3120 2530 3288 2564
rect 2026 2104 2060 2480
rect 2284 2104 2318 2480
rect 2542 2104 2576 2480
rect 2800 2104 2834 2480
rect 3058 2104 3092 2480
rect 3316 2104 3350 2480
rect 2088 2020 2256 2054
rect 2346 2020 2514 2054
rect 2604 2020 2772 2054
rect 2862 2020 3030 2054
rect 3120 2020 3288 2054
rect 2088 1912 2256 1946
rect 2346 1912 2514 1946
rect 2604 1912 2772 1946
rect 2862 1912 3030 1946
rect 3120 1912 3288 1946
rect 2026 1486 2060 1862
rect 2284 1486 2318 1862
rect 2542 1486 2576 1862
rect 2800 1486 2834 1862
rect 3058 1486 3092 1862
rect 3316 1486 3350 1862
rect 2088 1402 2256 1436
rect 2346 1402 2514 1436
rect 2604 1402 2772 1436
rect 2862 1402 3030 1436
rect 3120 1402 3288 1436
rect 2088 1294 2256 1328
rect 2346 1294 2514 1328
rect 2604 1294 2772 1328
rect 2862 1294 3030 1328
rect 3120 1294 3288 1328
rect 2026 868 2060 1244
rect 2284 868 2318 1244
rect 2542 868 2576 1244
rect 2800 868 2834 1244
rect 3058 868 3092 1244
rect 3316 868 3350 1244
rect 2088 784 2256 818
rect 2346 784 2514 818
rect 2604 784 2772 818
rect 2862 784 3030 818
rect 3120 784 3288 818
rect 2088 676 2256 710
rect 2346 676 2514 710
rect 2604 676 2772 710
rect 2862 676 3030 710
rect 3120 676 3288 710
rect 2026 250 2060 626
rect 2284 250 2318 626
rect 2542 250 2576 626
rect 2800 250 2834 626
rect 3058 250 3092 626
rect 3316 250 3350 626
rect 2088 166 2256 200
rect 2346 166 2514 200
rect 2604 166 2772 200
rect 2862 166 3030 200
rect 3120 166 3288 200
rect 3512 64 3692 276
rect 3888 3766 4056 3800
rect 4146 3766 4314 3800
rect 4404 3766 4572 3800
rect 4662 3766 4830 3800
rect 4920 3766 5088 3800
rect 3826 3340 3860 3716
rect 4084 3340 4118 3716
rect 4342 3340 4376 3716
rect 4600 3340 4634 3716
rect 4858 3340 4892 3716
rect 5116 3340 5150 3716
rect 3888 3256 4056 3290
rect 4146 3256 4314 3290
rect 4404 3256 4572 3290
rect 4662 3256 4830 3290
rect 4920 3256 5088 3290
rect 3888 3148 4056 3182
rect 4146 3148 4314 3182
rect 4404 3148 4572 3182
rect 4662 3148 4830 3182
rect 4920 3148 5088 3182
rect 3826 2722 3860 3098
rect 4084 2722 4118 3098
rect 4342 2722 4376 3098
rect 4600 2722 4634 3098
rect 4858 2722 4892 3098
rect 5116 2722 5150 3098
rect 3888 2638 4056 2672
rect 4146 2638 4314 2672
rect 4404 2638 4572 2672
rect 4662 2638 4830 2672
rect 4920 2638 5088 2672
rect 3888 2530 4056 2564
rect 4146 2530 4314 2564
rect 4404 2530 4572 2564
rect 4662 2530 4830 2564
rect 4920 2530 5088 2564
rect 3826 2104 3860 2480
rect 4084 2104 4118 2480
rect 4342 2104 4376 2480
rect 4600 2104 4634 2480
rect 4858 2104 4892 2480
rect 5116 2104 5150 2480
rect 3888 2020 4056 2054
rect 4146 2020 4314 2054
rect 4404 2020 4572 2054
rect 4662 2020 4830 2054
rect 4920 2020 5088 2054
rect 3888 1912 4056 1946
rect 4146 1912 4314 1946
rect 4404 1912 4572 1946
rect 4662 1912 4830 1946
rect 4920 1912 5088 1946
rect 3826 1486 3860 1862
rect 4084 1486 4118 1862
rect 4342 1486 4376 1862
rect 4600 1486 4634 1862
rect 4858 1486 4892 1862
rect 5116 1486 5150 1862
rect 3888 1402 4056 1436
rect 4146 1402 4314 1436
rect 4404 1402 4572 1436
rect 4662 1402 4830 1436
rect 4920 1402 5088 1436
rect 3888 1294 4056 1328
rect 4146 1294 4314 1328
rect 4404 1294 4572 1328
rect 4662 1294 4830 1328
rect 4920 1294 5088 1328
rect 3826 868 3860 1244
rect 4084 868 4118 1244
rect 4342 868 4376 1244
rect 4600 868 4634 1244
rect 4858 868 4892 1244
rect 5116 868 5150 1244
rect 3888 784 4056 818
rect 4146 784 4314 818
rect 4404 784 4572 818
rect 4662 784 4830 818
rect 4920 784 5088 818
rect 3888 676 4056 710
rect 4146 676 4314 710
rect 4404 676 4572 710
rect 4662 676 4830 710
rect 4920 676 5088 710
rect 3826 250 3860 626
rect 4084 250 4118 626
rect 4342 250 4376 626
rect 4600 250 4634 626
rect 4858 250 4892 626
rect 5116 250 5150 626
rect 3888 166 4056 200
rect 4146 166 4314 200
rect 4404 166 4572 200
rect 4662 166 4830 200
rect 4920 166 5088 200
rect 5288 64 5468 276
rect 5688 3766 5856 3800
rect 5946 3766 6114 3800
rect 6204 3766 6372 3800
rect 6462 3766 6630 3800
rect 6720 3766 6888 3800
rect 5626 3340 5660 3716
rect 5884 3340 5918 3716
rect 6142 3340 6176 3716
rect 6400 3340 6434 3716
rect 6658 3340 6692 3716
rect 6916 3340 6950 3716
rect 5688 3256 5856 3290
rect 5946 3256 6114 3290
rect 6204 3256 6372 3290
rect 6462 3256 6630 3290
rect 6720 3256 6888 3290
rect 5688 3148 5856 3182
rect 5946 3148 6114 3182
rect 6204 3148 6372 3182
rect 6462 3148 6630 3182
rect 6720 3148 6888 3182
rect 5626 2722 5660 3098
rect 5884 2722 5918 3098
rect 6142 2722 6176 3098
rect 6400 2722 6434 3098
rect 6658 2722 6692 3098
rect 6916 2722 6950 3098
rect 5688 2638 5856 2672
rect 5946 2638 6114 2672
rect 6204 2638 6372 2672
rect 6462 2638 6630 2672
rect 6720 2638 6888 2672
rect 5688 2530 5856 2564
rect 5946 2530 6114 2564
rect 6204 2530 6372 2564
rect 6462 2530 6630 2564
rect 6720 2530 6888 2564
rect 5626 2104 5660 2480
rect 5884 2104 5918 2480
rect 6142 2104 6176 2480
rect 6400 2104 6434 2480
rect 6658 2104 6692 2480
rect 6916 2104 6950 2480
rect 5688 2020 5856 2054
rect 5946 2020 6114 2054
rect 6204 2020 6372 2054
rect 6462 2020 6630 2054
rect 6720 2020 6888 2054
rect 5688 1912 5856 1946
rect 5946 1912 6114 1946
rect 6204 1912 6372 1946
rect 6462 1912 6630 1946
rect 6720 1912 6888 1946
rect 5626 1486 5660 1862
rect 5884 1486 5918 1862
rect 6142 1486 6176 1862
rect 6400 1486 6434 1862
rect 6658 1486 6692 1862
rect 6916 1486 6950 1862
rect 5688 1402 5856 1436
rect 5946 1402 6114 1436
rect 6204 1402 6372 1436
rect 6462 1402 6630 1436
rect 6720 1402 6888 1436
rect 5688 1294 5856 1328
rect 5946 1294 6114 1328
rect 6204 1294 6372 1328
rect 6462 1294 6630 1328
rect 6720 1294 6888 1328
rect 5626 868 5660 1244
rect 5884 868 5918 1244
rect 6142 868 6176 1244
rect 6400 868 6434 1244
rect 6658 868 6692 1244
rect 6916 868 6950 1244
rect 5688 784 5856 818
rect 5946 784 6114 818
rect 6204 784 6372 818
rect 6462 784 6630 818
rect 6720 784 6888 818
rect 5688 676 5856 710
rect 5946 676 6114 710
rect 6204 676 6372 710
rect 6462 676 6630 710
rect 6720 676 6888 710
rect 5626 250 5660 626
rect 5884 250 5918 626
rect 6142 250 6176 626
rect 6400 250 6434 626
rect 6658 250 6692 626
rect 6916 250 6950 626
rect 5688 166 5856 200
rect 5946 166 6114 200
rect 6204 166 6372 200
rect 6462 166 6630 200
rect 6720 166 6888 200
rect 14688 3766 14856 3800
rect 14946 3766 15114 3800
rect 15204 3766 15372 3800
rect 15462 3766 15630 3800
rect 15720 3766 15888 3800
rect 14626 3340 14660 3716
rect 14884 3340 14918 3716
rect 15142 3340 15176 3716
rect 15400 3340 15434 3716
rect 15658 3340 15692 3716
rect 15916 3340 15950 3716
rect 14688 3256 14856 3290
rect 14946 3256 15114 3290
rect 15204 3256 15372 3290
rect 15462 3256 15630 3290
rect 15720 3256 15888 3290
rect 14688 3148 14856 3182
rect 14946 3148 15114 3182
rect 15204 3148 15372 3182
rect 15462 3148 15630 3182
rect 15720 3148 15888 3182
rect 14626 2722 14660 3098
rect 14884 2722 14918 3098
rect 15142 2722 15176 3098
rect 15400 2722 15434 3098
rect 15658 2722 15692 3098
rect 15916 2722 15950 3098
rect 14688 2638 14856 2672
rect 14946 2638 15114 2672
rect 15204 2638 15372 2672
rect 15462 2638 15630 2672
rect 15720 2638 15888 2672
rect 14688 2530 14856 2564
rect 14946 2530 15114 2564
rect 15204 2530 15372 2564
rect 15462 2530 15630 2564
rect 15720 2530 15888 2564
rect 14626 2104 14660 2480
rect 14884 2104 14918 2480
rect 15142 2104 15176 2480
rect 15400 2104 15434 2480
rect 15658 2104 15692 2480
rect 15916 2104 15950 2480
rect 14688 2020 14856 2054
rect 14946 2020 15114 2054
rect 15204 2020 15372 2054
rect 15462 2020 15630 2054
rect 15720 2020 15888 2054
rect 14688 1912 14856 1946
rect 14946 1912 15114 1946
rect 15204 1912 15372 1946
rect 15462 1912 15630 1946
rect 15720 1912 15888 1946
rect 14626 1486 14660 1862
rect 14884 1486 14918 1862
rect 15142 1486 15176 1862
rect 15400 1486 15434 1862
rect 15658 1486 15692 1862
rect 15916 1486 15950 1862
rect 14688 1402 14856 1436
rect 14946 1402 15114 1436
rect 15204 1402 15372 1436
rect 15462 1402 15630 1436
rect 15720 1402 15888 1436
rect 14688 1294 14856 1328
rect 14946 1294 15114 1328
rect 15204 1294 15372 1328
rect 15462 1294 15630 1328
rect 15720 1294 15888 1328
rect 14626 868 14660 1244
rect 14884 868 14918 1244
rect 15142 868 15176 1244
rect 15400 868 15434 1244
rect 15658 868 15692 1244
rect 15916 868 15950 1244
rect 14688 784 14856 818
rect 14946 784 15114 818
rect 15204 784 15372 818
rect 15462 784 15630 818
rect 15720 784 15888 818
rect 14688 676 14856 710
rect 14946 676 15114 710
rect 15204 676 15372 710
rect 15462 676 15630 710
rect 15720 676 15888 710
rect 14626 250 14660 626
rect 14884 250 14918 626
rect 15142 250 15176 626
rect 15400 250 15434 626
rect 15658 250 15692 626
rect 15916 250 15950 626
rect 14688 166 14856 200
rect 14946 166 15114 200
rect 15204 166 15372 200
rect 15462 166 15630 200
rect 15720 166 15888 200
rect 16096 68 16276 268
rect 16488 3766 16656 3800
rect 16746 3766 16914 3800
rect 17004 3766 17172 3800
rect 17262 3766 17430 3800
rect 17520 3766 17688 3800
rect 16426 3340 16460 3716
rect 16684 3340 16718 3716
rect 16942 3340 16976 3716
rect 17200 3340 17234 3716
rect 17458 3340 17492 3716
rect 17716 3340 17750 3716
rect 16488 3256 16656 3290
rect 16746 3256 16914 3290
rect 17004 3256 17172 3290
rect 17262 3256 17430 3290
rect 17520 3256 17688 3290
rect 16488 3148 16656 3182
rect 16746 3148 16914 3182
rect 17004 3148 17172 3182
rect 17262 3148 17430 3182
rect 17520 3148 17688 3182
rect 16426 2722 16460 3098
rect 16684 2722 16718 3098
rect 16942 2722 16976 3098
rect 17200 2722 17234 3098
rect 17458 2722 17492 3098
rect 17716 2722 17750 3098
rect 16488 2638 16656 2672
rect 16746 2638 16914 2672
rect 17004 2638 17172 2672
rect 17262 2638 17430 2672
rect 17520 2638 17688 2672
rect 16488 2530 16656 2564
rect 16746 2530 16914 2564
rect 17004 2530 17172 2564
rect 17262 2530 17430 2564
rect 17520 2530 17688 2564
rect 16426 2104 16460 2480
rect 16684 2104 16718 2480
rect 16942 2104 16976 2480
rect 17200 2104 17234 2480
rect 17458 2104 17492 2480
rect 17716 2104 17750 2480
rect 16488 2020 16656 2054
rect 16746 2020 16914 2054
rect 17004 2020 17172 2054
rect 17262 2020 17430 2054
rect 17520 2020 17688 2054
rect 16488 1912 16656 1946
rect 16746 1912 16914 1946
rect 17004 1912 17172 1946
rect 17262 1912 17430 1946
rect 17520 1912 17688 1946
rect 16426 1486 16460 1862
rect 16684 1486 16718 1862
rect 16942 1486 16976 1862
rect 17200 1486 17234 1862
rect 17458 1486 17492 1862
rect 17716 1486 17750 1862
rect 16488 1402 16656 1436
rect 16746 1402 16914 1436
rect 17004 1402 17172 1436
rect 17262 1402 17430 1436
rect 17520 1402 17688 1436
rect 16488 1294 16656 1328
rect 16746 1294 16914 1328
rect 17004 1294 17172 1328
rect 17262 1294 17430 1328
rect 17520 1294 17688 1328
rect 16426 868 16460 1244
rect 16684 868 16718 1244
rect 16942 868 16976 1244
rect 17200 868 17234 1244
rect 17458 868 17492 1244
rect 17716 868 17750 1244
rect 16488 784 16656 818
rect 16746 784 16914 818
rect 17004 784 17172 818
rect 17262 784 17430 818
rect 17520 784 17688 818
rect 16488 676 16656 710
rect 16746 676 16914 710
rect 17004 676 17172 710
rect 17262 676 17430 710
rect 17520 676 17688 710
rect 16426 250 16460 626
rect 16684 250 16718 626
rect 16942 250 16976 626
rect 17200 250 17234 626
rect 17458 250 17492 626
rect 17716 250 17750 626
rect 16488 166 16656 200
rect 16746 166 16914 200
rect 17004 166 17172 200
rect 17262 166 17430 200
rect 17520 166 17688 200
rect 17912 64 18092 276
rect 18288 3766 18456 3800
rect 18546 3766 18714 3800
rect 18804 3766 18972 3800
rect 19062 3766 19230 3800
rect 19320 3766 19488 3800
rect 18226 3340 18260 3716
rect 18484 3340 18518 3716
rect 18742 3340 18776 3716
rect 19000 3340 19034 3716
rect 19258 3340 19292 3716
rect 19516 3340 19550 3716
rect 18288 3256 18456 3290
rect 18546 3256 18714 3290
rect 18804 3256 18972 3290
rect 19062 3256 19230 3290
rect 19320 3256 19488 3290
rect 18288 3148 18456 3182
rect 18546 3148 18714 3182
rect 18804 3148 18972 3182
rect 19062 3148 19230 3182
rect 19320 3148 19488 3182
rect 18226 2722 18260 3098
rect 18484 2722 18518 3098
rect 18742 2722 18776 3098
rect 19000 2722 19034 3098
rect 19258 2722 19292 3098
rect 19516 2722 19550 3098
rect 18288 2638 18456 2672
rect 18546 2638 18714 2672
rect 18804 2638 18972 2672
rect 19062 2638 19230 2672
rect 19320 2638 19488 2672
rect 18288 2530 18456 2564
rect 18546 2530 18714 2564
rect 18804 2530 18972 2564
rect 19062 2530 19230 2564
rect 19320 2530 19488 2564
rect 18226 2104 18260 2480
rect 18484 2104 18518 2480
rect 18742 2104 18776 2480
rect 19000 2104 19034 2480
rect 19258 2104 19292 2480
rect 19516 2104 19550 2480
rect 18288 2020 18456 2054
rect 18546 2020 18714 2054
rect 18804 2020 18972 2054
rect 19062 2020 19230 2054
rect 19320 2020 19488 2054
rect 18288 1912 18456 1946
rect 18546 1912 18714 1946
rect 18804 1912 18972 1946
rect 19062 1912 19230 1946
rect 19320 1912 19488 1946
rect 18226 1486 18260 1862
rect 18484 1486 18518 1862
rect 18742 1486 18776 1862
rect 19000 1486 19034 1862
rect 19258 1486 19292 1862
rect 19516 1486 19550 1862
rect 18288 1402 18456 1436
rect 18546 1402 18714 1436
rect 18804 1402 18972 1436
rect 19062 1402 19230 1436
rect 19320 1402 19488 1436
rect 18288 1294 18456 1328
rect 18546 1294 18714 1328
rect 18804 1294 18972 1328
rect 19062 1294 19230 1328
rect 19320 1294 19488 1328
rect 18226 868 18260 1244
rect 18484 868 18518 1244
rect 18742 868 18776 1244
rect 19000 868 19034 1244
rect 19258 868 19292 1244
rect 19516 868 19550 1244
rect 18288 784 18456 818
rect 18546 784 18714 818
rect 18804 784 18972 818
rect 19062 784 19230 818
rect 19320 784 19488 818
rect 18288 676 18456 710
rect 18546 676 18714 710
rect 18804 676 18972 710
rect 19062 676 19230 710
rect 19320 676 19488 710
rect 18226 250 18260 626
rect 18484 250 18518 626
rect 18742 250 18776 626
rect 19000 250 19034 626
rect 19258 250 19292 626
rect 19516 250 19550 626
rect 18288 166 18456 200
rect 18546 166 18714 200
rect 18804 166 18972 200
rect 19062 166 19230 200
rect 19320 166 19488 200
rect 19688 64 19868 276
rect 20088 3766 20256 3800
rect 20346 3766 20514 3800
rect 20604 3766 20772 3800
rect 20862 3766 21030 3800
rect 21120 3766 21288 3800
rect 20026 3340 20060 3716
rect 20284 3340 20318 3716
rect 20542 3340 20576 3716
rect 20800 3340 20834 3716
rect 21058 3340 21092 3716
rect 21316 3340 21350 3716
rect 20088 3256 20256 3290
rect 20346 3256 20514 3290
rect 20604 3256 20772 3290
rect 20862 3256 21030 3290
rect 21120 3256 21288 3290
rect 20088 3148 20256 3182
rect 20346 3148 20514 3182
rect 20604 3148 20772 3182
rect 20862 3148 21030 3182
rect 21120 3148 21288 3182
rect 20026 2722 20060 3098
rect 20284 2722 20318 3098
rect 20542 2722 20576 3098
rect 20800 2722 20834 3098
rect 21058 2722 21092 3098
rect 21316 2722 21350 3098
rect 20088 2638 20256 2672
rect 20346 2638 20514 2672
rect 20604 2638 20772 2672
rect 20862 2638 21030 2672
rect 21120 2638 21288 2672
rect 20088 2530 20256 2564
rect 20346 2530 20514 2564
rect 20604 2530 20772 2564
rect 20862 2530 21030 2564
rect 21120 2530 21288 2564
rect 20026 2104 20060 2480
rect 20284 2104 20318 2480
rect 20542 2104 20576 2480
rect 20800 2104 20834 2480
rect 21058 2104 21092 2480
rect 21316 2104 21350 2480
rect 20088 2020 20256 2054
rect 20346 2020 20514 2054
rect 20604 2020 20772 2054
rect 20862 2020 21030 2054
rect 21120 2020 21288 2054
rect 20088 1912 20256 1946
rect 20346 1912 20514 1946
rect 20604 1912 20772 1946
rect 20862 1912 21030 1946
rect 21120 1912 21288 1946
rect 20026 1486 20060 1862
rect 20284 1486 20318 1862
rect 20542 1486 20576 1862
rect 20800 1486 20834 1862
rect 21058 1486 21092 1862
rect 21316 1486 21350 1862
rect 20088 1402 20256 1436
rect 20346 1402 20514 1436
rect 20604 1402 20772 1436
rect 20862 1402 21030 1436
rect 21120 1402 21288 1436
rect 20088 1294 20256 1328
rect 20346 1294 20514 1328
rect 20604 1294 20772 1328
rect 20862 1294 21030 1328
rect 21120 1294 21288 1328
rect 20026 868 20060 1244
rect 20284 868 20318 1244
rect 20542 868 20576 1244
rect 20800 868 20834 1244
rect 21058 868 21092 1244
rect 21316 868 21350 1244
rect 20088 784 20256 818
rect 20346 784 20514 818
rect 20604 784 20772 818
rect 20862 784 21030 818
rect 21120 784 21288 818
rect 20088 676 20256 710
rect 20346 676 20514 710
rect 20604 676 20772 710
rect 20862 676 21030 710
rect 21120 676 21288 710
rect 20026 250 20060 626
rect 20284 250 20318 626
rect 20542 250 20576 626
rect 20800 250 20834 626
rect 21058 250 21092 626
rect 21316 250 21350 626
rect 20088 166 20256 200
rect 20346 166 20514 200
rect 20604 166 20772 200
rect 20862 166 21030 200
rect 21120 166 21288 200
<< metal1 >>
rect 7428 27436 7552 27442
rect 7428 27336 7440 27436
rect 7540 27336 7552 27436
rect 7428 27330 7552 27336
rect 6488 27168 8364 27232
rect 6488 27134 6552 27168
rect 6620 27134 6710 27168
rect 6778 27134 6868 27168
rect 6936 27134 7026 27168
rect 7094 27134 7184 27168
rect 7252 27134 7342 27168
rect 7410 27134 7500 27168
rect 7568 27134 7658 27168
rect 7726 27134 7816 27168
rect 7884 27134 7974 27168
rect 8042 27134 8364 27168
rect 6488 27124 8364 27134
rect 8708 27168 10584 27232
rect 8708 27134 8772 27168
rect 8840 27134 8930 27168
rect 8998 27134 9088 27168
rect 9156 27134 9246 27168
rect 9314 27134 9404 27168
rect 9472 27134 9562 27168
rect 9630 27134 9720 27168
rect 9788 27134 9878 27168
rect 9946 27134 10036 27168
rect 10104 27134 10194 27168
rect 10262 27134 10584 27168
rect 8708 27124 10584 27134
rect 10888 27168 12764 27232
rect 10888 27134 10952 27168
rect 11020 27134 11110 27168
rect 11178 27134 11268 27168
rect 11336 27134 11426 27168
rect 11494 27134 11584 27168
rect 11652 27134 11742 27168
rect 11810 27134 11900 27168
rect 11968 27134 12058 27168
rect 12126 27134 12216 27168
rect 12284 27134 12374 27168
rect 12442 27134 12764 27168
rect 10888 27124 12764 27134
rect 13068 27168 14944 27232
rect 13068 27134 13132 27168
rect 13200 27134 13290 27168
rect 13358 27134 13448 27168
rect 13516 27134 13606 27168
rect 13674 27134 13764 27168
rect 13832 27134 13922 27168
rect 13990 27134 14080 27168
rect 14148 27134 14238 27168
rect 14306 27134 14396 27168
rect 14464 27134 14554 27168
rect 14622 27134 14944 27168
rect 13068 27124 14944 27134
rect 15268 27168 17144 27232
rect 15268 27134 15332 27168
rect 15400 27134 15490 27168
rect 15558 27134 15648 27168
rect 15716 27134 15806 27168
rect 15874 27134 15964 27168
rect 16032 27134 16122 27168
rect 16190 27134 16280 27168
rect 16348 27134 16438 27168
rect 16506 27134 16596 27168
rect 16664 27134 16754 27168
rect 16822 27134 17144 27168
rect 15268 27124 17144 27134
rect 6484 27075 6530 27087
rect 6484 26868 6490 27075
rect 6524 26868 6530 27075
rect 6622 26912 6632 27092
rect 6696 26912 6706 27092
rect 6800 27075 6846 27087
rect 6466 26688 6476 26868
rect 6540 26688 6550 26868
rect 6642 26699 6648 26912
rect 6682 26699 6688 26912
rect 6800 26868 6806 27075
rect 6840 26868 6846 27075
rect 6938 26912 6948 27092
rect 7012 26912 7022 27092
rect 7116 27075 7162 27087
rect 6484 26687 6530 26688
rect 6642 26687 6688 26699
rect 6782 26688 6792 26868
rect 6856 26688 6866 26868
rect 6958 26699 6964 26912
rect 6998 26699 7004 26912
rect 7116 26868 7122 27075
rect 7156 26868 7162 27075
rect 7254 26912 7264 27092
rect 7328 26912 7338 27092
rect 7432 27075 7478 27087
rect 6800 26687 6846 26688
rect 6958 26687 7004 26699
rect 7098 26688 7108 26868
rect 7172 26688 7182 26868
rect 7274 26699 7280 26912
rect 7314 26699 7320 26912
rect 7432 26868 7438 27075
rect 7472 26868 7478 27075
rect 7570 26912 7580 27092
rect 7644 26912 7654 27092
rect 7748 27075 7794 27087
rect 7116 26687 7162 26688
rect 7274 26687 7320 26699
rect 7414 26688 7424 26868
rect 7488 26688 7498 26868
rect 7590 26699 7596 26912
rect 7630 26699 7636 26912
rect 7748 26868 7754 27075
rect 7788 26868 7794 27075
rect 7886 26912 7896 27092
rect 7960 26912 7970 27092
rect 8064 27075 8110 27087
rect 7432 26687 7478 26688
rect 7590 26687 7636 26699
rect 7730 26688 7740 26868
rect 7804 26688 7814 26868
rect 7906 26699 7912 26912
rect 7946 26699 7952 26912
rect 8064 26868 8070 27075
rect 8104 26868 8110 27075
rect 7748 26687 7794 26688
rect 7906 26687 7952 26699
rect 8046 26688 8056 26868
rect 8120 26688 8130 26868
rect 8064 26687 8110 26688
rect 8160 26656 8364 27124
rect 8704 27075 8750 27087
rect 8704 26868 8710 27075
rect 8744 26868 8750 27075
rect 8842 26912 8852 27092
rect 8916 26912 8926 27092
rect 9020 27075 9066 27087
rect 8686 26688 8696 26868
rect 8760 26688 8770 26868
rect 8862 26699 8868 26912
rect 8902 26699 8908 26912
rect 9020 26868 9026 27075
rect 9060 26868 9066 27075
rect 9158 26912 9168 27092
rect 9232 26912 9242 27092
rect 9336 27075 9382 27087
rect 8704 26687 8750 26688
rect 8862 26687 8908 26699
rect 9002 26688 9012 26868
rect 9076 26688 9086 26868
rect 9178 26699 9184 26912
rect 9218 26699 9224 26912
rect 9336 26868 9342 27075
rect 9376 26868 9382 27075
rect 9474 26912 9484 27092
rect 9548 26912 9558 27092
rect 9652 27075 9698 27087
rect 9020 26687 9066 26688
rect 9178 26687 9224 26699
rect 9318 26688 9328 26868
rect 9392 26688 9402 26868
rect 9494 26699 9500 26912
rect 9534 26699 9540 26912
rect 9652 26868 9658 27075
rect 9692 26868 9698 27075
rect 9790 26912 9800 27092
rect 9864 26912 9874 27092
rect 9968 27075 10014 27087
rect 9336 26687 9382 26688
rect 9494 26687 9540 26699
rect 9634 26688 9644 26868
rect 9708 26688 9718 26868
rect 9810 26699 9816 26912
rect 9850 26699 9856 26912
rect 9968 26868 9974 27075
rect 10008 26868 10014 27075
rect 10106 26912 10116 27092
rect 10180 26912 10190 27092
rect 10284 27075 10330 27087
rect 9652 26687 9698 26688
rect 9810 26687 9856 26699
rect 9950 26688 9960 26868
rect 10024 26688 10034 26868
rect 10126 26699 10132 26912
rect 10166 26699 10172 26912
rect 10284 26868 10290 27075
rect 10324 26868 10330 27075
rect 9968 26687 10014 26688
rect 10126 26687 10172 26699
rect 10266 26688 10276 26868
rect 10340 26688 10350 26868
rect 10284 26687 10330 26688
rect 10380 26656 10584 27124
rect 10884 27075 10930 27087
rect 10884 26868 10890 27075
rect 10924 26868 10930 27075
rect 11022 26912 11032 27092
rect 11096 26912 11106 27092
rect 11200 27075 11246 27087
rect 10866 26688 10876 26868
rect 10940 26688 10950 26868
rect 11042 26699 11048 26912
rect 11082 26699 11088 26912
rect 11200 26868 11206 27075
rect 11240 26868 11246 27075
rect 11338 26912 11348 27092
rect 11412 26912 11422 27092
rect 11516 27075 11562 27087
rect 10884 26687 10930 26688
rect 11042 26687 11088 26699
rect 11182 26688 11192 26868
rect 11256 26688 11266 26868
rect 11358 26699 11364 26912
rect 11398 26699 11404 26912
rect 11516 26868 11522 27075
rect 11556 26868 11562 27075
rect 11654 26912 11664 27092
rect 11728 26912 11738 27092
rect 11832 27075 11878 27087
rect 11200 26687 11246 26688
rect 11358 26687 11404 26699
rect 11498 26688 11508 26868
rect 11572 26688 11582 26868
rect 11674 26699 11680 26912
rect 11714 26699 11720 26912
rect 11832 26868 11838 27075
rect 11872 26868 11878 27075
rect 11970 26912 11980 27092
rect 12044 26912 12054 27092
rect 12148 27075 12194 27087
rect 11516 26687 11562 26688
rect 11674 26687 11720 26699
rect 11814 26688 11824 26868
rect 11888 26688 11898 26868
rect 11990 26699 11996 26912
rect 12030 26699 12036 26912
rect 12148 26868 12154 27075
rect 12188 26868 12194 27075
rect 12286 26912 12296 27092
rect 12360 26912 12370 27092
rect 12464 27075 12510 27087
rect 11832 26687 11878 26688
rect 11990 26687 12036 26699
rect 12130 26688 12140 26868
rect 12204 26688 12214 26868
rect 12306 26699 12312 26912
rect 12346 26699 12352 26912
rect 12464 26868 12470 27075
rect 12504 26868 12510 27075
rect 12148 26687 12194 26688
rect 12306 26687 12352 26699
rect 12446 26688 12456 26868
rect 12520 26688 12530 26868
rect 12464 26687 12510 26688
rect 12560 26656 12764 27124
rect 13064 27075 13110 27087
rect 13064 26868 13070 27075
rect 13104 26868 13110 27075
rect 13202 26912 13212 27092
rect 13276 26912 13286 27092
rect 13380 27075 13426 27087
rect 13046 26688 13056 26868
rect 13120 26688 13130 26868
rect 13222 26699 13228 26912
rect 13262 26699 13268 26912
rect 13380 26868 13386 27075
rect 13420 26868 13426 27075
rect 13518 26912 13528 27092
rect 13592 26912 13602 27092
rect 13696 27075 13742 27087
rect 13064 26687 13110 26688
rect 13222 26687 13268 26699
rect 13362 26688 13372 26868
rect 13436 26688 13446 26868
rect 13538 26699 13544 26912
rect 13578 26699 13584 26912
rect 13696 26868 13702 27075
rect 13736 26868 13742 27075
rect 13834 26912 13844 27092
rect 13908 26912 13918 27092
rect 14012 27075 14058 27087
rect 13380 26687 13426 26688
rect 13538 26687 13584 26699
rect 13678 26688 13688 26868
rect 13752 26688 13762 26868
rect 13854 26699 13860 26912
rect 13894 26699 13900 26912
rect 14012 26868 14018 27075
rect 14052 26868 14058 27075
rect 14150 26912 14160 27092
rect 14224 26912 14234 27092
rect 14328 27075 14374 27087
rect 13696 26687 13742 26688
rect 13854 26687 13900 26699
rect 13994 26688 14004 26868
rect 14068 26688 14078 26868
rect 14170 26699 14176 26912
rect 14210 26699 14216 26912
rect 14328 26868 14334 27075
rect 14368 26868 14374 27075
rect 14466 26912 14476 27092
rect 14540 26912 14550 27092
rect 14644 27075 14690 27087
rect 14012 26687 14058 26688
rect 14170 26687 14216 26699
rect 14310 26688 14320 26868
rect 14384 26688 14394 26868
rect 14486 26699 14492 26912
rect 14526 26699 14532 26912
rect 14644 26868 14650 27075
rect 14684 26868 14690 27075
rect 14328 26687 14374 26688
rect 14486 26687 14532 26699
rect 14626 26688 14636 26868
rect 14700 26688 14710 26868
rect 14644 26687 14690 26688
rect 14740 26656 14944 27124
rect 15264 27075 15310 27087
rect 15264 26868 15270 27075
rect 15304 26868 15310 27075
rect 15402 26912 15412 27092
rect 15476 26912 15486 27092
rect 15580 27075 15626 27087
rect 15246 26688 15256 26868
rect 15320 26688 15330 26868
rect 15422 26699 15428 26912
rect 15462 26699 15468 26912
rect 15580 26868 15586 27075
rect 15620 26868 15626 27075
rect 15718 26912 15728 27092
rect 15792 26912 15802 27092
rect 15896 27075 15942 27087
rect 15264 26687 15310 26688
rect 15422 26687 15468 26699
rect 15562 26688 15572 26868
rect 15636 26688 15646 26868
rect 15738 26699 15744 26912
rect 15778 26699 15784 26912
rect 15896 26868 15902 27075
rect 15936 26868 15942 27075
rect 16034 26912 16044 27092
rect 16108 26912 16118 27092
rect 16212 27075 16258 27087
rect 15580 26687 15626 26688
rect 15738 26687 15784 26699
rect 15878 26688 15888 26868
rect 15952 26688 15962 26868
rect 16054 26699 16060 26912
rect 16094 26699 16100 26912
rect 16212 26868 16218 27075
rect 16252 26868 16258 27075
rect 16350 26912 16360 27092
rect 16424 26912 16434 27092
rect 16528 27075 16574 27087
rect 15896 26687 15942 26688
rect 16054 26687 16100 26699
rect 16194 26688 16204 26868
rect 16268 26688 16278 26868
rect 16370 26699 16376 26912
rect 16410 26699 16416 26912
rect 16528 26868 16534 27075
rect 16568 26868 16574 27075
rect 16666 26912 16676 27092
rect 16740 26912 16750 27092
rect 16844 27075 16890 27087
rect 16212 26687 16258 26688
rect 16370 26687 16416 26699
rect 16510 26688 16520 26868
rect 16584 26688 16594 26868
rect 16686 26699 16692 26912
rect 16726 26699 16732 26912
rect 16844 26868 16850 27075
rect 16884 26868 16890 27075
rect 16528 26687 16574 26688
rect 16686 26687 16732 26699
rect 16826 26688 16836 26868
rect 16900 26688 16910 26868
rect 16844 26687 16890 26688
rect 16940 26656 17144 27124
rect 6488 26640 8364 26656
rect 6488 26606 6552 26640
rect 6620 26606 6710 26640
rect 6778 26606 6868 26640
rect 6936 26606 7026 26640
rect 7094 26606 7184 26640
rect 7252 26606 7342 26640
rect 7410 26606 7500 26640
rect 7568 26606 7658 26640
rect 7726 26606 7816 26640
rect 7884 26606 7974 26640
rect 8042 26606 8364 26640
rect 6488 26532 8364 26606
rect 6488 26498 6552 26532
rect 6620 26498 6710 26532
rect 6778 26498 6868 26532
rect 6936 26498 7026 26532
rect 7094 26498 7184 26532
rect 7252 26498 7342 26532
rect 7410 26498 7500 26532
rect 7568 26498 7658 26532
rect 7726 26498 7816 26532
rect 7884 26498 7974 26532
rect 8042 26498 8364 26532
rect 6488 26488 8364 26498
rect 8708 26640 10584 26656
rect 8708 26606 8772 26640
rect 8840 26606 8930 26640
rect 8998 26606 9088 26640
rect 9156 26606 9246 26640
rect 9314 26606 9404 26640
rect 9472 26606 9562 26640
rect 9630 26606 9720 26640
rect 9788 26606 9878 26640
rect 9946 26606 10036 26640
rect 10104 26606 10194 26640
rect 10262 26606 10584 26640
rect 8708 26532 10584 26606
rect 8708 26498 8772 26532
rect 8840 26498 8930 26532
rect 8998 26498 9088 26532
rect 9156 26498 9246 26532
rect 9314 26498 9404 26532
rect 9472 26498 9562 26532
rect 9630 26498 9720 26532
rect 9788 26498 9878 26532
rect 9946 26498 10036 26532
rect 10104 26498 10194 26532
rect 10262 26498 10584 26532
rect 8708 26488 10584 26498
rect 10888 26640 12764 26656
rect 10888 26606 10952 26640
rect 11020 26606 11110 26640
rect 11178 26606 11268 26640
rect 11336 26606 11426 26640
rect 11494 26606 11584 26640
rect 11652 26606 11742 26640
rect 11810 26606 11900 26640
rect 11968 26606 12058 26640
rect 12126 26606 12216 26640
rect 12284 26606 12374 26640
rect 12442 26606 12764 26640
rect 10888 26532 12764 26606
rect 10888 26498 10952 26532
rect 11020 26498 11110 26532
rect 11178 26498 11268 26532
rect 11336 26498 11426 26532
rect 11494 26498 11584 26532
rect 11652 26498 11742 26532
rect 11810 26498 11900 26532
rect 11968 26498 12058 26532
rect 12126 26498 12216 26532
rect 12284 26498 12374 26532
rect 12442 26498 12764 26532
rect 10888 26488 12764 26498
rect 13068 26640 14944 26656
rect 13068 26606 13132 26640
rect 13200 26606 13290 26640
rect 13358 26606 13448 26640
rect 13516 26606 13606 26640
rect 13674 26606 13764 26640
rect 13832 26606 13922 26640
rect 13990 26606 14080 26640
rect 14148 26606 14238 26640
rect 14306 26606 14396 26640
rect 14464 26606 14554 26640
rect 14622 26606 14944 26640
rect 13068 26532 14944 26606
rect 13068 26498 13132 26532
rect 13200 26498 13290 26532
rect 13358 26498 13448 26532
rect 13516 26498 13606 26532
rect 13674 26498 13764 26532
rect 13832 26498 13922 26532
rect 13990 26498 14080 26532
rect 14148 26498 14238 26532
rect 14306 26498 14396 26532
rect 14464 26498 14554 26532
rect 14622 26498 14944 26532
rect 13068 26488 14944 26498
rect 15268 26640 17144 26656
rect 15268 26606 15332 26640
rect 15400 26606 15490 26640
rect 15558 26606 15648 26640
rect 15716 26606 15806 26640
rect 15874 26606 15964 26640
rect 16032 26606 16122 26640
rect 16190 26606 16280 26640
rect 16348 26606 16438 26640
rect 16506 26606 16596 26640
rect 16664 26606 16754 26640
rect 16822 26606 17144 26640
rect 15268 26532 17144 26606
rect 15268 26498 15332 26532
rect 15400 26498 15490 26532
rect 15558 26498 15648 26532
rect 15716 26498 15806 26532
rect 15874 26498 15964 26532
rect 16032 26498 16122 26532
rect 16190 26498 16280 26532
rect 16348 26498 16438 26532
rect 16506 26498 16596 26532
rect 16664 26498 16754 26532
rect 16822 26498 17144 26532
rect 15268 26488 17144 26498
rect 6484 26439 6530 26451
rect 6484 26232 6490 26439
rect 6524 26232 6530 26439
rect 6622 26276 6632 26456
rect 6696 26276 6706 26456
rect 6800 26439 6846 26451
rect 6466 26052 6476 26232
rect 6540 26052 6550 26232
rect 6642 26063 6648 26276
rect 6682 26063 6688 26276
rect 6800 26232 6806 26439
rect 6840 26232 6846 26439
rect 6938 26276 6948 26456
rect 7012 26276 7022 26456
rect 7116 26439 7162 26451
rect 6484 26051 6530 26052
rect 6642 26051 6688 26063
rect 6782 26052 6792 26232
rect 6856 26052 6866 26232
rect 6958 26063 6964 26276
rect 6998 26063 7004 26276
rect 7116 26232 7122 26439
rect 7156 26232 7162 26439
rect 7254 26276 7264 26456
rect 7328 26276 7338 26456
rect 7432 26439 7478 26451
rect 6800 26051 6846 26052
rect 6958 26051 7004 26063
rect 7098 26052 7108 26232
rect 7172 26052 7182 26232
rect 7274 26063 7280 26276
rect 7314 26063 7320 26276
rect 7432 26232 7438 26439
rect 7472 26232 7478 26439
rect 7570 26276 7580 26456
rect 7644 26276 7654 26456
rect 7748 26439 7794 26451
rect 7116 26051 7162 26052
rect 7274 26051 7320 26063
rect 7414 26052 7424 26232
rect 7488 26052 7498 26232
rect 7590 26063 7596 26276
rect 7630 26063 7636 26276
rect 7748 26232 7754 26439
rect 7788 26232 7794 26439
rect 7886 26276 7896 26456
rect 7960 26276 7970 26456
rect 8064 26439 8110 26451
rect 7432 26051 7478 26052
rect 7590 26051 7636 26063
rect 7730 26052 7740 26232
rect 7804 26052 7814 26232
rect 7906 26063 7912 26276
rect 7946 26063 7952 26276
rect 8064 26232 8070 26439
rect 8104 26232 8110 26439
rect 7748 26051 7794 26052
rect 7906 26051 7952 26063
rect 8046 26052 8056 26232
rect 8120 26052 8130 26232
rect 8064 26051 8110 26052
rect 8160 26016 8364 26488
rect 8704 26439 8750 26451
rect 8704 26232 8710 26439
rect 8744 26232 8750 26439
rect 8842 26276 8852 26456
rect 8916 26276 8926 26456
rect 9020 26439 9066 26451
rect 8686 26052 8696 26232
rect 8760 26052 8770 26232
rect 8862 26063 8868 26276
rect 8902 26063 8908 26276
rect 9020 26232 9026 26439
rect 9060 26232 9066 26439
rect 9158 26276 9168 26456
rect 9232 26276 9242 26456
rect 9336 26439 9382 26451
rect 8704 26051 8750 26052
rect 8862 26051 8908 26063
rect 9002 26052 9012 26232
rect 9076 26052 9086 26232
rect 9178 26063 9184 26276
rect 9218 26063 9224 26276
rect 9336 26232 9342 26439
rect 9376 26232 9382 26439
rect 9474 26276 9484 26456
rect 9548 26276 9558 26456
rect 9652 26439 9698 26451
rect 9020 26051 9066 26052
rect 9178 26051 9224 26063
rect 9318 26052 9328 26232
rect 9392 26052 9402 26232
rect 9494 26063 9500 26276
rect 9534 26063 9540 26276
rect 9652 26232 9658 26439
rect 9692 26232 9698 26439
rect 9790 26276 9800 26456
rect 9864 26276 9874 26456
rect 9968 26439 10014 26451
rect 9336 26051 9382 26052
rect 9494 26051 9540 26063
rect 9634 26052 9644 26232
rect 9708 26052 9718 26232
rect 9810 26063 9816 26276
rect 9850 26063 9856 26276
rect 9968 26232 9974 26439
rect 10008 26232 10014 26439
rect 10106 26276 10116 26456
rect 10180 26276 10190 26456
rect 10284 26439 10330 26451
rect 9652 26051 9698 26052
rect 9810 26051 9856 26063
rect 9950 26052 9960 26232
rect 10024 26052 10034 26232
rect 10126 26063 10132 26276
rect 10166 26063 10172 26276
rect 10284 26232 10290 26439
rect 10324 26232 10330 26439
rect 9968 26051 10014 26052
rect 10126 26051 10172 26063
rect 10266 26052 10276 26232
rect 10340 26052 10350 26232
rect 10284 26051 10330 26052
rect 10380 26016 10584 26488
rect 10884 26439 10930 26451
rect 10884 26232 10890 26439
rect 10924 26232 10930 26439
rect 11022 26276 11032 26456
rect 11096 26276 11106 26456
rect 11200 26439 11246 26451
rect 10866 26052 10876 26232
rect 10940 26052 10950 26232
rect 11042 26063 11048 26276
rect 11082 26063 11088 26276
rect 11200 26232 11206 26439
rect 11240 26232 11246 26439
rect 11338 26276 11348 26456
rect 11412 26276 11422 26456
rect 11516 26439 11562 26451
rect 10884 26051 10930 26052
rect 11042 26051 11088 26063
rect 11182 26052 11192 26232
rect 11256 26052 11266 26232
rect 11358 26063 11364 26276
rect 11398 26063 11404 26276
rect 11516 26232 11522 26439
rect 11556 26232 11562 26439
rect 11654 26276 11664 26456
rect 11728 26276 11738 26456
rect 11832 26439 11878 26451
rect 11200 26051 11246 26052
rect 11358 26051 11404 26063
rect 11498 26052 11508 26232
rect 11572 26052 11582 26232
rect 11674 26063 11680 26276
rect 11714 26063 11720 26276
rect 11832 26232 11838 26439
rect 11872 26232 11878 26439
rect 11970 26276 11980 26456
rect 12044 26276 12054 26456
rect 12148 26439 12194 26451
rect 11516 26051 11562 26052
rect 11674 26051 11720 26063
rect 11814 26052 11824 26232
rect 11888 26052 11898 26232
rect 11990 26063 11996 26276
rect 12030 26063 12036 26276
rect 12148 26232 12154 26439
rect 12188 26232 12194 26439
rect 12286 26276 12296 26456
rect 12360 26276 12370 26456
rect 12464 26439 12510 26451
rect 11832 26051 11878 26052
rect 11990 26051 12036 26063
rect 12130 26052 12140 26232
rect 12204 26052 12214 26232
rect 12306 26063 12312 26276
rect 12346 26063 12352 26276
rect 12464 26232 12470 26439
rect 12504 26232 12510 26439
rect 12148 26051 12194 26052
rect 12306 26051 12352 26063
rect 12446 26052 12456 26232
rect 12520 26052 12530 26232
rect 12464 26051 12510 26052
rect 12560 26016 12764 26488
rect 13064 26439 13110 26451
rect 13064 26232 13070 26439
rect 13104 26232 13110 26439
rect 13202 26276 13212 26456
rect 13276 26276 13286 26456
rect 13380 26439 13426 26451
rect 13046 26052 13056 26232
rect 13120 26052 13130 26232
rect 13222 26063 13228 26276
rect 13262 26063 13268 26276
rect 13380 26232 13386 26439
rect 13420 26232 13426 26439
rect 13518 26276 13528 26456
rect 13592 26276 13602 26456
rect 13696 26439 13742 26451
rect 13064 26051 13110 26052
rect 13222 26051 13268 26063
rect 13362 26052 13372 26232
rect 13436 26052 13446 26232
rect 13538 26063 13544 26276
rect 13578 26063 13584 26276
rect 13696 26232 13702 26439
rect 13736 26232 13742 26439
rect 13834 26276 13844 26456
rect 13908 26276 13918 26456
rect 14012 26439 14058 26451
rect 13380 26051 13426 26052
rect 13538 26051 13584 26063
rect 13678 26052 13688 26232
rect 13752 26052 13762 26232
rect 13854 26063 13860 26276
rect 13894 26063 13900 26276
rect 14012 26232 14018 26439
rect 14052 26232 14058 26439
rect 14150 26276 14160 26456
rect 14224 26276 14234 26456
rect 14328 26439 14374 26451
rect 13696 26051 13742 26052
rect 13854 26051 13900 26063
rect 13994 26052 14004 26232
rect 14068 26052 14078 26232
rect 14170 26063 14176 26276
rect 14210 26063 14216 26276
rect 14328 26232 14334 26439
rect 14368 26232 14374 26439
rect 14466 26276 14476 26456
rect 14540 26276 14550 26456
rect 14644 26439 14690 26451
rect 14012 26051 14058 26052
rect 14170 26051 14216 26063
rect 14310 26052 14320 26232
rect 14384 26052 14394 26232
rect 14486 26063 14492 26276
rect 14526 26063 14532 26276
rect 14644 26232 14650 26439
rect 14684 26232 14690 26439
rect 14328 26051 14374 26052
rect 14486 26051 14532 26063
rect 14626 26052 14636 26232
rect 14700 26052 14710 26232
rect 14644 26051 14690 26052
rect 14740 26016 14944 26488
rect 15264 26439 15310 26451
rect 15264 26232 15270 26439
rect 15304 26232 15310 26439
rect 15402 26276 15412 26456
rect 15476 26276 15486 26456
rect 15580 26439 15626 26451
rect 15246 26052 15256 26232
rect 15320 26052 15330 26232
rect 15422 26063 15428 26276
rect 15462 26063 15468 26276
rect 15580 26232 15586 26439
rect 15620 26232 15626 26439
rect 15718 26276 15728 26456
rect 15792 26276 15802 26456
rect 15896 26439 15942 26451
rect 15264 26051 15310 26052
rect 15422 26051 15468 26063
rect 15562 26052 15572 26232
rect 15636 26052 15646 26232
rect 15738 26063 15744 26276
rect 15778 26063 15784 26276
rect 15896 26232 15902 26439
rect 15936 26232 15942 26439
rect 16034 26276 16044 26456
rect 16108 26276 16118 26456
rect 16212 26439 16258 26451
rect 15580 26051 15626 26052
rect 15738 26051 15784 26063
rect 15878 26052 15888 26232
rect 15952 26052 15962 26232
rect 16054 26063 16060 26276
rect 16094 26063 16100 26276
rect 16212 26232 16218 26439
rect 16252 26232 16258 26439
rect 16350 26276 16360 26456
rect 16424 26276 16434 26456
rect 16528 26439 16574 26451
rect 15896 26051 15942 26052
rect 16054 26051 16100 26063
rect 16194 26052 16204 26232
rect 16268 26052 16278 26232
rect 16370 26063 16376 26276
rect 16410 26063 16416 26276
rect 16528 26232 16534 26439
rect 16568 26232 16574 26439
rect 16666 26276 16676 26456
rect 16740 26276 16750 26456
rect 16844 26439 16890 26451
rect 16212 26051 16258 26052
rect 16370 26051 16416 26063
rect 16510 26052 16520 26232
rect 16584 26052 16594 26232
rect 16686 26063 16692 26276
rect 16726 26063 16732 26276
rect 16844 26232 16850 26439
rect 16884 26232 16890 26439
rect 16528 26051 16574 26052
rect 16686 26051 16732 26063
rect 16826 26052 16836 26232
rect 16900 26052 16910 26232
rect 16844 26051 16890 26052
rect 16940 26016 17144 26488
rect 6488 26004 8364 26016
rect 6488 25970 6552 26004
rect 6620 25970 6710 26004
rect 6778 25970 6868 26004
rect 6936 25970 7026 26004
rect 7094 25970 7184 26004
rect 7252 25970 7342 26004
rect 7410 25970 7500 26004
rect 7568 25970 7658 26004
rect 7726 25970 7816 26004
rect 7884 25970 7974 26004
rect 8042 25970 8364 26004
rect 6488 25896 8364 25970
rect 6488 25862 6552 25896
rect 6620 25862 6710 25896
rect 6778 25862 6868 25896
rect 6936 25862 7026 25896
rect 7094 25862 7184 25896
rect 7252 25862 7342 25896
rect 7410 25862 7500 25896
rect 7568 25862 7658 25896
rect 7726 25862 7816 25896
rect 7884 25862 7974 25896
rect 8042 25862 8364 25896
rect 6488 25848 8364 25862
rect 8708 26004 10584 26016
rect 8708 25970 8772 26004
rect 8840 25970 8930 26004
rect 8998 25970 9088 26004
rect 9156 25970 9246 26004
rect 9314 25970 9404 26004
rect 9472 25970 9562 26004
rect 9630 25970 9720 26004
rect 9788 25970 9878 26004
rect 9946 25970 10036 26004
rect 10104 25970 10194 26004
rect 10262 25970 10584 26004
rect 8708 25896 10584 25970
rect 8708 25862 8772 25896
rect 8840 25862 8930 25896
rect 8998 25862 9088 25896
rect 9156 25862 9246 25896
rect 9314 25862 9404 25896
rect 9472 25862 9562 25896
rect 9630 25862 9720 25896
rect 9788 25862 9878 25896
rect 9946 25862 10036 25896
rect 10104 25862 10194 25896
rect 10262 25862 10584 25896
rect 8708 25848 10584 25862
rect 10888 26004 12764 26016
rect 10888 25970 10952 26004
rect 11020 25970 11110 26004
rect 11178 25970 11268 26004
rect 11336 25970 11426 26004
rect 11494 25970 11584 26004
rect 11652 25970 11742 26004
rect 11810 25970 11900 26004
rect 11968 25970 12058 26004
rect 12126 25970 12216 26004
rect 12284 25970 12374 26004
rect 12442 25970 12764 26004
rect 10888 25896 12764 25970
rect 10888 25862 10952 25896
rect 11020 25862 11110 25896
rect 11178 25862 11268 25896
rect 11336 25862 11426 25896
rect 11494 25862 11584 25896
rect 11652 25862 11742 25896
rect 11810 25862 11900 25896
rect 11968 25862 12058 25896
rect 12126 25862 12216 25896
rect 12284 25862 12374 25896
rect 12442 25862 12764 25896
rect 10888 25848 12764 25862
rect 13068 26004 14944 26016
rect 13068 25970 13132 26004
rect 13200 25970 13290 26004
rect 13358 25970 13448 26004
rect 13516 25970 13606 26004
rect 13674 25970 13764 26004
rect 13832 25970 13922 26004
rect 13990 25970 14080 26004
rect 14148 25970 14238 26004
rect 14306 25970 14396 26004
rect 14464 25970 14554 26004
rect 14622 25970 14944 26004
rect 13068 25896 14944 25970
rect 13068 25862 13132 25896
rect 13200 25862 13290 25896
rect 13358 25862 13448 25896
rect 13516 25862 13606 25896
rect 13674 25862 13764 25896
rect 13832 25862 13922 25896
rect 13990 25862 14080 25896
rect 14148 25862 14238 25896
rect 14306 25862 14396 25896
rect 14464 25862 14554 25896
rect 14622 25862 14944 25896
rect 13068 25848 14944 25862
rect 15268 26004 17144 26016
rect 15268 25970 15332 26004
rect 15400 25970 15490 26004
rect 15558 25970 15648 26004
rect 15716 25970 15806 26004
rect 15874 25970 15964 26004
rect 16032 25970 16122 26004
rect 16190 25970 16280 26004
rect 16348 25970 16438 26004
rect 16506 25970 16596 26004
rect 16664 25970 16754 26004
rect 16822 25970 17144 26004
rect 15268 25896 17144 25970
rect 15268 25862 15332 25896
rect 15400 25862 15490 25896
rect 15558 25862 15648 25896
rect 15716 25862 15806 25896
rect 15874 25862 15964 25896
rect 16032 25862 16122 25896
rect 16190 25862 16280 25896
rect 16348 25862 16438 25896
rect 16506 25862 16596 25896
rect 16664 25862 16754 25896
rect 16822 25862 17144 25896
rect 15268 25848 17144 25862
rect 6484 25803 6530 25815
rect 6484 25592 6490 25803
rect 6524 25592 6530 25803
rect 6622 25636 6632 25816
rect 6696 25636 6706 25816
rect 6800 25803 6846 25815
rect 6466 25412 6476 25592
rect 6540 25412 6550 25592
rect 6642 25427 6648 25636
rect 6682 25427 6688 25636
rect 6800 25592 6806 25803
rect 6840 25592 6846 25803
rect 6938 25636 6948 25816
rect 7012 25636 7022 25816
rect 7116 25803 7162 25815
rect 6642 25415 6688 25427
rect 6782 25412 6792 25592
rect 6856 25412 6866 25592
rect 6958 25427 6964 25636
rect 6998 25427 7004 25636
rect 7116 25592 7122 25803
rect 7156 25592 7162 25803
rect 7254 25636 7264 25816
rect 7328 25636 7338 25816
rect 7432 25803 7478 25815
rect 6958 25415 7004 25427
rect 7098 25412 7108 25592
rect 7172 25412 7182 25592
rect 7274 25427 7280 25636
rect 7314 25427 7320 25636
rect 7432 25592 7438 25803
rect 7472 25592 7478 25803
rect 7570 25636 7580 25816
rect 7644 25636 7654 25816
rect 7748 25803 7794 25815
rect 7274 25415 7320 25427
rect 7414 25412 7424 25592
rect 7488 25412 7498 25592
rect 7590 25427 7596 25636
rect 7630 25427 7636 25636
rect 7748 25592 7754 25803
rect 7788 25592 7794 25803
rect 7886 25636 7896 25816
rect 7960 25636 7970 25816
rect 8064 25803 8110 25815
rect 7590 25415 7636 25427
rect 7730 25412 7740 25592
rect 7804 25412 7814 25592
rect 7906 25427 7912 25636
rect 7946 25427 7952 25636
rect 8064 25592 8070 25803
rect 8104 25592 8110 25803
rect 7906 25415 7952 25427
rect 8046 25412 8056 25592
rect 8120 25412 8130 25592
rect 8160 25376 8364 25848
rect 8704 25803 8750 25815
rect 8704 25592 8710 25803
rect 8744 25592 8750 25803
rect 8842 25636 8852 25816
rect 8916 25636 8926 25816
rect 9020 25803 9066 25815
rect 8686 25412 8696 25592
rect 8760 25412 8770 25592
rect 8862 25427 8868 25636
rect 8902 25427 8908 25636
rect 9020 25592 9026 25803
rect 9060 25592 9066 25803
rect 9158 25636 9168 25816
rect 9232 25636 9242 25816
rect 9336 25803 9382 25815
rect 8862 25415 8908 25427
rect 9002 25412 9012 25592
rect 9076 25412 9086 25592
rect 9178 25427 9184 25636
rect 9218 25427 9224 25636
rect 9336 25592 9342 25803
rect 9376 25592 9382 25803
rect 9474 25636 9484 25816
rect 9548 25636 9558 25816
rect 9652 25803 9698 25815
rect 9178 25415 9224 25427
rect 9318 25412 9328 25592
rect 9392 25412 9402 25592
rect 9494 25427 9500 25636
rect 9534 25427 9540 25636
rect 9652 25592 9658 25803
rect 9692 25592 9698 25803
rect 9790 25636 9800 25816
rect 9864 25636 9874 25816
rect 9968 25803 10014 25815
rect 9494 25415 9540 25427
rect 9634 25412 9644 25592
rect 9708 25412 9718 25592
rect 9810 25427 9816 25636
rect 9850 25427 9856 25636
rect 9968 25592 9974 25803
rect 10008 25592 10014 25803
rect 10106 25636 10116 25816
rect 10180 25636 10190 25816
rect 10284 25803 10330 25815
rect 9810 25415 9856 25427
rect 9950 25412 9960 25592
rect 10024 25412 10034 25592
rect 10126 25427 10132 25636
rect 10166 25427 10172 25636
rect 10284 25592 10290 25803
rect 10324 25592 10330 25803
rect 10126 25415 10172 25427
rect 10266 25412 10276 25592
rect 10340 25412 10350 25592
rect 10380 25376 10584 25848
rect 10884 25803 10930 25815
rect 10884 25592 10890 25803
rect 10924 25592 10930 25803
rect 11022 25636 11032 25816
rect 11096 25636 11106 25816
rect 11200 25803 11246 25815
rect 10866 25412 10876 25592
rect 10940 25412 10950 25592
rect 11042 25427 11048 25636
rect 11082 25427 11088 25636
rect 11200 25592 11206 25803
rect 11240 25592 11246 25803
rect 11338 25636 11348 25816
rect 11412 25636 11422 25816
rect 11516 25803 11562 25815
rect 11042 25415 11088 25427
rect 11182 25412 11192 25592
rect 11256 25412 11266 25592
rect 11358 25427 11364 25636
rect 11398 25427 11404 25636
rect 11516 25592 11522 25803
rect 11556 25592 11562 25803
rect 11654 25636 11664 25816
rect 11728 25636 11738 25816
rect 11832 25803 11878 25815
rect 11358 25415 11404 25427
rect 11498 25412 11508 25592
rect 11572 25412 11582 25592
rect 11674 25427 11680 25636
rect 11714 25427 11720 25636
rect 11832 25592 11838 25803
rect 11872 25592 11878 25803
rect 11970 25636 11980 25816
rect 12044 25636 12054 25816
rect 12148 25803 12194 25815
rect 11674 25415 11720 25427
rect 11814 25412 11824 25592
rect 11888 25412 11898 25592
rect 11990 25427 11996 25636
rect 12030 25427 12036 25636
rect 12148 25592 12154 25803
rect 12188 25592 12194 25803
rect 12286 25636 12296 25816
rect 12360 25636 12370 25816
rect 12464 25803 12510 25815
rect 11990 25415 12036 25427
rect 12130 25412 12140 25592
rect 12204 25412 12214 25592
rect 12306 25427 12312 25636
rect 12346 25427 12352 25636
rect 12464 25592 12470 25803
rect 12504 25592 12510 25803
rect 12306 25415 12352 25427
rect 12446 25412 12456 25592
rect 12520 25412 12530 25592
rect 12560 25376 12764 25848
rect 13064 25803 13110 25815
rect 13064 25592 13070 25803
rect 13104 25592 13110 25803
rect 13202 25636 13212 25816
rect 13276 25636 13286 25816
rect 13380 25803 13426 25815
rect 13046 25412 13056 25592
rect 13120 25412 13130 25592
rect 13222 25427 13228 25636
rect 13262 25427 13268 25636
rect 13380 25592 13386 25803
rect 13420 25592 13426 25803
rect 13518 25636 13528 25816
rect 13592 25636 13602 25816
rect 13696 25803 13742 25815
rect 13222 25415 13268 25427
rect 13362 25412 13372 25592
rect 13436 25412 13446 25592
rect 13538 25427 13544 25636
rect 13578 25427 13584 25636
rect 13696 25592 13702 25803
rect 13736 25592 13742 25803
rect 13834 25636 13844 25816
rect 13908 25636 13918 25816
rect 14012 25803 14058 25815
rect 13538 25415 13584 25427
rect 13678 25412 13688 25592
rect 13752 25412 13762 25592
rect 13854 25427 13860 25636
rect 13894 25427 13900 25636
rect 14012 25592 14018 25803
rect 14052 25592 14058 25803
rect 14150 25636 14160 25816
rect 14224 25636 14234 25816
rect 14328 25803 14374 25815
rect 13854 25415 13900 25427
rect 13994 25412 14004 25592
rect 14068 25412 14078 25592
rect 14170 25427 14176 25636
rect 14210 25427 14216 25636
rect 14328 25592 14334 25803
rect 14368 25592 14374 25803
rect 14466 25636 14476 25816
rect 14540 25636 14550 25816
rect 14644 25803 14690 25815
rect 14170 25415 14216 25427
rect 14310 25412 14320 25592
rect 14384 25412 14394 25592
rect 14486 25427 14492 25636
rect 14526 25427 14532 25636
rect 14644 25592 14650 25803
rect 14684 25592 14690 25803
rect 14486 25415 14532 25427
rect 14626 25412 14636 25592
rect 14700 25412 14710 25592
rect 14740 25376 14944 25848
rect 15264 25803 15310 25815
rect 15264 25592 15270 25803
rect 15304 25592 15310 25803
rect 15402 25636 15412 25816
rect 15476 25636 15486 25816
rect 15580 25803 15626 25815
rect 15246 25412 15256 25592
rect 15320 25412 15330 25592
rect 15422 25427 15428 25636
rect 15462 25427 15468 25636
rect 15580 25592 15586 25803
rect 15620 25592 15626 25803
rect 15718 25636 15728 25816
rect 15792 25636 15802 25816
rect 15896 25803 15942 25815
rect 15422 25415 15468 25427
rect 15562 25412 15572 25592
rect 15636 25412 15646 25592
rect 15738 25427 15744 25636
rect 15778 25427 15784 25636
rect 15896 25592 15902 25803
rect 15936 25592 15942 25803
rect 16034 25636 16044 25816
rect 16108 25636 16118 25816
rect 16212 25803 16258 25815
rect 15738 25415 15784 25427
rect 15878 25412 15888 25592
rect 15952 25412 15962 25592
rect 16054 25427 16060 25636
rect 16094 25427 16100 25636
rect 16212 25592 16218 25803
rect 16252 25592 16258 25803
rect 16350 25636 16360 25816
rect 16424 25636 16434 25816
rect 16528 25803 16574 25815
rect 16054 25415 16100 25427
rect 16194 25412 16204 25592
rect 16268 25412 16278 25592
rect 16370 25427 16376 25636
rect 16410 25427 16416 25636
rect 16528 25592 16534 25803
rect 16568 25592 16574 25803
rect 16666 25636 16676 25816
rect 16740 25636 16750 25816
rect 16844 25803 16890 25815
rect 16370 25415 16416 25427
rect 16510 25412 16520 25592
rect 16584 25412 16594 25592
rect 16686 25427 16692 25636
rect 16726 25427 16732 25636
rect 16844 25592 16850 25803
rect 16884 25592 16890 25803
rect 16686 25415 16732 25427
rect 16826 25412 16836 25592
rect 16900 25412 16910 25592
rect 16940 25376 17144 25848
rect 19048 25436 19232 25442
rect 6488 25368 8364 25376
rect 6488 25334 6552 25368
rect 6620 25334 6710 25368
rect 6778 25334 6868 25368
rect 6936 25334 7026 25368
rect 7094 25334 7184 25368
rect 7252 25334 7342 25368
rect 7410 25334 7500 25368
rect 7568 25334 7658 25368
rect 7726 25334 7816 25368
rect 7884 25334 7974 25368
rect 8042 25334 8364 25368
rect 6488 25320 8364 25334
rect 8708 25368 10584 25376
rect 8708 25334 8772 25368
rect 8840 25334 8930 25368
rect 8998 25334 9088 25368
rect 9156 25334 9246 25368
rect 9314 25334 9404 25368
rect 9472 25334 9562 25368
rect 9630 25334 9720 25368
rect 9788 25334 9878 25368
rect 9946 25334 10036 25368
rect 10104 25334 10194 25368
rect 10262 25334 10584 25368
rect 8708 25320 10584 25334
rect 10888 25368 12764 25376
rect 10888 25334 10952 25368
rect 11020 25334 11110 25368
rect 11178 25334 11268 25368
rect 11336 25334 11426 25368
rect 11494 25334 11584 25368
rect 11652 25334 11742 25368
rect 11810 25334 11900 25368
rect 11968 25334 12058 25368
rect 12126 25334 12216 25368
rect 12284 25334 12374 25368
rect 12442 25334 12764 25368
rect 10888 25320 12764 25334
rect 13068 25368 14944 25376
rect 13068 25334 13132 25368
rect 13200 25334 13290 25368
rect 13358 25334 13448 25368
rect 13516 25334 13606 25368
rect 13674 25334 13764 25368
rect 13832 25334 13922 25368
rect 13990 25334 14080 25368
rect 14148 25334 14238 25368
rect 14306 25334 14396 25368
rect 14464 25334 14554 25368
rect 14622 25334 14944 25368
rect 13068 25320 14944 25334
rect 15268 25368 17144 25376
rect 15268 25334 15332 25368
rect 15400 25334 15490 25368
rect 15558 25334 15648 25368
rect 15716 25334 15806 25368
rect 15874 25334 15964 25368
rect 16032 25334 16122 25368
rect 16190 25334 16280 25368
rect 16348 25334 16438 25368
rect 16506 25334 16596 25368
rect 16664 25334 16754 25368
rect 16822 25334 17144 25368
rect 15268 25320 17144 25334
rect 6488 25272 17144 25320
rect 18340 25296 19060 25436
rect 19220 25296 19232 25436
rect 8020 25116 17004 25272
rect 18340 25120 18580 25296
rect 19048 25290 19232 25296
rect 6520 25096 17004 25116
rect 6520 25072 8224 25096
rect 6520 25038 6538 25072
rect 6572 25038 6730 25072
rect 6764 25038 6922 25072
rect 6956 25038 7114 25072
rect 7148 25038 7306 25072
rect 7340 25038 7498 25072
rect 7532 25038 7690 25072
rect 7724 25038 7882 25072
rect 7916 25038 8224 25072
rect 6520 25032 8224 25038
rect 8740 25072 10444 25096
rect 8740 25038 8758 25072
rect 8792 25038 8950 25072
rect 8984 25038 9142 25072
rect 9176 25038 9334 25072
rect 9368 25038 9526 25072
rect 9560 25038 9718 25072
rect 9752 25038 9910 25072
rect 9944 25038 10102 25072
rect 10136 25038 10444 25072
rect 8740 25032 10444 25038
rect 10920 25072 12624 25096
rect 10920 25038 10938 25072
rect 10972 25038 11130 25072
rect 11164 25038 11322 25072
rect 11356 25038 11514 25072
rect 11548 25038 11706 25072
rect 11740 25038 11898 25072
rect 11932 25038 12090 25072
rect 12124 25038 12282 25072
rect 12316 25038 12624 25072
rect 10920 25032 12624 25038
rect 13100 25072 14804 25096
rect 13100 25038 13118 25072
rect 13152 25038 13310 25072
rect 13344 25038 13502 25072
rect 13536 25038 13694 25072
rect 13728 25038 13886 25072
rect 13920 25038 14078 25072
rect 14112 25038 14270 25072
rect 14304 25038 14462 25072
rect 14496 25038 14804 25072
rect 13100 25032 14804 25038
rect 15300 25072 17004 25096
rect 15300 25038 15318 25072
rect 15352 25038 15510 25072
rect 15544 25038 15702 25072
rect 15736 25038 15894 25072
rect 15928 25038 16086 25072
rect 16120 25038 16278 25072
rect 16312 25038 16470 25072
rect 16504 25038 16662 25072
rect 16696 25038 17004 25072
rect 15300 25032 17004 25038
rect 6484 24979 6530 24991
rect 6484 24768 6490 24979
rect 6524 24768 6530 24979
rect 6562 24812 6572 24992
rect 6636 24812 6646 24992
rect 6676 24979 6722 24991
rect 6466 24588 6476 24768
rect 6540 24588 6550 24768
rect 6580 24603 6586 24812
rect 6620 24603 6626 24812
rect 6676 24768 6682 24979
rect 6716 24768 6722 24979
rect 6754 24812 6764 24992
rect 6828 24812 6838 24992
rect 6868 24979 6914 24991
rect 6580 24591 6626 24603
rect 6654 24588 6664 24768
rect 6728 24588 6738 24768
rect 6772 24603 6778 24812
rect 6812 24603 6818 24812
rect 6868 24768 6874 24979
rect 6908 24768 6914 24979
rect 6946 24812 6956 24992
rect 7020 24812 7030 24992
rect 7060 24979 7106 24991
rect 6772 24591 6818 24603
rect 6846 24588 6856 24768
rect 6920 24588 6930 24768
rect 6964 24603 6970 24812
rect 7004 24603 7010 24812
rect 7060 24768 7066 24979
rect 7100 24768 7106 24979
rect 7138 24812 7148 24992
rect 7212 24812 7222 24992
rect 7252 24979 7298 24991
rect 6964 24591 7010 24603
rect 7042 24588 7052 24768
rect 7116 24588 7126 24768
rect 7156 24603 7162 24812
rect 7196 24603 7202 24812
rect 7252 24768 7258 24979
rect 7292 24768 7298 24979
rect 7330 24812 7340 24992
rect 7404 24812 7414 24992
rect 7444 24979 7490 24991
rect 7156 24591 7202 24603
rect 7234 24588 7244 24768
rect 7308 24588 7318 24768
rect 7348 24603 7354 24812
rect 7388 24603 7394 24812
rect 7444 24768 7450 24979
rect 7484 24768 7490 24979
rect 7522 24812 7532 24992
rect 7596 24812 7606 24992
rect 7636 24979 7682 24991
rect 7348 24591 7394 24603
rect 7426 24588 7436 24768
rect 7500 24588 7510 24768
rect 7540 24603 7546 24812
rect 7580 24603 7586 24812
rect 7636 24768 7642 24979
rect 7676 24768 7682 24979
rect 7714 24812 7724 24992
rect 7788 24812 7798 24992
rect 7828 24979 7874 24991
rect 7540 24591 7586 24603
rect 7618 24588 7628 24768
rect 7692 24588 7702 24768
rect 7732 24603 7738 24812
rect 7772 24603 7778 24812
rect 7828 24768 7834 24979
rect 7868 24768 7874 24979
rect 7906 24812 7916 24992
rect 7980 24812 7990 24992
rect 7732 24591 7778 24603
rect 7810 24588 7820 24768
rect 7884 24588 7894 24768
rect 7924 24603 7930 24812
rect 7964 24603 7970 24812
rect 7924 24591 7970 24603
rect 8020 24552 8224 25032
rect 8704 24979 8750 24991
rect 8704 24768 8710 24979
rect 8744 24768 8750 24979
rect 8782 24812 8792 24992
rect 8856 24812 8866 24992
rect 8896 24979 8942 24991
rect 8686 24588 8696 24768
rect 8760 24588 8770 24768
rect 8800 24603 8806 24812
rect 8840 24603 8846 24812
rect 8896 24768 8902 24979
rect 8936 24768 8942 24979
rect 8974 24812 8984 24992
rect 9048 24812 9058 24992
rect 9088 24979 9134 24991
rect 8800 24591 8846 24603
rect 8874 24588 8884 24768
rect 8948 24588 8958 24768
rect 8992 24603 8998 24812
rect 9032 24603 9038 24812
rect 9088 24768 9094 24979
rect 9128 24768 9134 24979
rect 9166 24812 9176 24992
rect 9240 24812 9250 24992
rect 9280 24979 9326 24991
rect 8992 24591 9038 24603
rect 9066 24588 9076 24768
rect 9140 24588 9150 24768
rect 9184 24603 9190 24812
rect 9224 24603 9230 24812
rect 9280 24768 9286 24979
rect 9320 24768 9326 24979
rect 9358 24812 9368 24992
rect 9432 24812 9442 24992
rect 9472 24979 9518 24991
rect 9184 24591 9230 24603
rect 9262 24588 9272 24768
rect 9336 24588 9346 24768
rect 9376 24603 9382 24812
rect 9416 24603 9422 24812
rect 9472 24768 9478 24979
rect 9512 24768 9518 24979
rect 9550 24812 9560 24992
rect 9624 24812 9634 24992
rect 9664 24979 9710 24991
rect 9376 24591 9422 24603
rect 9454 24588 9464 24768
rect 9528 24588 9538 24768
rect 9568 24603 9574 24812
rect 9608 24603 9614 24812
rect 9664 24768 9670 24979
rect 9704 24768 9710 24979
rect 9742 24812 9752 24992
rect 9816 24812 9826 24992
rect 9856 24979 9902 24991
rect 9568 24591 9614 24603
rect 9646 24588 9656 24768
rect 9720 24588 9730 24768
rect 9760 24603 9766 24812
rect 9800 24603 9806 24812
rect 9856 24768 9862 24979
rect 9896 24768 9902 24979
rect 9934 24812 9944 24992
rect 10008 24812 10018 24992
rect 10048 24979 10094 24991
rect 9760 24591 9806 24603
rect 9838 24588 9848 24768
rect 9912 24588 9922 24768
rect 9952 24603 9958 24812
rect 9992 24603 9998 24812
rect 10048 24768 10054 24979
rect 10088 24768 10094 24979
rect 10126 24812 10136 24992
rect 10200 24812 10210 24992
rect 9952 24591 9998 24603
rect 10030 24588 10040 24768
rect 10104 24588 10114 24768
rect 10144 24603 10150 24812
rect 10184 24603 10190 24812
rect 10144 24591 10190 24603
rect 10240 24552 10444 25032
rect 10884 24979 10930 24991
rect 10884 24768 10890 24979
rect 10924 24768 10930 24979
rect 10962 24812 10972 24992
rect 11036 24812 11046 24992
rect 11076 24979 11122 24991
rect 10866 24588 10876 24768
rect 10940 24588 10950 24768
rect 10980 24603 10986 24812
rect 11020 24603 11026 24812
rect 11076 24768 11082 24979
rect 11116 24768 11122 24979
rect 11154 24812 11164 24992
rect 11228 24812 11238 24992
rect 11268 24979 11314 24991
rect 10980 24591 11026 24603
rect 11054 24588 11064 24768
rect 11128 24588 11138 24768
rect 11172 24603 11178 24812
rect 11212 24603 11218 24812
rect 11268 24768 11274 24979
rect 11308 24768 11314 24979
rect 11346 24812 11356 24992
rect 11420 24812 11430 24992
rect 11460 24979 11506 24991
rect 11172 24591 11218 24603
rect 11246 24588 11256 24768
rect 11320 24588 11330 24768
rect 11364 24603 11370 24812
rect 11404 24603 11410 24812
rect 11460 24768 11466 24979
rect 11500 24768 11506 24979
rect 11538 24812 11548 24992
rect 11612 24812 11622 24992
rect 11652 24979 11698 24991
rect 11364 24591 11410 24603
rect 11442 24588 11452 24768
rect 11516 24588 11526 24768
rect 11556 24603 11562 24812
rect 11596 24603 11602 24812
rect 11652 24768 11658 24979
rect 11692 24768 11698 24979
rect 11730 24812 11740 24992
rect 11804 24812 11814 24992
rect 11844 24979 11890 24991
rect 11556 24591 11602 24603
rect 11634 24588 11644 24768
rect 11708 24588 11718 24768
rect 11748 24603 11754 24812
rect 11788 24603 11794 24812
rect 11844 24768 11850 24979
rect 11884 24768 11890 24979
rect 11922 24812 11932 24992
rect 11996 24812 12006 24992
rect 12036 24979 12082 24991
rect 11748 24591 11794 24603
rect 11826 24588 11836 24768
rect 11900 24588 11910 24768
rect 11940 24603 11946 24812
rect 11980 24603 11986 24812
rect 12036 24768 12042 24979
rect 12076 24768 12082 24979
rect 12114 24812 12124 24992
rect 12188 24812 12198 24992
rect 12228 24979 12274 24991
rect 11940 24591 11986 24603
rect 12018 24588 12028 24768
rect 12092 24588 12102 24768
rect 12132 24603 12138 24812
rect 12172 24603 12178 24812
rect 12228 24768 12234 24979
rect 12268 24768 12274 24979
rect 12306 24812 12316 24992
rect 12380 24812 12390 24992
rect 12132 24591 12178 24603
rect 12210 24588 12220 24768
rect 12284 24588 12294 24768
rect 12324 24603 12330 24812
rect 12364 24603 12370 24812
rect 12324 24591 12370 24603
rect 12420 24552 12624 25032
rect 13064 24979 13110 24991
rect 13064 24768 13070 24979
rect 13104 24768 13110 24979
rect 13142 24812 13152 24992
rect 13216 24812 13226 24992
rect 13256 24979 13302 24991
rect 13046 24588 13056 24768
rect 13120 24588 13130 24768
rect 13160 24603 13166 24812
rect 13200 24603 13206 24812
rect 13256 24768 13262 24979
rect 13296 24768 13302 24979
rect 13334 24812 13344 24992
rect 13408 24812 13418 24992
rect 13448 24979 13494 24991
rect 13160 24591 13206 24603
rect 13234 24588 13244 24768
rect 13308 24588 13318 24768
rect 13352 24603 13358 24812
rect 13392 24603 13398 24812
rect 13448 24768 13454 24979
rect 13488 24768 13494 24979
rect 13526 24812 13536 24992
rect 13600 24812 13610 24992
rect 13640 24979 13686 24991
rect 13352 24591 13398 24603
rect 13426 24588 13436 24768
rect 13500 24588 13510 24768
rect 13544 24603 13550 24812
rect 13584 24603 13590 24812
rect 13640 24768 13646 24979
rect 13680 24768 13686 24979
rect 13718 24812 13728 24992
rect 13792 24812 13802 24992
rect 13832 24979 13878 24991
rect 13544 24591 13590 24603
rect 13622 24588 13632 24768
rect 13696 24588 13706 24768
rect 13736 24603 13742 24812
rect 13776 24603 13782 24812
rect 13832 24768 13838 24979
rect 13872 24768 13878 24979
rect 13910 24812 13920 24992
rect 13984 24812 13994 24992
rect 14024 24979 14070 24991
rect 13736 24591 13782 24603
rect 13814 24588 13824 24768
rect 13888 24588 13898 24768
rect 13928 24603 13934 24812
rect 13968 24603 13974 24812
rect 14024 24768 14030 24979
rect 14064 24768 14070 24979
rect 14102 24812 14112 24992
rect 14176 24812 14186 24992
rect 14216 24979 14262 24991
rect 13928 24591 13974 24603
rect 14006 24588 14016 24768
rect 14080 24588 14090 24768
rect 14120 24603 14126 24812
rect 14160 24603 14166 24812
rect 14216 24768 14222 24979
rect 14256 24768 14262 24979
rect 14294 24812 14304 24992
rect 14368 24812 14378 24992
rect 14408 24979 14454 24991
rect 14120 24591 14166 24603
rect 14198 24588 14208 24768
rect 14272 24588 14282 24768
rect 14312 24603 14318 24812
rect 14352 24603 14358 24812
rect 14408 24768 14414 24979
rect 14448 24768 14454 24979
rect 14486 24812 14496 24992
rect 14560 24812 14570 24992
rect 14312 24591 14358 24603
rect 14390 24588 14400 24768
rect 14464 24588 14474 24768
rect 14504 24603 14510 24812
rect 14544 24603 14550 24812
rect 14504 24591 14550 24603
rect 14600 24552 14804 25032
rect 15264 24979 15310 24991
rect 15264 24768 15270 24979
rect 15304 24768 15310 24979
rect 15342 24812 15352 24992
rect 15416 24812 15426 24992
rect 15456 24979 15502 24991
rect 15246 24588 15256 24768
rect 15320 24588 15330 24768
rect 15360 24603 15366 24812
rect 15400 24603 15406 24812
rect 15456 24768 15462 24979
rect 15496 24768 15502 24979
rect 15534 24812 15544 24992
rect 15608 24812 15618 24992
rect 15648 24979 15694 24991
rect 15360 24591 15406 24603
rect 15434 24588 15444 24768
rect 15508 24588 15518 24768
rect 15552 24603 15558 24812
rect 15592 24603 15598 24812
rect 15648 24768 15654 24979
rect 15688 24768 15694 24979
rect 15726 24812 15736 24992
rect 15800 24812 15810 24992
rect 15840 24979 15886 24991
rect 15552 24591 15598 24603
rect 15626 24588 15636 24768
rect 15700 24588 15710 24768
rect 15744 24603 15750 24812
rect 15784 24603 15790 24812
rect 15840 24768 15846 24979
rect 15880 24768 15886 24979
rect 15918 24812 15928 24992
rect 15992 24812 16002 24992
rect 16032 24979 16078 24991
rect 15744 24591 15790 24603
rect 15822 24588 15832 24768
rect 15896 24588 15906 24768
rect 15936 24603 15942 24812
rect 15976 24603 15982 24812
rect 16032 24768 16038 24979
rect 16072 24768 16078 24979
rect 16110 24812 16120 24992
rect 16184 24812 16194 24992
rect 16224 24979 16270 24991
rect 15936 24591 15982 24603
rect 16014 24588 16024 24768
rect 16088 24588 16098 24768
rect 16128 24603 16134 24812
rect 16168 24603 16174 24812
rect 16224 24768 16230 24979
rect 16264 24768 16270 24979
rect 16302 24812 16312 24992
rect 16376 24812 16386 24992
rect 16416 24979 16462 24991
rect 16128 24591 16174 24603
rect 16206 24588 16216 24768
rect 16280 24588 16290 24768
rect 16320 24603 16326 24812
rect 16360 24603 16366 24812
rect 16416 24768 16422 24979
rect 16456 24768 16462 24979
rect 16494 24812 16504 24992
rect 16568 24812 16578 24992
rect 16608 24979 16654 24991
rect 16320 24591 16366 24603
rect 16398 24588 16408 24768
rect 16472 24588 16482 24768
rect 16512 24603 16518 24812
rect 16552 24603 16558 24812
rect 16608 24768 16614 24979
rect 16648 24768 16654 24979
rect 16686 24812 16696 24992
rect 16760 24812 16770 24992
rect 16512 24591 16558 24603
rect 16590 24588 16600 24768
rect 16664 24588 16674 24768
rect 16704 24603 16710 24812
rect 16744 24603 16750 24812
rect 16704 24591 16750 24603
rect 16800 24552 17004 25032
rect 18270 24600 18280 25120
rect 18640 24600 18650 25120
rect 19030 25040 19040 25260
rect 19240 25040 19250 25260
rect 18904 25020 19000 25036
rect 6616 24544 8224 24552
rect 6616 24510 6634 24544
rect 6668 24510 6826 24544
rect 6860 24510 7018 24544
rect 7052 24510 7210 24544
rect 7244 24510 7402 24544
rect 7436 24510 7594 24544
rect 7628 24510 7786 24544
rect 7820 24510 8224 24544
rect 6616 24436 8224 24510
rect 8836 24544 10444 24552
rect 8836 24510 8854 24544
rect 8888 24510 9046 24544
rect 9080 24510 9238 24544
rect 9272 24510 9430 24544
rect 9464 24510 9622 24544
rect 9656 24510 9814 24544
rect 9848 24510 10006 24544
rect 10040 24510 10444 24544
rect 8836 24436 10444 24510
rect 6616 24402 6634 24436
rect 6668 24402 6826 24436
rect 6860 24402 7018 24436
rect 7052 24402 7210 24436
rect 7244 24402 7402 24436
rect 7436 24402 7594 24436
rect 7628 24402 7786 24436
rect 7820 24402 8156 24436
rect 6616 24396 8156 24402
rect 6484 24343 6530 24355
rect 6484 24132 6490 24343
rect 6524 24132 6530 24343
rect 6562 24176 6572 24356
rect 6636 24176 6646 24356
rect 6676 24343 6722 24355
rect 6466 23952 6476 24132
rect 6540 23952 6550 24132
rect 6580 23967 6586 24176
rect 6620 23967 6626 24176
rect 6676 24132 6682 24343
rect 6716 24132 6722 24343
rect 6754 24176 6764 24356
rect 6828 24176 6838 24356
rect 6868 24343 6914 24355
rect 6580 23955 6626 23967
rect 6654 23952 6664 24132
rect 6728 23952 6738 24132
rect 6772 23967 6778 24176
rect 6812 23967 6818 24176
rect 6868 24132 6874 24343
rect 6908 24132 6914 24343
rect 6946 24176 6956 24356
rect 7020 24176 7030 24356
rect 7060 24343 7106 24355
rect 6772 23955 6818 23967
rect 6846 23952 6856 24132
rect 6920 23952 6930 24132
rect 6964 23967 6970 24176
rect 7004 23967 7010 24176
rect 7060 24132 7066 24343
rect 7100 24132 7106 24343
rect 7138 24176 7148 24356
rect 7212 24176 7222 24356
rect 7252 24343 7298 24355
rect 6964 23955 7010 23967
rect 7042 23952 7052 24132
rect 7116 23952 7126 24132
rect 7156 23967 7162 24176
rect 7196 23967 7202 24176
rect 7252 24132 7258 24343
rect 7292 24132 7298 24343
rect 7330 24176 7340 24356
rect 7404 24176 7414 24356
rect 7444 24343 7490 24355
rect 7156 23955 7202 23967
rect 7234 23952 7244 24132
rect 7308 23952 7318 24132
rect 7348 23967 7354 24176
rect 7388 23967 7394 24176
rect 7444 24132 7450 24343
rect 7484 24132 7490 24343
rect 7522 24176 7532 24356
rect 7596 24176 7606 24356
rect 7636 24343 7682 24355
rect 7348 23955 7394 23967
rect 7426 23952 7436 24132
rect 7500 23952 7510 24132
rect 7540 23967 7546 24176
rect 7580 23967 7586 24176
rect 7636 24132 7642 24343
rect 7676 24132 7682 24343
rect 7714 24176 7724 24356
rect 7788 24176 7798 24356
rect 7828 24343 7874 24355
rect 7540 23955 7586 23967
rect 7618 23952 7628 24132
rect 7692 23952 7702 24132
rect 7732 23967 7738 24176
rect 7772 23967 7778 24176
rect 7828 24132 7834 24343
rect 7868 24132 7874 24343
rect 7906 24176 7916 24356
rect 7980 24176 7990 24356
rect 8020 24212 8156 24396
rect 8328 24212 8338 24436
rect 8836 24402 8854 24436
rect 8888 24402 9046 24436
rect 9080 24402 9238 24436
rect 9272 24402 9430 24436
rect 9464 24402 9622 24436
rect 9656 24402 9814 24436
rect 9848 24402 10006 24436
rect 10040 24402 10444 24436
rect 8836 24396 10444 24402
rect 11016 24544 12624 24552
rect 11016 24510 11034 24544
rect 11068 24510 11226 24544
rect 11260 24510 11418 24544
rect 11452 24510 11610 24544
rect 11644 24510 11802 24544
rect 11836 24510 11994 24544
rect 12028 24510 12186 24544
rect 12220 24510 12624 24544
rect 11016 24436 12624 24510
rect 11016 24402 11034 24436
rect 11068 24402 11226 24436
rect 11260 24402 11418 24436
rect 11452 24402 11610 24436
rect 11644 24402 11802 24436
rect 11836 24402 11994 24436
rect 12028 24402 12186 24436
rect 12220 24402 12624 24436
rect 11016 24396 12624 24402
rect 13196 24544 14804 24552
rect 13196 24510 13214 24544
rect 13248 24510 13406 24544
rect 13440 24510 13598 24544
rect 13632 24510 13790 24544
rect 13824 24510 13982 24544
rect 14016 24510 14174 24544
rect 14208 24510 14366 24544
rect 14400 24510 14804 24544
rect 13196 24436 14804 24510
rect 13196 24402 13214 24436
rect 13248 24402 13406 24436
rect 13440 24402 13598 24436
rect 13632 24402 13790 24436
rect 13824 24402 13982 24436
rect 14016 24402 14174 24436
rect 14208 24402 14366 24436
rect 14400 24402 14804 24436
rect 13196 24396 14804 24402
rect 15396 24544 17004 24552
rect 15396 24510 15414 24544
rect 15448 24510 15606 24544
rect 15640 24510 15798 24544
rect 15832 24510 15990 24544
rect 16024 24510 16182 24544
rect 16216 24510 16374 24544
rect 16408 24510 16566 24544
rect 16600 24510 17004 24544
rect 15396 24436 17004 24510
rect 15396 24402 15414 24436
rect 15448 24402 15606 24436
rect 15640 24402 15798 24436
rect 15832 24402 15990 24436
rect 16024 24402 16182 24436
rect 16216 24402 16374 24436
rect 16408 24402 16566 24436
rect 16600 24402 17004 24436
rect 15396 24396 17004 24402
rect 8704 24343 8750 24355
rect 7732 23955 7778 23967
rect 7810 23952 7820 24132
rect 7884 23952 7894 24132
rect 7924 23967 7930 24176
rect 7964 23967 7970 24176
rect 7924 23955 7970 23967
rect 8020 23916 8224 24212
rect 8704 24132 8710 24343
rect 8744 24132 8750 24343
rect 8782 24176 8792 24356
rect 8856 24176 8866 24356
rect 8896 24343 8942 24355
rect 8686 23952 8696 24132
rect 8760 23952 8770 24132
rect 8800 23967 8806 24176
rect 8840 23967 8846 24176
rect 8896 24132 8902 24343
rect 8936 24132 8942 24343
rect 8974 24176 8984 24356
rect 9048 24176 9058 24356
rect 9088 24343 9134 24355
rect 8800 23955 8846 23967
rect 8874 23952 8884 24132
rect 8948 23952 8958 24132
rect 8992 23967 8998 24176
rect 9032 23967 9038 24176
rect 9088 24132 9094 24343
rect 9128 24132 9134 24343
rect 9166 24176 9176 24356
rect 9240 24176 9250 24356
rect 9280 24343 9326 24355
rect 8992 23955 9038 23967
rect 9066 23952 9076 24132
rect 9140 23952 9150 24132
rect 9184 23967 9190 24176
rect 9224 23967 9230 24176
rect 9280 24132 9286 24343
rect 9320 24132 9326 24343
rect 9358 24176 9368 24356
rect 9432 24176 9442 24356
rect 9472 24343 9518 24355
rect 9184 23955 9230 23967
rect 9262 23952 9272 24132
rect 9336 23952 9346 24132
rect 9376 23967 9382 24176
rect 9416 23967 9422 24176
rect 9472 24132 9478 24343
rect 9512 24132 9518 24343
rect 9550 24176 9560 24356
rect 9624 24176 9634 24356
rect 9664 24343 9710 24355
rect 9376 23955 9422 23967
rect 9454 23952 9464 24132
rect 9528 23952 9538 24132
rect 9568 23967 9574 24176
rect 9608 23967 9614 24176
rect 9664 24132 9670 24343
rect 9704 24132 9710 24343
rect 9742 24176 9752 24356
rect 9816 24176 9826 24356
rect 9856 24343 9902 24355
rect 9568 23955 9614 23967
rect 9646 23952 9656 24132
rect 9720 23952 9730 24132
rect 9760 23967 9766 24176
rect 9800 23967 9806 24176
rect 9856 24132 9862 24343
rect 9896 24132 9902 24343
rect 9934 24176 9944 24356
rect 10008 24176 10018 24356
rect 10048 24343 10094 24355
rect 9760 23955 9806 23967
rect 9838 23952 9848 24132
rect 9912 23952 9922 24132
rect 9952 23967 9958 24176
rect 9992 23967 9998 24176
rect 10048 24132 10054 24343
rect 10088 24132 10094 24343
rect 10126 24176 10136 24356
rect 10200 24176 10210 24356
rect 9952 23955 9998 23967
rect 10030 23952 10040 24132
rect 10104 23952 10114 24132
rect 10144 23967 10150 24176
rect 10184 23967 10190 24176
rect 10144 23955 10190 23967
rect 10240 23916 10444 24396
rect 10884 24343 10930 24355
rect 10884 24132 10890 24343
rect 10924 24132 10930 24343
rect 10962 24176 10972 24356
rect 11036 24176 11046 24356
rect 11076 24343 11122 24355
rect 10866 23952 10876 24132
rect 10940 23952 10950 24132
rect 10980 23967 10986 24176
rect 11020 23967 11026 24176
rect 11076 24132 11082 24343
rect 11116 24132 11122 24343
rect 11154 24176 11164 24356
rect 11228 24176 11238 24356
rect 11268 24343 11314 24355
rect 10980 23955 11026 23967
rect 11054 23952 11064 24132
rect 11128 23952 11138 24132
rect 11172 23967 11178 24176
rect 11212 23967 11218 24176
rect 11268 24132 11274 24343
rect 11308 24132 11314 24343
rect 11346 24176 11356 24356
rect 11420 24176 11430 24356
rect 11460 24343 11506 24355
rect 11172 23955 11218 23967
rect 11246 23952 11256 24132
rect 11320 23952 11330 24132
rect 11364 23967 11370 24176
rect 11404 23967 11410 24176
rect 11460 24132 11466 24343
rect 11500 24132 11506 24343
rect 11538 24176 11548 24356
rect 11612 24176 11622 24356
rect 11652 24343 11698 24355
rect 11364 23955 11410 23967
rect 11442 23952 11452 24132
rect 11516 23952 11526 24132
rect 11556 23967 11562 24176
rect 11596 23967 11602 24176
rect 11652 24132 11658 24343
rect 11692 24132 11698 24343
rect 11730 24176 11740 24356
rect 11804 24176 11814 24356
rect 11844 24343 11890 24355
rect 11556 23955 11602 23967
rect 11634 23952 11644 24132
rect 11708 23952 11718 24132
rect 11748 23967 11754 24176
rect 11788 23967 11794 24176
rect 11844 24132 11850 24343
rect 11884 24132 11890 24343
rect 11922 24176 11932 24356
rect 11996 24176 12006 24356
rect 12036 24343 12082 24355
rect 11748 23955 11794 23967
rect 11826 23952 11836 24132
rect 11900 23952 11910 24132
rect 11940 23967 11946 24176
rect 11980 23967 11986 24176
rect 12036 24132 12042 24343
rect 12076 24132 12082 24343
rect 12114 24176 12124 24356
rect 12188 24176 12198 24356
rect 12228 24343 12274 24355
rect 11940 23955 11986 23967
rect 12018 23952 12028 24132
rect 12092 23952 12102 24132
rect 12132 23967 12138 24176
rect 12172 23967 12178 24176
rect 12228 24132 12234 24343
rect 12268 24132 12274 24343
rect 12306 24176 12316 24356
rect 12380 24176 12390 24356
rect 12132 23955 12178 23967
rect 12210 23952 12220 24132
rect 12284 23952 12294 24132
rect 12324 23967 12330 24176
rect 12364 23967 12370 24176
rect 12324 23955 12370 23967
rect 12420 23916 12624 24396
rect 13064 24343 13110 24355
rect 13064 24132 13070 24343
rect 13104 24132 13110 24343
rect 13142 24176 13152 24356
rect 13216 24176 13226 24356
rect 13256 24343 13302 24355
rect 13046 23952 13056 24132
rect 13120 23952 13130 24132
rect 13160 23967 13166 24176
rect 13200 23967 13206 24176
rect 13256 24132 13262 24343
rect 13296 24132 13302 24343
rect 13334 24176 13344 24356
rect 13408 24176 13418 24356
rect 13448 24343 13494 24355
rect 13160 23955 13206 23967
rect 13234 23952 13244 24132
rect 13308 23952 13318 24132
rect 13352 23967 13358 24176
rect 13392 23967 13398 24176
rect 13448 24132 13454 24343
rect 13488 24132 13494 24343
rect 13526 24176 13536 24356
rect 13600 24176 13610 24356
rect 13640 24343 13686 24355
rect 13352 23955 13398 23967
rect 13426 23952 13436 24132
rect 13500 23952 13510 24132
rect 13544 23967 13550 24176
rect 13584 23967 13590 24176
rect 13640 24132 13646 24343
rect 13680 24132 13686 24343
rect 13718 24176 13728 24356
rect 13792 24176 13802 24356
rect 13832 24343 13878 24355
rect 13544 23955 13590 23967
rect 13622 23952 13632 24132
rect 13696 23952 13706 24132
rect 13736 23967 13742 24176
rect 13776 23967 13782 24176
rect 13832 24132 13838 24343
rect 13872 24132 13878 24343
rect 13910 24176 13920 24356
rect 13984 24176 13994 24356
rect 14024 24343 14070 24355
rect 13736 23955 13782 23967
rect 13814 23952 13824 24132
rect 13888 23952 13898 24132
rect 13928 23967 13934 24176
rect 13968 23967 13974 24176
rect 14024 24132 14030 24343
rect 14064 24132 14070 24343
rect 14102 24176 14112 24356
rect 14176 24176 14186 24356
rect 14216 24343 14262 24355
rect 13928 23955 13974 23967
rect 14006 23952 14016 24132
rect 14080 23952 14090 24132
rect 14120 23967 14126 24176
rect 14160 23967 14166 24176
rect 14216 24132 14222 24343
rect 14256 24132 14262 24343
rect 14294 24176 14304 24356
rect 14368 24176 14378 24356
rect 14408 24343 14454 24355
rect 14120 23955 14166 23967
rect 14198 23952 14208 24132
rect 14272 23952 14282 24132
rect 14312 23967 14318 24176
rect 14352 23967 14358 24176
rect 14408 24132 14414 24343
rect 14448 24132 14454 24343
rect 14486 24176 14496 24356
rect 14560 24176 14570 24356
rect 14312 23955 14358 23967
rect 14390 23952 14400 24132
rect 14464 23952 14474 24132
rect 14504 23967 14510 24176
rect 14544 23967 14550 24176
rect 14504 23955 14550 23967
rect 14600 23916 14804 24396
rect 15264 24343 15310 24355
rect 15264 24132 15270 24343
rect 15304 24132 15310 24343
rect 15342 24176 15352 24356
rect 15416 24176 15426 24356
rect 15456 24343 15502 24355
rect 15246 23952 15256 24132
rect 15320 23952 15330 24132
rect 15360 23967 15366 24176
rect 15400 23967 15406 24176
rect 15456 24132 15462 24343
rect 15496 24132 15502 24343
rect 15534 24176 15544 24356
rect 15608 24176 15618 24356
rect 15648 24343 15694 24355
rect 15360 23955 15406 23967
rect 15434 23952 15444 24132
rect 15508 23952 15518 24132
rect 15552 23967 15558 24176
rect 15592 23967 15598 24176
rect 15648 24132 15654 24343
rect 15688 24132 15694 24343
rect 15726 24176 15736 24356
rect 15800 24176 15810 24356
rect 15840 24343 15886 24355
rect 15552 23955 15598 23967
rect 15626 23952 15636 24132
rect 15700 23952 15710 24132
rect 15744 23967 15750 24176
rect 15784 23967 15790 24176
rect 15840 24132 15846 24343
rect 15880 24132 15886 24343
rect 15918 24176 15928 24356
rect 15992 24176 16002 24356
rect 16032 24343 16078 24355
rect 15744 23955 15790 23967
rect 15822 23952 15832 24132
rect 15896 23952 15906 24132
rect 15936 23967 15942 24176
rect 15976 23967 15982 24176
rect 16032 24132 16038 24343
rect 16072 24132 16078 24343
rect 16110 24176 16120 24356
rect 16184 24176 16194 24356
rect 16224 24343 16270 24355
rect 15936 23955 15982 23967
rect 16014 23952 16024 24132
rect 16088 23952 16098 24132
rect 16128 23967 16134 24176
rect 16168 23967 16174 24176
rect 16224 24132 16230 24343
rect 16264 24132 16270 24343
rect 16302 24176 16312 24356
rect 16376 24176 16386 24356
rect 16416 24343 16462 24355
rect 16128 23955 16174 23967
rect 16206 23952 16216 24132
rect 16280 23952 16290 24132
rect 16320 23967 16326 24176
rect 16360 23967 16366 24176
rect 16416 24132 16422 24343
rect 16456 24132 16462 24343
rect 16494 24176 16504 24356
rect 16568 24176 16578 24356
rect 16608 24343 16654 24355
rect 16320 23955 16366 23967
rect 16398 23952 16408 24132
rect 16472 23952 16482 24132
rect 16512 23967 16518 24176
rect 16552 23967 16558 24176
rect 16608 24132 16614 24343
rect 16648 24132 16654 24343
rect 16686 24176 16696 24356
rect 16760 24176 16770 24356
rect 16512 23955 16558 23967
rect 16590 23952 16600 24132
rect 16664 23952 16674 24132
rect 16704 23967 16710 24176
rect 16744 23967 16750 24176
rect 16704 23955 16750 23967
rect 16800 23916 17004 24396
rect 6520 23908 8224 23916
rect 6520 23874 6538 23908
rect 6572 23874 6730 23908
rect 6764 23874 6922 23908
rect 6956 23874 7114 23908
rect 7148 23874 7306 23908
rect 7340 23874 7498 23908
rect 7532 23874 7690 23908
rect 7724 23874 7882 23908
rect 7916 23874 8224 23908
rect 6520 23820 8224 23874
rect 8740 23908 10444 23916
rect 8740 23874 8758 23908
rect 8792 23874 8950 23908
rect 8984 23874 9142 23908
rect 9176 23874 9334 23908
rect 9368 23874 9526 23908
rect 9560 23874 9718 23908
rect 9752 23874 9910 23908
rect 9944 23874 10102 23908
rect 10136 23874 10444 23908
rect 8740 23820 10444 23874
rect 10920 23908 12624 23916
rect 10920 23874 10938 23908
rect 10972 23874 11130 23908
rect 11164 23874 11322 23908
rect 11356 23874 11514 23908
rect 11548 23874 11706 23908
rect 11740 23874 11898 23908
rect 11932 23874 12090 23908
rect 12124 23874 12282 23908
rect 12316 23874 12624 23908
rect 10920 23820 12624 23874
rect 13100 23908 14804 23916
rect 13100 23874 13118 23908
rect 13152 23874 13310 23908
rect 13344 23874 13502 23908
rect 13536 23874 13694 23908
rect 13728 23874 13886 23908
rect 13920 23874 14078 23908
rect 14112 23874 14270 23908
rect 14304 23874 14462 23908
rect 14496 23874 14804 23908
rect 13100 23820 14804 23874
rect 15300 23908 17004 23916
rect 15300 23874 15318 23908
rect 15352 23874 15510 23908
rect 15544 23874 15702 23908
rect 15736 23874 15894 23908
rect 15928 23874 16086 23908
rect 16120 23874 16278 23908
rect 16312 23874 16470 23908
rect 16504 23874 16662 23908
rect 16696 23874 17004 23908
rect 15300 23820 17004 23874
rect 6600 23494 7752 23536
rect 6600 23460 6754 23494
rect 6788 23460 6946 23494
rect 6980 23460 7138 23494
rect 7172 23460 7330 23494
rect 7364 23460 7522 23494
rect 7556 23460 7752 23494
rect 6600 23456 7752 23460
rect 8320 23494 9472 23536
rect 8320 23460 8474 23494
rect 8508 23460 8666 23494
rect 8700 23460 8858 23494
rect 8892 23460 9050 23494
rect 9084 23460 9242 23494
rect 9276 23460 9472 23494
rect 8320 23456 9472 23460
rect 6742 23454 6800 23456
rect 6934 23454 6992 23456
rect 7126 23454 7184 23456
rect 7318 23454 7376 23456
rect 7510 23454 7568 23456
rect 6604 23410 6650 23422
rect 6604 23200 6610 23410
rect 6644 23200 6650 23410
rect 6686 23244 6696 23424
rect 6748 23244 6758 23424
rect 6796 23410 6842 23422
rect 6590 23020 6600 23200
rect 6652 23020 6662 23200
rect 6700 23034 6706 23244
rect 6740 23034 6746 23244
rect 6796 23200 6802 23410
rect 6836 23200 6842 23410
rect 6878 23244 6888 23424
rect 6940 23244 6950 23424
rect 6988 23410 7034 23422
rect 6700 23022 6746 23034
rect 6782 23020 6792 23200
rect 6844 23020 6854 23200
rect 6892 23034 6898 23244
rect 6932 23034 6938 23244
rect 6988 23200 6994 23410
rect 7028 23200 7034 23410
rect 7070 23244 7080 23424
rect 7132 23244 7142 23424
rect 7180 23410 7226 23422
rect 6892 23022 6938 23034
rect 6974 23020 6984 23200
rect 7036 23020 7046 23200
rect 7084 23034 7090 23244
rect 7124 23034 7130 23244
rect 7180 23200 7186 23410
rect 7220 23200 7226 23410
rect 7262 23244 7272 23424
rect 7324 23244 7334 23424
rect 7372 23410 7418 23422
rect 7084 23022 7130 23034
rect 7166 23020 7176 23200
rect 7228 23020 7238 23200
rect 7276 23034 7282 23244
rect 7316 23034 7322 23244
rect 7372 23200 7378 23410
rect 7412 23200 7418 23410
rect 7454 23244 7464 23424
rect 7516 23244 7526 23424
rect 7564 23410 7610 23422
rect 7276 23022 7322 23034
rect 7358 23020 7368 23200
rect 7420 23020 7430 23200
rect 7468 23034 7474 23244
rect 7508 23034 7514 23244
rect 7564 23200 7570 23410
rect 7604 23200 7610 23410
rect 7468 23022 7514 23034
rect 7550 23020 7560 23200
rect 7612 23020 7622 23200
rect 6646 22984 6704 22990
rect 6838 22984 6896 22990
rect 7030 22984 7088 22990
rect 7222 22984 7280 22990
rect 7414 22984 7472 22990
rect 7652 22984 7752 23456
rect 8462 23454 8520 23456
rect 8654 23454 8712 23456
rect 8846 23454 8904 23456
rect 9038 23454 9096 23456
rect 9230 23454 9288 23456
rect 8324 23410 8370 23422
rect 8324 23200 8330 23410
rect 8364 23200 8370 23410
rect 8406 23244 8416 23424
rect 8468 23244 8478 23424
rect 8516 23410 8562 23422
rect 8310 23020 8320 23200
rect 8372 23020 8382 23200
rect 8420 23034 8426 23244
rect 8460 23034 8466 23244
rect 8516 23200 8522 23410
rect 8556 23200 8562 23410
rect 8598 23244 8608 23424
rect 8660 23244 8670 23424
rect 8708 23410 8754 23422
rect 8420 23022 8466 23034
rect 8502 23020 8512 23200
rect 8564 23020 8574 23200
rect 8612 23034 8618 23244
rect 8652 23034 8658 23244
rect 8708 23200 8714 23410
rect 8748 23200 8754 23410
rect 8790 23244 8800 23424
rect 8852 23244 8862 23424
rect 8900 23410 8946 23422
rect 8612 23022 8658 23034
rect 8694 23020 8704 23200
rect 8756 23020 8766 23200
rect 8804 23034 8810 23244
rect 8844 23034 8850 23244
rect 8900 23200 8906 23410
rect 8940 23200 8946 23410
rect 8982 23244 8992 23424
rect 9044 23244 9054 23424
rect 9092 23410 9138 23422
rect 8804 23022 8850 23034
rect 8886 23020 8896 23200
rect 8948 23020 8958 23200
rect 8996 23034 9002 23244
rect 9036 23034 9042 23244
rect 9092 23200 9098 23410
rect 9132 23200 9138 23410
rect 9174 23244 9184 23424
rect 9236 23244 9246 23424
rect 9284 23410 9330 23422
rect 8996 23022 9042 23034
rect 9078 23020 9088 23200
rect 9140 23020 9150 23200
rect 9188 23034 9194 23244
rect 9228 23034 9234 23244
rect 9284 23200 9290 23410
rect 9324 23200 9330 23410
rect 9188 23022 9234 23034
rect 9270 23020 9280 23200
rect 9332 23020 9342 23200
rect 8366 22984 8424 22990
rect 8558 22984 8616 22990
rect 8750 22984 8808 22990
rect 8942 22984 9000 22990
rect 9134 22984 9192 22990
rect 9372 22984 9472 23456
rect 18318 23420 18328 23852
rect 18688 23420 18698 23852
rect 18904 23452 18958 25020
rect 18992 23452 19000 25020
rect 18904 23156 19000 23452
rect 19280 25020 19376 25032
rect 19280 23452 19286 25020
rect 19320 23452 19376 25020
rect 19034 23364 19044 23448
rect 19232 23364 19242 23448
rect 18892 23148 19000 23156
rect 19280 23148 19376 23452
rect 6636 22950 6658 22984
rect 6692 22950 6850 22984
rect 6884 22950 7042 22984
rect 7076 22950 7234 22984
rect 7268 22950 7426 22984
rect 7460 22950 7752 22984
rect 6636 22876 7752 22950
rect 6636 22842 6658 22876
rect 6692 22842 6850 22876
rect 6884 22842 7042 22876
rect 7076 22842 7234 22876
rect 7268 22842 7426 22876
rect 7460 22842 7752 22876
rect 6636 22840 7752 22842
rect 8356 22950 8378 22984
rect 8412 22950 8570 22984
rect 8604 22950 8762 22984
rect 8796 22950 8954 22984
rect 8988 22950 9146 22984
rect 9180 22950 9472 22984
rect 8356 22876 9472 22950
rect 8356 22842 8378 22876
rect 8412 22842 8570 22876
rect 8604 22842 8762 22876
rect 8796 22842 8954 22876
rect 8988 22842 9146 22876
rect 9180 22842 9472 22876
rect 8356 22840 9472 22842
rect 6646 22836 6704 22840
rect 6838 22836 6896 22840
rect 7030 22836 7088 22840
rect 7222 22836 7280 22840
rect 7414 22836 7472 22840
rect 6604 22792 6650 22804
rect 6604 22584 6610 22792
rect 6644 22584 6650 22792
rect 6686 22628 6696 22808
rect 6748 22628 6758 22808
rect 6796 22792 6842 22804
rect 6590 22404 6600 22584
rect 6652 22404 6662 22584
rect 6700 22416 6706 22628
rect 6740 22416 6746 22628
rect 6796 22584 6802 22792
rect 6836 22584 6842 22792
rect 6878 22628 6888 22808
rect 6940 22628 6950 22808
rect 6988 22792 7034 22804
rect 6700 22404 6746 22416
rect 6782 22404 6792 22584
rect 6844 22404 6854 22584
rect 6892 22416 6898 22628
rect 6932 22416 6938 22628
rect 6988 22584 6994 22792
rect 7028 22584 7034 22792
rect 7070 22628 7080 22808
rect 7132 22628 7142 22808
rect 7180 22792 7226 22804
rect 6892 22404 6938 22416
rect 6974 22404 6984 22584
rect 7036 22404 7046 22584
rect 7084 22416 7090 22628
rect 7124 22416 7130 22628
rect 7180 22584 7186 22792
rect 7220 22584 7226 22792
rect 7262 22628 7272 22808
rect 7324 22628 7334 22808
rect 7372 22792 7418 22804
rect 7084 22404 7130 22416
rect 7166 22404 7176 22584
rect 7228 22404 7238 22584
rect 7276 22416 7282 22628
rect 7316 22416 7322 22628
rect 7372 22584 7378 22792
rect 7412 22584 7418 22792
rect 7454 22628 7464 22808
rect 7516 22628 7526 22808
rect 7564 22792 7610 22804
rect 7276 22404 7322 22416
rect 7358 22404 7368 22584
rect 7420 22404 7430 22584
rect 7468 22416 7474 22628
rect 7508 22416 7514 22628
rect 7564 22584 7570 22792
rect 7604 22584 7610 22792
rect 7468 22404 7514 22416
rect 7550 22404 7560 22584
rect 7612 22404 7622 22584
rect 6742 22368 6800 22372
rect 6934 22368 6992 22372
rect 7126 22368 7184 22372
rect 7318 22368 7376 22372
rect 7510 22368 7568 22372
rect 7652 22368 7752 22840
rect 8366 22836 8424 22840
rect 8558 22836 8616 22840
rect 8750 22836 8808 22840
rect 8942 22836 9000 22840
rect 9134 22836 9192 22840
rect 8324 22792 8370 22804
rect 8324 22584 8330 22792
rect 8364 22584 8370 22792
rect 8406 22628 8416 22808
rect 8468 22628 8478 22808
rect 8516 22792 8562 22804
rect 8310 22404 8320 22584
rect 8372 22404 8382 22584
rect 8420 22416 8426 22628
rect 8460 22416 8466 22628
rect 8516 22584 8522 22792
rect 8556 22584 8562 22792
rect 8598 22628 8608 22808
rect 8660 22628 8670 22808
rect 8708 22792 8754 22804
rect 8420 22404 8466 22416
rect 8502 22404 8512 22584
rect 8564 22404 8574 22584
rect 8612 22416 8618 22628
rect 8652 22416 8658 22628
rect 8708 22584 8714 22792
rect 8748 22584 8754 22792
rect 8790 22628 8800 22808
rect 8852 22628 8862 22808
rect 8900 22792 8946 22804
rect 8612 22404 8658 22416
rect 8694 22404 8704 22584
rect 8756 22404 8766 22584
rect 8804 22416 8810 22628
rect 8844 22416 8850 22628
rect 8900 22584 8906 22792
rect 8940 22584 8946 22792
rect 8982 22628 8992 22808
rect 9044 22628 9054 22808
rect 9092 22792 9138 22804
rect 8804 22404 8850 22416
rect 8886 22404 8896 22584
rect 8948 22404 8958 22584
rect 8996 22416 9002 22628
rect 9036 22416 9042 22628
rect 9092 22584 9098 22792
rect 9132 22584 9138 22792
rect 9174 22628 9184 22808
rect 9236 22628 9246 22808
rect 9284 22792 9330 22804
rect 8996 22404 9042 22416
rect 9078 22404 9088 22584
rect 9140 22404 9150 22584
rect 9188 22416 9194 22628
rect 9228 22416 9234 22628
rect 9284 22584 9290 22792
rect 9324 22584 9330 22792
rect 9188 22404 9234 22416
rect 9270 22404 9280 22584
rect 9332 22404 9342 22584
rect 8462 22368 8520 22372
rect 8654 22368 8712 22372
rect 8846 22368 8904 22372
rect 9038 22368 9096 22372
rect 9230 22368 9288 22372
rect 9372 22368 9472 22840
rect 18188 23104 19412 23148
rect 18188 23070 18454 23104
rect 18488 23070 18646 23104
rect 18680 23070 18838 23104
rect 18872 23070 19030 23104
rect 19064 23070 19222 23104
rect 19256 23070 19412 23104
rect 18188 23068 19412 23070
rect 18188 22580 18260 23068
rect 18442 23064 18500 23068
rect 18634 23064 18692 23068
rect 18826 23064 18884 23068
rect 19018 23064 19076 23068
rect 19210 23064 19268 23068
rect 18304 23011 18350 23023
rect 18304 22800 18310 23011
rect 18344 22800 18350 23011
rect 18386 22844 18396 23024
rect 18448 22844 18458 23024
rect 18496 23011 18542 23023
rect 18290 22620 18300 22800
rect 18352 22620 18362 22800
rect 18400 22635 18406 22844
rect 18440 22635 18446 22844
rect 18496 22800 18502 23011
rect 18536 22800 18542 23011
rect 18578 22844 18588 23024
rect 18640 22844 18650 23024
rect 18688 23011 18734 23023
rect 18400 22623 18446 22635
rect 18482 22620 18492 22800
rect 18544 22620 18554 22800
rect 18592 22635 18598 22844
rect 18632 22635 18638 22844
rect 18688 22800 18694 23011
rect 18728 22800 18734 23011
rect 18770 22844 18780 23024
rect 18832 22844 18842 23024
rect 18880 23011 18926 23023
rect 18592 22623 18638 22635
rect 18674 22620 18684 22800
rect 18736 22620 18746 22800
rect 18784 22635 18790 22844
rect 18824 22635 18830 22844
rect 18880 22800 18886 23011
rect 18920 22800 18926 23011
rect 18962 22844 18972 23024
rect 19024 22844 19034 23024
rect 19072 23011 19118 23023
rect 18784 22623 18830 22635
rect 18866 22620 18876 22800
rect 18928 22620 18938 22800
rect 18976 22635 18982 22844
rect 19016 22635 19022 22844
rect 19072 22800 19078 23011
rect 19112 22800 19118 23011
rect 19154 22844 19164 23024
rect 19216 22844 19226 23024
rect 19264 23011 19310 23023
rect 18976 22623 19022 22635
rect 19058 22620 19068 22800
rect 19120 22620 19130 22800
rect 19168 22635 19174 22844
rect 19208 22635 19214 22844
rect 19264 22800 19270 23011
rect 19304 22800 19310 23011
rect 19168 22623 19214 22635
rect 19250 22620 19260 22800
rect 19312 22620 19322 22800
rect 18346 22580 18404 22582
rect 18538 22580 18596 22582
rect 18730 22580 18788 22582
rect 18922 22580 18980 22582
rect 19114 22580 19172 22582
rect 18188 22576 19176 22580
rect 18188 22572 18358 22576
rect 18392 22572 18550 22576
rect 18584 22572 18742 22576
rect 18776 22572 18934 22576
rect 18188 22472 18272 22572
rect 18860 22542 18934 22572
rect 18968 22542 19126 22576
rect 19160 22542 19176 22576
rect 18860 22500 19176 22542
rect 18860 22472 18920 22500
rect 18188 22460 18920 22472
rect 6736 22366 7752 22368
rect 6736 22332 6754 22366
rect 6788 22332 6946 22366
rect 6980 22332 7138 22366
rect 7172 22332 7330 22366
rect 7364 22332 7522 22366
rect 7556 22332 7752 22366
rect 6736 22258 7752 22332
rect 6736 22224 6754 22258
rect 6788 22224 6946 22258
rect 6980 22224 7138 22258
rect 7172 22224 7330 22258
rect 7364 22224 7522 22258
rect 7556 22224 7752 22258
rect 8456 22366 9472 22368
rect 8456 22332 8474 22366
rect 8508 22332 8666 22366
rect 8700 22332 8858 22366
rect 8892 22332 9050 22366
rect 9084 22332 9242 22366
rect 9276 22332 9472 22366
rect 8456 22258 9472 22332
rect 8456 22224 8474 22258
rect 8508 22224 8666 22258
rect 8700 22224 8858 22258
rect 8892 22224 9050 22258
rect 9084 22224 9242 22258
rect 9276 22224 9472 22258
rect 6742 22218 6800 22224
rect 6934 22218 6992 22224
rect 7126 22218 7184 22224
rect 7318 22218 7376 22224
rect 7510 22218 7568 22224
rect 6604 22174 6650 22186
rect 6604 21964 6610 22174
rect 6644 21964 6650 22174
rect 6686 22008 6696 22188
rect 6748 22008 6758 22188
rect 6796 22174 6842 22186
rect 6590 21784 6600 21964
rect 6652 21784 6662 21964
rect 6700 21798 6706 22008
rect 6740 21798 6746 22008
rect 6796 21964 6802 22174
rect 6836 21964 6842 22174
rect 6878 22008 6888 22188
rect 6940 22008 6950 22188
rect 6988 22174 7034 22186
rect 6700 21786 6746 21798
rect 6782 21784 6792 21964
rect 6844 21784 6854 21964
rect 6892 21798 6898 22008
rect 6932 21798 6938 22008
rect 6988 21964 6994 22174
rect 7028 21964 7034 22174
rect 7070 22008 7080 22188
rect 7132 22008 7142 22188
rect 7180 22174 7226 22186
rect 6892 21786 6938 21798
rect 6974 21784 6984 21964
rect 7036 21784 7046 21964
rect 7084 21798 7090 22008
rect 7124 21798 7130 22008
rect 7180 21964 7186 22174
rect 7220 21964 7226 22174
rect 7262 22008 7272 22188
rect 7324 22008 7334 22188
rect 7372 22174 7418 22186
rect 7084 21786 7130 21798
rect 7166 21784 7176 21964
rect 7228 21784 7238 21964
rect 7276 21798 7282 22008
rect 7316 21798 7322 22008
rect 7372 21964 7378 22174
rect 7412 21964 7418 22174
rect 7454 22008 7464 22188
rect 7516 22008 7526 22188
rect 7564 22174 7610 22186
rect 7276 21786 7322 21798
rect 7358 21784 7368 21964
rect 7420 21784 7430 21964
rect 7468 21798 7474 22008
rect 7508 21798 7514 22008
rect 7564 21964 7570 22174
rect 7604 21964 7610 22174
rect 7468 21786 7514 21798
rect 7550 21784 7560 21964
rect 7612 21784 7622 21964
rect 6646 21748 6704 21754
rect 6838 21748 6896 21754
rect 7030 21748 7088 21754
rect 7222 21748 7280 21754
rect 7414 21748 7472 21754
rect 7652 21748 7752 22224
rect 8462 22218 8520 22224
rect 8654 22218 8712 22224
rect 8846 22218 8904 22224
rect 9038 22218 9096 22224
rect 9230 22218 9288 22224
rect 8324 22174 8370 22186
rect 8324 21964 8330 22174
rect 8364 21964 8370 22174
rect 8406 22008 8416 22188
rect 8468 22008 8478 22188
rect 8516 22174 8562 22186
rect 8310 21784 8320 21964
rect 8372 21784 8382 21964
rect 8420 21798 8426 22008
rect 8460 21798 8466 22008
rect 8516 21964 8522 22174
rect 8556 21964 8562 22174
rect 8598 22008 8608 22188
rect 8660 22008 8670 22188
rect 8708 22174 8754 22186
rect 8420 21786 8466 21798
rect 8502 21784 8512 21964
rect 8564 21784 8574 21964
rect 8612 21798 8618 22008
rect 8652 21798 8658 22008
rect 8708 21964 8714 22174
rect 8748 21964 8754 22174
rect 8790 22008 8800 22188
rect 8852 22008 8862 22188
rect 8900 22174 8946 22186
rect 8612 21786 8658 21798
rect 8694 21784 8704 21964
rect 8756 21784 8766 21964
rect 8804 21798 8810 22008
rect 8844 21798 8850 22008
rect 8900 21964 8906 22174
rect 8940 21964 8946 22174
rect 8982 22008 8992 22188
rect 9044 22008 9054 22188
rect 9092 22174 9138 22186
rect 8804 21786 8850 21798
rect 8886 21784 8896 21964
rect 8948 21784 8958 21964
rect 8996 21798 9002 22008
rect 9036 21798 9042 22008
rect 9092 21964 9098 22174
rect 9132 21964 9138 22174
rect 9174 22008 9184 22188
rect 9236 22008 9246 22188
rect 9284 22174 9330 22186
rect 8996 21786 9042 21798
rect 9078 21784 9088 21964
rect 9140 21784 9150 21964
rect 9188 21798 9194 22008
rect 9228 21798 9234 22008
rect 9284 21964 9290 22174
rect 9324 21964 9330 22174
rect 9188 21786 9234 21798
rect 9270 21784 9280 21964
rect 9332 21784 9342 21964
rect 8366 21748 8424 21754
rect 8558 21748 8616 21754
rect 8750 21748 8808 21754
rect 8942 21748 9000 21754
rect 9134 21748 9192 21754
rect 9372 21748 9472 22224
rect 6640 21714 6658 21748
rect 6692 21714 6850 21748
rect 6884 21714 7042 21748
rect 7076 21714 7234 21748
rect 7268 21714 7426 21748
rect 7460 21714 7752 21748
rect 6640 21616 7752 21714
rect 8360 21714 8378 21748
rect 8412 21714 8570 21748
rect 8604 21714 8762 21748
rect 8796 21714 8954 21748
rect 8988 21714 9146 21748
rect 9180 21714 9472 21748
rect 8360 21688 9472 21714
rect 18164 22236 19268 22336
rect 18164 22202 18454 22236
rect 18488 22202 18646 22236
rect 18680 22202 18838 22236
rect 18872 22202 19030 22236
rect 19064 22202 19222 22236
rect 19256 22202 19268 22236
rect 18164 22200 19268 22202
rect 18164 21728 18260 22200
rect 18442 22196 18500 22200
rect 18634 22196 18692 22200
rect 18826 22196 18884 22200
rect 19018 22196 19076 22200
rect 19210 22196 19268 22200
rect 18304 22152 18350 22164
rect 18304 21944 18310 22152
rect 18344 21944 18350 22152
rect 18382 21988 18392 22168
rect 18444 21988 18454 22168
rect 18496 22152 18542 22164
rect 18290 21764 18300 21944
rect 18352 21764 18362 21944
rect 18400 21776 18406 21988
rect 18440 21776 18446 21988
rect 18496 21944 18502 22152
rect 18536 21944 18542 22152
rect 18574 21988 18584 22168
rect 18636 21988 18646 22168
rect 18688 22152 18734 22164
rect 18400 21764 18446 21776
rect 18478 21764 18488 21944
rect 18540 21764 18550 21944
rect 18592 21776 18598 21988
rect 18632 21776 18638 21988
rect 18688 21944 18694 22152
rect 18728 21944 18734 22152
rect 18766 21988 18776 22168
rect 18828 21988 18838 22168
rect 18880 22152 18926 22164
rect 18592 21764 18638 21776
rect 18670 21764 18680 21944
rect 18732 21764 18742 21944
rect 18784 21776 18790 21988
rect 18824 21776 18830 21988
rect 18880 21944 18886 22152
rect 18920 21944 18926 22152
rect 18958 21988 18968 22168
rect 19020 21988 19030 22168
rect 19072 22152 19118 22164
rect 18784 21764 18830 21776
rect 18862 21764 18872 21944
rect 18924 21764 18934 21944
rect 18976 21776 18982 21988
rect 19016 21776 19022 21988
rect 19072 21944 19078 22152
rect 19112 21944 19118 22152
rect 19150 21988 19160 22168
rect 19212 21988 19222 22168
rect 19264 22152 19310 22164
rect 18976 21764 19022 21776
rect 19054 21764 19064 21944
rect 19116 21764 19126 21944
rect 19168 21776 19174 21988
rect 19208 21776 19214 21988
rect 19264 21944 19270 22152
rect 19304 21944 19310 22152
rect 19168 21764 19214 21776
rect 19246 21764 19256 21944
rect 19308 21764 19318 21944
rect 18346 21728 18404 21732
rect 18538 21728 18596 21732
rect 18730 21728 18788 21732
rect 18922 21728 18980 21732
rect 19114 21728 19172 21732
rect 18164 21726 19176 21728
rect 18164 21692 18358 21726
rect 18392 21692 18550 21726
rect 18584 21692 18742 21726
rect 18776 21692 18934 21726
rect 18968 21692 19126 21726
rect 19160 21692 19176 21726
rect 18164 21688 19176 21692
rect 8360 21618 19176 21688
rect 8360 21616 18358 21618
rect 7200 21556 7344 21616
rect 8920 21584 18358 21616
rect 18392 21584 18550 21618
rect 18584 21584 18742 21618
rect 18776 21584 18934 21618
rect 18968 21584 19126 21618
rect 19160 21584 19176 21618
rect 8920 21580 19176 21584
rect 8920 21556 18260 21580
rect 18346 21578 18404 21580
rect 18538 21578 18596 21580
rect 18730 21578 18788 21580
rect 18922 21578 18980 21580
rect 19114 21578 19172 21580
rect 7200 21460 18260 21556
rect 7200 21396 9064 21460
rect 7200 21368 7344 21396
rect 8920 21368 9064 21396
rect 6648 21348 7888 21368
rect 6648 21314 6672 21348
rect 6840 21314 6930 21348
rect 7098 21314 7188 21348
rect 7356 21314 7446 21348
rect 7614 21314 7704 21348
rect 7872 21314 7888 21348
rect 6648 21308 7888 21314
rect 8368 21348 9608 21368
rect 8368 21314 8392 21348
rect 8560 21314 8650 21348
rect 8818 21314 8908 21348
rect 9076 21314 9166 21348
rect 9334 21314 9424 21348
rect 9592 21314 9608 21348
rect 8368 21308 9608 21314
rect 6590 21096 6600 21276
rect 6652 21096 6662 21276
rect 6862 21264 6908 21276
rect 6604 20888 6610 21096
rect 6644 20888 6650 21096
rect 6862 21056 6868 21264
rect 6902 21056 6908 21264
rect 6604 20876 6650 20888
rect 6850 20876 6860 21056
rect 6912 20876 6922 21056
rect 6952 20844 7072 21308
rect 7106 21096 7116 21276
rect 7168 21096 7178 21276
rect 7120 20888 7126 21096
rect 7160 20888 7166 21096
rect 7120 20876 7166 20888
rect 7212 20844 7332 21308
rect 7378 21264 7424 21276
rect 7378 21056 7384 21264
rect 7418 21056 7424 21264
rect 7366 20876 7376 21056
rect 7428 20876 7438 21056
rect 7472 20844 7592 21308
rect 7622 21096 7632 21276
rect 7684 21096 7694 21276
rect 7894 21264 7940 21276
rect 7636 20888 7642 21096
rect 7676 20888 7682 21096
rect 7894 21056 7900 21264
rect 7934 21056 7940 21264
rect 8310 21096 8320 21276
rect 8372 21096 8382 21276
rect 8582 21264 8628 21276
rect 7636 20876 7682 20888
rect 7882 20876 7892 21056
rect 7944 20876 7954 21056
rect 8324 20888 8330 21096
rect 8364 20888 8370 21096
rect 8582 21056 8588 21264
rect 8622 21056 8628 21264
rect 8324 20876 8370 20888
rect 8570 20876 8580 21056
rect 8632 20876 8642 21056
rect 8672 20844 8792 21308
rect 8826 21096 8836 21276
rect 8888 21096 8898 21276
rect 8840 20888 8846 21096
rect 8880 20888 8886 21096
rect 8840 20876 8886 20888
rect 8932 20844 9052 21308
rect 9098 21264 9144 21276
rect 9098 21056 9104 21264
rect 9138 21056 9144 21264
rect 9086 20876 9096 21056
rect 9148 20876 9158 21056
rect 9192 20844 9312 21308
rect 9342 21096 9352 21276
rect 9404 21096 9414 21276
rect 9614 21264 9660 21276
rect 9356 20888 9362 21096
rect 9396 20888 9402 21096
rect 9614 21056 9620 21264
rect 9654 21056 9660 21264
rect 10320 21220 11900 21300
rect 9356 20876 9402 20888
rect 9602 20876 9612 21056
rect 9664 20876 9674 21056
rect 10320 20860 10380 21220
rect 10840 20860 11900 21220
rect 6648 20840 7888 20844
rect 8368 20840 9608 20844
rect 6644 20838 7888 20840
rect 6644 20804 6672 20838
rect 6840 20804 6930 20838
rect 7098 20804 7188 20838
rect 7356 20804 7446 20838
rect 7614 20804 7704 20838
rect 7872 20804 7888 20838
rect 6644 20730 7888 20804
rect 6644 20696 6672 20730
rect 6840 20696 6930 20730
rect 7098 20696 7188 20730
rect 7356 20696 7446 20730
rect 7614 20696 7704 20730
rect 7872 20696 7888 20730
rect 6644 20692 7888 20696
rect 8364 20838 9608 20840
rect 8364 20804 8392 20838
rect 8560 20804 8650 20838
rect 8818 20804 8908 20838
rect 9076 20804 9166 20838
rect 9334 20804 9424 20838
rect 9592 20804 9608 20838
rect 8364 20730 9608 20804
rect 10320 20780 11900 20860
rect 8364 20696 8392 20730
rect 8560 20696 8650 20730
rect 8818 20696 8908 20730
rect 9076 20696 9166 20730
rect 9334 20696 9424 20730
rect 9592 20696 9608 20730
rect 8364 20692 9608 20696
rect 6660 20690 6852 20692
rect 6918 20690 7110 20692
rect 7176 20690 7368 20692
rect 7434 20690 7626 20692
rect 7692 20690 7884 20692
rect 8380 20690 8572 20692
rect 8638 20690 8830 20692
rect 8896 20690 9088 20692
rect 9154 20690 9346 20692
rect 9412 20690 9604 20692
rect 6590 20480 6600 20660
rect 6652 20480 6662 20660
rect 6862 20646 6908 20658
rect 6604 20270 6610 20480
rect 6644 20270 6650 20480
rect 6862 20440 6868 20646
rect 6902 20440 6908 20646
rect 6604 20258 6650 20270
rect 6850 20260 6860 20440
rect 6912 20260 6922 20440
rect 6862 20258 6908 20260
rect 6952 20226 7072 20690
rect 7106 20480 7116 20660
rect 7168 20480 7178 20660
rect 7120 20270 7126 20480
rect 7160 20270 7166 20480
rect 7120 20258 7166 20270
rect 7212 20228 7332 20690
rect 7378 20646 7424 20658
rect 7378 20440 7384 20646
rect 7418 20440 7424 20646
rect 7366 20260 7376 20440
rect 7428 20260 7438 20440
rect 7378 20258 7424 20260
rect 7200 20226 7344 20228
rect 7472 20226 7592 20690
rect 7622 20480 7632 20660
rect 7684 20480 7694 20660
rect 7894 20646 7940 20658
rect 7636 20270 7642 20480
rect 7676 20270 7682 20480
rect 7894 20440 7900 20646
rect 7934 20440 7940 20646
rect 8310 20480 8320 20660
rect 8372 20480 8382 20660
rect 8582 20646 8628 20658
rect 7636 20258 7682 20270
rect 7882 20260 7892 20440
rect 7944 20260 7954 20440
rect 8324 20270 8330 20480
rect 8364 20270 8370 20480
rect 8582 20440 8588 20646
rect 8622 20440 8628 20646
rect 7894 20258 7940 20260
rect 8324 20258 8370 20270
rect 8570 20260 8580 20440
rect 8632 20260 8642 20440
rect 8582 20258 8628 20260
rect 8672 20226 8792 20690
rect 8826 20480 8836 20660
rect 8888 20480 8898 20660
rect 8840 20270 8846 20480
rect 8880 20270 8886 20480
rect 8840 20258 8886 20270
rect 8932 20228 9052 20690
rect 9098 20646 9144 20658
rect 9098 20440 9104 20646
rect 9138 20440 9144 20646
rect 9086 20260 9096 20440
rect 9148 20260 9158 20440
rect 9098 20258 9144 20260
rect 8920 20226 9064 20228
rect 9192 20226 9312 20690
rect 9342 20480 9352 20660
rect 9404 20480 9414 20660
rect 9614 20646 9660 20658
rect 9356 20270 9362 20480
rect 9396 20270 9402 20480
rect 9614 20440 9620 20646
rect 9654 20440 9660 20646
rect 9356 20258 9402 20270
rect 9602 20260 9612 20440
rect 9664 20260 9674 20440
rect 9614 20258 9660 20260
rect 6660 20224 6852 20226
rect 6918 20224 7110 20226
rect 7176 20224 7368 20226
rect 7434 20224 7626 20226
rect 7692 20224 7884 20226
rect 8380 20224 8572 20226
rect 8638 20224 8830 20226
rect 8896 20224 9088 20226
rect 9154 20224 9346 20226
rect 9412 20224 9604 20226
rect 6648 20220 7888 20224
rect 8368 20220 9608 20224
rect 6648 20186 6672 20220
rect 6840 20186 6930 20220
rect 7098 20186 7188 20220
rect 7356 20186 7446 20220
rect 7614 20186 7704 20220
rect 7872 20186 7892 20220
rect 6648 20112 7892 20186
rect 6648 20078 6672 20112
rect 6840 20078 6930 20112
rect 7098 20078 7188 20112
rect 7356 20078 7446 20112
rect 7614 20078 7704 20112
rect 7872 20078 7892 20112
rect 6648 20072 7892 20078
rect 8368 20186 8392 20220
rect 8560 20186 8650 20220
rect 8818 20186 8908 20220
rect 9076 20186 9166 20220
rect 9334 20186 9424 20220
rect 9592 20186 9612 20220
rect 8368 20112 9612 20186
rect 8368 20078 8392 20112
rect 8560 20078 8650 20112
rect 8818 20078 8908 20112
rect 9076 20078 9166 20112
rect 9334 20078 9424 20112
rect 9592 20078 9612 20112
rect 8368 20072 9612 20078
rect 6590 19860 6600 20040
rect 6652 19860 6662 20040
rect 6862 20028 6908 20040
rect 6604 19652 6610 19860
rect 6644 19652 6650 19860
rect 6862 19820 6868 20028
rect 6902 19820 6908 20028
rect 6604 19640 6650 19652
rect 6850 19640 6860 19820
rect 6912 19640 6922 19820
rect 6952 19608 7072 20072
rect 7106 19860 7116 20040
rect 7168 19860 7178 20040
rect 7120 19652 7126 19860
rect 7160 19652 7166 19860
rect 7120 19640 7166 19652
rect 7212 19608 7332 20072
rect 7378 20028 7424 20040
rect 7378 19820 7384 20028
rect 7418 19820 7424 20028
rect 7366 19640 7376 19820
rect 7428 19640 7438 19820
rect 7472 19608 7592 20072
rect 7622 19860 7632 20040
rect 7684 19860 7694 20040
rect 7894 20028 7940 20040
rect 7636 19652 7642 19860
rect 7676 19652 7682 19860
rect 7894 19820 7900 20028
rect 7934 19820 7940 20028
rect 8310 19860 8320 20040
rect 8372 19860 8382 20040
rect 8582 20028 8628 20040
rect 7636 19640 7682 19652
rect 7882 19640 7892 19820
rect 7944 19640 7954 19820
rect 8324 19652 8330 19860
rect 8364 19652 8370 19860
rect 8582 19820 8588 20028
rect 8622 19820 8628 20028
rect 8324 19640 8370 19652
rect 8570 19640 8580 19820
rect 8632 19640 8642 19820
rect 8672 19608 8792 20072
rect 8826 19860 8836 20040
rect 8888 19860 8898 20040
rect 8840 19652 8846 19860
rect 8880 19652 8886 19860
rect 8840 19640 8886 19652
rect 8932 19608 9052 20072
rect 9098 20028 9144 20040
rect 9098 19820 9104 20028
rect 9138 19820 9144 20028
rect 9086 19640 9096 19820
rect 9148 19640 9158 19820
rect 9192 19608 9312 20072
rect 9342 19860 9352 20040
rect 9404 19860 9414 20040
rect 9614 20028 9660 20040
rect 9356 19652 9362 19860
rect 9396 19652 9402 19860
rect 9614 19820 9620 20028
rect 9654 19820 9660 20028
rect 10024 19836 10752 19844
rect 9356 19640 9402 19652
rect 9602 19640 9612 19820
rect 9664 19640 9674 19820
rect 10024 19768 10188 19836
rect 10260 19798 10752 19836
rect 10260 19768 10314 19798
rect 10024 19764 10314 19768
rect 10348 19764 10506 19798
rect 10540 19764 10698 19798
rect 10732 19764 10752 19798
rect 10024 19756 10752 19764
rect 6648 19604 6852 19608
rect 6644 19602 6852 19604
rect 6644 19568 6672 19602
rect 6840 19572 6852 19602
rect 6918 19602 7368 19608
rect 6918 19572 6930 19602
rect 6840 19568 6930 19572
rect 7098 19568 7188 19602
rect 7356 19572 7368 19602
rect 7434 19602 7884 19608
rect 8368 19604 8572 19608
rect 7434 19572 7446 19602
rect 7356 19568 7446 19572
rect 7614 19568 7704 19602
rect 7872 19572 7884 19602
rect 8364 19602 8572 19604
rect 7872 19568 7888 19572
rect 6644 19494 7888 19568
rect 6644 19460 6672 19494
rect 6840 19460 6930 19494
rect 7098 19460 7188 19494
rect 7356 19460 7446 19494
rect 7614 19460 7704 19494
rect 7872 19460 7888 19494
rect 6644 19456 7888 19460
rect 8364 19568 8392 19602
rect 8560 19572 8572 19602
rect 8638 19602 9088 19608
rect 8638 19572 8650 19602
rect 8560 19568 8650 19572
rect 8818 19568 8908 19602
rect 9076 19572 9088 19602
rect 9154 19602 9604 19608
rect 9154 19572 9166 19602
rect 9076 19568 9166 19572
rect 9334 19568 9424 19602
rect 9592 19572 9604 19602
rect 9592 19568 9608 19572
rect 8364 19494 9608 19568
rect 8364 19460 8392 19494
rect 8560 19460 8650 19494
rect 8818 19460 8908 19494
rect 9076 19460 9166 19494
rect 9334 19460 9424 19494
rect 9592 19460 9608 19494
rect 8364 19456 9608 19460
rect 6660 19454 6852 19456
rect 6918 19454 7110 19456
rect 7176 19454 7368 19456
rect 7434 19454 7626 19456
rect 7692 19454 7884 19456
rect 8380 19454 8572 19456
rect 8638 19454 8830 19456
rect 8896 19454 9088 19456
rect 9154 19454 9346 19456
rect 9412 19454 9604 19456
rect 6590 19244 6600 19424
rect 6652 19244 6662 19424
rect 6862 19410 6908 19422
rect 6604 19034 6610 19244
rect 6644 19034 6650 19244
rect 6862 19204 6868 19410
rect 6902 19204 6908 19410
rect 6604 19022 6650 19034
rect 6850 19024 6860 19204
rect 6912 19024 6922 19204
rect 6862 19022 6908 19024
rect 6952 18990 7072 19454
rect 7200 19452 7344 19454
rect 7106 19244 7116 19424
rect 7168 19244 7178 19424
rect 7120 19034 7126 19244
rect 7160 19034 7166 19244
rect 7120 19022 7166 19034
rect 7212 18990 7332 19452
rect 7378 19410 7424 19422
rect 7378 19204 7384 19410
rect 7418 19204 7424 19410
rect 7366 19024 7376 19204
rect 7428 19024 7438 19204
rect 7378 19022 7424 19024
rect 7472 18990 7592 19454
rect 7622 19244 7632 19424
rect 7684 19244 7694 19424
rect 7894 19410 7940 19422
rect 7636 19034 7642 19244
rect 7676 19034 7682 19244
rect 7894 19204 7900 19410
rect 7934 19204 7940 19410
rect 8310 19244 8320 19424
rect 8372 19244 8382 19424
rect 8582 19410 8628 19422
rect 7636 19022 7682 19034
rect 7882 19024 7892 19204
rect 7944 19024 7954 19204
rect 8324 19034 8330 19244
rect 8364 19034 8370 19244
rect 8582 19204 8588 19410
rect 8622 19204 8628 19410
rect 7894 19022 7940 19024
rect 8324 19022 8370 19034
rect 8570 19024 8580 19204
rect 8632 19024 8642 19204
rect 8582 19022 8628 19024
rect 8672 18990 8792 19454
rect 8920 19452 9064 19454
rect 8826 19244 8836 19424
rect 8888 19244 8898 19424
rect 8840 19034 8846 19244
rect 8880 19034 8886 19244
rect 8840 19022 8886 19034
rect 8932 18990 9052 19452
rect 9098 19410 9144 19422
rect 9098 19204 9104 19410
rect 9138 19204 9144 19410
rect 9086 19024 9096 19204
rect 9148 19024 9158 19204
rect 9098 19022 9144 19024
rect 9192 18990 9312 19454
rect 9342 19244 9352 19424
rect 9404 19244 9414 19424
rect 9614 19410 9660 19422
rect 9356 19034 9362 19244
rect 9396 19034 9402 19244
rect 9614 19204 9620 19410
rect 9654 19204 9660 19410
rect 10024 19296 10120 19756
rect 10164 19714 10210 19726
rect 10164 19504 10170 19714
rect 10204 19504 10210 19714
rect 10242 19548 10252 19728
rect 10312 19548 10322 19728
rect 10356 19714 10402 19726
rect 10150 19324 10160 19504
rect 10220 19324 10230 19504
rect 10260 19338 10266 19548
rect 10300 19338 10306 19548
rect 10356 19504 10362 19714
rect 10396 19504 10402 19714
rect 10434 19548 10444 19728
rect 10504 19548 10514 19728
rect 10548 19714 10594 19726
rect 10260 19326 10306 19338
rect 10338 19324 10348 19504
rect 10408 19324 10418 19504
rect 10452 19338 10458 19548
rect 10492 19338 10498 19548
rect 10548 19504 10554 19714
rect 10588 19504 10594 19714
rect 10626 19548 10636 19728
rect 10696 19548 10706 19728
rect 10740 19714 10786 19726
rect 10452 19326 10498 19338
rect 10530 19324 10540 19504
rect 10600 19324 10610 19504
rect 10644 19338 10650 19548
rect 10684 19338 10690 19548
rect 10740 19504 10746 19714
rect 10780 19504 10786 19714
rect 10818 19548 10828 19728
rect 10888 19548 10898 19728
rect 10644 19326 10690 19338
rect 10722 19324 10732 19504
rect 10792 19324 10802 19504
rect 10836 19338 10842 19548
rect 10876 19338 10882 19548
rect 10836 19326 10882 19338
rect 10024 19288 10844 19296
rect 10024 19254 10218 19288
rect 10252 19254 10410 19288
rect 10444 19254 10602 19288
rect 10636 19254 10794 19288
rect 10828 19254 10844 19288
rect 10024 19216 10844 19254
rect 9356 19022 9402 19034
rect 9602 19024 9612 19204
rect 9664 19024 9674 19204
rect 9614 19022 9660 19024
rect 6660 18988 6852 18990
rect 6918 18988 7110 18990
rect 7176 18988 7368 18990
rect 7434 18988 7626 18990
rect 7692 18988 7884 18990
rect 8380 18988 8572 18990
rect 8638 18988 8830 18990
rect 8896 18988 9088 18990
rect 9154 18988 9346 18990
rect 9412 18988 9604 18990
rect 6648 18984 7888 18988
rect 8368 18984 9608 18988
rect 6648 18950 6672 18984
rect 6840 18950 6930 18984
rect 7098 18950 7188 18984
rect 7356 18950 7446 18984
rect 7614 18950 7704 18984
rect 7872 18950 7892 18984
rect 6648 18876 7892 18950
rect 6648 18842 6672 18876
rect 6840 18842 6930 18876
rect 7098 18842 7188 18876
rect 7356 18842 7446 18876
rect 7614 18842 7704 18876
rect 7872 18842 7892 18876
rect 6648 18836 7892 18842
rect 8368 18950 8392 18984
rect 8560 18950 8650 18984
rect 8818 18950 8908 18984
rect 9076 18950 9166 18984
rect 9334 18950 9424 18984
rect 9592 18950 9612 18984
rect 8368 18876 9612 18950
rect 8368 18842 8392 18876
rect 8560 18842 8650 18876
rect 8818 18842 8908 18876
rect 9076 18842 9166 18876
rect 9334 18842 9424 18876
rect 9592 18842 9612 18876
rect 8368 18836 9612 18842
rect 10024 18876 11044 18924
rect 10024 18842 10218 18876
rect 10252 18842 10410 18876
rect 10444 18842 10602 18876
rect 10636 18842 10794 18876
rect 10828 18842 10986 18876
rect 11020 18842 11044 18876
rect 10024 18836 11044 18842
rect 6590 18624 6600 18804
rect 6652 18624 6662 18804
rect 6862 18792 6908 18804
rect 6604 18416 6610 18624
rect 6644 18416 6650 18624
rect 6862 18584 6868 18792
rect 6902 18584 6908 18792
rect 6604 18404 6650 18416
rect 6850 18404 6860 18584
rect 6912 18404 6922 18584
rect 6952 18372 7072 18836
rect 7106 18624 7116 18804
rect 7168 18624 7178 18804
rect 7120 18416 7126 18624
rect 7160 18416 7166 18624
rect 7120 18404 7166 18416
rect 7212 18372 7332 18836
rect 7378 18792 7424 18804
rect 7378 18584 7384 18792
rect 7418 18584 7424 18792
rect 7366 18404 7376 18584
rect 7428 18404 7438 18584
rect 7472 18372 7592 18836
rect 7622 18624 7632 18804
rect 7684 18624 7694 18804
rect 7894 18792 7940 18804
rect 7636 18416 7642 18624
rect 7676 18416 7682 18624
rect 7894 18584 7900 18792
rect 7934 18584 7940 18792
rect 8310 18624 8320 18804
rect 8372 18624 8382 18804
rect 8582 18792 8628 18804
rect 7636 18404 7682 18416
rect 7882 18404 7892 18584
rect 7944 18404 7954 18584
rect 8324 18416 8330 18624
rect 8364 18416 8370 18624
rect 8582 18584 8588 18792
rect 8622 18584 8628 18792
rect 8324 18404 8370 18416
rect 8570 18404 8580 18584
rect 8632 18404 8642 18584
rect 8672 18372 8792 18836
rect 8826 18624 8836 18804
rect 8888 18624 8898 18804
rect 8840 18416 8846 18624
rect 8880 18416 8886 18624
rect 8840 18404 8886 18416
rect 8932 18372 9052 18836
rect 9098 18792 9144 18804
rect 9098 18584 9104 18792
rect 9138 18584 9144 18792
rect 9086 18404 9096 18584
rect 9148 18404 9158 18584
rect 9192 18372 9312 18836
rect 9342 18624 9352 18804
rect 9404 18624 9414 18804
rect 9614 18792 9660 18804
rect 9356 18416 9362 18624
rect 9396 18416 9402 18624
rect 9614 18584 9620 18792
rect 9654 18584 9660 18792
rect 9356 18404 9402 18416
rect 9602 18404 9612 18584
rect 9664 18404 9674 18584
rect 10024 18372 10120 18836
rect 10164 18792 10210 18804
rect 10164 18584 10170 18792
rect 10204 18584 10210 18792
rect 10242 18624 10252 18804
rect 10312 18624 10322 18804
rect 10356 18792 10402 18804
rect 10150 18404 10160 18584
rect 10220 18404 10230 18584
rect 10260 18416 10266 18624
rect 10300 18416 10306 18624
rect 10356 18584 10362 18792
rect 10396 18584 10402 18792
rect 10434 18624 10444 18804
rect 10504 18624 10514 18804
rect 10548 18792 10594 18804
rect 10260 18404 10306 18416
rect 10338 18404 10348 18584
rect 10408 18404 10418 18584
rect 10452 18416 10458 18624
rect 10492 18416 10498 18624
rect 10548 18584 10554 18792
rect 10588 18584 10594 18792
rect 10626 18624 10636 18804
rect 10696 18624 10706 18804
rect 10740 18792 10786 18804
rect 10452 18404 10498 18416
rect 10530 18404 10540 18584
rect 10600 18404 10610 18584
rect 10644 18416 10650 18624
rect 10684 18416 10690 18624
rect 10740 18584 10746 18792
rect 10780 18584 10786 18792
rect 10818 18624 10828 18804
rect 10888 18624 10898 18804
rect 10932 18792 10978 18804
rect 10644 18404 10690 18416
rect 10722 18404 10732 18584
rect 10792 18404 10802 18584
rect 10836 18416 10842 18624
rect 10876 18416 10882 18624
rect 10932 18584 10938 18792
rect 10972 18584 10978 18792
rect 11010 18624 11020 18804
rect 11080 18624 11090 18804
rect 11124 18792 11170 18804
rect 10836 18404 10882 18416
rect 10914 18404 10924 18584
rect 10984 18404 10994 18584
rect 11028 18416 11034 18624
rect 11068 18416 11074 18624
rect 11124 18584 11130 18792
rect 11164 18584 11170 18792
rect 11028 18404 11074 18416
rect 11106 18404 11116 18584
rect 11176 18404 11186 18584
rect 6648 18366 6852 18372
rect 6648 18332 6672 18366
rect 6840 18356 6852 18366
rect 6918 18366 7368 18372
rect 6918 18356 6930 18366
rect 6840 18332 6930 18356
rect 7098 18332 7188 18366
rect 7356 18356 7368 18366
rect 7434 18366 7884 18372
rect 7434 18356 7446 18366
rect 7356 18332 7446 18356
rect 7614 18332 7704 18366
rect 7872 18356 7884 18366
rect 8368 18366 8572 18372
rect 7872 18332 7892 18356
rect 6648 18258 7892 18332
rect 6648 18224 6672 18258
rect 6840 18224 6930 18258
rect 7098 18224 7188 18258
rect 7356 18224 7446 18258
rect 7614 18224 7704 18258
rect 7872 18224 7892 18258
rect 6648 18220 7892 18224
rect 8368 18332 8392 18366
rect 8560 18356 8572 18366
rect 8638 18366 9088 18372
rect 8638 18356 8650 18366
rect 8560 18332 8650 18356
rect 8818 18332 8908 18366
rect 9076 18356 9088 18366
rect 9154 18366 9604 18372
rect 9154 18356 9166 18366
rect 9076 18332 9166 18356
rect 9334 18332 9424 18366
rect 9592 18356 9604 18366
rect 10024 18366 11140 18372
rect 9592 18332 9612 18356
rect 8368 18258 9612 18332
rect 8368 18224 8392 18258
rect 8560 18224 8650 18258
rect 8818 18224 8908 18258
rect 9076 18224 9166 18258
rect 9334 18224 9424 18258
rect 9592 18224 9612 18258
rect 8368 18220 9612 18224
rect 10024 18332 10314 18366
rect 10348 18332 10506 18366
rect 10540 18332 10698 18366
rect 10732 18332 10890 18366
rect 10924 18332 11082 18366
rect 11116 18332 11140 18366
rect 10024 18258 11140 18332
rect 10024 18224 10314 18258
rect 10348 18224 10506 18258
rect 10540 18224 10698 18258
rect 10732 18224 10890 18258
rect 10924 18224 11082 18258
rect 11116 18224 11140 18258
rect 6660 18218 6852 18220
rect 6918 18218 7110 18220
rect 7176 18218 7368 18220
rect 7434 18218 7626 18220
rect 7692 18218 7884 18220
rect 8380 18218 8572 18220
rect 8638 18218 8830 18220
rect 8896 18218 9088 18220
rect 9154 18218 9346 18220
rect 9412 18218 9604 18220
rect 6590 18008 6600 18188
rect 6652 18008 6662 18188
rect 6862 18174 6908 18186
rect 6604 17798 6610 18008
rect 6644 17798 6650 18008
rect 6862 17968 6868 18174
rect 6902 17968 6908 18174
rect 6604 17786 6650 17798
rect 6850 17788 6860 17968
rect 6912 17788 6922 17968
rect 6862 17786 6908 17788
rect 6952 17756 7072 18218
rect 7106 18008 7116 18188
rect 7168 18008 7178 18188
rect 7120 17798 7126 18008
rect 7160 17798 7166 18008
rect 7120 17786 7166 17798
rect 7212 17756 7332 18218
rect 7378 18174 7424 18186
rect 7378 17968 7384 18174
rect 7418 17968 7424 18174
rect 7366 17788 7376 17968
rect 7428 17788 7438 17968
rect 7378 17786 7424 17788
rect 7472 17756 7592 18218
rect 7622 18008 7632 18188
rect 7684 18008 7694 18188
rect 7894 18174 7940 18186
rect 7636 17798 7642 18008
rect 7676 17798 7682 18008
rect 7894 17968 7900 18174
rect 7934 17968 7940 18174
rect 8310 18008 8320 18188
rect 8372 18008 8382 18188
rect 8582 18174 8628 18186
rect 7636 17786 7682 17798
rect 7882 17788 7892 17968
rect 7944 17788 7954 17968
rect 8324 17798 8330 18008
rect 8364 17798 8370 18008
rect 8582 17968 8588 18174
rect 8622 17968 8628 18174
rect 7894 17786 7940 17788
rect 8324 17786 8370 17798
rect 8570 17788 8580 17968
rect 8632 17788 8642 17968
rect 8582 17786 8628 17788
rect 8028 17776 8232 17782
rect 6648 17748 7888 17756
rect 6648 17714 6672 17748
rect 6840 17714 6930 17748
rect 7098 17714 7188 17748
rect 7356 17714 7446 17748
rect 7614 17714 7704 17748
rect 7872 17714 7888 17748
rect 6648 17696 7888 17714
rect 8028 17616 8040 17776
rect 8220 17616 8232 17776
rect 8672 17756 8792 18218
rect 8826 18008 8836 18188
rect 8888 18008 8898 18188
rect 8840 17798 8846 18008
rect 8880 17798 8886 18008
rect 8840 17786 8886 17798
rect 8932 17756 9052 18218
rect 9098 18174 9144 18186
rect 9098 17968 9104 18174
rect 9138 17968 9144 18174
rect 9086 17788 9096 17968
rect 9148 17788 9158 17968
rect 9098 17786 9144 17788
rect 9192 17756 9312 18218
rect 10024 18216 11140 18224
rect 9342 18008 9352 18188
rect 9404 18008 9414 18188
rect 9614 18174 9660 18186
rect 9356 17798 9362 18008
rect 9396 17798 9402 18008
rect 9614 17968 9620 18174
rect 9654 17968 9660 18174
rect 9356 17786 9402 17798
rect 9602 17788 9612 17968
rect 9664 17788 9674 17968
rect 9614 17786 9660 17788
rect 10024 17756 10120 18216
rect 10164 18174 10210 18186
rect 10164 17964 10170 18174
rect 10204 17964 10210 18174
rect 10242 18008 10252 18188
rect 10312 18008 10322 18188
rect 10356 18174 10402 18186
rect 10150 17784 10160 17964
rect 10220 17784 10230 17964
rect 10260 17798 10266 18008
rect 10300 17798 10306 18008
rect 10356 17964 10362 18174
rect 10396 17964 10402 18174
rect 10434 18008 10444 18188
rect 10504 18008 10514 18188
rect 10548 18174 10594 18186
rect 10260 17786 10306 17798
rect 10338 17784 10348 17964
rect 10408 17784 10418 17964
rect 10452 17798 10458 18008
rect 10492 17798 10498 18008
rect 10548 17964 10554 18174
rect 10588 17964 10594 18174
rect 10626 18008 10636 18188
rect 10696 18008 10706 18188
rect 10740 18174 10786 18186
rect 10452 17786 10498 17798
rect 10530 17784 10540 17964
rect 10600 17784 10610 17964
rect 10644 17798 10650 18008
rect 10684 17798 10690 18008
rect 10740 17964 10746 18174
rect 10780 17964 10786 18174
rect 10818 18008 10828 18188
rect 10888 18008 10898 18188
rect 10932 18174 10978 18186
rect 10644 17786 10690 17798
rect 10722 17784 10732 17964
rect 10792 17784 10802 17964
rect 10836 17798 10842 18008
rect 10876 17798 10882 18008
rect 10932 17964 10938 18174
rect 10972 17964 10978 18174
rect 11010 18008 11020 18188
rect 11080 18008 11090 18188
rect 11124 18174 11170 18186
rect 10836 17786 10882 17798
rect 10914 17784 10924 17964
rect 10984 17784 10994 17964
rect 11028 17798 11034 18008
rect 11068 17798 11074 18008
rect 11124 17964 11130 18174
rect 11164 17964 11170 18174
rect 11028 17786 11074 17798
rect 11106 17784 11116 17964
rect 11176 17784 11186 17964
rect 8368 17748 9608 17756
rect 8368 17714 8392 17748
rect 8560 17714 8650 17748
rect 8818 17714 8908 17748
rect 9076 17714 9166 17748
rect 9334 17714 9424 17748
rect 9592 17714 9608 17748
rect 8368 17696 9608 17714
rect 10024 17748 11044 17756
rect 10024 17714 10218 17748
rect 10252 17714 10410 17748
rect 10444 17714 10602 17748
rect 10636 17714 10794 17748
rect 10828 17714 10986 17748
rect 11020 17714 11044 17748
rect 10024 17712 11044 17714
rect 8028 17610 8232 17616
rect 9400 17280 9600 17696
rect 10024 17652 11300 17712
rect 9400 16980 10160 17280
rect 1288 10768 1580 10774
rect 1288 10532 1300 10768
rect 1568 10532 1580 10768
rect 2578 10660 2588 11148
rect 4792 10660 4802 11148
rect 6090 10808 6282 10820
rect 6086 10608 6096 10808
rect 6276 10608 6286 10808
rect 6090 10596 6282 10608
rect 1288 10526 1580 10532
rect 6724 10428 7576 10436
rect 5156 10388 7576 10428
rect 5156 10364 9548 10388
rect 5156 10330 5174 10364
rect 5208 10330 5366 10364
rect 5400 10330 5558 10364
rect 5592 10330 5750 10364
rect 5784 10330 5942 10364
rect 5976 10330 6134 10364
rect 6168 10330 6326 10364
rect 6360 10330 6518 10364
rect 6552 10330 6710 10364
rect 6744 10330 6902 10364
rect 6936 10334 9548 10364
rect 6936 10330 7770 10334
rect 5156 10324 7770 10330
rect 7156 10300 7770 10324
rect 7804 10300 7962 10334
rect 7996 10300 8154 10334
rect 8188 10300 8346 10334
rect 8380 10300 8538 10334
rect 8572 10300 8730 10334
rect 8764 10300 8922 10334
rect 8956 10300 9114 10334
rect 9148 10300 9306 10334
rect 9340 10300 9498 10334
rect 9532 10300 9548 10334
rect 7156 10292 9548 10300
rect 5120 10271 5166 10283
rect 5120 10060 5126 10271
rect 5160 10060 5166 10271
rect 5202 10104 5212 10284
rect 5268 10104 5278 10284
rect 5312 10271 5358 10283
rect 2578 9440 2588 9908
rect 4780 9440 4790 9908
rect 5106 9880 5116 10060
rect 5172 9880 5182 10060
rect 5216 9895 5222 10104
rect 5256 9895 5262 10104
rect 5312 10060 5318 10271
rect 5352 10060 5358 10271
rect 5394 10104 5404 10284
rect 5460 10104 5470 10284
rect 5504 10271 5550 10283
rect 5216 9883 5262 9895
rect 5298 9880 5308 10060
rect 5364 9880 5374 10060
rect 5408 9895 5414 10104
rect 5448 9895 5454 10104
rect 5504 10060 5510 10271
rect 5544 10060 5550 10271
rect 5586 10104 5596 10284
rect 5652 10104 5662 10284
rect 5696 10271 5742 10283
rect 5408 9883 5454 9895
rect 5490 9880 5500 10060
rect 5556 9880 5566 10060
rect 5600 9895 5606 10104
rect 5640 9895 5646 10104
rect 5696 10060 5702 10271
rect 5736 10060 5742 10271
rect 5778 10104 5788 10284
rect 5844 10104 5854 10284
rect 5888 10271 5934 10283
rect 5600 9883 5646 9895
rect 5682 9880 5692 10060
rect 5748 9880 5758 10060
rect 5792 9895 5798 10104
rect 5832 9895 5838 10104
rect 5888 10060 5894 10271
rect 5928 10060 5934 10271
rect 5970 10104 5980 10284
rect 6036 10104 6046 10284
rect 6080 10271 6126 10283
rect 5792 9883 5838 9895
rect 5874 9880 5884 10060
rect 5940 9880 5950 10060
rect 5984 9895 5990 10104
rect 6024 9895 6030 10104
rect 6080 10060 6086 10271
rect 6120 10060 6126 10271
rect 6162 10104 6172 10284
rect 6228 10104 6238 10284
rect 6272 10271 6318 10283
rect 5984 9883 6030 9895
rect 6066 9880 6076 10060
rect 6132 9880 6142 10060
rect 6176 9895 6182 10104
rect 6216 9895 6222 10104
rect 6272 10060 6278 10271
rect 6312 10060 6318 10271
rect 6354 10104 6364 10284
rect 6420 10104 6430 10284
rect 6464 10271 6510 10283
rect 6176 9883 6222 9895
rect 6258 9880 6268 10060
rect 6324 9880 6334 10060
rect 6368 9895 6374 10104
rect 6408 9895 6414 10104
rect 6464 10060 6470 10271
rect 6504 10060 6510 10271
rect 6546 10104 6556 10284
rect 6612 10104 6622 10284
rect 6656 10271 6702 10283
rect 6368 9883 6414 9895
rect 6450 9880 6460 10060
rect 6516 9880 6526 10060
rect 6560 9895 6566 10104
rect 6600 9895 6606 10104
rect 6656 10060 6662 10271
rect 6696 10060 6702 10271
rect 6738 10104 6748 10284
rect 6804 10104 6814 10284
rect 6848 10271 6894 10283
rect 6560 9883 6606 9895
rect 6642 9880 6652 10060
rect 6708 9880 6718 10060
rect 6752 9895 6758 10104
rect 6792 9895 6798 10104
rect 6848 10060 6854 10271
rect 6888 10060 6894 10271
rect 6930 10104 6940 10284
rect 6996 10104 7006 10284
rect 7040 10271 7086 10283
rect 6752 9883 6798 9895
rect 6834 9880 6844 10060
rect 6900 9880 6910 10060
rect 6944 9895 6950 10104
rect 6984 9895 6990 10104
rect 7040 10060 7046 10271
rect 7080 10060 7086 10271
rect 6944 9883 6990 9895
rect 7026 9880 7036 10060
rect 7092 9880 7102 10060
rect 7156 9844 7576 10292
rect 7620 10250 7666 10262
rect 7620 10044 7626 10250
rect 7660 10044 7666 10250
rect 7702 10080 7712 10264
rect 7768 10080 7778 10264
rect 7812 10250 7858 10262
rect 7606 9860 7616 10044
rect 7672 9860 7682 10044
rect 7716 9874 7722 10080
rect 7756 9874 7762 10080
rect 7812 10044 7818 10250
rect 7852 10044 7858 10250
rect 7894 10080 7904 10264
rect 7960 10080 7970 10264
rect 8004 10250 8050 10262
rect 7716 9862 7762 9874
rect 7798 9860 7808 10044
rect 7864 9860 7874 10044
rect 7908 9874 7914 10080
rect 7948 9874 7954 10080
rect 8004 10044 8010 10250
rect 8044 10044 8050 10250
rect 8086 10080 8096 10264
rect 8152 10080 8162 10264
rect 8196 10250 8242 10262
rect 7908 9862 7954 9874
rect 7990 9860 8000 10044
rect 8056 9860 8066 10044
rect 8100 9874 8106 10080
rect 8140 9874 8146 10080
rect 8196 10044 8202 10250
rect 8236 10044 8242 10250
rect 8278 10080 8288 10264
rect 8344 10080 8354 10264
rect 8388 10250 8434 10262
rect 8100 9862 8146 9874
rect 8182 9860 8192 10044
rect 8248 9860 8258 10044
rect 8292 9874 8298 10080
rect 8332 9874 8338 10080
rect 8388 10044 8394 10250
rect 8428 10044 8434 10250
rect 8470 10080 8480 10264
rect 8536 10080 8546 10264
rect 8580 10250 8626 10262
rect 8292 9862 8338 9874
rect 8374 9860 8384 10044
rect 8440 9860 8450 10044
rect 8484 9874 8490 10080
rect 8524 9874 8530 10080
rect 8580 10044 8586 10250
rect 8620 10044 8626 10250
rect 8662 10080 8672 10264
rect 8728 10080 8738 10264
rect 8772 10250 8818 10262
rect 8484 9862 8530 9874
rect 8566 9860 8576 10044
rect 8632 9860 8642 10044
rect 8676 9874 8682 10080
rect 8716 9874 8722 10080
rect 8772 10044 8778 10250
rect 8812 10044 8818 10250
rect 8854 10080 8864 10264
rect 8920 10080 8930 10264
rect 8964 10250 9010 10262
rect 8676 9862 8722 9874
rect 8758 9860 8768 10044
rect 8824 9860 8834 10044
rect 8868 9874 8874 10080
rect 8908 9874 8914 10080
rect 8964 10044 8970 10250
rect 9004 10044 9010 10250
rect 9046 10080 9056 10264
rect 9112 10080 9122 10264
rect 9156 10250 9202 10262
rect 8868 9862 8914 9874
rect 8950 9860 8960 10044
rect 9016 9860 9026 10044
rect 9060 9874 9066 10080
rect 9100 9874 9106 10080
rect 9156 10044 9162 10250
rect 9196 10044 9202 10250
rect 9238 10080 9248 10264
rect 9304 10080 9314 10264
rect 9348 10250 9394 10262
rect 9060 9862 9106 9874
rect 9142 9860 9152 10044
rect 9208 9860 9218 10044
rect 9252 9874 9258 10080
rect 9292 9874 9298 10080
rect 9348 10044 9354 10250
rect 9388 10044 9394 10250
rect 9430 10080 9440 10264
rect 9496 10080 9506 10264
rect 9540 10250 9586 10262
rect 9252 9862 9298 9874
rect 9334 9860 9344 10044
rect 9400 9860 9410 10044
rect 9444 9874 9450 10080
rect 9484 9874 9490 10080
rect 9540 10044 9546 10250
rect 9580 10044 9586 10250
rect 9444 9862 9490 9874
rect 9526 9860 9536 10044
rect 9592 9860 9602 10044
rect 5252 9836 7576 9844
rect 5252 9802 5270 9836
rect 5304 9802 5462 9836
rect 5496 9802 5654 9836
rect 5688 9802 5846 9836
rect 5880 9802 6038 9836
rect 6072 9802 6230 9836
rect 6264 9802 6422 9836
rect 6456 9802 6614 9836
rect 6648 9802 6806 9836
rect 6840 9802 6998 9836
rect 7032 9832 7576 9836
rect 7032 9824 9452 9832
rect 7032 9802 7674 9824
rect 5252 9790 7674 9802
rect 7708 9790 7866 9824
rect 7900 9790 8058 9824
rect 8092 9790 8250 9824
rect 8284 9790 8442 9824
rect 8476 9790 8634 9824
rect 8668 9790 8826 9824
rect 8860 9790 9018 9824
rect 9052 9790 9210 9824
rect 9244 9790 9402 9824
rect 9436 9790 9452 9824
rect 5252 9728 9452 9790
rect 5252 9694 5270 9728
rect 5304 9694 5462 9728
rect 5496 9694 5654 9728
rect 5688 9694 5846 9728
rect 5880 9694 6038 9728
rect 6072 9694 6230 9728
rect 6264 9694 6422 9728
rect 6456 9694 6614 9728
rect 6648 9694 6806 9728
rect 6840 9694 6998 9728
rect 7032 9716 9452 9728
rect 7032 9694 7674 9716
rect 5252 9688 7674 9694
rect 7156 9682 7674 9688
rect 7708 9682 7866 9716
rect 7900 9682 8058 9716
rect 8092 9682 8250 9716
rect 8284 9682 8442 9716
rect 8476 9682 8634 9716
rect 8668 9682 8826 9716
rect 8860 9682 9018 9716
rect 9052 9682 9210 9716
rect 9244 9682 9402 9716
rect 9436 9682 9452 9716
rect 7156 9676 9452 9682
rect 5120 9635 5166 9647
rect 5120 9428 5126 9635
rect 5160 9428 5166 9635
rect 5202 9472 5212 9652
rect 5268 9472 5278 9652
rect 5312 9635 5358 9647
rect 5106 9248 5116 9428
rect 5172 9248 5182 9428
rect 5216 9259 5222 9472
rect 5256 9259 5262 9472
rect 5312 9428 5318 9635
rect 5352 9428 5358 9635
rect 5394 9472 5404 9652
rect 5460 9472 5470 9652
rect 5504 9635 5550 9647
rect 5120 9247 5166 9248
rect 5216 9247 5262 9259
rect 5298 9248 5308 9428
rect 5364 9248 5374 9428
rect 5408 9259 5414 9472
rect 5448 9259 5454 9472
rect 5504 9428 5510 9635
rect 5544 9428 5550 9635
rect 5586 9472 5596 9652
rect 5652 9472 5662 9652
rect 5696 9635 5742 9647
rect 5312 9247 5358 9248
rect 5408 9247 5454 9259
rect 5490 9248 5500 9428
rect 5556 9248 5566 9428
rect 5600 9259 5606 9472
rect 5640 9259 5646 9472
rect 5696 9428 5702 9635
rect 5736 9428 5742 9635
rect 5778 9472 5788 9652
rect 5844 9472 5854 9652
rect 5888 9635 5934 9647
rect 5504 9247 5550 9248
rect 5600 9247 5646 9259
rect 5682 9248 5692 9428
rect 5748 9248 5758 9428
rect 5792 9259 5798 9472
rect 5832 9259 5838 9472
rect 5888 9428 5894 9635
rect 5928 9428 5934 9635
rect 5970 9472 5980 9652
rect 6036 9472 6046 9652
rect 6080 9635 6126 9647
rect 5696 9247 5742 9248
rect 5792 9247 5838 9259
rect 5874 9248 5884 9428
rect 5940 9248 5950 9428
rect 5984 9259 5990 9472
rect 6024 9259 6030 9472
rect 6080 9428 6086 9635
rect 6120 9428 6126 9635
rect 6162 9472 6172 9652
rect 6228 9472 6238 9652
rect 6272 9635 6318 9647
rect 5888 9247 5934 9248
rect 5984 9247 6030 9259
rect 6066 9248 6076 9428
rect 6132 9248 6142 9428
rect 6176 9259 6182 9472
rect 6216 9259 6222 9472
rect 6272 9428 6278 9635
rect 6312 9428 6318 9635
rect 6354 9472 6364 9652
rect 6420 9472 6430 9652
rect 6464 9635 6510 9647
rect 6080 9247 6126 9248
rect 6176 9247 6222 9259
rect 6258 9248 6268 9428
rect 6324 9248 6334 9428
rect 6368 9259 6374 9472
rect 6408 9259 6414 9472
rect 6464 9428 6470 9635
rect 6504 9428 6510 9635
rect 6546 9472 6556 9652
rect 6612 9472 6622 9652
rect 6656 9635 6702 9647
rect 6272 9247 6318 9248
rect 6368 9247 6414 9259
rect 6450 9248 6460 9428
rect 6516 9248 6526 9428
rect 6560 9259 6566 9472
rect 6600 9259 6606 9472
rect 6656 9428 6662 9635
rect 6696 9428 6702 9635
rect 6738 9472 6748 9652
rect 6804 9472 6814 9652
rect 6848 9635 6894 9647
rect 6464 9247 6510 9248
rect 6560 9247 6606 9259
rect 6642 9248 6652 9428
rect 6708 9248 6718 9428
rect 6752 9259 6758 9472
rect 6792 9259 6798 9472
rect 6848 9428 6854 9635
rect 6888 9428 6894 9635
rect 6930 9472 6940 9652
rect 6996 9472 7006 9652
rect 7040 9635 7086 9647
rect 6656 9247 6702 9248
rect 6752 9247 6798 9259
rect 6834 9248 6844 9428
rect 6900 9248 6910 9428
rect 6944 9259 6950 9472
rect 6984 9259 6990 9472
rect 7040 9428 7046 9635
rect 7080 9428 7086 9635
rect 6848 9247 6894 9248
rect 6944 9247 6990 9259
rect 7026 9248 7036 9428
rect 7092 9248 7102 9428
rect 7040 9247 7086 9248
rect 7156 9212 7576 9676
rect 7620 9632 7666 9644
rect 7620 9428 7626 9632
rect 7660 9428 7666 9632
rect 7702 9464 7712 9648
rect 7768 9464 7778 9648
rect 7812 9632 7858 9644
rect 7606 9244 7616 9428
rect 7672 9244 7682 9428
rect 7716 9256 7722 9464
rect 7756 9256 7762 9464
rect 7812 9428 7818 9632
rect 7852 9428 7858 9632
rect 7894 9464 7904 9648
rect 7960 9464 7970 9648
rect 8004 9632 8050 9644
rect 7716 9244 7762 9256
rect 7798 9244 7808 9428
rect 7864 9244 7874 9428
rect 7908 9256 7914 9464
rect 7948 9256 7954 9464
rect 8004 9428 8010 9632
rect 8044 9428 8050 9632
rect 8086 9464 8096 9648
rect 8152 9464 8162 9648
rect 8196 9632 8242 9644
rect 7908 9244 7954 9256
rect 7990 9244 8000 9428
rect 8056 9244 8066 9428
rect 8100 9256 8106 9464
rect 8140 9256 8146 9464
rect 8196 9428 8202 9632
rect 8236 9428 8242 9632
rect 8278 9464 8288 9648
rect 8344 9464 8354 9648
rect 8388 9632 8434 9644
rect 8100 9244 8146 9256
rect 8182 9244 8192 9428
rect 8248 9244 8258 9428
rect 8292 9256 8298 9464
rect 8332 9256 8338 9464
rect 8388 9428 8394 9632
rect 8428 9428 8434 9632
rect 8470 9464 8480 9648
rect 8536 9464 8546 9648
rect 8580 9632 8626 9644
rect 8292 9244 8338 9256
rect 8374 9244 8384 9428
rect 8440 9244 8450 9428
rect 8484 9256 8490 9464
rect 8524 9256 8530 9464
rect 8580 9428 8586 9632
rect 8620 9428 8626 9632
rect 8662 9464 8672 9648
rect 8728 9464 8738 9648
rect 8772 9632 8818 9644
rect 8484 9244 8530 9256
rect 8566 9244 8576 9428
rect 8632 9244 8642 9428
rect 8676 9256 8682 9464
rect 8716 9256 8722 9464
rect 8772 9428 8778 9632
rect 8812 9428 8818 9632
rect 8854 9464 8864 9648
rect 8920 9464 8930 9648
rect 8964 9632 9010 9644
rect 8676 9244 8722 9256
rect 8758 9244 8768 9428
rect 8824 9244 8834 9428
rect 8868 9256 8874 9464
rect 8908 9256 8914 9464
rect 8964 9428 8970 9632
rect 9004 9428 9010 9632
rect 9046 9464 9056 9648
rect 9112 9464 9122 9648
rect 9156 9632 9202 9644
rect 8868 9244 8914 9256
rect 8950 9244 8960 9428
rect 9016 9244 9026 9428
rect 9060 9256 9066 9464
rect 9100 9256 9106 9464
rect 9156 9428 9162 9632
rect 9196 9428 9202 9632
rect 9238 9464 9248 9648
rect 9304 9464 9314 9648
rect 9348 9632 9394 9644
rect 9060 9244 9106 9256
rect 9142 9244 9152 9428
rect 9208 9244 9218 9428
rect 9252 9256 9258 9464
rect 9292 9256 9298 9464
rect 9348 9428 9354 9632
rect 9388 9428 9394 9632
rect 9430 9464 9440 9648
rect 9496 9464 9506 9648
rect 9540 9632 9586 9644
rect 9252 9244 9298 9256
rect 9334 9244 9344 9428
rect 9400 9244 9410 9428
rect 9444 9256 9450 9464
rect 9484 9256 9490 9464
rect 9540 9428 9546 9632
rect 9580 9428 9586 9632
rect 9444 9244 9490 9256
rect 9526 9244 9536 9428
rect 9592 9244 9602 9428
rect 7156 9208 9548 9212
rect 5156 9206 9548 9208
rect 5156 9200 7770 9206
rect 5156 9166 5174 9200
rect 5208 9166 5366 9200
rect 5400 9166 5558 9200
rect 5592 9166 5750 9200
rect 5784 9166 5942 9200
rect 5976 9166 6134 9200
rect 6168 9166 6326 9200
rect 6360 9166 6518 9200
rect 6552 9166 6710 9200
rect 6744 9166 6902 9200
rect 6936 9172 7770 9200
rect 7804 9172 7962 9206
rect 7996 9172 8154 9206
rect 8188 9172 8346 9206
rect 8380 9172 8538 9206
rect 8572 9172 8730 9206
rect 8764 9172 8922 9206
rect 8956 9172 9114 9206
rect 9148 9172 9306 9206
rect 9340 9172 9498 9206
rect 9532 9172 9548 9206
rect 6936 9166 9548 9172
rect 5156 9104 9548 9166
rect 7156 9098 9548 9104
rect 7156 9064 7770 9098
rect 7804 9064 7962 9098
rect 7996 9064 8154 9098
rect 8188 9064 8346 9098
rect 8380 9064 8538 9098
rect 8572 9064 8730 9098
rect 8764 9064 8922 9098
rect 8956 9064 9114 9098
rect 9148 9064 9306 9098
rect 9340 9064 9498 9098
rect 9532 9064 9548 9098
rect 7156 9056 9548 9064
rect 1532 8970 1736 8972
rect 1532 8968 1976 8970
rect 1520 8964 1976 8968
rect 2528 8964 2844 8970
rect 1520 8904 1672 8964
rect 2056 8904 2066 8964
rect 2528 8904 2540 8964
rect 2832 8904 2844 8964
rect 1520 8898 1976 8904
rect 2528 8898 2844 8904
rect 3464 8964 3780 8970
rect 3464 8904 3476 8964
rect 3768 8904 3780 8964
rect 3464 8898 3780 8904
rect 1520 8896 1736 8898
rect 1520 8704 1604 8896
rect 4578 8868 4588 8984
rect 1816 8802 4588 8868
rect 1816 8768 1834 8802
rect 1868 8768 2026 8802
rect 2060 8768 2218 8802
rect 2252 8768 2410 8802
rect 2444 8768 2602 8802
rect 2636 8768 2794 8802
rect 2828 8768 2986 8802
rect 3020 8768 3178 8802
rect 3212 8768 3370 8802
rect 3404 8768 3562 8802
rect 3596 8768 4588 8802
rect 1816 8760 4588 8768
rect -9928 8356 -8884 8364
rect -9928 8306 -9044 8356
rect -9928 8272 -9906 8306
rect -9872 8272 -9714 8306
rect -9680 8272 -9522 8306
rect -9488 8272 -9330 8306
rect -9296 8272 -9138 8306
rect -9104 8280 -9044 8306
rect -8904 8280 -8884 8356
rect 1520 8356 1540 8704
rect 1596 8356 1604 8704
rect 1684 8718 1730 8730
rect 1684 8508 1690 8718
rect 1724 8508 1730 8718
rect 1766 8552 1776 8732
rect 1828 8552 1838 8732
rect 1876 8718 1922 8730
rect -9104 8272 -8884 8280
rect -9928 8264 -8884 8272
rect -10056 8222 -10010 8234
rect -10056 8012 -10050 8222
rect -10016 8012 -10010 8222
rect -9974 8056 -9964 8236
rect -9912 8056 -9902 8236
rect -9864 8222 -9818 8234
rect -10070 7832 -10060 8012
rect -10008 7832 -9998 8012
rect -9960 7846 -9954 8056
rect -9920 7846 -9914 8056
rect -9864 8012 -9858 8222
rect -9824 8012 -9818 8222
rect -9782 8056 -9772 8236
rect -9720 8056 -9710 8236
rect -9672 8222 -9626 8234
rect -9960 7834 -9914 7846
rect -9878 7832 -9868 8012
rect -9816 7832 -9806 8012
rect -9768 7846 -9762 8056
rect -9728 7846 -9722 8056
rect -9672 8012 -9666 8222
rect -9632 8012 -9626 8222
rect -9590 8056 -9580 8236
rect -9528 8056 -9518 8236
rect -9480 8222 -9434 8234
rect -9768 7834 -9722 7846
rect -9686 7832 -9676 8012
rect -9624 7832 -9614 8012
rect -9576 7846 -9570 8056
rect -9536 7846 -9530 8056
rect -9480 8012 -9474 8222
rect -9440 8012 -9434 8222
rect -9398 8056 -9388 8236
rect -9336 8056 -9326 8236
rect -9288 8222 -9242 8234
rect -9576 7834 -9530 7846
rect -9494 7832 -9484 8012
rect -9432 7832 -9422 8012
rect -9384 7846 -9378 8056
rect -9344 7846 -9338 8056
rect -9288 8012 -9282 8222
rect -9248 8012 -9242 8222
rect -9206 8056 -9196 8236
rect -9144 8056 -9134 8236
rect -9096 8222 -9050 8234
rect -9384 7834 -9338 7846
rect -9302 7832 -9292 8012
rect -9240 7832 -9230 8012
rect -9192 7846 -9186 8056
rect -9152 7846 -9146 8056
rect -9096 8012 -9090 8222
rect -9056 8012 -9050 8222
rect -9192 7834 -9146 7846
rect -9110 7832 -9100 8012
rect -9048 7832 -9038 8012
rect -9004 7804 -8884 8264
rect -8670 8196 -8660 8296
rect -8480 8196 -8470 8296
rect -8670 8190 -8470 8196
rect -10020 7796 -8884 7804
rect -10020 7762 -10002 7796
rect -9968 7762 -9810 7796
rect -9776 7762 -9618 7796
rect -9584 7762 -9426 7796
rect -9392 7762 -9234 7796
rect -9200 7762 -8884 7796
rect -10020 7688 -8884 7762
rect -10020 7654 -10002 7688
rect -9968 7654 -9810 7688
rect -9776 7654 -9618 7688
rect -9584 7654 -9426 7688
rect -9392 7654 -9234 7688
rect -9200 7654 -8884 7688
rect -10020 7648 -8884 7654
rect -10056 7604 -10010 7616
rect -10056 7396 -10050 7604
rect -10016 7396 -10010 7604
rect -9974 7440 -9964 7620
rect -9912 7440 -9902 7620
rect -9864 7604 -9818 7616
rect -10070 7216 -10060 7396
rect -10008 7216 -9998 7396
rect -9960 7228 -9954 7440
rect -9920 7228 -9914 7440
rect -9864 7396 -9858 7604
rect -9824 7396 -9818 7604
rect -9782 7440 -9772 7620
rect -9720 7440 -9710 7620
rect -9672 7604 -9626 7616
rect -9960 7216 -9914 7228
rect -9878 7216 -9868 7396
rect -9816 7216 -9806 7396
rect -9768 7228 -9762 7440
rect -9728 7228 -9722 7440
rect -9672 7396 -9666 7604
rect -9632 7396 -9626 7604
rect -9590 7440 -9580 7620
rect -9528 7440 -9518 7620
rect -9480 7604 -9434 7616
rect -9768 7216 -9722 7228
rect -9686 7216 -9676 7396
rect -9624 7216 -9614 7396
rect -9576 7228 -9570 7440
rect -9536 7228 -9530 7440
rect -9480 7396 -9474 7604
rect -9440 7396 -9434 7604
rect -9398 7440 -9388 7620
rect -9336 7440 -9326 7620
rect -9288 7604 -9242 7616
rect -9576 7216 -9530 7228
rect -9494 7216 -9484 7396
rect -9432 7216 -9422 7396
rect -9384 7228 -9378 7440
rect -9344 7228 -9338 7440
rect -9288 7396 -9282 7604
rect -9248 7396 -9242 7604
rect -9206 7440 -9196 7620
rect -9144 7440 -9134 7620
rect -9096 7604 -9050 7616
rect -9384 7216 -9338 7228
rect -9302 7216 -9292 7396
rect -9240 7216 -9230 7396
rect -9192 7228 -9186 7440
rect -9152 7228 -9146 7440
rect -9096 7396 -9090 7604
rect -9056 7396 -9050 7604
rect -9192 7216 -9146 7228
rect -9110 7216 -9100 7396
rect -9048 7216 -9038 7396
rect -9004 7184 -8884 7648
rect -9924 7178 -8884 7184
rect -9924 7144 -9906 7178
rect -9872 7144 -9714 7178
rect -9680 7144 -9522 7178
rect -9488 7144 -9330 7178
rect -9296 7144 -9138 7178
rect -9104 7144 -8884 7178
rect -9924 7070 -8884 7144
rect -9924 7036 -9906 7070
rect -9872 7036 -9714 7070
rect -9680 7036 -9522 7070
rect -9488 7036 -9330 7070
rect -9296 7036 -9138 7070
rect -9104 7036 -8884 7070
rect -8748 8168 -8702 8180
rect -8748 7040 -8742 8168
rect -8708 7040 -8702 8168
rect -8438 8168 -8392 8180
rect -8438 7044 -8432 8168
rect -8398 7044 -8392 8168
rect 1520 8160 1604 8356
rect 1670 8328 1680 8508
rect 1732 8328 1742 8508
rect 1780 8342 1786 8552
rect 1820 8342 1826 8552
rect 1876 8508 1882 8718
rect 1916 8508 1922 8718
rect 1958 8552 1968 8732
rect 2020 8552 2030 8732
rect 2068 8718 2114 8730
rect 1780 8330 1826 8342
rect 1862 8328 1872 8508
rect 1924 8328 1934 8508
rect 1972 8342 1978 8552
rect 2012 8342 2018 8552
rect 2068 8508 2074 8718
rect 2108 8508 2114 8718
rect 2150 8552 2160 8732
rect 2212 8552 2222 8732
rect 2260 8718 2306 8730
rect 1972 8330 2018 8342
rect 2054 8328 2064 8508
rect 2116 8328 2126 8508
rect 2164 8342 2170 8552
rect 2204 8342 2210 8552
rect 2260 8508 2266 8718
rect 2300 8508 2306 8718
rect 2342 8552 2352 8732
rect 2404 8552 2414 8732
rect 2452 8718 2498 8730
rect 2164 8330 2210 8342
rect 2246 8328 2256 8508
rect 2308 8328 2318 8508
rect 2356 8342 2362 8552
rect 2396 8342 2402 8552
rect 2452 8508 2458 8718
rect 2492 8508 2498 8718
rect 2534 8552 2544 8732
rect 2596 8552 2606 8732
rect 2644 8718 2690 8730
rect 2356 8330 2402 8342
rect 2438 8328 2448 8508
rect 2500 8328 2510 8508
rect 2548 8342 2554 8552
rect 2588 8342 2594 8552
rect 2644 8508 2650 8718
rect 2684 8508 2690 8718
rect 2726 8552 2736 8732
rect 2788 8552 2798 8732
rect 2836 8718 2882 8730
rect 2548 8330 2594 8342
rect 2630 8328 2640 8508
rect 2692 8328 2702 8508
rect 2740 8342 2746 8552
rect 2780 8342 2786 8552
rect 2836 8508 2842 8718
rect 2876 8508 2882 8718
rect 2918 8552 2928 8732
rect 2980 8552 2990 8732
rect 3028 8718 3074 8730
rect 2740 8330 2786 8342
rect 2822 8328 2832 8508
rect 2884 8328 2894 8508
rect 2932 8342 2938 8552
rect 2972 8342 2978 8552
rect 3028 8508 3034 8718
rect 3068 8508 3074 8718
rect 3110 8552 3120 8732
rect 3172 8552 3182 8732
rect 3220 8718 3266 8730
rect 2932 8330 2978 8342
rect 3014 8328 3024 8508
rect 3076 8328 3086 8508
rect 3124 8342 3130 8552
rect 3164 8342 3170 8552
rect 3220 8508 3226 8718
rect 3260 8508 3266 8718
rect 3302 8552 3312 8732
rect 3364 8552 3374 8732
rect 3412 8718 3458 8730
rect 3124 8330 3170 8342
rect 3206 8328 3216 8508
rect 3268 8328 3278 8508
rect 3316 8342 3322 8552
rect 3356 8342 3362 8552
rect 3412 8508 3418 8718
rect 3452 8508 3458 8718
rect 3494 8552 3504 8732
rect 3556 8552 3566 8732
rect 3604 8718 3650 8730
rect 3316 8330 3362 8342
rect 3398 8328 3408 8508
rect 3460 8328 3470 8508
rect 3508 8342 3514 8552
rect 3548 8342 3554 8552
rect 3604 8508 3610 8718
rect 3644 8508 3650 8718
rect 3734 8672 3806 8684
rect 3508 8330 3554 8342
rect 3590 8328 3600 8508
rect 3652 8328 3662 8508
rect 3730 8416 3740 8672
rect 3800 8416 3810 8672
rect 3928 8432 4588 8760
rect 5008 8432 5018 8984
rect 7156 8980 7576 9056
rect 5152 8768 7296 8816
rect 5152 8734 5174 8768
rect 5208 8734 5366 8768
rect 5400 8734 5558 8768
rect 5592 8734 5750 8768
rect 5784 8734 5942 8768
rect 5976 8734 6134 8768
rect 6168 8734 6326 8768
rect 6360 8734 6518 8768
rect 6552 8734 6710 8768
rect 6744 8734 6902 8768
rect 6936 8734 7296 8768
rect 5152 8728 7296 8734
rect 5120 8684 5166 8696
rect 5120 8476 5126 8684
rect 5160 8476 5166 8684
rect 5202 8520 5212 8700
rect 5268 8520 5278 8700
rect 5312 8684 5358 8696
rect 3734 8404 3806 8416
rect 3928 8300 4212 8432
rect 1724 8292 4212 8300
rect 5106 8296 5116 8476
rect 5172 8296 5182 8476
rect 5216 8308 5222 8520
rect 5256 8308 5262 8520
rect 5312 8476 5318 8684
rect 5352 8476 5358 8684
rect 5394 8520 5404 8700
rect 5460 8520 5470 8700
rect 5504 8684 5550 8696
rect 5216 8296 5262 8308
rect 5298 8296 5308 8476
rect 5364 8296 5374 8476
rect 5408 8308 5414 8520
rect 5448 8308 5454 8520
rect 5504 8476 5510 8684
rect 5544 8476 5550 8684
rect 5586 8520 5596 8700
rect 5652 8520 5662 8700
rect 5696 8684 5742 8696
rect 5408 8296 5454 8308
rect 5490 8296 5500 8476
rect 5556 8296 5566 8476
rect 5600 8308 5606 8520
rect 5640 8308 5646 8520
rect 5696 8476 5702 8684
rect 5736 8476 5742 8684
rect 5778 8520 5788 8700
rect 5844 8520 5854 8700
rect 5888 8684 5934 8696
rect 5600 8296 5646 8308
rect 5682 8296 5692 8476
rect 5748 8296 5758 8476
rect 5792 8308 5798 8520
rect 5832 8308 5838 8520
rect 5888 8476 5894 8684
rect 5928 8476 5934 8684
rect 5970 8520 5980 8700
rect 6036 8520 6046 8700
rect 6080 8684 6126 8696
rect 5792 8296 5838 8308
rect 5874 8296 5884 8476
rect 5940 8296 5950 8476
rect 5984 8308 5990 8520
rect 6024 8308 6030 8520
rect 6080 8476 6086 8684
rect 6120 8476 6126 8684
rect 6162 8520 6172 8700
rect 6228 8520 6238 8700
rect 6272 8684 6318 8696
rect 5984 8296 6030 8308
rect 6066 8296 6076 8476
rect 6132 8296 6142 8476
rect 6176 8308 6182 8520
rect 6216 8308 6222 8520
rect 6272 8476 6278 8684
rect 6312 8476 6318 8684
rect 6354 8520 6364 8700
rect 6420 8520 6430 8700
rect 6464 8684 6510 8696
rect 6176 8296 6222 8308
rect 6258 8296 6268 8476
rect 6324 8296 6334 8476
rect 6368 8308 6374 8520
rect 6408 8308 6414 8520
rect 6464 8476 6470 8684
rect 6504 8476 6510 8684
rect 6546 8520 6556 8700
rect 6612 8520 6622 8700
rect 6656 8684 6702 8696
rect 6368 8296 6414 8308
rect 6450 8296 6460 8476
rect 6516 8296 6526 8476
rect 6560 8308 6566 8520
rect 6600 8308 6606 8520
rect 6656 8476 6662 8684
rect 6696 8476 6702 8684
rect 6738 8520 6748 8700
rect 6804 8520 6814 8700
rect 6848 8684 6894 8696
rect 6560 8296 6606 8308
rect 6642 8296 6652 8476
rect 6708 8296 6718 8476
rect 6752 8308 6758 8520
rect 6792 8308 6798 8520
rect 6848 8476 6854 8684
rect 6888 8476 6894 8684
rect 6930 8520 6940 8700
rect 6996 8520 7006 8700
rect 7040 8684 7086 8696
rect 6752 8296 6798 8308
rect 6834 8296 6844 8476
rect 6900 8296 6910 8476
rect 6944 8308 6950 8520
rect 6984 8308 6990 8520
rect 7040 8476 7046 8684
rect 7080 8476 7086 8684
rect 6944 8296 6990 8308
rect 7026 8296 7036 8476
rect 7092 8296 7100 8476
rect 1724 8258 1738 8292
rect 1772 8258 1930 8292
rect 1964 8258 2122 8292
rect 2156 8258 2314 8292
rect 2348 8258 2506 8292
rect 2540 8258 2698 8292
rect 2732 8258 2890 8292
rect 2924 8258 3082 8292
rect 3116 8258 3274 8292
rect 3308 8258 3466 8292
rect 3500 8258 4212 8292
rect 7128 8264 7296 8728
rect 1724 8192 4212 8258
rect 1520 8154 1752 8160
rect 1520 8152 1976 8154
rect 2528 8152 2872 8154
rect 1520 8148 1764 8152
rect 1520 8088 1672 8148
rect 2056 8088 2066 8152
rect 2528 8088 2540 8152
rect 2860 8088 2872 8152
rect 1520 8084 1976 8088
rect 1520 7856 1604 8084
rect 1660 8082 1976 8084
rect 2528 8082 2872 8088
rect 3464 8152 3780 8158
rect 3464 8092 3476 8152
rect 3768 8092 3780 8152
rect 3464 8086 3780 8092
rect 3928 8044 4212 8192
rect 5252 8258 7296 8264
rect 5252 8224 5270 8258
rect 5304 8224 5462 8258
rect 5496 8224 5654 8258
rect 5688 8224 5846 8258
rect 5880 8224 6038 8258
rect 6072 8224 6230 8258
rect 6264 8224 6422 8258
rect 6456 8224 6614 8258
rect 6648 8224 6806 8258
rect 6840 8224 6998 8258
rect 7032 8224 7296 8258
rect 5252 8150 7296 8224
rect 5252 8116 5270 8150
rect 5304 8116 5462 8150
rect 5496 8116 5654 8150
rect 5688 8116 5846 8150
rect 5880 8116 6038 8150
rect 6072 8116 6230 8150
rect 6264 8116 6422 8150
rect 6456 8116 6614 8150
rect 6648 8116 6806 8150
rect 6840 8116 6998 8150
rect 7032 8116 7296 8150
rect 5252 8108 7296 8116
rect 1820 7982 4212 8044
rect 1820 7948 1834 7982
rect 1868 7948 2026 7982
rect 2060 7948 2218 7982
rect 2252 7948 2410 7982
rect 2444 7948 2602 7982
rect 2636 7948 2794 7982
rect 2828 7948 2986 7982
rect 3020 7948 3178 7982
rect 3212 7948 3370 7982
rect 3404 7948 3562 7982
rect 3596 7948 4212 7982
rect 1820 7940 4212 7948
rect 1684 7898 1730 7910
rect 1520 7844 1606 7856
rect 1520 7588 1540 7844
rect 1600 7588 1606 7844
rect 1684 7688 1690 7898
rect 1724 7688 1730 7898
rect 1766 7732 1776 7912
rect 1828 7732 1838 7912
rect 1876 7898 1922 7910
rect 1520 7576 1606 7588
rect 1520 7336 1604 7576
rect 1670 7508 1680 7688
rect 1732 7508 1742 7688
rect 1780 7522 1786 7732
rect 1820 7522 1826 7732
rect 1876 7688 1882 7898
rect 1916 7688 1922 7898
rect 1958 7732 1968 7912
rect 2020 7732 2030 7912
rect 2068 7898 2114 7910
rect 1780 7510 1826 7522
rect 1862 7508 1872 7688
rect 1924 7508 1934 7688
rect 1972 7522 1978 7732
rect 2012 7522 2018 7732
rect 2068 7688 2074 7898
rect 2108 7688 2114 7898
rect 2150 7732 2160 7912
rect 2212 7732 2222 7912
rect 2260 7898 2306 7910
rect 1972 7510 2018 7522
rect 2054 7508 2064 7688
rect 2116 7508 2126 7688
rect 2164 7522 2170 7732
rect 2204 7522 2210 7732
rect 2260 7688 2266 7898
rect 2300 7688 2306 7898
rect 2342 7732 2352 7912
rect 2404 7732 2414 7912
rect 2452 7898 2498 7910
rect 2164 7510 2210 7522
rect 2246 7508 2256 7688
rect 2308 7508 2318 7688
rect 2356 7522 2362 7732
rect 2396 7522 2402 7732
rect 2452 7688 2458 7898
rect 2492 7688 2498 7898
rect 2534 7732 2544 7912
rect 2596 7732 2606 7912
rect 2644 7898 2690 7910
rect 2356 7510 2402 7522
rect 2438 7508 2448 7688
rect 2500 7508 2510 7688
rect 2548 7522 2554 7732
rect 2588 7522 2594 7732
rect 2644 7688 2650 7898
rect 2684 7688 2690 7898
rect 2726 7732 2736 7912
rect 2788 7732 2798 7912
rect 2836 7898 2882 7910
rect 2548 7510 2594 7522
rect 2630 7508 2640 7688
rect 2692 7508 2702 7688
rect 2740 7522 2746 7732
rect 2780 7522 2786 7732
rect 2836 7688 2842 7898
rect 2876 7688 2882 7898
rect 2918 7732 2928 7912
rect 2980 7732 2990 7912
rect 3028 7898 3074 7910
rect 2740 7510 2786 7522
rect 2822 7508 2832 7688
rect 2884 7508 2894 7688
rect 2932 7522 2938 7732
rect 2972 7522 2978 7732
rect 3028 7688 3034 7898
rect 3068 7688 3074 7898
rect 3110 7732 3120 7912
rect 3172 7732 3182 7912
rect 3220 7898 3266 7910
rect 2932 7510 2978 7522
rect 3014 7508 3024 7688
rect 3076 7508 3086 7688
rect 3124 7522 3130 7732
rect 3164 7522 3170 7732
rect 3220 7688 3226 7898
rect 3260 7688 3266 7898
rect 3302 7732 3312 7912
rect 3364 7732 3374 7912
rect 3412 7898 3458 7910
rect 3124 7510 3170 7522
rect 3206 7508 3216 7688
rect 3268 7508 3278 7688
rect 3316 7522 3322 7732
rect 3356 7522 3362 7732
rect 3412 7688 3418 7898
rect 3452 7688 3458 7898
rect 3494 7732 3504 7912
rect 3556 7732 3566 7912
rect 3604 7898 3650 7910
rect 3316 7510 3362 7522
rect 3398 7508 3408 7688
rect 3460 7508 3470 7688
rect 3508 7522 3514 7732
rect 3548 7522 3554 7732
rect 3604 7688 3610 7898
rect 3644 7688 3650 7898
rect 3734 7824 3806 7836
rect 3508 7510 3554 7522
rect 3590 7508 3600 7688
rect 3652 7508 3662 7688
rect 3730 7568 3740 7824
rect 3800 7568 3810 7824
rect 3734 7556 3806 7568
rect 3928 7480 4212 7940
rect 5120 8066 5166 8078
rect 5120 7856 5126 8066
rect 5160 7856 5166 8066
rect 5202 7900 5212 8080
rect 5268 7900 5278 8080
rect 5312 8066 5358 8078
rect 5106 7676 5116 7856
rect 5172 7676 5182 7856
rect 5216 7690 5222 7900
rect 5256 7690 5262 7900
rect 5312 7856 5318 8066
rect 5352 7856 5358 8066
rect 5394 7900 5404 8080
rect 5460 7900 5470 8080
rect 5504 8066 5550 8078
rect 5216 7678 5262 7690
rect 5298 7676 5308 7856
rect 5364 7676 5374 7856
rect 5408 7690 5414 7900
rect 5448 7690 5454 7900
rect 5504 7856 5510 8066
rect 5544 7856 5550 8066
rect 5586 7900 5596 8080
rect 5652 7900 5662 8080
rect 5696 8066 5742 8078
rect 5408 7678 5454 7690
rect 5490 7676 5500 7856
rect 5556 7676 5566 7856
rect 5600 7690 5606 7900
rect 5640 7690 5646 7900
rect 5696 7856 5702 8066
rect 5736 7856 5742 8066
rect 5778 7900 5788 8080
rect 5844 7900 5854 8080
rect 5888 8066 5934 8078
rect 5600 7678 5646 7690
rect 5682 7676 5692 7856
rect 5748 7676 5758 7856
rect 5792 7690 5798 7900
rect 5832 7690 5838 7900
rect 5888 7856 5894 8066
rect 5928 7856 5934 8066
rect 5970 7900 5980 8080
rect 6036 7900 6046 8080
rect 6080 8066 6126 8078
rect 5792 7678 5838 7690
rect 5874 7676 5884 7856
rect 5940 7676 5950 7856
rect 5984 7690 5990 7900
rect 6024 7690 6030 7900
rect 6080 7856 6086 8066
rect 6120 7856 6126 8066
rect 6162 7900 6172 8080
rect 6228 7900 6238 8080
rect 6272 8066 6318 8078
rect 5984 7678 6030 7690
rect 6066 7676 6076 7856
rect 6132 7676 6142 7856
rect 6176 7690 6182 7900
rect 6216 7690 6222 7900
rect 6272 7856 6278 8066
rect 6312 7856 6318 8066
rect 6354 7900 6364 8080
rect 6420 7900 6430 8080
rect 6464 8066 6510 8078
rect 6176 7678 6222 7690
rect 6258 7676 6268 7856
rect 6324 7676 6334 7856
rect 6368 7690 6374 7900
rect 6408 7690 6414 7900
rect 6464 7856 6470 8066
rect 6504 7856 6510 8066
rect 6546 7900 6556 8080
rect 6612 7900 6622 8080
rect 6656 8066 6702 8078
rect 6368 7678 6414 7690
rect 6450 7676 6460 7856
rect 6516 7676 6526 7856
rect 6560 7690 6566 7900
rect 6600 7690 6606 7900
rect 6656 7856 6662 8066
rect 6696 7856 6702 8066
rect 6738 7900 6748 8080
rect 6804 7900 6814 8080
rect 6848 8066 6894 8078
rect 6560 7678 6606 7690
rect 6642 7676 6652 7856
rect 6708 7676 6718 7856
rect 6752 7690 6758 7900
rect 6792 7690 6798 7900
rect 6848 7856 6854 8066
rect 6888 7856 6894 8066
rect 6930 7900 6940 8080
rect 6996 7900 7006 8080
rect 7040 8066 7086 8078
rect 6752 7678 6798 7690
rect 6834 7676 6844 7856
rect 6900 7676 6910 7856
rect 6944 7690 6950 7900
rect 6984 7690 6990 7900
rect 7040 7856 7046 8066
rect 7080 7856 7086 8066
rect 6944 7678 6990 7690
rect 7026 7676 7036 7856
rect 7092 7676 7100 7856
rect 7128 7648 7296 8108
rect 5156 7640 7296 7648
rect 5156 7606 5174 7640
rect 5208 7606 5366 7640
rect 5400 7606 5558 7640
rect 5592 7606 5750 7640
rect 5784 7606 5942 7640
rect 5976 7606 6134 7640
rect 6168 7606 6326 7640
rect 6360 7606 6518 7640
rect 6552 7606 6710 7640
rect 6744 7606 6902 7640
rect 6936 7606 7296 7640
rect 5156 7572 7296 7606
rect 5392 7552 7296 7572
rect 1720 7472 4212 7480
rect 1720 7438 1738 7472
rect 1772 7438 1930 7472
rect 1964 7438 2122 7472
rect 2156 7438 2314 7472
rect 2348 7438 2506 7472
rect 2540 7438 2698 7472
rect 2732 7438 2890 7472
rect 2924 7438 3082 7472
rect 3116 7438 3274 7472
rect 3308 7438 3466 7472
rect 3500 7438 4212 7472
rect 1720 7372 4212 7438
rect 6372 7512 6568 7552
rect 6920 7512 7296 7552
rect 6372 7384 6384 7512
rect 1520 7328 2068 7336
rect 2528 7328 2844 7334
rect 1520 7268 1672 7328
rect 2056 7268 2068 7328
rect 2526 7268 2536 7328
rect 2832 7268 2844 7328
rect 1520 7260 2068 7268
rect 2528 7262 2844 7268
rect 3464 7328 3780 7334
rect 3464 7268 3476 7328
rect 3768 7268 3780 7328
rect 3464 7262 3780 7268
rect -9924 7028 -8884 7036
rect -10056 6986 -10010 6998
rect -10056 6776 -10050 6986
rect -10016 6776 -10010 6986
rect -9974 6820 -9964 7000
rect -9912 6820 -9902 7000
rect -9864 6986 -9818 6998
rect -10070 6596 -10060 6776
rect -10008 6596 -9998 6776
rect -9960 6610 -9954 6820
rect -9920 6610 -9914 6820
rect -9864 6776 -9858 6986
rect -9824 6776 -9818 6986
rect -9782 6820 -9772 7000
rect -9720 6820 -9710 7000
rect -9672 6986 -9626 6998
rect -9960 6598 -9914 6610
rect -9878 6596 -9868 6776
rect -9816 6596 -9806 6776
rect -9768 6610 -9762 6820
rect -9728 6610 -9722 6820
rect -9672 6776 -9666 6986
rect -9632 6776 -9626 6986
rect -9590 6820 -9580 7000
rect -9528 6820 -9518 7000
rect -9480 6986 -9434 6998
rect -9768 6598 -9722 6610
rect -9686 6596 -9676 6776
rect -9624 6596 -9614 6776
rect -9576 6610 -9570 6820
rect -9536 6610 -9530 6820
rect -9480 6776 -9474 6986
rect -9440 6776 -9434 6986
rect -9398 6820 -9388 7000
rect -9336 6820 -9326 7000
rect -9288 6986 -9242 6998
rect -9576 6598 -9530 6610
rect -9494 6596 -9484 6776
rect -9432 6596 -9422 6776
rect -9384 6610 -9378 6820
rect -9344 6610 -9338 6820
rect -9288 6776 -9282 6986
rect -9248 6776 -9242 6986
rect -9206 6820 -9196 7000
rect -9144 6820 -9134 7000
rect -9096 6986 -9050 6998
rect -9384 6598 -9338 6610
rect -9302 6596 -9292 6776
rect -9240 6596 -9230 6776
rect -9192 6610 -9186 6820
rect -9152 6610 -9146 6820
rect -9096 6776 -9090 6986
rect -9056 6776 -9050 6986
rect -9192 6598 -9146 6610
rect -9110 6596 -9100 6776
rect -9048 6596 -9038 6776
rect -9004 6568 -8884 7028
rect -8766 6828 -8756 7040
rect -8680 6828 -8670 7040
rect -8466 6832 -8456 7044
rect -8380 6832 -8370 7044
rect 1520 7004 1604 7260
rect 3928 7228 4212 7372
rect 1816 7162 4212 7228
rect 1816 7128 1834 7162
rect 1868 7128 2026 7162
rect 2060 7128 2218 7162
rect 2252 7128 2410 7162
rect 2444 7128 2602 7162
rect 2636 7128 2794 7162
rect 2828 7128 2986 7162
rect 3020 7128 3178 7162
rect 3212 7128 3370 7162
rect 3404 7128 3562 7162
rect 3596 7128 4212 7162
rect 1816 7120 4212 7128
rect -8748 6600 -8742 6828
rect -8708 6600 -8702 6828
rect -8748 6588 -8702 6600
rect -8438 6600 -8432 6832
rect -8398 6600 -8392 6832
rect -8438 6588 -8392 6600
rect 1520 6748 1536 7004
rect 1596 6748 1604 7004
rect 1684 7078 1730 7090
rect 1684 6868 1690 7078
rect 1724 6868 1730 7078
rect 1766 6912 1776 7092
rect 1828 6912 1838 7092
rect 1876 7078 1922 7090
rect -10020 6560 -8884 6568
rect -10020 6526 -10002 6560
rect -9968 6526 -9810 6560
rect -9776 6526 -9618 6560
rect -9584 6526 -9426 6560
rect -9392 6526 -9234 6560
rect -9200 6526 -8884 6560
rect -10020 6468 -8884 6526
rect -8670 6572 -8470 6578
rect -8670 6492 -8660 6572
rect -8480 6492 -8470 6572
rect 1520 6520 1604 6748
rect 1670 6688 1680 6868
rect 1732 6688 1742 6868
rect 1780 6702 1786 6912
rect 1820 6702 1826 6912
rect 1876 6868 1882 7078
rect 1916 6868 1922 7078
rect 1958 6912 1968 7092
rect 2020 6912 2030 7092
rect 2068 7078 2114 7090
rect 1780 6690 1826 6702
rect 1862 6688 1872 6868
rect 1924 6688 1934 6868
rect 1972 6702 1978 6912
rect 2012 6702 2018 6912
rect 2068 6868 2074 7078
rect 2108 6868 2114 7078
rect 2150 6912 2160 7092
rect 2212 6912 2222 7092
rect 2260 7078 2306 7090
rect 1972 6690 2018 6702
rect 2054 6688 2064 6868
rect 2116 6688 2126 6868
rect 2164 6702 2170 6912
rect 2204 6702 2210 6912
rect 2260 6868 2266 7078
rect 2300 6868 2306 7078
rect 2342 6912 2352 7092
rect 2404 6912 2414 7092
rect 2452 7078 2498 7090
rect 2164 6690 2210 6702
rect 2246 6688 2256 6868
rect 2308 6688 2318 6868
rect 2356 6702 2362 6912
rect 2396 6702 2402 6912
rect 2452 6868 2458 7078
rect 2492 6868 2498 7078
rect 2534 6912 2544 7092
rect 2596 6912 2606 7092
rect 2644 7078 2690 7090
rect 2356 6690 2402 6702
rect 2438 6688 2448 6868
rect 2500 6688 2510 6868
rect 2548 6702 2554 6912
rect 2588 6702 2594 6912
rect 2644 6868 2650 7078
rect 2684 6868 2690 7078
rect 2726 6912 2736 7092
rect 2788 6912 2798 7092
rect 2836 7078 2882 7090
rect 2548 6690 2594 6702
rect 2630 6688 2640 6868
rect 2692 6688 2702 6868
rect 2740 6702 2746 6912
rect 2780 6702 2786 6912
rect 2836 6868 2842 7078
rect 2876 6868 2882 7078
rect 2918 6912 2928 7092
rect 2980 6912 2990 7092
rect 3028 7078 3074 7090
rect 2740 6690 2786 6702
rect 2822 6688 2832 6868
rect 2884 6688 2894 6868
rect 2932 6702 2938 6912
rect 2972 6702 2978 6912
rect 3028 6868 3034 7078
rect 3068 6868 3074 7078
rect 3110 6912 3120 7092
rect 3172 6912 3182 7092
rect 3220 7078 3266 7090
rect 2932 6690 2978 6702
rect 3014 6688 3024 6868
rect 3076 6688 3086 6868
rect 3124 6702 3130 6912
rect 3164 6702 3170 6912
rect 3220 6868 3226 7078
rect 3260 6868 3266 7078
rect 3302 6912 3312 7092
rect 3364 6912 3374 7092
rect 3412 7078 3458 7090
rect 3124 6690 3170 6702
rect 3206 6688 3216 6868
rect 3268 6688 3278 6868
rect 3316 6702 3322 6912
rect 3356 6702 3362 6912
rect 3412 6868 3418 7078
rect 3452 6868 3458 7078
rect 3494 6912 3504 7092
rect 3556 6912 3566 7092
rect 3604 7078 3650 7090
rect 3316 6690 3362 6702
rect 3398 6688 3408 6868
rect 3460 6688 3470 6868
rect 3508 6702 3514 6912
rect 3548 6702 3554 6912
rect 3604 6868 3610 7078
rect 3644 6868 3650 7078
rect 3734 7012 3806 7024
rect 3508 6690 3554 6702
rect 3590 6688 3600 6868
rect 3652 6688 3662 6868
rect 3730 6756 3740 7012
rect 3800 6756 3810 7012
rect 3734 6744 3806 6756
rect 3928 6660 4212 7120
rect 6374 7000 6384 7384
rect 7076 7392 7296 7512
rect 7324 8596 7576 8980
rect 7620 9014 7666 9026
rect 7620 8808 7626 9014
rect 7660 8808 7666 9014
rect 7702 8844 7712 9028
rect 7768 8844 7778 9028
rect 7812 9014 7858 9026
rect 7606 8624 7616 8808
rect 7672 8624 7682 8808
rect 7716 8638 7722 8844
rect 7756 8638 7762 8844
rect 7812 8808 7818 9014
rect 7852 8808 7858 9014
rect 7894 8844 7904 9028
rect 7960 8844 7970 9028
rect 8004 9014 8050 9026
rect 7716 8626 7762 8638
rect 7798 8624 7808 8808
rect 7864 8624 7874 8808
rect 7908 8638 7914 8844
rect 7948 8638 7954 8844
rect 8004 8808 8010 9014
rect 8044 8808 8050 9014
rect 8086 8844 8096 9028
rect 8152 8844 8162 9028
rect 8196 9014 8242 9026
rect 7908 8626 7954 8638
rect 7990 8624 8000 8808
rect 8056 8624 8066 8808
rect 8100 8638 8106 8844
rect 8140 8638 8146 8844
rect 8196 8808 8202 9014
rect 8236 8808 8242 9014
rect 8278 8844 8288 9028
rect 8344 8844 8354 9028
rect 8388 9014 8434 9026
rect 8100 8626 8146 8638
rect 8182 8624 8192 8808
rect 8248 8624 8258 8808
rect 8292 8638 8298 8844
rect 8332 8638 8338 8844
rect 8388 8808 8394 9014
rect 8428 8808 8434 9014
rect 8470 8844 8480 9028
rect 8536 8844 8546 9028
rect 8580 9014 8626 9026
rect 8292 8626 8338 8638
rect 8374 8624 8384 8808
rect 8440 8624 8450 8808
rect 8484 8638 8490 8844
rect 8524 8638 8530 8844
rect 8580 8808 8586 9014
rect 8620 8808 8626 9014
rect 8662 8844 8672 9028
rect 8728 8844 8738 9028
rect 8772 9014 8818 9026
rect 8484 8626 8530 8638
rect 8566 8624 8576 8808
rect 8632 8624 8642 8808
rect 8676 8638 8682 8844
rect 8716 8638 8722 8844
rect 8772 8808 8778 9014
rect 8812 8808 8818 9014
rect 8854 8844 8864 9028
rect 8920 8844 8930 9028
rect 8964 9014 9010 9026
rect 8676 8626 8722 8638
rect 8758 8624 8768 8808
rect 8824 8624 8834 8808
rect 8868 8638 8874 8844
rect 8908 8638 8914 8844
rect 8964 8808 8970 9014
rect 9004 8808 9010 9014
rect 9046 8844 9056 9028
rect 9112 8844 9122 9028
rect 9156 9014 9202 9026
rect 8868 8626 8914 8638
rect 8950 8624 8960 8808
rect 9016 8624 9026 8808
rect 9060 8638 9066 8844
rect 9100 8638 9106 8844
rect 9156 8808 9162 9014
rect 9196 8808 9202 9014
rect 9238 8844 9248 9028
rect 9304 8844 9314 9028
rect 9348 9014 9394 9026
rect 9060 8626 9106 8638
rect 9142 8624 9152 8808
rect 9208 8624 9218 8808
rect 9252 8638 9258 8844
rect 9292 8638 9298 8844
rect 9348 8808 9354 9014
rect 9388 8808 9394 9014
rect 9430 8844 9440 9028
rect 9496 8844 9506 9028
rect 9540 9014 9586 9026
rect 9252 8626 9298 8638
rect 9334 8624 9344 8808
rect 9400 8624 9410 8808
rect 9444 8638 9450 8844
rect 9484 8638 9490 8844
rect 9540 8808 9546 9014
rect 9580 8808 9586 9014
rect 9444 8626 9490 8638
rect 9526 8624 9536 8808
rect 9592 8624 9602 8808
rect 7324 8588 9452 8596
rect 7324 8554 7674 8588
rect 7708 8554 7866 8588
rect 7900 8554 8058 8588
rect 8092 8554 8250 8588
rect 8284 8554 8442 8588
rect 8476 8554 8634 8588
rect 8668 8554 8826 8588
rect 8860 8554 9018 8588
rect 9052 8554 9210 8588
rect 9244 8554 9402 8588
rect 9436 8554 9452 8588
rect 7324 8480 9452 8554
rect 7324 8446 7674 8480
rect 7708 8446 7866 8480
rect 7900 8446 8058 8480
rect 8092 8446 8250 8480
rect 8284 8446 8442 8480
rect 8476 8446 8634 8480
rect 8668 8446 8826 8480
rect 8860 8446 9018 8480
rect 9052 8446 9210 8480
rect 9244 8446 9402 8480
rect 9436 8446 9452 8480
rect 7324 8440 9452 8446
rect 7324 7976 7576 8440
rect 7620 8396 7666 8408
rect 7620 8192 7626 8396
rect 7660 8192 7666 8396
rect 7702 8228 7712 8412
rect 7768 8228 7778 8412
rect 7812 8396 7858 8408
rect 7606 8008 7616 8192
rect 7672 8008 7682 8192
rect 7716 8020 7722 8228
rect 7756 8020 7762 8228
rect 7812 8192 7818 8396
rect 7852 8192 7858 8396
rect 7894 8228 7904 8412
rect 7960 8228 7970 8412
rect 8004 8396 8050 8408
rect 7716 8008 7762 8020
rect 7798 8008 7808 8192
rect 7864 8008 7874 8192
rect 7908 8020 7914 8228
rect 7948 8020 7954 8228
rect 8004 8192 8010 8396
rect 8044 8192 8050 8396
rect 8086 8228 8096 8412
rect 8152 8228 8162 8412
rect 8196 8396 8242 8408
rect 7908 8008 7954 8020
rect 7990 8008 8000 8192
rect 8056 8008 8066 8192
rect 8100 8020 8106 8228
rect 8140 8020 8146 8228
rect 8196 8192 8202 8396
rect 8236 8192 8242 8396
rect 8278 8228 8288 8412
rect 8344 8228 8354 8412
rect 8388 8396 8434 8408
rect 8100 8008 8146 8020
rect 8182 8008 8192 8192
rect 8248 8008 8258 8192
rect 8292 8020 8298 8228
rect 8332 8020 8338 8228
rect 8388 8192 8394 8396
rect 8428 8192 8434 8396
rect 8470 8228 8480 8412
rect 8536 8228 8546 8412
rect 8580 8396 8626 8408
rect 8292 8008 8338 8020
rect 8374 8008 8384 8192
rect 8440 8008 8450 8192
rect 8484 8020 8490 8228
rect 8524 8020 8530 8228
rect 8580 8192 8586 8396
rect 8620 8192 8626 8396
rect 8662 8228 8672 8412
rect 8728 8228 8738 8412
rect 8772 8396 8818 8408
rect 8484 8008 8530 8020
rect 8566 8008 8576 8192
rect 8632 8008 8642 8192
rect 8676 8020 8682 8228
rect 8716 8020 8722 8228
rect 8772 8192 8778 8396
rect 8812 8192 8818 8396
rect 8854 8228 8864 8412
rect 8920 8228 8930 8412
rect 8964 8396 9010 8408
rect 8676 8008 8722 8020
rect 8758 8008 8768 8192
rect 8824 8008 8834 8192
rect 8868 8020 8874 8228
rect 8908 8020 8914 8228
rect 8964 8192 8970 8396
rect 9004 8192 9010 8396
rect 9046 8228 9056 8412
rect 9112 8228 9122 8412
rect 9156 8396 9202 8408
rect 8868 8008 8914 8020
rect 8950 8008 8960 8192
rect 9016 8008 9026 8192
rect 9060 8020 9066 8228
rect 9100 8020 9106 8228
rect 9156 8192 9162 8396
rect 9196 8192 9202 8396
rect 9238 8228 9248 8412
rect 9304 8228 9314 8412
rect 9348 8396 9394 8408
rect 9060 8008 9106 8020
rect 9142 8008 9152 8192
rect 9208 8008 9218 8192
rect 9252 8020 9258 8228
rect 9292 8020 9298 8228
rect 9348 8192 9354 8396
rect 9388 8192 9394 8396
rect 9430 8228 9440 8412
rect 9496 8228 9506 8412
rect 9540 8396 9586 8408
rect 9252 8008 9298 8020
rect 9334 8008 9344 8192
rect 9400 8008 9410 8192
rect 9444 8020 9450 8228
rect 9484 8020 9490 8228
rect 9540 8192 9546 8396
rect 9580 8192 9586 8396
rect 9444 8008 9490 8020
rect 9526 8008 9536 8192
rect 9592 8008 9602 8192
rect 7324 7970 9548 7976
rect 7324 7936 7770 7970
rect 7804 7936 7962 7970
rect 7996 7936 8154 7970
rect 8188 7936 8346 7970
rect 8380 7936 8538 7970
rect 8572 7936 8730 7970
rect 8764 7936 8922 7970
rect 8956 7936 9114 7970
rect 9148 7936 9306 7970
rect 9340 7936 9498 7970
rect 9532 7936 9548 7970
rect 7324 7862 9548 7936
rect 7324 7828 7770 7862
rect 7804 7828 7962 7862
rect 7996 7828 8154 7862
rect 8188 7828 8346 7862
rect 8380 7828 8538 7862
rect 8572 7828 8730 7862
rect 8764 7828 8922 7862
rect 8956 7828 9114 7862
rect 9148 7828 9306 7862
rect 9340 7828 9498 7862
rect 9532 7828 9548 7862
rect 7324 7820 9548 7828
rect 7076 7000 7086 7392
rect 7324 7360 7576 7820
rect 7620 7778 7666 7790
rect 7620 7572 7626 7778
rect 7660 7572 7666 7778
rect 7702 7608 7712 7792
rect 7768 7608 7778 7792
rect 7812 7778 7858 7790
rect 7606 7388 7616 7572
rect 7672 7388 7682 7572
rect 7716 7402 7722 7608
rect 7756 7402 7762 7608
rect 7812 7572 7818 7778
rect 7852 7572 7858 7778
rect 7894 7608 7904 7792
rect 7960 7608 7970 7792
rect 8004 7778 8050 7790
rect 7716 7390 7762 7402
rect 7798 7388 7808 7572
rect 7864 7388 7874 7572
rect 7908 7402 7914 7608
rect 7948 7402 7954 7608
rect 8004 7572 8010 7778
rect 8044 7572 8050 7778
rect 8086 7608 8096 7792
rect 8152 7608 8162 7792
rect 8196 7778 8242 7790
rect 7908 7390 7954 7402
rect 7990 7388 8000 7572
rect 8056 7388 8066 7572
rect 8100 7402 8106 7608
rect 8140 7402 8146 7608
rect 8196 7572 8202 7778
rect 8236 7572 8242 7778
rect 8278 7608 8288 7792
rect 8344 7608 8354 7792
rect 8388 7778 8434 7790
rect 8100 7390 8146 7402
rect 8182 7388 8192 7572
rect 8248 7388 8258 7572
rect 8292 7402 8298 7608
rect 8332 7402 8338 7608
rect 8388 7572 8394 7778
rect 8428 7572 8434 7778
rect 8470 7608 8480 7792
rect 8536 7608 8546 7792
rect 8580 7778 8626 7790
rect 8292 7390 8338 7402
rect 8374 7388 8384 7572
rect 8440 7388 8450 7572
rect 8484 7402 8490 7608
rect 8524 7402 8530 7608
rect 8580 7572 8586 7778
rect 8620 7572 8626 7778
rect 8662 7608 8672 7792
rect 8728 7608 8738 7792
rect 8772 7778 8818 7790
rect 8484 7390 8530 7402
rect 8566 7388 8576 7572
rect 8632 7388 8642 7572
rect 8676 7402 8682 7608
rect 8716 7402 8722 7608
rect 8772 7572 8778 7778
rect 8812 7572 8818 7778
rect 8854 7608 8864 7792
rect 8920 7608 8930 7792
rect 8964 7778 9010 7790
rect 8676 7390 8722 7402
rect 8758 7388 8768 7572
rect 8824 7388 8834 7572
rect 8868 7402 8874 7608
rect 8908 7402 8914 7608
rect 8964 7572 8970 7778
rect 9004 7572 9010 7778
rect 9046 7608 9056 7792
rect 9112 7608 9122 7792
rect 9156 7778 9202 7790
rect 8868 7390 8914 7402
rect 8950 7388 8960 7572
rect 9016 7388 9026 7572
rect 9060 7402 9066 7608
rect 9100 7402 9106 7608
rect 9156 7572 9162 7778
rect 9196 7572 9202 7778
rect 9238 7608 9248 7792
rect 9304 7608 9314 7792
rect 9348 7778 9394 7790
rect 9060 7390 9106 7402
rect 9142 7388 9152 7572
rect 9208 7388 9218 7572
rect 9252 7402 9258 7608
rect 9292 7402 9298 7608
rect 9348 7572 9354 7778
rect 9388 7572 9394 7778
rect 9430 7608 9440 7792
rect 9496 7608 9506 7792
rect 9540 7778 9586 7790
rect 9252 7390 9298 7402
rect 9334 7388 9344 7572
rect 9400 7388 9410 7572
rect 9444 7402 9450 7608
rect 9484 7402 9490 7608
rect 9540 7572 9546 7778
rect 9580 7572 9586 7778
rect 9444 7390 9490 7402
rect 9526 7388 9536 7572
rect 9592 7388 9602 7572
rect 7156 7352 9452 7360
rect 7156 7318 7674 7352
rect 7708 7318 7866 7352
rect 7900 7318 8058 7352
rect 8092 7318 8250 7352
rect 8284 7318 8442 7352
rect 8476 7318 8634 7352
rect 8668 7318 8826 7352
rect 8860 7318 9018 7352
rect 9052 7318 9210 7352
rect 9244 7318 9402 7352
rect 9436 7318 9452 7352
rect 7156 7244 9452 7318
rect 7156 7210 7674 7244
rect 7708 7210 7866 7244
rect 7900 7210 8058 7244
rect 8092 7210 8250 7244
rect 8284 7210 8442 7244
rect 8476 7210 8634 7244
rect 8668 7210 8826 7244
rect 8860 7210 9018 7244
rect 9052 7210 9210 7244
rect 9244 7210 9402 7244
rect 9436 7210 9452 7244
rect 7156 7204 9452 7210
rect 7156 6928 7576 7204
rect 7620 7160 7666 7172
rect 7620 6956 7626 7160
rect 7660 6956 7666 7160
rect 7702 6992 7712 7176
rect 7768 6992 7778 7176
rect 7812 7160 7858 7172
rect 1724 6652 4212 6660
rect 1724 6618 1738 6652
rect 1772 6618 1930 6652
rect 1964 6618 2122 6652
rect 2156 6618 2314 6652
rect 2348 6618 2506 6652
rect 2540 6618 2698 6652
rect 2732 6618 2890 6652
rect 2924 6618 3082 6652
rect 3116 6618 3274 6652
rect 3308 6618 3466 6652
rect 3500 6618 4212 6652
rect 1724 6552 4212 6618
rect 6990 6600 7000 6928
rect 7528 6740 7576 6928
rect 7606 6772 7616 6956
rect 7672 6772 7682 6956
rect 7716 6784 7722 6992
rect 7756 6784 7762 6992
rect 7812 6956 7818 7160
rect 7852 6956 7858 7160
rect 7894 6992 7904 7176
rect 7960 6992 7970 7176
rect 8004 7160 8050 7172
rect 7716 6772 7762 6784
rect 7798 6772 7808 6956
rect 7864 6772 7874 6956
rect 7908 6784 7914 6992
rect 7948 6784 7954 6992
rect 8004 6956 8010 7160
rect 8044 6956 8050 7160
rect 8086 6992 8096 7176
rect 8152 6992 8162 7176
rect 8196 7160 8242 7172
rect 7908 6772 7954 6784
rect 7990 6772 8000 6956
rect 8056 6772 8066 6956
rect 8100 6784 8106 6992
rect 8140 6784 8146 6992
rect 8196 6956 8202 7160
rect 8236 6956 8242 7160
rect 8278 6992 8288 7176
rect 8344 6992 8354 7176
rect 8388 7160 8434 7172
rect 8100 6772 8146 6784
rect 8182 6772 8192 6956
rect 8248 6772 8258 6956
rect 8292 6784 8298 6992
rect 8332 6784 8338 6992
rect 8388 6956 8394 7160
rect 8428 6956 8434 7160
rect 8470 6992 8480 7176
rect 8536 6992 8546 7176
rect 8580 7160 8626 7172
rect 8292 6772 8338 6784
rect 8374 6772 8384 6956
rect 8440 6772 8450 6956
rect 8484 6784 8490 6992
rect 8524 6784 8530 6992
rect 8580 6956 8586 7160
rect 8620 6956 8626 7160
rect 8662 6992 8672 7176
rect 8728 6992 8738 7176
rect 8772 7160 8818 7172
rect 8484 6772 8530 6784
rect 8566 6772 8576 6956
rect 8632 6772 8642 6956
rect 8676 6784 8682 6992
rect 8716 6784 8722 6992
rect 8772 6956 8778 7160
rect 8812 6956 8818 7160
rect 8854 6992 8864 7176
rect 8920 6992 8930 7176
rect 8964 7160 9010 7172
rect 8676 6772 8722 6784
rect 8758 6772 8768 6956
rect 8824 6772 8834 6956
rect 8868 6784 8874 6992
rect 8908 6784 8914 6992
rect 8964 6956 8970 7160
rect 9004 6956 9010 7160
rect 9046 6992 9056 7176
rect 9112 6992 9122 7176
rect 9156 7160 9202 7172
rect 8868 6772 8914 6784
rect 8950 6772 8960 6956
rect 9016 6772 9026 6956
rect 9060 6784 9066 6992
rect 9100 6784 9106 6992
rect 9156 6956 9162 7160
rect 9196 6956 9202 7160
rect 9238 6992 9248 7176
rect 9304 6992 9314 7176
rect 9348 7160 9394 7172
rect 9060 6772 9106 6784
rect 9142 6772 9152 6956
rect 9208 6772 9218 6956
rect 9252 6784 9258 6992
rect 9292 6784 9298 6992
rect 9348 6956 9354 7160
rect 9388 6956 9394 7160
rect 9430 6992 9440 7176
rect 9496 6992 9506 7176
rect 9540 7160 9586 7172
rect 9252 6772 9298 6784
rect 9334 6772 9344 6956
rect 9400 6772 9410 6956
rect 9444 6784 9450 6992
rect 9484 6784 9490 6992
rect 9540 6956 9546 7160
rect 9580 6956 9586 7160
rect 9444 6772 9490 6784
rect 9526 6772 9536 6956
rect 9592 6772 9602 6956
rect 7528 6734 9548 6740
rect 7528 6700 7770 6734
rect 7804 6700 7962 6734
rect 7996 6700 8154 6734
rect 8188 6700 8346 6734
rect 8380 6700 8538 6734
rect 8572 6700 8730 6734
rect 8764 6700 8922 6734
rect 8956 6700 9114 6734
rect 9148 6700 9306 6734
rect 9340 6700 9498 6734
rect 9532 6700 9548 6734
rect 7528 6626 9548 6700
rect 7528 6600 7770 6626
rect 7156 6592 7770 6600
rect 7804 6592 7962 6626
rect 7996 6592 8154 6626
rect 8188 6592 8346 6626
rect 8380 6592 8538 6626
rect 8572 6592 8730 6626
rect 8764 6592 8922 6626
rect 8956 6592 9114 6626
rect 9148 6592 9306 6626
rect 9340 6592 9498 6626
rect 9532 6592 9548 6626
rect 7156 6584 9548 6592
rect 1660 6520 1976 6522
rect 1520 6516 1976 6520
rect 1520 6456 1672 6516
rect 1964 6456 1976 6516
rect 1520 6448 1976 6456
rect 2528 6516 2844 6522
rect 2528 6456 2540 6516
rect 2832 6456 2844 6516
rect 2528 6450 2844 6456
rect 3464 6512 3780 6518
rect 3464 6452 3476 6512
rect 3768 6452 3780 6512
rect 7156 6472 7576 6584
rect 3464 6446 3780 6452
rect -10060 6226 -8908 6268
rect -10060 6192 -9906 6226
rect -9872 6192 -9714 6226
rect -9680 6192 -9522 6226
rect -9488 6192 -9330 6226
rect -9296 6192 -9138 6226
rect -9104 6192 -8908 6226
rect -10060 6188 -8908 6192
rect -9918 6186 -9860 6188
rect -9726 6186 -9668 6188
rect -9534 6186 -9476 6188
rect -9342 6186 -9284 6188
rect -9150 6186 -9092 6188
rect -9008 6164 -8908 6188
rect -10056 6142 -10010 6154
rect -10056 5932 -10050 6142
rect -10016 5932 -10010 6142
rect -9974 5976 -9964 6156
rect -9912 5976 -9902 6156
rect -9864 6142 -9818 6154
rect -10070 5752 -10060 5932
rect -10008 5752 -9998 5932
rect -9960 5766 -9954 5976
rect -9920 5766 -9914 5976
rect -9864 5932 -9858 6142
rect -9824 5932 -9818 6142
rect -9782 5976 -9772 6156
rect -9720 5976 -9710 6156
rect -9672 6142 -9626 6154
rect -9960 5754 -9914 5766
rect -9878 5752 -9868 5932
rect -9816 5752 -9806 5932
rect -9768 5766 -9762 5976
rect -9728 5766 -9722 5976
rect -9672 5932 -9666 6142
rect -9632 5932 -9626 6142
rect -9590 5976 -9580 6156
rect -9528 5976 -9518 6156
rect -9480 6142 -9434 6154
rect -9768 5754 -9722 5766
rect -9686 5752 -9676 5932
rect -9624 5752 -9614 5932
rect -9576 5766 -9570 5976
rect -9536 5766 -9530 5976
rect -9480 5932 -9474 6142
rect -9440 5932 -9434 6142
rect -9398 5976 -9388 6156
rect -9336 5976 -9326 6156
rect -9288 6142 -9242 6154
rect -9576 5754 -9530 5766
rect -9494 5752 -9484 5932
rect -9432 5752 -9422 5932
rect -9384 5766 -9378 5976
rect -9344 5766 -9338 5976
rect -9288 5932 -9282 6142
rect -9248 5932 -9242 6142
rect -9206 5976 -9196 6156
rect -9144 5976 -9134 6156
rect -9096 6142 -9050 6154
rect -9384 5754 -9338 5766
rect -9302 5752 -9292 5932
rect -9240 5752 -9230 5932
rect -9192 5766 -9186 5976
rect -9152 5766 -9146 5976
rect -9096 5932 -9090 6142
rect -9056 5932 -9050 6142
rect -9008 5988 -8992 6164
rect -8824 5988 -8814 6164
rect 6950 6156 6960 6472
rect 7456 6156 7576 6472
rect 7620 6542 7666 6554
rect 7620 6336 7626 6542
rect 7660 6336 7666 6542
rect 7702 6372 7712 6556
rect 7768 6372 7778 6556
rect 7812 6542 7858 6554
rect 7156 6124 7576 6156
rect 7606 6152 7616 6336
rect 7672 6152 7682 6336
rect 7716 6166 7722 6372
rect 7756 6166 7762 6372
rect 7812 6336 7818 6542
rect 7852 6336 7858 6542
rect 7894 6372 7904 6556
rect 7960 6372 7970 6556
rect 8004 6542 8050 6554
rect 7716 6154 7762 6166
rect 7798 6152 7808 6336
rect 7864 6152 7874 6336
rect 7908 6166 7914 6372
rect 7948 6166 7954 6372
rect 8004 6336 8010 6542
rect 8044 6336 8050 6542
rect 8086 6372 8096 6556
rect 8152 6372 8162 6556
rect 8196 6542 8242 6554
rect 7908 6154 7954 6166
rect 7990 6152 8000 6336
rect 8056 6152 8066 6336
rect 8100 6166 8106 6372
rect 8140 6166 8146 6372
rect 8196 6336 8202 6542
rect 8236 6336 8242 6542
rect 8278 6372 8288 6556
rect 8344 6372 8354 6556
rect 8388 6542 8434 6554
rect 8100 6154 8146 6166
rect 8182 6152 8192 6336
rect 8248 6152 8258 6336
rect 8292 6166 8298 6372
rect 8332 6166 8338 6372
rect 8388 6336 8394 6542
rect 8428 6336 8434 6542
rect 8470 6372 8480 6556
rect 8536 6372 8546 6556
rect 8580 6542 8626 6554
rect 8292 6154 8338 6166
rect 8374 6152 8384 6336
rect 8440 6152 8450 6336
rect 8484 6166 8490 6372
rect 8524 6166 8530 6372
rect 8580 6336 8586 6542
rect 8620 6336 8626 6542
rect 8662 6372 8672 6556
rect 8728 6372 8738 6556
rect 8772 6542 8818 6554
rect 8484 6154 8530 6166
rect 8566 6152 8576 6336
rect 8632 6152 8642 6336
rect 8676 6166 8682 6372
rect 8716 6166 8722 6372
rect 8772 6336 8778 6542
rect 8812 6336 8818 6542
rect 8854 6372 8864 6556
rect 8920 6372 8930 6556
rect 8964 6542 9010 6554
rect 8676 6154 8722 6166
rect 8758 6152 8768 6336
rect 8824 6152 8834 6336
rect 8868 6166 8874 6372
rect 8908 6166 8914 6372
rect 8964 6336 8970 6542
rect 9004 6336 9010 6542
rect 9046 6372 9056 6556
rect 9112 6372 9122 6556
rect 9156 6542 9202 6554
rect 8868 6154 8914 6166
rect 8950 6152 8960 6336
rect 9016 6152 9026 6336
rect 9060 6166 9066 6372
rect 9100 6166 9106 6372
rect 9156 6336 9162 6542
rect 9196 6336 9202 6542
rect 9238 6372 9248 6556
rect 9304 6372 9314 6556
rect 9348 6542 9394 6554
rect 9060 6154 9106 6166
rect 9142 6152 9152 6336
rect 9208 6152 9218 6336
rect 9252 6166 9258 6372
rect 9292 6166 9298 6372
rect 9348 6336 9354 6542
rect 9388 6336 9394 6542
rect 9430 6372 9440 6556
rect 9496 6372 9506 6556
rect 9540 6542 9586 6554
rect 9252 6154 9298 6166
rect 9334 6152 9344 6336
rect 9400 6152 9410 6336
rect 9444 6166 9450 6372
rect 9484 6166 9490 6372
rect 9540 6336 9546 6542
rect 9580 6336 9586 6542
rect 9444 6154 9490 6166
rect 9526 6152 9536 6336
rect 9592 6152 9602 6336
rect 7156 6116 9452 6124
rect 7156 6082 7674 6116
rect 7708 6082 7866 6116
rect 7900 6082 8058 6116
rect 8092 6082 8250 6116
rect 8284 6082 8442 6116
rect 8476 6082 8634 6116
rect 8668 6082 8826 6116
rect 8860 6082 9018 6116
rect 9052 6082 9210 6116
rect 9244 6082 9402 6116
rect 9436 6082 9452 6116
rect 7156 6080 9452 6082
rect -396 5988 6664 6052
rect -9192 5754 -9146 5766
rect -9110 5752 -9100 5932
rect -9048 5752 -9038 5932
rect -10014 5716 -9956 5722
rect -9822 5716 -9764 5722
rect -9630 5716 -9572 5722
rect -9438 5716 -9380 5722
rect -9246 5716 -9188 5722
rect -9008 5716 -8908 5988
rect -10024 5682 -10002 5716
rect -9968 5682 -9810 5716
rect -9776 5682 -9618 5716
rect -9584 5682 -9426 5716
rect -9392 5682 -9234 5716
rect -9200 5682 -8908 5716
rect -10024 5608 -8908 5682
rect -10024 5574 -10002 5608
rect -9968 5574 -9810 5608
rect -9776 5574 -9618 5608
rect -9584 5574 -9426 5608
rect -9392 5574 -9234 5608
rect -9200 5574 -8908 5608
rect -10024 5572 -8908 5574
rect -10014 5568 -9956 5572
rect -9822 5568 -9764 5572
rect -9630 5568 -9572 5572
rect -9438 5568 -9380 5572
rect -9246 5568 -9188 5572
rect -10056 5524 -10010 5536
rect -10056 5316 -10050 5524
rect -10016 5316 -10010 5524
rect -9974 5360 -9964 5540
rect -9912 5360 -9902 5540
rect -9864 5524 -9818 5536
rect -10070 5136 -10060 5316
rect -10008 5136 -9998 5316
rect -9960 5148 -9954 5360
rect -9920 5148 -9914 5360
rect -9864 5316 -9858 5524
rect -9824 5316 -9818 5524
rect -9782 5360 -9772 5540
rect -9720 5360 -9710 5540
rect -9672 5524 -9626 5536
rect -9960 5136 -9914 5148
rect -9878 5136 -9868 5316
rect -9816 5136 -9806 5316
rect -9768 5148 -9762 5360
rect -9728 5148 -9722 5360
rect -9672 5316 -9666 5524
rect -9632 5316 -9626 5524
rect -9590 5360 -9580 5540
rect -9528 5360 -9518 5540
rect -9480 5524 -9434 5536
rect -9768 5136 -9722 5148
rect -9686 5136 -9676 5316
rect -9624 5136 -9614 5316
rect -9576 5148 -9570 5360
rect -9536 5148 -9530 5360
rect -9480 5316 -9474 5524
rect -9440 5316 -9434 5524
rect -9398 5360 -9388 5540
rect -9336 5360 -9326 5540
rect -9288 5524 -9242 5536
rect -9576 5136 -9530 5148
rect -9494 5136 -9484 5316
rect -9432 5136 -9422 5316
rect -9384 5148 -9378 5360
rect -9344 5148 -9338 5360
rect -9288 5316 -9282 5524
rect -9248 5316 -9242 5524
rect -9206 5360 -9196 5540
rect -9144 5360 -9134 5540
rect -9096 5524 -9050 5536
rect -9384 5136 -9338 5148
rect -9302 5136 -9292 5316
rect -9240 5136 -9230 5316
rect -9192 5148 -9186 5360
rect -9152 5148 -9146 5360
rect -9096 5316 -9090 5524
rect -9056 5316 -9050 5524
rect -9192 5136 -9146 5148
rect -9110 5136 -9100 5316
rect -9048 5136 -9038 5316
rect -9918 5100 -9860 5104
rect -9726 5100 -9668 5104
rect -9534 5100 -9476 5104
rect -9342 5100 -9284 5104
rect -9150 5100 -9092 5104
rect -9008 5100 -8908 5572
rect -9924 5098 -8908 5100
rect -9924 5064 -9906 5098
rect -9872 5064 -9714 5098
rect -9680 5064 -9522 5098
rect -9488 5064 -9330 5098
rect -9296 5064 -9138 5098
rect -9104 5064 -8908 5098
rect -396 5984 6768 5988
rect -396 5946 6904 5984
rect -396 5912 370 5946
rect 404 5912 562 5946
rect 596 5912 754 5946
rect 788 5912 946 5946
rect 980 5912 1138 5946
rect 1172 5912 2170 5946
rect 2204 5912 2362 5946
rect 2396 5912 2554 5946
rect 2588 5912 2746 5946
rect 2780 5912 2938 5946
rect 2972 5912 3970 5946
rect 4004 5912 4162 5946
rect 4196 5912 4354 5946
rect 4388 5912 4546 5946
rect 4580 5912 4738 5946
rect 4772 5912 5770 5946
rect 5804 5912 5962 5946
rect 5996 5912 6154 5946
rect 6188 5912 6346 5946
rect 6380 5912 6538 5946
rect 6572 5912 6904 5946
rect -396 5908 6904 5912
rect -396 5436 84 5908
rect 358 5906 416 5908
rect 550 5906 608 5908
rect 742 5906 800 5908
rect 934 5906 992 5908
rect 1126 5906 1184 5908
rect 220 5862 266 5874
rect 220 5652 226 5862
rect 260 5652 266 5862
rect 302 5696 312 5876
rect 364 5696 374 5876
rect 412 5862 458 5874
rect 206 5472 216 5652
rect 268 5472 278 5652
rect 316 5486 322 5696
rect 356 5486 362 5696
rect 412 5652 418 5862
rect 452 5652 458 5862
rect 494 5696 504 5876
rect 556 5696 566 5876
rect 604 5862 650 5874
rect 316 5474 362 5486
rect 398 5472 408 5652
rect 460 5472 470 5652
rect 508 5486 514 5696
rect 548 5486 554 5696
rect 604 5652 610 5862
rect 644 5652 650 5862
rect 686 5696 696 5876
rect 748 5696 758 5876
rect 796 5862 842 5874
rect 508 5474 554 5486
rect 590 5472 600 5652
rect 652 5472 662 5652
rect 700 5486 706 5696
rect 740 5486 746 5696
rect 796 5652 802 5862
rect 836 5652 842 5862
rect 878 5696 888 5876
rect 940 5696 950 5876
rect 988 5862 1034 5874
rect 700 5474 746 5486
rect 782 5472 792 5652
rect 844 5472 854 5652
rect 892 5486 898 5696
rect 932 5486 938 5696
rect 988 5652 994 5862
rect 1028 5652 1034 5862
rect 1070 5696 1080 5876
rect 1132 5696 1142 5876
rect 1180 5862 1226 5874
rect 892 5474 938 5486
rect 974 5472 984 5652
rect 1036 5472 1046 5652
rect 1084 5486 1090 5696
rect 1124 5486 1130 5696
rect 1180 5652 1186 5862
rect 1220 5652 1226 5862
rect 1084 5474 1130 5486
rect 1166 5472 1176 5652
rect 1228 5472 1238 5652
rect 262 5436 320 5442
rect 454 5436 512 5442
rect 646 5436 704 5442
rect 838 5436 896 5442
rect 1030 5436 1088 5442
rect 1268 5436 1500 5908
rect 2158 5906 2216 5908
rect 2350 5906 2408 5908
rect 2542 5906 2600 5908
rect 2734 5906 2792 5908
rect 2926 5906 2984 5908
rect 2020 5862 2066 5874
rect 2020 5652 2026 5862
rect 2060 5652 2066 5862
rect 2102 5696 2112 5876
rect 2164 5696 2174 5876
rect 2212 5862 2258 5874
rect 2006 5472 2016 5652
rect 2068 5472 2078 5652
rect 2116 5486 2122 5696
rect 2156 5486 2162 5696
rect 2212 5652 2218 5862
rect 2252 5652 2258 5862
rect 2294 5696 2304 5876
rect 2356 5696 2366 5876
rect 2404 5862 2450 5874
rect 2116 5474 2162 5486
rect 2198 5472 2208 5652
rect 2260 5472 2270 5652
rect 2308 5486 2314 5696
rect 2348 5486 2354 5696
rect 2404 5652 2410 5862
rect 2444 5652 2450 5862
rect 2486 5696 2496 5876
rect 2548 5696 2558 5876
rect 2596 5862 2642 5874
rect 2308 5474 2354 5486
rect 2390 5472 2400 5652
rect 2452 5472 2462 5652
rect 2500 5486 2506 5696
rect 2540 5486 2546 5696
rect 2596 5652 2602 5862
rect 2636 5652 2642 5862
rect 2678 5696 2688 5876
rect 2740 5696 2750 5876
rect 2788 5862 2834 5874
rect 2500 5474 2546 5486
rect 2582 5472 2592 5652
rect 2644 5472 2654 5652
rect 2692 5486 2698 5696
rect 2732 5486 2738 5696
rect 2788 5652 2794 5862
rect 2828 5652 2834 5862
rect 2870 5696 2880 5876
rect 2932 5696 2942 5876
rect 2980 5862 3026 5874
rect 2692 5474 2738 5486
rect 2774 5472 2784 5652
rect 2836 5472 2846 5652
rect 2884 5486 2890 5696
rect 2924 5486 2930 5696
rect 2980 5652 2986 5862
rect 3020 5652 3026 5862
rect 2884 5474 2930 5486
rect 2966 5472 2976 5652
rect 3028 5472 3038 5652
rect 2062 5436 2120 5442
rect 2254 5436 2312 5442
rect 2446 5436 2504 5442
rect 2638 5436 2696 5442
rect 2830 5436 2888 5442
rect 3068 5436 3304 5908
rect 3958 5906 4016 5908
rect 4150 5906 4208 5908
rect 4342 5906 4400 5908
rect 4534 5906 4592 5908
rect 4726 5906 4784 5908
rect 3820 5862 3866 5874
rect 3820 5652 3826 5862
rect 3860 5652 3866 5862
rect 3902 5696 3912 5876
rect 3964 5696 3974 5876
rect 4012 5862 4058 5874
rect 3806 5472 3816 5652
rect 3868 5472 3878 5652
rect 3916 5486 3922 5696
rect 3956 5486 3962 5696
rect 4012 5652 4018 5862
rect 4052 5652 4058 5862
rect 4094 5696 4104 5876
rect 4156 5696 4166 5876
rect 4204 5862 4250 5874
rect 3916 5474 3962 5486
rect 3998 5472 4008 5652
rect 4060 5472 4070 5652
rect 4108 5486 4114 5696
rect 4148 5486 4154 5696
rect 4204 5652 4210 5862
rect 4244 5652 4250 5862
rect 4286 5696 4296 5876
rect 4348 5696 4358 5876
rect 4396 5862 4442 5874
rect 4108 5474 4154 5486
rect 4190 5472 4200 5652
rect 4252 5472 4262 5652
rect 4300 5486 4306 5696
rect 4340 5486 4346 5696
rect 4396 5652 4402 5862
rect 4436 5652 4442 5862
rect 4478 5696 4488 5876
rect 4540 5696 4550 5876
rect 4588 5862 4634 5874
rect 4300 5474 4346 5486
rect 4382 5472 4392 5652
rect 4444 5472 4454 5652
rect 4492 5486 4498 5696
rect 4532 5486 4538 5696
rect 4588 5652 4594 5862
rect 4628 5652 4634 5862
rect 4670 5696 4680 5876
rect 4732 5696 4742 5876
rect 4780 5862 4826 5874
rect 4492 5474 4538 5486
rect 4574 5472 4584 5652
rect 4636 5472 4646 5652
rect 4684 5486 4690 5696
rect 4724 5486 4730 5696
rect 4780 5652 4786 5862
rect 4820 5652 4826 5862
rect 4684 5474 4730 5486
rect 4766 5472 4776 5652
rect 4828 5472 4838 5652
rect 3862 5436 3920 5442
rect 4054 5436 4112 5442
rect 4246 5436 4304 5442
rect 4438 5436 4496 5442
rect 4630 5436 4688 5442
rect 4868 5436 5104 5908
rect 5758 5906 5816 5908
rect 5950 5906 6008 5908
rect 6142 5906 6200 5908
rect 6334 5906 6392 5908
rect 6526 5906 6584 5908
rect 5620 5862 5666 5874
rect 5620 5652 5626 5862
rect 5660 5652 5666 5862
rect 5702 5696 5712 5876
rect 5764 5696 5774 5876
rect 5812 5862 5858 5874
rect 5606 5472 5616 5652
rect 5668 5472 5678 5652
rect 5716 5486 5722 5696
rect 5756 5486 5762 5696
rect 5812 5652 5818 5862
rect 5852 5652 5858 5862
rect 5894 5696 5904 5876
rect 5956 5696 5966 5876
rect 6004 5862 6050 5874
rect 5716 5474 5762 5486
rect 5798 5472 5808 5652
rect 5860 5472 5870 5652
rect 5908 5486 5914 5696
rect 5948 5486 5954 5696
rect 6004 5652 6010 5862
rect 6044 5652 6050 5862
rect 6086 5696 6096 5876
rect 6148 5696 6158 5876
rect 6196 5862 6242 5874
rect 5908 5474 5954 5486
rect 5990 5472 6000 5652
rect 6052 5472 6062 5652
rect 6100 5486 6106 5696
rect 6140 5486 6146 5696
rect 6196 5652 6202 5862
rect 6236 5652 6242 5862
rect 6278 5696 6288 5876
rect 6340 5696 6350 5876
rect 6388 5862 6434 5874
rect 6100 5474 6146 5486
rect 6182 5472 6192 5652
rect 6244 5472 6254 5652
rect 6292 5486 6298 5696
rect 6332 5486 6338 5696
rect 6388 5652 6394 5862
rect 6428 5652 6434 5862
rect 6470 5696 6480 5876
rect 6532 5696 6542 5876
rect 6580 5862 6626 5874
rect 6292 5474 6338 5486
rect 6374 5472 6384 5652
rect 6436 5472 6446 5652
rect 6484 5486 6490 5696
rect 6524 5486 6530 5696
rect 6580 5652 6586 5862
rect 6620 5652 6626 5862
rect 6484 5474 6530 5486
rect 6566 5472 6576 5652
rect 6628 5472 6638 5652
rect 5662 5436 5720 5442
rect 5854 5436 5912 5442
rect 6046 5436 6104 5442
rect 6238 5436 6296 5442
rect 6430 5436 6488 5442
rect 6668 5436 6904 5908
rect 7078 5580 7088 6080
rect 7372 6008 9452 6080
rect 7372 5974 7674 6008
rect 7708 5974 7866 6008
rect 7900 5974 8058 6008
rect 8092 5974 8250 6008
rect 8284 5974 8442 6008
rect 8476 5974 8634 6008
rect 8668 5974 8826 6008
rect 8860 5974 9018 6008
rect 9052 5974 9210 6008
rect 9244 5974 9402 6008
rect 9436 5974 9452 6008
rect 7372 5968 9452 5974
rect 7372 5580 7576 5968
rect 7620 5924 7666 5936
rect 7620 5720 7626 5924
rect 7660 5720 7666 5924
rect 7702 5756 7712 5940
rect 7768 5756 7778 5940
rect 7812 5924 7858 5936
rect -396 5402 274 5436
rect 308 5402 466 5436
rect 500 5402 658 5436
rect 692 5402 850 5436
rect 884 5402 1042 5436
rect 1076 5402 2074 5436
rect 2108 5402 2266 5436
rect 2300 5402 2458 5436
rect 2492 5402 2650 5436
rect 2684 5402 2842 5436
rect 2876 5402 3874 5436
rect 3908 5402 4066 5436
rect 4100 5402 4258 5436
rect 4292 5402 4450 5436
rect 4484 5402 4642 5436
rect 4676 5402 5674 5436
rect 5708 5402 5866 5436
rect 5900 5402 6058 5436
rect 6092 5402 6250 5436
rect 6284 5402 6442 5436
rect 6476 5402 6904 5436
rect -396 5328 6904 5402
rect -396 5294 274 5328
rect 308 5294 466 5328
rect 500 5294 658 5328
rect 692 5294 850 5328
rect 884 5294 1042 5328
rect 1076 5294 2074 5328
rect 2108 5294 2266 5328
rect 2300 5294 2458 5328
rect 2492 5294 2650 5328
rect 2684 5294 2842 5328
rect 2876 5294 3874 5328
rect 3908 5294 4066 5328
rect 4100 5294 4258 5328
rect 4292 5294 4450 5328
rect 4484 5294 4642 5328
rect 4676 5294 5674 5328
rect 5708 5294 5866 5328
rect 5900 5294 6058 5328
rect 6092 5294 6250 5328
rect 6284 5294 6442 5328
rect 6476 5294 6904 5328
rect -396 5292 6904 5294
rect -396 5092 84 5292
rect 262 5288 320 5292
rect 454 5288 512 5292
rect 646 5288 704 5292
rect 838 5288 896 5292
rect 1030 5288 1088 5292
rect -9924 4990 -8908 5064
rect -9924 4956 -9906 4990
rect -9872 4956 -9714 4990
rect -9680 4956 -9522 4990
rect -9488 4956 -9330 4990
rect -9296 4956 -9138 4990
rect -9104 4956 -8908 4990
rect -9918 4950 -9860 4956
rect -9726 4950 -9668 4956
rect -9534 4950 -9476 4956
rect -9342 4950 -9284 4956
rect -9150 4950 -9092 4956
rect -10056 4906 -10010 4918
rect -10056 4696 -10050 4906
rect -10016 4696 -10010 4906
rect -9974 4740 -9964 4920
rect -9912 4740 -9902 4920
rect -9864 4906 -9818 4918
rect -10070 4516 -10060 4696
rect -10008 4516 -9998 4696
rect -9960 4530 -9954 4740
rect -9920 4530 -9914 4740
rect -9864 4696 -9858 4906
rect -9824 4696 -9818 4906
rect -9782 4740 -9772 4920
rect -9720 4740 -9710 4920
rect -9672 4906 -9626 4918
rect -9960 4518 -9914 4530
rect -9878 4516 -9868 4696
rect -9816 4516 -9806 4696
rect -9768 4530 -9762 4740
rect -9728 4530 -9722 4740
rect -9672 4696 -9666 4906
rect -9632 4696 -9626 4906
rect -9590 4740 -9580 4920
rect -9528 4740 -9518 4920
rect -9480 4906 -9434 4918
rect -9768 4518 -9722 4530
rect -9686 4516 -9676 4696
rect -9624 4516 -9614 4696
rect -9576 4530 -9570 4740
rect -9536 4530 -9530 4740
rect -9480 4696 -9474 4906
rect -9440 4696 -9434 4906
rect -9398 4740 -9388 4920
rect -9336 4740 -9326 4920
rect -9288 4906 -9242 4918
rect -9576 4518 -9530 4530
rect -9494 4516 -9484 4696
rect -9432 4516 -9422 4696
rect -9384 4530 -9378 4740
rect -9344 4530 -9338 4740
rect -9288 4696 -9282 4906
rect -9248 4696 -9242 4906
rect -9206 4740 -9196 4920
rect -9144 4740 -9134 4920
rect -9096 4906 -9050 4918
rect -9384 4518 -9338 4530
rect -9302 4516 -9292 4696
rect -9240 4516 -9230 4696
rect -9192 4530 -9186 4740
rect -9152 4530 -9146 4740
rect -9096 4696 -9090 4906
rect -9056 4696 -9050 4906
rect -9192 4518 -9146 4530
rect -9110 4516 -9100 4696
rect -9048 4516 -9038 4696
rect -10014 4480 -9956 4486
rect -9822 4480 -9764 4486
rect -9630 4480 -9572 4486
rect -9438 4480 -9380 4486
rect -9246 4480 -9188 4486
rect -9008 4480 -8908 4956
rect -10020 4446 -10002 4480
rect -9968 4446 -9810 4480
rect -9776 4446 -9618 4480
rect -9584 4446 -9426 4480
rect -9392 4446 -9234 4480
rect -9200 4446 -8908 4480
rect -10020 4348 -8908 4446
rect -3192 4532 -3008 4568
rect -3192 4420 -3172 4532
rect -3028 4420 -3008 4532
rect -9460 4100 -9316 4348
rect -3192 4200 -3008 4420
rect -414 4400 -404 5092
rect 28 4820 84 5092
rect 220 5244 266 5256
rect 220 5036 226 5244
rect 260 5036 266 5244
rect 302 5080 312 5260
rect 364 5080 374 5260
rect 412 5244 458 5256
rect 206 4856 216 5036
rect 268 4856 278 5036
rect 316 4868 322 5080
rect 356 4868 362 5080
rect 412 5036 418 5244
rect 452 5036 458 5244
rect 494 5080 504 5260
rect 556 5080 566 5260
rect 604 5244 650 5256
rect 316 4856 362 4868
rect 398 4856 408 5036
rect 460 4856 470 5036
rect 508 4868 514 5080
rect 548 4868 554 5080
rect 604 5036 610 5244
rect 644 5036 650 5244
rect 686 5080 696 5260
rect 748 5080 758 5260
rect 796 5244 842 5256
rect 508 4856 554 4868
rect 590 4856 600 5036
rect 652 4856 662 5036
rect 700 4868 706 5080
rect 740 4868 746 5080
rect 796 5036 802 5244
rect 836 5036 842 5244
rect 878 5080 888 5260
rect 940 5080 950 5260
rect 988 5244 1034 5256
rect 700 4856 746 4868
rect 782 4856 792 5036
rect 844 4856 854 5036
rect 892 4868 898 5080
rect 932 4868 938 5080
rect 988 5036 994 5244
rect 1028 5036 1034 5244
rect 1070 5080 1080 5260
rect 1132 5080 1142 5260
rect 1180 5244 1226 5256
rect 892 4856 938 4868
rect 974 4856 984 5036
rect 1036 4856 1046 5036
rect 1084 4868 1090 5080
rect 1124 4868 1130 5080
rect 1180 5036 1186 5244
rect 1220 5036 1226 5244
rect 1084 4856 1130 4868
rect 1166 4856 1176 5036
rect 1228 4856 1238 5036
rect 358 4820 416 4824
rect 550 4820 608 4824
rect 742 4820 800 4824
rect 934 4820 992 4824
rect 1126 4820 1184 4824
rect 1268 4820 1500 5292
rect 2062 5288 2120 5292
rect 2254 5288 2312 5292
rect 2446 5288 2504 5292
rect 2638 5288 2696 5292
rect 2830 5288 2888 5292
rect 2020 5244 2066 5256
rect 2020 5036 2026 5244
rect 2060 5036 2066 5244
rect 2102 5080 2112 5260
rect 2164 5080 2174 5260
rect 2212 5244 2258 5256
rect 2006 4856 2016 5036
rect 2068 4856 2078 5036
rect 2116 4868 2122 5080
rect 2156 4868 2162 5080
rect 2212 5036 2218 5244
rect 2252 5036 2258 5244
rect 2294 5080 2304 5260
rect 2356 5080 2366 5260
rect 2404 5244 2450 5256
rect 2116 4856 2162 4868
rect 2198 4856 2208 5036
rect 2260 4856 2270 5036
rect 2308 4868 2314 5080
rect 2348 4868 2354 5080
rect 2404 5036 2410 5244
rect 2444 5036 2450 5244
rect 2486 5080 2496 5260
rect 2548 5080 2558 5260
rect 2596 5244 2642 5256
rect 2308 4856 2354 4868
rect 2390 4856 2400 5036
rect 2452 4856 2462 5036
rect 2500 4868 2506 5080
rect 2540 4868 2546 5080
rect 2596 5036 2602 5244
rect 2636 5036 2642 5244
rect 2678 5080 2688 5260
rect 2740 5080 2750 5260
rect 2788 5244 2834 5256
rect 2500 4856 2546 4868
rect 2582 4856 2592 5036
rect 2644 4856 2654 5036
rect 2692 4868 2698 5080
rect 2732 4868 2738 5080
rect 2788 5036 2794 5244
rect 2828 5036 2834 5244
rect 2870 5080 2880 5260
rect 2932 5080 2942 5260
rect 2980 5244 3026 5256
rect 2692 4856 2738 4868
rect 2774 4856 2784 5036
rect 2836 4856 2846 5036
rect 2884 4868 2890 5080
rect 2924 4868 2930 5080
rect 2980 5036 2986 5244
rect 3020 5036 3026 5244
rect 2884 4856 2930 4868
rect 2966 4856 2976 5036
rect 3028 4856 3038 5036
rect 2158 4820 2216 4824
rect 2350 4820 2408 4824
rect 2542 4820 2600 4824
rect 2734 4820 2792 4824
rect 2926 4820 2984 4824
rect 3068 4820 3304 5292
rect 3862 5288 3920 5292
rect 4054 5288 4112 5292
rect 4246 5288 4304 5292
rect 4438 5288 4496 5292
rect 4630 5288 4688 5292
rect 3820 5244 3866 5256
rect 3820 5036 3826 5244
rect 3860 5036 3866 5244
rect 3902 5080 3912 5260
rect 3964 5080 3974 5260
rect 4012 5244 4058 5256
rect 3806 4856 3816 5036
rect 3868 4856 3878 5036
rect 3916 4868 3922 5080
rect 3956 4868 3962 5080
rect 4012 5036 4018 5244
rect 4052 5036 4058 5244
rect 4094 5080 4104 5260
rect 4156 5080 4166 5260
rect 4204 5244 4250 5256
rect 3916 4856 3962 4868
rect 3998 4856 4008 5036
rect 4060 4856 4070 5036
rect 4108 4868 4114 5080
rect 4148 4868 4154 5080
rect 4204 5036 4210 5244
rect 4244 5036 4250 5244
rect 4286 5080 4296 5260
rect 4348 5080 4358 5260
rect 4396 5244 4442 5256
rect 4108 4856 4154 4868
rect 4190 4856 4200 5036
rect 4252 4856 4262 5036
rect 4300 4868 4306 5080
rect 4340 4868 4346 5080
rect 4396 5036 4402 5244
rect 4436 5036 4442 5244
rect 4478 5080 4488 5260
rect 4540 5080 4550 5260
rect 4588 5244 4634 5256
rect 4300 4856 4346 4868
rect 4382 4856 4392 5036
rect 4444 4856 4454 5036
rect 4492 4868 4498 5080
rect 4532 4868 4538 5080
rect 4588 5036 4594 5244
rect 4628 5036 4634 5244
rect 4670 5080 4680 5260
rect 4732 5080 4742 5260
rect 4780 5244 4826 5256
rect 4492 4856 4538 4868
rect 4574 4856 4584 5036
rect 4636 4856 4646 5036
rect 4684 4868 4690 5080
rect 4724 4868 4730 5080
rect 4780 5036 4786 5244
rect 4820 5036 4826 5244
rect 4684 4856 4730 4868
rect 4766 4856 4776 5036
rect 4828 4856 4838 5036
rect 3958 4820 4016 4824
rect 4150 4820 4208 4824
rect 4342 4820 4400 4824
rect 4534 4820 4592 4824
rect 4726 4820 4784 4824
rect 4868 4820 5104 5292
rect 5662 5288 5720 5292
rect 5854 5288 5912 5292
rect 6046 5288 6104 5292
rect 6238 5288 6296 5292
rect 6430 5288 6488 5292
rect 5620 5244 5666 5256
rect 5620 5036 5626 5244
rect 5660 5036 5666 5244
rect 5702 5080 5712 5260
rect 5764 5080 5774 5260
rect 5812 5244 5858 5256
rect 5606 4856 5616 5036
rect 5668 4856 5678 5036
rect 5716 4868 5722 5080
rect 5756 4868 5762 5080
rect 5812 5036 5818 5244
rect 5852 5036 5858 5244
rect 5894 5080 5904 5260
rect 5956 5080 5966 5260
rect 6004 5244 6050 5256
rect 5716 4856 5762 4868
rect 5798 4856 5808 5036
rect 5860 4856 5870 5036
rect 5908 4868 5914 5080
rect 5948 4868 5954 5080
rect 6004 5036 6010 5244
rect 6044 5036 6050 5244
rect 6086 5080 6096 5260
rect 6148 5080 6158 5260
rect 6196 5244 6242 5256
rect 5908 4856 5954 4868
rect 5990 4856 6000 5036
rect 6052 4856 6062 5036
rect 6100 4868 6106 5080
rect 6140 4868 6146 5080
rect 6196 5036 6202 5244
rect 6236 5036 6242 5244
rect 6278 5080 6288 5260
rect 6340 5080 6350 5260
rect 6388 5244 6434 5256
rect 6100 4856 6146 4868
rect 6182 4856 6192 5036
rect 6244 4856 6254 5036
rect 6292 4868 6298 5080
rect 6332 4868 6338 5080
rect 6388 5036 6394 5244
rect 6428 5036 6434 5244
rect 6470 5080 6480 5260
rect 6532 5080 6542 5260
rect 6580 5244 6626 5256
rect 6292 4856 6338 4868
rect 6374 4856 6384 5036
rect 6436 4856 6446 5036
rect 6484 4868 6490 5080
rect 6524 4868 6530 5080
rect 6580 5036 6586 5244
rect 6620 5036 6626 5244
rect 6484 4856 6530 4868
rect 6566 4856 6576 5036
rect 6628 4856 6638 5036
rect 5758 4820 5816 4824
rect 5950 4820 6008 4824
rect 6142 4820 6200 4824
rect 6334 4820 6392 4824
rect 6526 4820 6584 4824
rect 6668 4820 6904 5292
rect 28 4818 6904 4820
rect 28 4784 370 4818
rect 404 4784 562 4818
rect 596 4784 754 4818
rect 788 4784 946 4818
rect 980 4784 1138 4818
rect 1172 4784 2170 4818
rect 2204 4784 2362 4818
rect 2396 4784 2554 4818
rect 2588 4784 2746 4818
rect 2780 4784 2938 4818
rect 2972 4784 3970 4818
rect 4004 4784 4162 4818
rect 4196 4784 4354 4818
rect 4388 4784 4546 4818
rect 4580 4784 4738 4818
rect 4772 4784 5770 4818
rect 5804 4784 5962 4818
rect 5996 4784 6154 4818
rect 6188 4784 6346 4818
rect 6380 4784 6538 4818
rect 6572 4784 6904 4818
rect 7156 5504 7576 5580
rect 7606 5536 7616 5720
rect 7672 5536 7682 5720
rect 7716 5548 7722 5756
rect 7756 5548 7762 5756
rect 7812 5720 7818 5924
rect 7852 5720 7858 5924
rect 7894 5756 7904 5940
rect 7960 5756 7970 5940
rect 8004 5924 8050 5936
rect 7716 5536 7762 5548
rect 7798 5536 7808 5720
rect 7864 5536 7874 5720
rect 7908 5548 7914 5756
rect 7948 5548 7954 5756
rect 8004 5720 8010 5924
rect 8044 5720 8050 5924
rect 8086 5756 8096 5940
rect 8152 5756 8162 5940
rect 8196 5924 8242 5936
rect 7908 5536 7954 5548
rect 7990 5536 8000 5720
rect 8056 5536 8066 5720
rect 8100 5548 8106 5756
rect 8140 5548 8146 5756
rect 8196 5720 8202 5924
rect 8236 5720 8242 5924
rect 8278 5756 8288 5940
rect 8344 5756 8354 5940
rect 8388 5924 8434 5936
rect 8100 5536 8146 5548
rect 8182 5536 8192 5720
rect 8248 5536 8258 5720
rect 8292 5548 8298 5756
rect 8332 5548 8338 5756
rect 8388 5720 8394 5924
rect 8428 5720 8434 5924
rect 8470 5756 8480 5940
rect 8536 5756 8546 5940
rect 8580 5924 8626 5936
rect 8292 5536 8338 5548
rect 8374 5536 8384 5720
rect 8440 5536 8450 5720
rect 8484 5548 8490 5756
rect 8524 5548 8530 5756
rect 8580 5720 8586 5924
rect 8620 5720 8626 5924
rect 8662 5756 8672 5940
rect 8728 5756 8738 5940
rect 8772 5924 8818 5936
rect 8484 5536 8530 5548
rect 8566 5536 8576 5720
rect 8632 5536 8642 5720
rect 8676 5548 8682 5756
rect 8716 5548 8722 5756
rect 8772 5720 8778 5924
rect 8812 5720 8818 5924
rect 8854 5756 8864 5940
rect 8920 5756 8930 5940
rect 8964 5924 9010 5936
rect 8676 5536 8722 5548
rect 8758 5536 8768 5720
rect 8824 5536 8834 5720
rect 8868 5548 8874 5756
rect 8908 5548 8914 5756
rect 8964 5720 8970 5924
rect 9004 5720 9010 5924
rect 9046 5756 9056 5940
rect 9112 5756 9122 5940
rect 9156 5924 9202 5936
rect 8868 5536 8914 5548
rect 8950 5536 8960 5720
rect 9016 5536 9026 5720
rect 9060 5548 9066 5756
rect 9100 5548 9106 5756
rect 9156 5720 9162 5924
rect 9196 5720 9202 5924
rect 9238 5756 9248 5940
rect 9304 5756 9314 5940
rect 9348 5924 9394 5936
rect 9060 5536 9106 5548
rect 9142 5536 9152 5720
rect 9208 5536 9218 5720
rect 9252 5548 9258 5756
rect 9292 5548 9298 5756
rect 9348 5720 9354 5924
rect 9388 5720 9394 5924
rect 9430 5756 9440 5940
rect 9496 5756 9506 5940
rect 9540 5924 9586 5936
rect 9252 5536 9298 5548
rect 9334 5536 9344 5720
rect 9400 5536 9410 5720
rect 9444 5548 9450 5756
rect 9484 5548 9490 5756
rect 9540 5720 9546 5924
rect 9580 5720 9586 5924
rect 9444 5536 9490 5548
rect 9526 5536 9536 5720
rect 9592 5536 9602 5720
rect 7156 5498 9548 5504
rect 7156 5464 7770 5498
rect 7804 5464 7962 5498
rect 7996 5464 8154 5498
rect 8188 5464 8346 5498
rect 8380 5464 8538 5498
rect 8572 5464 8730 5498
rect 8764 5464 8922 5498
rect 8956 5464 9114 5498
rect 9148 5464 9306 5498
rect 9340 5464 9498 5498
rect 9532 5464 9548 5498
rect 7156 5390 9548 5464
rect 7156 5356 7770 5390
rect 7804 5356 7962 5390
rect 7996 5356 8154 5390
rect 8188 5356 8346 5390
rect 8380 5356 8538 5390
rect 8572 5356 8730 5390
rect 8764 5356 8922 5390
rect 8956 5356 9114 5390
rect 9148 5356 9306 5390
rect 9340 5356 9498 5390
rect 9532 5356 9548 5390
rect 7156 5348 9548 5356
rect 7156 4888 7576 5348
rect 7620 5306 7666 5318
rect 7620 5100 7626 5306
rect 7660 5100 7666 5306
rect 7702 5136 7712 5320
rect 7768 5136 7778 5320
rect 7812 5306 7858 5318
rect 7606 4916 7616 5100
rect 7672 4916 7682 5100
rect 7716 4930 7722 5136
rect 7756 4930 7762 5136
rect 7812 5100 7818 5306
rect 7852 5100 7858 5306
rect 7894 5136 7904 5320
rect 7960 5136 7970 5320
rect 8004 5306 8050 5318
rect 7716 4918 7762 4930
rect 7798 4916 7808 5100
rect 7864 4916 7874 5100
rect 7908 4930 7914 5136
rect 7948 4930 7954 5136
rect 8004 5100 8010 5306
rect 8044 5100 8050 5306
rect 8086 5136 8096 5320
rect 8152 5136 8162 5320
rect 8196 5306 8242 5318
rect 7908 4918 7954 4930
rect 7990 4916 8000 5100
rect 8056 4916 8066 5100
rect 8100 4930 8106 5136
rect 8140 4930 8146 5136
rect 8196 5100 8202 5306
rect 8236 5100 8242 5306
rect 8278 5136 8288 5320
rect 8344 5136 8354 5320
rect 8388 5306 8434 5318
rect 8100 4918 8146 4930
rect 8182 4916 8192 5100
rect 8248 4916 8258 5100
rect 8292 4930 8298 5136
rect 8332 4930 8338 5136
rect 8388 5100 8394 5306
rect 8428 5100 8434 5306
rect 8470 5136 8480 5320
rect 8536 5136 8546 5320
rect 8580 5306 8626 5318
rect 8292 4918 8338 4930
rect 8374 4916 8384 5100
rect 8440 4916 8450 5100
rect 8484 4930 8490 5136
rect 8524 4930 8530 5136
rect 8580 5100 8586 5306
rect 8620 5100 8626 5306
rect 8662 5136 8672 5320
rect 8728 5136 8738 5320
rect 8772 5306 8818 5318
rect 8484 4918 8530 4930
rect 8566 4916 8576 5100
rect 8632 4916 8642 5100
rect 8676 4930 8682 5136
rect 8716 4930 8722 5136
rect 8772 5100 8778 5306
rect 8812 5100 8818 5306
rect 8854 5136 8864 5320
rect 8920 5136 8930 5320
rect 8964 5306 9010 5318
rect 8676 4918 8722 4930
rect 8758 4916 8768 5100
rect 8824 4916 8834 5100
rect 8868 4930 8874 5136
rect 8908 4930 8914 5136
rect 8964 5100 8970 5306
rect 9004 5100 9010 5306
rect 9046 5136 9056 5320
rect 9112 5136 9122 5320
rect 9156 5306 9202 5318
rect 8868 4918 8914 4930
rect 8950 4916 8960 5100
rect 9016 4916 9026 5100
rect 9060 4930 9066 5136
rect 9100 4930 9106 5136
rect 9156 5100 9162 5306
rect 9196 5100 9202 5306
rect 9238 5136 9248 5320
rect 9304 5136 9314 5320
rect 9348 5306 9394 5318
rect 9060 4918 9106 4930
rect 9142 4916 9152 5100
rect 9208 4916 9218 5100
rect 9252 4930 9258 5136
rect 9292 4930 9298 5136
rect 9348 5100 9354 5306
rect 9388 5100 9394 5306
rect 9430 5136 9440 5320
rect 9496 5136 9506 5320
rect 9540 5306 9586 5318
rect 9252 4918 9298 4930
rect 9334 4916 9344 5100
rect 9400 4916 9410 5100
rect 9444 4930 9450 5136
rect 9484 4930 9490 5136
rect 9540 5100 9546 5306
rect 9580 5100 9586 5306
rect 9444 4918 9490 4930
rect 9526 4916 9536 5100
rect 9592 4916 9602 5100
rect 7156 4880 9452 4888
rect 7156 4846 7674 4880
rect 7708 4846 7866 4880
rect 7900 4846 8058 4880
rect 8092 4846 8250 4880
rect 8284 4846 8442 4880
rect 8476 4846 8634 4880
rect 8668 4846 8826 4880
rect 8860 4846 9018 4880
rect 9052 4846 9210 4880
rect 9244 4846 9402 4880
rect 9436 4846 9452 4880
rect 7156 4792 9452 4846
rect 28 4710 6904 4784
rect 28 4676 370 4710
rect 404 4676 562 4710
rect 596 4676 754 4710
rect 788 4676 946 4710
rect 980 4676 1138 4710
rect 1172 4676 2170 4710
rect 2204 4676 2362 4710
rect 2396 4676 2554 4710
rect 2588 4676 2746 4710
rect 2780 4676 2938 4710
rect 2972 4676 3970 4710
rect 4004 4676 4162 4710
rect 4196 4676 4354 4710
rect 4388 4676 4546 4710
rect 4580 4676 4738 4710
rect 4772 4676 5770 4710
rect 5804 4676 5962 4710
rect 5996 4676 6154 4710
rect 6188 4676 6346 4710
rect 6380 4676 6538 4710
rect 6572 4676 6904 4710
rect 28 4400 84 4676
rect 358 4670 416 4676
rect 550 4670 608 4676
rect 742 4670 800 4676
rect 934 4670 992 4676
rect 1126 4670 1184 4676
rect 220 4626 266 4638
rect 220 4416 226 4626
rect 260 4416 266 4626
rect 302 4460 312 4640
rect 364 4460 374 4640
rect 412 4626 458 4638
rect -396 4200 84 4400
rect 206 4236 216 4416
rect 268 4236 278 4416
rect 316 4250 322 4460
rect 356 4250 362 4460
rect 412 4416 418 4626
rect 452 4416 458 4626
rect 494 4460 504 4640
rect 556 4460 566 4640
rect 604 4626 650 4638
rect 316 4238 362 4250
rect 398 4236 408 4416
rect 460 4236 470 4416
rect 508 4250 514 4460
rect 548 4250 554 4460
rect 604 4416 610 4626
rect 644 4416 650 4626
rect 686 4460 696 4640
rect 748 4460 758 4640
rect 796 4626 842 4638
rect 508 4238 554 4250
rect 590 4236 600 4416
rect 652 4236 662 4416
rect 700 4250 706 4460
rect 740 4250 746 4460
rect 796 4416 802 4626
rect 836 4416 842 4626
rect 878 4460 888 4640
rect 940 4460 950 4640
rect 988 4626 1034 4638
rect 700 4238 746 4250
rect 782 4236 792 4416
rect 844 4236 854 4416
rect 892 4250 898 4460
rect 932 4250 938 4460
rect 988 4416 994 4626
rect 1028 4416 1034 4626
rect 1070 4460 1080 4640
rect 1132 4460 1142 4640
rect 1180 4626 1226 4638
rect 892 4238 938 4250
rect 974 4236 984 4416
rect 1036 4236 1046 4416
rect 1084 4250 1090 4460
rect 1124 4250 1130 4460
rect 1180 4416 1186 4626
rect 1220 4416 1226 4626
rect 1084 4238 1130 4250
rect 1166 4236 1176 4416
rect 1228 4236 1238 4416
rect 262 4200 320 4206
rect 454 4200 512 4206
rect 646 4200 704 4206
rect 838 4200 896 4206
rect 1030 4200 1088 4206
rect 1268 4200 1500 4676
rect 2158 4670 2216 4676
rect 2350 4670 2408 4676
rect 2542 4670 2600 4676
rect 2734 4670 2792 4676
rect 2926 4670 2984 4676
rect 2020 4626 2066 4638
rect 2020 4416 2026 4626
rect 2060 4416 2066 4626
rect 2102 4460 2112 4640
rect 2164 4460 2174 4640
rect 2212 4626 2258 4638
rect 2006 4236 2016 4416
rect 2068 4236 2078 4416
rect 2116 4250 2122 4460
rect 2156 4250 2162 4460
rect 2212 4416 2218 4626
rect 2252 4416 2258 4626
rect 2294 4460 2304 4640
rect 2356 4460 2366 4640
rect 2404 4626 2450 4638
rect 2116 4238 2162 4250
rect 2198 4236 2208 4416
rect 2260 4236 2270 4416
rect 2308 4250 2314 4460
rect 2348 4250 2354 4460
rect 2404 4416 2410 4626
rect 2444 4416 2450 4626
rect 2486 4460 2496 4640
rect 2548 4460 2558 4640
rect 2596 4626 2642 4638
rect 2308 4238 2354 4250
rect 2390 4236 2400 4416
rect 2452 4236 2462 4416
rect 2500 4250 2506 4460
rect 2540 4250 2546 4460
rect 2596 4416 2602 4626
rect 2636 4416 2642 4626
rect 2678 4460 2688 4640
rect 2740 4460 2750 4640
rect 2788 4626 2834 4638
rect 2500 4238 2546 4250
rect 2582 4236 2592 4416
rect 2644 4236 2654 4416
rect 2692 4250 2698 4460
rect 2732 4250 2738 4460
rect 2788 4416 2794 4626
rect 2828 4416 2834 4626
rect 2870 4460 2880 4640
rect 2932 4460 2942 4640
rect 2980 4626 3026 4638
rect 2692 4238 2738 4250
rect 2774 4236 2784 4416
rect 2836 4236 2846 4416
rect 2884 4250 2890 4460
rect 2924 4250 2930 4460
rect 2980 4416 2986 4626
rect 3020 4416 3026 4626
rect 2884 4238 2930 4250
rect 2966 4236 2976 4416
rect 3028 4236 3038 4416
rect 2062 4200 2120 4206
rect 2254 4200 2312 4206
rect 2446 4200 2504 4206
rect 2638 4200 2696 4206
rect 2830 4200 2888 4206
rect 3068 4200 3304 4676
rect 3958 4670 4016 4676
rect 4150 4670 4208 4676
rect 4342 4670 4400 4676
rect 4534 4670 4592 4676
rect 4726 4670 4784 4676
rect 3820 4626 3866 4638
rect 3820 4416 3826 4626
rect 3860 4416 3866 4626
rect 3902 4460 3912 4640
rect 3964 4460 3974 4640
rect 4012 4626 4058 4638
rect 3806 4236 3816 4416
rect 3868 4236 3878 4416
rect 3916 4250 3922 4460
rect 3956 4250 3962 4460
rect 4012 4416 4018 4626
rect 4052 4416 4058 4626
rect 4094 4460 4104 4640
rect 4156 4460 4166 4640
rect 4204 4626 4250 4638
rect 3916 4238 3962 4250
rect 3998 4236 4008 4416
rect 4060 4236 4070 4416
rect 4108 4250 4114 4460
rect 4148 4250 4154 4460
rect 4204 4416 4210 4626
rect 4244 4416 4250 4626
rect 4286 4460 4296 4640
rect 4348 4460 4358 4640
rect 4396 4626 4442 4638
rect 4108 4238 4154 4250
rect 4190 4236 4200 4416
rect 4252 4236 4262 4416
rect 4300 4250 4306 4460
rect 4340 4250 4346 4460
rect 4396 4416 4402 4626
rect 4436 4416 4442 4626
rect 4478 4460 4488 4640
rect 4540 4460 4550 4640
rect 4588 4626 4634 4638
rect 4300 4238 4346 4250
rect 4382 4236 4392 4416
rect 4444 4236 4454 4416
rect 4492 4250 4498 4460
rect 4532 4250 4538 4460
rect 4588 4416 4594 4626
rect 4628 4416 4634 4626
rect 4670 4460 4680 4640
rect 4732 4460 4742 4640
rect 4780 4626 4826 4638
rect 4492 4238 4538 4250
rect 4574 4236 4584 4416
rect 4636 4236 4646 4416
rect 4684 4250 4690 4460
rect 4724 4250 4730 4460
rect 4780 4416 4786 4626
rect 4820 4416 4826 4626
rect 4684 4238 4730 4250
rect 4766 4236 4776 4416
rect 4828 4236 4838 4416
rect 3862 4200 3920 4206
rect 4054 4200 4112 4206
rect 4246 4200 4304 4206
rect 4438 4200 4496 4206
rect 4630 4200 4688 4206
rect 4868 4200 5104 4676
rect 5758 4670 5816 4676
rect 5950 4670 6008 4676
rect 6142 4670 6200 4676
rect 6334 4670 6392 4676
rect 6526 4670 6584 4676
rect 5620 4626 5666 4638
rect 5620 4416 5626 4626
rect 5660 4416 5666 4626
rect 5702 4460 5712 4640
rect 5764 4460 5774 4640
rect 5812 4626 5858 4638
rect 5606 4236 5616 4416
rect 5668 4236 5678 4416
rect 5716 4250 5722 4460
rect 5756 4250 5762 4460
rect 5812 4416 5818 4626
rect 5852 4416 5858 4626
rect 5894 4460 5904 4640
rect 5956 4460 5966 4640
rect 6004 4626 6050 4638
rect 5716 4238 5762 4250
rect 5798 4236 5808 4416
rect 5860 4236 5870 4416
rect 5908 4250 5914 4460
rect 5948 4250 5954 4460
rect 6004 4416 6010 4626
rect 6044 4416 6050 4626
rect 6086 4460 6096 4640
rect 6148 4460 6158 4640
rect 6196 4626 6242 4638
rect 5908 4238 5954 4250
rect 5990 4236 6000 4416
rect 6052 4236 6062 4416
rect 6100 4250 6106 4460
rect 6140 4250 6146 4460
rect 6196 4416 6202 4626
rect 6236 4416 6242 4626
rect 6278 4460 6288 4640
rect 6340 4460 6350 4640
rect 6388 4626 6434 4638
rect 6100 4238 6146 4250
rect 6182 4236 6192 4416
rect 6244 4236 6254 4416
rect 6292 4250 6298 4460
rect 6332 4250 6338 4460
rect 6388 4416 6394 4626
rect 6428 4416 6434 4626
rect 6470 4460 6480 4640
rect 6532 4460 6542 4640
rect 6580 4626 6626 4638
rect 6292 4238 6338 4250
rect 6374 4236 6384 4416
rect 6436 4236 6446 4416
rect 6484 4250 6490 4460
rect 6524 4250 6530 4460
rect 6580 4416 6586 4626
rect 6620 4416 6626 4626
rect 6484 4238 6530 4250
rect 6566 4236 6576 4416
rect 6628 4236 6638 4416
rect 5662 4200 5720 4206
rect 5854 4200 5912 4206
rect 6046 4200 6104 4206
rect 6238 4200 6296 4206
rect 6430 4200 6488 4206
rect 6668 4200 6904 4676
rect 9840 4200 10160 16980
rect 10800 7928 11300 17652
rect 11480 11940 11900 20780
rect 18164 21108 18260 21460
rect 18304 21534 18350 21546
rect 18304 21324 18310 21534
rect 18344 21324 18350 21534
rect 18386 21368 18396 21548
rect 18448 21368 18458 21548
rect 18496 21534 18542 21546
rect 18294 21144 18304 21324
rect 18356 21144 18366 21324
rect 18400 21158 18406 21368
rect 18440 21158 18446 21368
rect 18496 21324 18502 21534
rect 18536 21324 18542 21534
rect 18578 21368 18588 21548
rect 18640 21368 18650 21548
rect 18688 21534 18734 21546
rect 18400 21146 18446 21158
rect 18482 21144 18492 21324
rect 18544 21144 18554 21324
rect 18592 21158 18598 21368
rect 18632 21158 18638 21368
rect 18688 21324 18694 21534
rect 18728 21324 18734 21534
rect 18770 21368 18780 21548
rect 18832 21368 18842 21548
rect 18880 21534 18926 21546
rect 18592 21146 18638 21158
rect 18674 21144 18684 21324
rect 18736 21144 18746 21324
rect 18784 21158 18790 21368
rect 18824 21158 18830 21368
rect 18880 21324 18886 21534
rect 18920 21324 18926 21534
rect 18962 21368 18972 21548
rect 19024 21368 19034 21548
rect 19072 21534 19118 21546
rect 18784 21146 18830 21158
rect 18866 21144 18876 21324
rect 18928 21144 18938 21324
rect 18976 21158 18982 21368
rect 19016 21158 19022 21368
rect 19072 21324 19078 21534
rect 19112 21324 19118 21534
rect 19154 21368 19164 21548
rect 19216 21368 19226 21548
rect 19264 21534 19310 21546
rect 18976 21146 19022 21158
rect 19058 21144 19068 21324
rect 19120 21144 19130 21324
rect 19168 21158 19174 21368
rect 19208 21158 19214 21368
rect 19264 21324 19270 21534
rect 19304 21324 19310 21534
rect 19168 21146 19214 21158
rect 19250 21144 19260 21324
rect 19312 21144 19322 21324
rect 18442 21108 18500 21114
rect 18634 21108 18692 21114
rect 18826 21108 18884 21114
rect 19018 21108 19076 21114
rect 19210 21108 19268 21114
rect 18164 21074 18454 21108
rect 18488 21074 18646 21108
rect 18680 21074 18838 21108
rect 18872 21074 19030 21108
rect 19064 21074 19222 21108
rect 19256 21074 19312 21108
rect 18164 20980 19312 21074
rect 18164 20868 18260 20980
rect 18164 20752 19588 20868
rect 18164 20718 18372 20752
rect 18540 20718 18630 20752
rect 18798 20718 18888 20752
rect 19056 20718 19146 20752
rect 19314 20718 19404 20752
rect 19572 20718 19588 20752
rect 18164 20712 19588 20718
rect 18164 20248 18260 20712
rect 18304 20668 18350 20680
rect 18304 20460 18310 20668
rect 18344 20460 18350 20668
rect 18550 20504 18560 20684
rect 18612 20504 18622 20684
rect 18820 20668 18866 20680
rect 18290 20280 18300 20460
rect 18352 20280 18362 20460
rect 18562 20292 18568 20504
rect 18602 20292 18608 20504
rect 18820 20460 18826 20668
rect 18860 20460 18866 20668
rect 19066 20504 19076 20684
rect 19128 20504 19138 20684
rect 19336 20668 19382 20680
rect 18562 20280 18608 20292
rect 18806 20280 18816 20460
rect 18868 20280 18878 20460
rect 19078 20292 19084 20504
rect 19118 20292 19124 20504
rect 19336 20460 19342 20668
rect 19376 20460 19382 20668
rect 19582 20504 19592 20684
rect 19644 20504 19654 20684
rect 19078 20280 19124 20292
rect 19322 20280 19332 20460
rect 19384 20280 19394 20460
rect 19594 20292 19600 20504
rect 19634 20292 19640 20504
rect 19594 20280 19640 20292
rect 18164 20242 19588 20248
rect 18164 20208 18372 20242
rect 18540 20208 18630 20242
rect 18798 20208 18888 20242
rect 19056 20208 19146 20242
rect 19314 20208 19404 20242
rect 19572 20208 19588 20242
rect 18164 20134 19588 20208
rect 18164 20100 18372 20134
rect 18540 20100 18630 20134
rect 18798 20100 18888 20134
rect 19056 20100 19146 20134
rect 19314 20100 19404 20134
rect 19572 20100 19588 20134
rect 18164 20092 19588 20100
rect 18164 19632 18260 20092
rect 18304 20050 18350 20062
rect 18304 19840 18310 20050
rect 18344 19840 18350 20050
rect 18550 19884 18560 20064
rect 18612 19884 18622 20064
rect 18820 20050 18866 20062
rect 18290 19660 18300 19840
rect 18352 19660 18362 19840
rect 18562 19674 18568 19884
rect 18602 19674 18608 19884
rect 18820 19840 18826 20050
rect 18860 19840 18866 20050
rect 19066 19884 19076 20064
rect 19128 19884 19138 20064
rect 19336 20050 19382 20062
rect 18562 19662 18608 19674
rect 18806 19660 18816 19840
rect 18868 19660 18878 19840
rect 19078 19674 19084 19884
rect 19118 19674 19124 19884
rect 19336 19840 19342 20050
rect 19376 19840 19382 20050
rect 19582 19884 19592 20064
rect 19644 19884 19654 20064
rect 19078 19662 19124 19674
rect 19322 19660 19332 19840
rect 19384 19660 19394 19840
rect 19594 19674 19600 19884
rect 19634 19674 19640 19884
rect 19594 19662 19640 19674
rect 18164 19624 19588 19632
rect 18164 19590 18372 19624
rect 18540 19590 18630 19624
rect 18798 19590 18888 19624
rect 19056 19590 19146 19624
rect 19314 19590 19404 19624
rect 19572 19590 19588 19624
rect 18164 19516 19588 19590
rect 18164 19482 18372 19516
rect 18540 19482 18630 19516
rect 18798 19482 18888 19516
rect 19056 19482 19146 19516
rect 19314 19482 19404 19516
rect 19572 19482 19588 19516
rect 18164 19476 19588 19482
rect 18164 19012 18260 19476
rect 18304 19432 18350 19444
rect 18304 19224 18310 19432
rect 18344 19224 18350 19432
rect 18550 19268 18560 19448
rect 18612 19268 18622 19448
rect 18820 19432 18866 19444
rect 18290 19044 18300 19224
rect 18352 19044 18362 19224
rect 18562 19056 18568 19268
rect 18602 19056 18608 19268
rect 18820 19224 18826 19432
rect 18860 19224 18866 19432
rect 19066 19268 19076 19448
rect 19128 19268 19138 19448
rect 19336 19432 19382 19444
rect 18562 19044 18608 19056
rect 18806 19044 18816 19224
rect 18868 19044 18878 19224
rect 19078 19056 19084 19268
rect 19118 19056 19124 19268
rect 19336 19224 19342 19432
rect 19376 19224 19382 19432
rect 19582 19268 19592 19448
rect 19644 19268 19654 19448
rect 19078 19044 19124 19056
rect 19322 19044 19332 19224
rect 19384 19044 19394 19224
rect 19594 19056 19600 19268
rect 19634 19056 19640 19268
rect 19594 19044 19640 19056
rect 18164 19006 19588 19012
rect 18164 18972 18372 19006
rect 18540 18972 18630 19006
rect 18798 18972 18888 19006
rect 19056 18972 19146 19006
rect 19314 18972 19404 19006
rect 19572 18972 19588 19006
rect 18164 18898 19588 18972
rect 18164 18864 18372 18898
rect 18540 18864 18630 18898
rect 18798 18864 18888 18898
rect 19056 18864 19146 18898
rect 19314 18864 19404 18898
rect 19572 18864 19588 18898
rect 18164 18856 19588 18864
rect 18164 18396 18260 18856
rect 18304 18814 18350 18826
rect 18304 18604 18310 18814
rect 18344 18604 18350 18814
rect 18550 18648 18560 18828
rect 18612 18648 18622 18828
rect 18820 18814 18866 18826
rect 18290 18424 18300 18604
rect 18352 18424 18362 18604
rect 18562 18438 18568 18648
rect 18602 18438 18608 18648
rect 18820 18604 18826 18814
rect 18860 18604 18866 18814
rect 19066 18648 19076 18828
rect 19128 18648 19138 18828
rect 19336 18814 19382 18826
rect 18562 18426 18608 18438
rect 18806 18424 18816 18604
rect 18868 18424 18878 18604
rect 19078 18438 19084 18648
rect 19118 18438 19124 18648
rect 19336 18604 19342 18814
rect 19376 18604 19382 18814
rect 19582 18648 19592 18828
rect 19644 18648 19654 18828
rect 19078 18426 19124 18438
rect 19322 18424 19332 18604
rect 19384 18424 19394 18604
rect 19594 18438 19600 18648
rect 19634 18438 19640 18648
rect 19594 18426 19640 18438
rect 18164 18388 19588 18396
rect 18164 18354 18372 18388
rect 18540 18354 18630 18388
rect 18798 18354 18888 18388
rect 19056 18354 19146 18388
rect 19314 18354 19404 18388
rect 19572 18354 19588 18388
rect 18164 18240 19588 18354
rect 18468 18156 18692 18162
rect 18468 18056 18480 18156
rect 18680 18056 18692 18156
rect 18468 18050 18692 18056
rect 11480 11500 24900 11940
rect 10790 7472 10800 7928
rect 11300 7472 11310 7928
rect 11480 4920 11900 11500
rect 15688 10768 15980 10774
rect 15688 10532 15700 10768
rect 15968 10532 15980 10768
rect 16978 10660 16988 11148
rect 19192 10660 19202 11148
rect 20490 10808 20682 10820
rect 20486 10608 20496 10808
rect 20676 10608 20686 10808
rect 20490 10596 20682 10608
rect 15688 10526 15980 10532
rect 21124 10428 21976 10436
rect 19556 10388 21976 10428
rect 19556 10364 23948 10388
rect 19556 10330 19574 10364
rect 19608 10330 19766 10364
rect 19800 10330 19958 10364
rect 19992 10330 20150 10364
rect 20184 10330 20342 10364
rect 20376 10330 20534 10364
rect 20568 10330 20726 10364
rect 20760 10330 20918 10364
rect 20952 10330 21110 10364
rect 21144 10330 21302 10364
rect 21336 10334 23948 10364
rect 21336 10330 22170 10334
rect 19556 10324 22170 10330
rect 21556 10300 22170 10324
rect 22204 10300 22362 10334
rect 22396 10300 22554 10334
rect 22588 10300 22746 10334
rect 22780 10300 22938 10334
rect 22972 10300 23130 10334
rect 23164 10300 23322 10334
rect 23356 10300 23514 10334
rect 23548 10300 23706 10334
rect 23740 10300 23898 10334
rect 23932 10300 23948 10334
rect 21556 10292 23948 10300
rect 19520 10271 19566 10283
rect 19520 10060 19526 10271
rect 19560 10060 19566 10271
rect 19602 10104 19612 10284
rect 19668 10104 19678 10284
rect 19712 10271 19758 10283
rect 16978 9440 16988 9908
rect 19180 9440 19190 9908
rect 19506 9880 19516 10060
rect 19572 9880 19582 10060
rect 19616 9895 19622 10104
rect 19656 9895 19662 10104
rect 19712 10060 19718 10271
rect 19752 10060 19758 10271
rect 19794 10104 19804 10284
rect 19860 10104 19870 10284
rect 19904 10271 19950 10283
rect 19616 9883 19662 9895
rect 19698 9880 19708 10060
rect 19764 9880 19774 10060
rect 19808 9895 19814 10104
rect 19848 9895 19854 10104
rect 19904 10060 19910 10271
rect 19944 10060 19950 10271
rect 19986 10104 19996 10284
rect 20052 10104 20062 10284
rect 20096 10271 20142 10283
rect 19808 9883 19854 9895
rect 19890 9880 19900 10060
rect 19956 9880 19966 10060
rect 20000 9895 20006 10104
rect 20040 9895 20046 10104
rect 20096 10060 20102 10271
rect 20136 10060 20142 10271
rect 20178 10104 20188 10284
rect 20244 10104 20254 10284
rect 20288 10271 20334 10283
rect 20000 9883 20046 9895
rect 20082 9880 20092 10060
rect 20148 9880 20158 10060
rect 20192 9895 20198 10104
rect 20232 9895 20238 10104
rect 20288 10060 20294 10271
rect 20328 10060 20334 10271
rect 20370 10104 20380 10284
rect 20436 10104 20446 10284
rect 20480 10271 20526 10283
rect 20192 9883 20238 9895
rect 20274 9880 20284 10060
rect 20340 9880 20350 10060
rect 20384 9895 20390 10104
rect 20424 9895 20430 10104
rect 20480 10060 20486 10271
rect 20520 10060 20526 10271
rect 20562 10104 20572 10284
rect 20628 10104 20638 10284
rect 20672 10271 20718 10283
rect 20384 9883 20430 9895
rect 20466 9880 20476 10060
rect 20532 9880 20542 10060
rect 20576 9895 20582 10104
rect 20616 9895 20622 10104
rect 20672 10060 20678 10271
rect 20712 10060 20718 10271
rect 20754 10104 20764 10284
rect 20820 10104 20830 10284
rect 20864 10271 20910 10283
rect 20576 9883 20622 9895
rect 20658 9880 20668 10060
rect 20724 9880 20734 10060
rect 20768 9895 20774 10104
rect 20808 9895 20814 10104
rect 20864 10060 20870 10271
rect 20904 10060 20910 10271
rect 20946 10104 20956 10284
rect 21012 10104 21022 10284
rect 21056 10271 21102 10283
rect 20768 9883 20814 9895
rect 20850 9880 20860 10060
rect 20916 9880 20926 10060
rect 20960 9895 20966 10104
rect 21000 9895 21006 10104
rect 21056 10060 21062 10271
rect 21096 10060 21102 10271
rect 21138 10104 21148 10284
rect 21204 10104 21214 10284
rect 21248 10271 21294 10283
rect 20960 9883 21006 9895
rect 21042 9880 21052 10060
rect 21108 9880 21118 10060
rect 21152 9895 21158 10104
rect 21192 9895 21198 10104
rect 21248 10060 21254 10271
rect 21288 10060 21294 10271
rect 21330 10104 21340 10284
rect 21396 10104 21406 10284
rect 21440 10271 21486 10283
rect 21152 9883 21198 9895
rect 21234 9880 21244 10060
rect 21300 9880 21310 10060
rect 21344 9895 21350 10104
rect 21384 9895 21390 10104
rect 21440 10060 21446 10271
rect 21480 10060 21486 10271
rect 21344 9883 21390 9895
rect 21426 9880 21436 10060
rect 21492 9880 21502 10060
rect 21556 9844 21976 10292
rect 22020 10250 22066 10262
rect 22020 10044 22026 10250
rect 22060 10044 22066 10250
rect 22102 10080 22112 10264
rect 22168 10080 22178 10264
rect 22212 10250 22258 10262
rect 22006 9860 22016 10044
rect 22072 9860 22082 10044
rect 22116 9874 22122 10080
rect 22156 9874 22162 10080
rect 22212 10044 22218 10250
rect 22252 10044 22258 10250
rect 22294 10080 22304 10264
rect 22360 10080 22370 10264
rect 22404 10250 22450 10262
rect 22116 9862 22162 9874
rect 22198 9860 22208 10044
rect 22264 9860 22274 10044
rect 22308 9874 22314 10080
rect 22348 9874 22354 10080
rect 22404 10044 22410 10250
rect 22444 10044 22450 10250
rect 22486 10080 22496 10264
rect 22552 10080 22562 10264
rect 22596 10250 22642 10262
rect 22308 9862 22354 9874
rect 22390 9860 22400 10044
rect 22456 9860 22466 10044
rect 22500 9874 22506 10080
rect 22540 9874 22546 10080
rect 22596 10044 22602 10250
rect 22636 10044 22642 10250
rect 22678 10080 22688 10264
rect 22744 10080 22754 10264
rect 22788 10250 22834 10262
rect 22500 9862 22546 9874
rect 22582 9860 22592 10044
rect 22648 9860 22658 10044
rect 22692 9874 22698 10080
rect 22732 9874 22738 10080
rect 22788 10044 22794 10250
rect 22828 10044 22834 10250
rect 22870 10080 22880 10264
rect 22936 10080 22946 10264
rect 22980 10250 23026 10262
rect 22692 9862 22738 9874
rect 22774 9860 22784 10044
rect 22840 9860 22850 10044
rect 22884 9874 22890 10080
rect 22924 9874 22930 10080
rect 22980 10044 22986 10250
rect 23020 10044 23026 10250
rect 23062 10080 23072 10264
rect 23128 10080 23138 10264
rect 23172 10250 23218 10262
rect 22884 9862 22930 9874
rect 22966 9860 22976 10044
rect 23032 9860 23042 10044
rect 23076 9874 23082 10080
rect 23116 9874 23122 10080
rect 23172 10044 23178 10250
rect 23212 10044 23218 10250
rect 23254 10080 23264 10264
rect 23320 10080 23330 10264
rect 23364 10250 23410 10262
rect 23076 9862 23122 9874
rect 23158 9860 23168 10044
rect 23224 9860 23234 10044
rect 23268 9874 23274 10080
rect 23308 9874 23314 10080
rect 23364 10044 23370 10250
rect 23404 10044 23410 10250
rect 23446 10080 23456 10264
rect 23512 10080 23522 10264
rect 23556 10250 23602 10262
rect 23268 9862 23314 9874
rect 23350 9860 23360 10044
rect 23416 9860 23426 10044
rect 23460 9874 23466 10080
rect 23500 9874 23506 10080
rect 23556 10044 23562 10250
rect 23596 10044 23602 10250
rect 23638 10080 23648 10264
rect 23704 10080 23714 10264
rect 23748 10250 23794 10262
rect 23460 9862 23506 9874
rect 23542 9860 23552 10044
rect 23608 9860 23618 10044
rect 23652 9874 23658 10080
rect 23692 9874 23698 10080
rect 23748 10044 23754 10250
rect 23788 10044 23794 10250
rect 23830 10080 23840 10264
rect 23896 10080 23906 10264
rect 23940 10250 23986 10262
rect 23652 9862 23698 9874
rect 23734 9860 23744 10044
rect 23800 9860 23810 10044
rect 23844 9874 23850 10080
rect 23884 9874 23890 10080
rect 23940 10044 23946 10250
rect 23980 10044 23986 10250
rect 23844 9862 23890 9874
rect 23926 9860 23936 10044
rect 23992 9860 24002 10044
rect 19652 9836 21976 9844
rect 19652 9802 19670 9836
rect 19704 9802 19862 9836
rect 19896 9802 20054 9836
rect 20088 9802 20246 9836
rect 20280 9802 20438 9836
rect 20472 9802 20630 9836
rect 20664 9802 20822 9836
rect 20856 9802 21014 9836
rect 21048 9802 21206 9836
rect 21240 9802 21398 9836
rect 21432 9832 21976 9836
rect 21432 9824 23852 9832
rect 21432 9802 22074 9824
rect 19652 9790 22074 9802
rect 22108 9790 22266 9824
rect 22300 9790 22458 9824
rect 22492 9790 22650 9824
rect 22684 9790 22842 9824
rect 22876 9790 23034 9824
rect 23068 9790 23226 9824
rect 23260 9790 23418 9824
rect 23452 9790 23610 9824
rect 23644 9790 23802 9824
rect 23836 9790 23852 9824
rect 19652 9728 23852 9790
rect 19652 9694 19670 9728
rect 19704 9694 19862 9728
rect 19896 9694 20054 9728
rect 20088 9694 20246 9728
rect 20280 9694 20438 9728
rect 20472 9694 20630 9728
rect 20664 9694 20822 9728
rect 20856 9694 21014 9728
rect 21048 9694 21206 9728
rect 21240 9694 21398 9728
rect 21432 9716 23852 9728
rect 21432 9694 22074 9716
rect 19652 9688 22074 9694
rect 21556 9682 22074 9688
rect 22108 9682 22266 9716
rect 22300 9682 22458 9716
rect 22492 9682 22650 9716
rect 22684 9682 22842 9716
rect 22876 9682 23034 9716
rect 23068 9682 23226 9716
rect 23260 9682 23418 9716
rect 23452 9682 23610 9716
rect 23644 9682 23802 9716
rect 23836 9682 23852 9716
rect 21556 9676 23852 9682
rect 19520 9635 19566 9647
rect 19520 9428 19526 9635
rect 19560 9428 19566 9635
rect 19602 9472 19612 9652
rect 19668 9472 19678 9652
rect 19712 9635 19758 9647
rect 19506 9248 19516 9428
rect 19572 9248 19582 9428
rect 19616 9259 19622 9472
rect 19656 9259 19662 9472
rect 19712 9428 19718 9635
rect 19752 9428 19758 9635
rect 19794 9472 19804 9652
rect 19860 9472 19870 9652
rect 19904 9635 19950 9647
rect 19520 9247 19566 9248
rect 19616 9247 19662 9259
rect 19698 9248 19708 9428
rect 19764 9248 19774 9428
rect 19808 9259 19814 9472
rect 19848 9259 19854 9472
rect 19904 9428 19910 9635
rect 19944 9428 19950 9635
rect 19986 9472 19996 9652
rect 20052 9472 20062 9652
rect 20096 9635 20142 9647
rect 19712 9247 19758 9248
rect 19808 9247 19854 9259
rect 19890 9248 19900 9428
rect 19956 9248 19966 9428
rect 20000 9259 20006 9472
rect 20040 9259 20046 9472
rect 20096 9428 20102 9635
rect 20136 9428 20142 9635
rect 20178 9472 20188 9652
rect 20244 9472 20254 9652
rect 20288 9635 20334 9647
rect 19904 9247 19950 9248
rect 20000 9247 20046 9259
rect 20082 9248 20092 9428
rect 20148 9248 20158 9428
rect 20192 9259 20198 9472
rect 20232 9259 20238 9472
rect 20288 9428 20294 9635
rect 20328 9428 20334 9635
rect 20370 9472 20380 9652
rect 20436 9472 20446 9652
rect 20480 9635 20526 9647
rect 20096 9247 20142 9248
rect 20192 9247 20238 9259
rect 20274 9248 20284 9428
rect 20340 9248 20350 9428
rect 20384 9259 20390 9472
rect 20424 9259 20430 9472
rect 20480 9428 20486 9635
rect 20520 9428 20526 9635
rect 20562 9472 20572 9652
rect 20628 9472 20638 9652
rect 20672 9635 20718 9647
rect 20288 9247 20334 9248
rect 20384 9247 20430 9259
rect 20466 9248 20476 9428
rect 20532 9248 20542 9428
rect 20576 9259 20582 9472
rect 20616 9259 20622 9472
rect 20672 9428 20678 9635
rect 20712 9428 20718 9635
rect 20754 9472 20764 9652
rect 20820 9472 20830 9652
rect 20864 9635 20910 9647
rect 20480 9247 20526 9248
rect 20576 9247 20622 9259
rect 20658 9248 20668 9428
rect 20724 9248 20734 9428
rect 20768 9259 20774 9472
rect 20808 9259 20814 9472
rect 20864 9428 20870 9635
rect 20904 9428 20910 9635
rect 20946 9472 20956 9652
rect 21012 9472 21022 9652
rect 21056 9635 21102 9647
rect 20672 9247 20718 9248
rect 20768 9247 20814 9259
rect 20850 9248 20860 9428
rect 20916 9248 20926 9428
rect 20960 9259 20966 9472
rect 21000 9259 21006 9472
rect 21056 9428 21062 9635
rect 21096 9428 21102 9635
rect 21138 9472 21148 9652
rect 21204 9472 21214 9652
rect 21248 9635 21294 9647
rect 20864 9247 20910 9248
rect 20960 9247 21006 9259
rect 21042 9248 21052 9428
rect 21108 9248 21118 9428
rect 21152 9259 21158 9472
rect 21192 9259 21198 9472
rect 21248 9428 21254 9635
rect 21288 9428 21294 9635
rect 21330 9472 21340 9652
rect 21396 9472 21406 9652
rect 21440 9635 21486 9647
rect 21056 9247 21102 9248
rect 21152 9247 21198 9259
rect 21234 9248 21244 9428
rect 21300 9248 21310 9428
rect 21344 9259 21350 9472
rect 21384 9259 21390 9472
rect 21440 9428 21446 9635
rect 21480 9428 21486 9635
rect 21248 9247 21294 9248
rect 21344 9247 21390 9259
rect 21426 9248 21436 9428
rect 21492 9248 21502 9428
rect 21440 9247 21486 9248
rect 21556 9212 21976 9676
rect 22020 9632 22066 9644
rect 22020 9428 22026 9632
rect 22060 9428 22066 9632
rect 22102 9464 22112 9648
rect 22168 9464 22178 9648
rect 22212 9632 22258 9644
rect 22006 9244 22016 9428
rect 22072 9244 22082 9428
rect 22116 9256 22122 9464
rect 22156 9256 22162 9464
rect 22212 9428 22218 9632
rect 22252 9428 22258 9632
rect 22294 9464 22304 9648
rect 22360 9464 22370 9648
rect 22404 9632 22450 9644
rect 22116 9244 22162 9256
rect 22198 9244 22208 9428
rect 22264 9244 22274 9428
rect 22308 9256 22314 9464
rect 22348 9256 22354 9464
rect 22404 9428 22410 9632
rect 22444 9428 22450 9632
rect 22486 9464 22496 9648
rect 22552 9464 22562 9648
rect 22596 9632 22642 9644
rect 22308 9244 22354 9256
rect 22390 9244 22400 9428
rect 22456 9244 22466 9428
rect 22500 9256 22506 9464
rect 22540 9256 22546 9464
rect 22596 9428 22602 9632
rect 22636 9428 22642 9632
rect 22678 9464 22688 9648
rect 22744 9464 22754 9648
rect 22788 9632 22834 9644
rect 22500 9244 22546 9256
rect 22582 9244 22592 9428
rect 22648 9244 22658 9428
rect 22692 9256 22698 9464
rect 22732 9256 22738 9464
rect 22788 9428 22794 9632
rect 22828 9428 22834 9632
rect 22870 9464 22880 9648
rect 22936 9464 22946 9648
rect 22980 9632 23026 9644
rect 22692 9244 22738 9256
rect 22774 9244 22784 9428
rect 22840 9244 22850 9428
rect 22884 9256 22890 9464
rect 22924 9256 22930 9464
rect 22980 9428 22986 9632
rect 23020 9428 23026 9632
rect 23062 9464 23072 9648
rect 23128 9464 23138 9648
rect 23172 9632 23218 9644
rect 22884 9244 22930 9256
rect 22966 9244 22976 9428
rect 23032 9244 23042 9428
rect 23076 9256 23082 9464
rect 23116 9256 23122 9464
rect 23172 9428 23178 9632
rect 23212 9428 23218 9632
rect 23254 9464 23264 9648
rect 23320 9464 23330 9648
rect 23364 9632 23410 9644
rect 23076 9244 23122 9256
rect 23158 9244 23168 9428
rect 23224 9244 23234 9428
rect 23268 9256 23274 9464
rect 23308 9256 23314 9464
rect 23364 9428 23370 9632
rect 23404 9428 23410 9632
rect 23446 9464 23456 9648
rect 23512 9464 23522 9648
rect 23556 9632 23602 9644
rect 23268 9244 23314 9256
rect 23350 9244 23360 9428
rect 23416 9244 23426 9428
rect 23460 9256 23466 9464
rect 23500 9256 23506 9464
rect 23556 9428 23562 9632
rect 23596 9428 23602 9632
rect 23638 9464 23648 9648
rect 23704 9464 23714 9648
rect 23748 9632 23794 9644
rect 23460 9244 23506 9256
rect 23542 9244 23552 9428
rect 23608 9244 23618 9428
rect 23652 9256 23658 9464
rect 23692 9256 23698 9464
rect 23748 9428 23754 9632
rect 23788 9428 23794 9632
rect 23830 9464 23840 9648
rect 23896 9464 23906 9648
rect 23940 9632 23986 9644
rect 23652 9244 23698 9256
rect 23734 9244 23744 9428
rect 23800 9244 23810 9428
rect 23844 9256 23850 9464
rect 23884 9256 23890 9464
rect 23940 9428 23946 9632
rect 23980 9428 23986 9632
rect 23844 9244 23890 9256
rect 23926 9244 23936 9428
rect 23992 9244 24002 9428
rect 21556 9208 23948 9212
rect 19556 9206 23948 9208
rect 19556 9200 22170 9206
rect 19556 9166 19574 9200
rect 19608 9166 19766 9200
rect 19800 9166 19958 9200
rect 19992 9166 20150 9200
rect 20184 9166 20342 9200
rect 20376 9166 20534 9200
rect 20568 9166 20726 9200
rect 20760 9166 20918 9200
rect 20952 9166 21110 9200
rect 21144 9166 21302 9200
rect 21336 9172 22170 9200
rect 22204 9172 22362 9206
rect 22396 9172 22554 9206
rect 22588 9172 22746 9206
rect 22780 9172 22938 9206
rect 22972 9172 23130 9206
rect 23164 9172 23322 9206
rect 23356 9172 23514 9206
rect 23548 9172 23706 9206
rect 23740 9172 23898 9206
rect 23932 9172 23948 9206
rect 21336 9166 23948 9172
rect 19556 9104 23948 9166
rect 21556 9098 23948 9104
rect 21556 9064 22170 9098
rect 22204 9064 22362 9098
rect 22396 9064 22554 9098
rect 22588 9064 22746 9098
rect 22780 9064 22938 9098
rect 22972 9064 23130 9098
rect 23164 9064 23322 9098
rect 23356 9064 23514 9098
rect 23548 9064 23706 9098
rect 23740 9064 23898 9098
rect 23932 9064 23948 9098
rect 21556 9056 23948 9064
rect 15932 8970 16136 8972
rect 15932 8968 16376 8970
rect 15920 8964 16376 8968
rect 16928 8964 17244 8970
rect 15920 8904 16072 8964
rect 16456 8904 16466 8964
rect 16928 8904 16940 8964
rect 17232 8904 17244 8964
rect 15920 8898 16376 8904
rect 16928 8898 17244 8904
rect 17864 8964 18180 8970
rect 17864 8904 17876 8964
rect 18168 8904 18180 8964
rect 17864 8898 18180 8904
rect 15920 8896 16136 8898
rect 15920 8704 16004 8896
rect 18978 8868 18988 8984
rect 16216 8802 18988 8868
rect 16216 8768 16234 8802
rect 16268 8768 16426 8802
rect 16460 8768 16618 8802
rect 16652 8768 16810 8802
rect 16844 8768 17002 8802
rect 17036 8768 17194 8802
rect 17228 8768 17386 8802
rect 17420 8768 17578 8802
rect 17612 8768 17770 8802
rect 17804 8768 17962 8802
rect 17996 8768 18988 8802
rect 16216 8760 18988 8768
rect 15920 8356 15940 8704
rect 15996 8356 16004 8704
rect 16084 8718 16130 8730
rect 16084 8508 16090 8718
rect 16124 8508 16130 8718
rect 16166 8552 16176 8732
rect 16228 8552 16238 8732
rect 16276 8718 16322 8730
rect 15920 8160 16004 8356
rect 16070 8328 16080 8508
rect 16132 8328 16142 8508
rect 16180 8342 16186 8552
rect 16220 8342 16226 8552
rect 16276 8508 16282 8718
rect 16316 8508 16322 8718
rect 16358 8552 16368 8732
rect 16420 8552 16430 8732
rect 16468 8718 16514 8730
rect 16180 8330 16226 8342
rect 16262 8328 16272 8508
rect 16324 8328 16334 8508
rect 16372 8342 16378 8552
rect 16412 8342 16418 8552
rect 16468 8508 16474 8718
rect 16508 8508 16514 8718
rect 16550 8552 16560 8732
rect 16612 8552 16622 8732
rect 16660 8718 16706 8730
rect 16372 8330 16418 8342
rect 16454 8328 16464 8508
rect 16516 8328 16526 8508
rect 16564 8342 16570 8552
rect 16604 8342 16610 8552
rect 16660 8508 16666 8718
rect 16700 8508 16706 8718
rect 16742 8552 16752 8732
rect 16804 8552 16814 8732
rect 16852 8718 16898 8730
rect 16564 8330 16610 8342
rect 16646 8328 16656 8508
rect 16708 8328 16718 8508
rect 16756 8342 16762 8552
rect 16796 8342 16802 8552
rect 16852 8508 16858 8718
rect 16892 8508 16898 8718
rect 16934 8552 16944 8732
rect 16996 8552 17006 8732
rect 17044 8718 17090 8730
rect 16756 8330 16802 8342
rect 16838 8328 16848 8508
rect 16900 8328 16910 8508
rect 16948 8342 16954 8552
rect 16988 8342 16994 8552
rect 17044 8508 17050 8718
rect 17084 8508 17090 8718
rect 17126 8552 17136 8732
rect 17188 8552 17198 8732
rect 17236 8718 17282 8730
rect 16948 8330 16994 8342
rect 17030 8328 17040 8508
rect 17092 8328 17102 8508
rect 17140 8342 17146 8552
rect 17180 8342 17186 8552
rect 17236 8508 17242 8718
rect 17276 8508 17282 8718
rect 17318 8552 17328 8732
rect 17380 8552 17390 8732
rect 17428 8718 17474 8730
rect 17140 8330 17186 8342
rect 17222 8328 17232 8508
rect 17284 8328 17294 8508
rect 17332 8342 17338 8552
rect 17372 8342 17378 8552
rect 17428 8508 17434 8718
rect 17468 8508 17474 8718
rect 17510 8552 17520 8732
rect 17572 8552 17582 8732
rect 17620 8718 17666 8730
rect 17332 8330 17378 8342
rect 17414 8328 17424 8508
rect 17476 8328 17486 8508
rect 17524 8342 17530 8552
rect 17564 8342 17570 8552
rect 17620 8508 17626 8718
rect 17660 8508 17666 8718
rect 17702 8552 17712 8732
rect 17764 8552 17774 8732
rect 17812 8718 17858 8730
rect 17524 8330 17570 8342
rect 17606 8328 17616 8508
rect 17668 8328 17678 8508
rect 17716 8342 17722 8552
rect 17756 8342 17762 8552
rect 17812 8508 17818 8718
rect 17852 8508 17858 8718
rect 17894 8552 17904 8732
rect 17956 8552 17966 8732
rect 18004 8718 18050 8730
rect 17716 8330 17762 8342
rect 17798 8328 17808 8508
rect 17860 8328 17870 8508
rect 17908 8342 17914 8552
rect 17948 8342 17954 8552
rect 18004 8508 18010 8718
rect 18044 8508 18050 8718
rect 18134 8672 18206 8684
rect 17908 8330 17954 8342
rect 17990 8328 18000 8508
rect 18052 8328 18062 8508
rect 18130 8416 18140 8672
rect 18200 8416 18210 8672
rect 18328 8432 18988 8760
rect 19408 8432 19418 8984
rect 21556 8980 21976 9056
rect 19552 8768 21696 8816
rect 19552 8734 19574 8768
rect 19608 8734 19766 8768
rect 19800 8734 19958 8768
rect 19992 8734 20150 8768
rect 20184 8734 20342 8768
rect 20376 8734 20534 8768
rect 20568 8734 20726 8768
rect 20760 8734 20918 8768
rect 20952 8734 21110 8768
rect 21144 8734 21302 8768
rect 21336 8734 21696 8768
rect 19552 8728 21696 8734
rect 19520 8684 19566 8696
rect 19520 8476 19526 8684
rect 19560 8476 19566 8684
rect 19602 8520 19612 8700
rect 19668 8520 19678 8700
rect 19712 8684 19758 8696
rect 18134 8404 18206 8416
rect 18328 8300 18612 8432
rect 16124 8292 18612 8300
rect 19506 8296 19516 8476
rect 19572 8296 19582 8476
rect 19616 8308 19622 8520
rect 19656 8308 19662 8520
rect 19712 8476 19718 8684
rect 19752 8476 19758 8684
rect 19794 8520 19804 8700
rect 19860 8520 19870 8700
rect 19904 8684 19950 8696
rect 19616 8296 19662 8308
rect 19698 8296 19708 8476
rect 19764 8296 19774 8476
rect 19808 8308 19814 8520
rect 19848 8308 19854 8520
rect 19904 8476 19910 8684
rect 19944 8476 19950 8684
rect 19986 8520 19996 8700
rect 20052 8520 20062 8700
rect 20096 8684 20142 8696
rect 19808 8296 19854 8308
rect 19890 8296 19900 8476
rect 19956 8296 19966 8476
rect 20000 8308 20006 8520
rect 20040 8308 20046 8520
rect 20096 8476 20102 8684
rect 20136 8476 20142 8684
rect 20178 8520 20188 8700
rect 20244 8520 20254 8700
rect 20288 8684 20334 8696
rect 20000 8296 20046 8308
rect 20082 8296 20092 8476
rect 20148 8296 20158 8476
rect 20192 8308 20198 8520
rect 20232 8308 20238 8520
rect 20288 8476 20294 8684
rect 20328 8476 20334 8684
rect 20370 8520 20380 8700
rect 20436 8520 20446 8700
rect 20480 8684 20526 8696
rect 20192 8296 20238 8308
rect 20274 8296 20284 8476
rect 20340 8296 20350 8476
rect 20384 8308 20390 8520
rect 20424 8308 20430 8520
rect 20480 8476 20486 8684
rect 20520 8476 20526 8684
rect 20562 8520 20572 8700
rect 20628 8520 20638 8700
rect 20672 8684 20718 8696
rect 20384 8296 20430 8308
rect 20466 8296 20476 8476
rect 20532 8296 20542 8476
rect 20576 8308 20582 8520
rect 20616 8308 20622 8520
rect 20672 8476 20678 8684
rect 20712 8476 20718 8684
rect 20754 8520 20764 8700
rect 20820 8520 20830 8700
rect 20864 8684 20910 8696
rect 20576 8296 20622 8308
rect 20658 8296 20668 8476
rect 20724 8296 20734 8476
rect 20768 8308 20774 8520
rect 20808 8308 20814 8520
rect 20864 8476 20870 8684
rect 20904 8476 20910 8684
rect 20946 8520 20956 8700
rect 21012 8520 21022 8700
rect 21056 8684 21102 8696
rect 20768 8296 20814 8308
rect 20850 8296 20860 8476
rect 20916 8296 20926 8476
rect 20960 8308 20966 8520
rect 21000 8308 21006 8520
rect 21056 8476 21062 8684
rect 21096 8476 21102 8684
rect 21138 8520 21148 8700
rect 21204 8520 21214 8700
rect 21248 8684 21294 8696
rect 20960 8296 21006 8308
rect 21042 8296 21052 8476
rect 21108 8296 21118 8476
rect 21152 8308 21158 8520
rect 21192 8308 21198 8520
rect 21248 8476 21254 8684
rect 21288 8476 21294 8684
rect 21330 8520 21340 8700
rect 21396 8520 21406 8700
rect 21440 8684 21486 8696
rect 21152 8296 21198 8308
rect 21234 8296 21244 8476
rect 21300 8296 21310 8476
rect 21344 8308 21350 8520
rect 21384 8308 21390 8520
rect 21440 8476 21446 8684
rect 21480 8476 21486 8684
rect 21344 8296 21390 8308
rect 21426 8296 21436 8476
rect 21492 8296 21500 8476
rect 16124 8258 16138 8292
rect 16172 8258 16330 8292
rect 16364 8258 16522 8292
rect 16556 8258 16714 8292
rect 16748 8258 16906 8292
rect 16940 8258 17098 8292
rect 17132 8258 17290 8292
rect 17324 8258 17482 8292
rect 17516 8258 17674 8292
rect 17708 8258 17866 8292
rect 17900 8258 18612 8292
rect 21528 8264 21696 8728
rect 16124 8192 18612 8258
rect 15920 8154 16152 8160
rect 15920 8152 16376 8154
rect 16928 8152 17272 8154
rect 15920 8148 16164 8152
rect 15920 8088 16072 8148
rect 16456 8088 16466 8152
rect 16928 8088 16940 8152
rect 17260 8088 17272 8152
rect 15920 8084 16376 8088
rect 15920 7856 16004 8084
rect 16060 8082 16376 8084
rect 16928 8082 17272 8088
rect 17864 8152 18180 8158
rect 17864 8092 17876 8152
rect 18168 8092 18180 8152
rect 17864 8086 18180 8092
rect 18328 8044 18612 8192
rect 19652 8258 21696 8264
rect 19652 8224 19670 8258
rect 19704 8224 19862 8258
rect 19896 8224 20054 8258
rect 20088 8224 20246 8258
rect 20280 8224 20438 8258
rect 20472 8224 20630 8258
rect 20664 8224 20822 8258
rect 20856 8224 21014 8258
rect 21048 8224 21206 8258
rect 21240 8224 21398 8258
rect 21432 8224 21696 8258
rect 19652 8150 21696 8224
rect 19652 8116 19670 8150
rect 19704 8116 19862 8150
rect 19896 8116 20054 8150
rect 20088 8116 20246 8150
rect 20280 8116 20438 8150
rect 20472 8116 20630 8150
rect 20664 8116 20822 8150
rect 20856 8116 21014 8150
rect 21048 8116 21206 8150
rect 21240 8116 21398 8150
rect 21432 8116 21696 8150
rect 19652 8108 21696 8116
rect 16220 7982 18612 8044
rect 16220 7948 16234 7982
rect 16268 7948 16426 7982
rect 16460 7948 16618 7982
rect 16652 7948 16810 7982
rect 16844 7948 17002 7982
rect 17036 7948 17194 7982
rect 17228 7948 17386 7982
rect 17420 7948 17578 7982
rect 17612 7948 17770 7982
rect 17804 7948 17962 7982
rect 17996 7948 18612 7982
rect 16220 7940 18612 7948
rect 16084 7898 16130 7910
rect 15920 7844 16006 7856
rect 15920 7588 15940 7844
rect 16000 7588 16006 7844
rect 16084 7688 16090 7898
rect 16124 7688 16130 7898
rect 16166 7732 16176 7912
rect 16228 7732 16238 7912
rect 16276 7898 16322 7910
rect 15920 7576 16006 7588
rect 15920 7336 16004 7576
rect 16070 7508 16080 7688
rect 16132 7508 16142 7688
rect 16180 7522 16186 7732
rect 16220 7522 16226 7732
rect 16276 7688 16282 7898
rect 16316 7688 16322 7898
rect 16358 7732 16368 7912
rect 16420 7732 16430 7912
rect 16468 7898 16514 7910
rect 16180 7510 16226 7522
rect 16262 7508 16272 7688
rect 16324 7508 16334 7688
rect 16372 7522 16378 7732
rect 16412 7522 16418 7732
rect 16468 7688 16474 7898
rect 16508 7688 16514 7898
rect 16550 7732 16560 7912
rect 16612 7732 16622 7912
rect 16660 7898 16706 7910
rect 16372 7510 16418 7522
rect 16454 7508 16464 7688
rect 16516 7508 16526 7688
rect 16564 7522 16570 7732
rect 16604 7522 16610 7732
rect 16660 7688 16666 7898
rect 16700 7688 16706 7898
rect 16742 7732 16752 7912
rect 16804 7732 16814 7912
rect 16852 7898 16898 7910
rect 16564 7510 16610 7522
rect 16646 7508 16656 7688
rect 16708 7508 16718 7688
rect 16756 7522 16762 7732
rect 16796 7522 16802 7732
rect 16852 7688 16858 7898
rect 16892 7688 16898 7898
rect 16934 7732 16944 7912
rect 16996 7732 17006 7912
rect 17044 7898 17090 7910
rect 16756 7510 16802 7522
rect 16838 7508 16848 7688
rect 16900 7508 16910 7688
rect 16948 7522 16954 7732
rect 16988 7522 16994 7732
rect 17044 7688 17050 7898
rect 17084 7688 17090 7898
rect 17126 7732 17136 7912
rect 17188 7732 17198 7912
rect 17236 7898 17282 7910
rect 16948 7510 16994 7522
rect 17030 7508 17040 7688
rect 17092 7508 17102 7688
rect 17140 7522 17146 7732
rect 17180 7522 17186 7732
rect 17236 7688 17242 7898
rect 17276 7688 17282 7898
rect 17318 7732 17328 7912
rect 17380 7732 17390 7912
rect 17428 7898 17474 7910
rect 17140 7510 17186 7522
rect 17222 7508 17232 7688
rect 17284 7508 17294 7688
rect 17332 7522 17338 7732
rect 17372 7522 17378 7732
rect 17428 7688 17434 7898
rect 17468 7688 17474 7898
rect 17510 7732 17520 7912
rect 17572 7732 17582 7912
rect 17620 7898 17666 7910
rect 17332 7510 17378 7522
rect 17414 7508 17424 7688
rect 17476 7508 17486 7688
rect 17524 7522 17530 7732
rect 17564 7522 17570 7732
rect 17620 7688 17626 7898
rect 17660 7688 17666 7898
rect 17702 7732 17712 7912
rect 17764 7732 17774 7912
rect 17812 7898 17858 7910
rect 17524 7510 17570 7522
rect 17606 7508 17616 7688
rect 17668 7508 17678 7688
rect 17716 7522 17722 7732
rect 17756 7522 17762 7732
rect 17812 7688 17818 7898
rect 17852 7688 17858 7898
rect 17894 7732 17904 7912
rect 17956 7732 17966 7912
rect 18004 7898 18050 7910
rect 17716 7510 17762 7522
rect 17798 7508 17808 7688
rect 17860 7508 17870 7688
rect 17908 7522 17914 7732
rect 17948 7522 17954 7732
rect 18004 7688 18010 7898
rect 18044 7688 18050 7898
rect 18134 7824 18206 7836
rect 17908 7510 17954 7522
rect 17990 7508 18000 7688
rect 18052 7508 18062 7688
rect 18130 7568 18140 7824
rect 18200 7568 18210 7824
rect 18134 7556 18206 7568
rect 18328 7480 18612 7940
rect 19520 8066 19566 8078
rect 19520 7856 19526 8066
rect 19560 7856 19566 8066
rect 19602 7900 19612 8080
rect 19668 7900 19678 8080
rect 19712 8066 19758 8078
rect 19506 7676 19516 7856
rect 19572 7676 19582 7856
rect 19616 7690 19622 7900
rect 19656 7690 19662 7900
rect 19712 7856 19718 8066
rect 19752 7856 19758 8066
rect 19794 7900 19804 8080
rect 19860 7900 19870 8080
rect 19904 8066 19950 8078
rect 19616 7678 19662 7690
rect 19698 7676 19708 7856
rect 19764 7676 19774 7856
rect 19808 7690 19814 7900
rect 19848 7690 19854 7900
rect 19904 7856 19910 8066
rect 19944 7856 19950 8066
rect 19986 7900 19996 8080
rect 20052 7900 20062 8080
rect 20096 8066 20142 8078
rect 19808 7678 19854 7690
rect 19890 7676 19900 7856
rect 19956 7676 19966 7856
rect 20000 7690 20006 7900
rect 20040 7690 20046 7900
rect 20096 7856 20102 8066
rect 20136 7856 20142 8066
rect 20178 7900 20188 8080
rect 20244 7900 20254 8080
rect 20288 8066 20334 8078
rect 20000 7678 20046 7690
rect 20082 7676 20092 7856
rect 20148 7676 20158 7856
rect 20192 7690 20198 7900
rect 20232 7690 20238 7900
rect 20288 7856 20294 8066
rect 20328 7856 20334 8066
rect 20370 7900 20380 8080
rect 20436 7900 20446 8080
rect 20480 8066 20526 8078
rect 20192 7678 20238 7690
rect 20274 7676 20284 7856
rect 20340 7676 20350 7856
rect 20384 7690 20390 7900
rect 20424 7690 20430 7900
rect 20480 7856 20486 8066
rect 20520 7856 20526 8066
rect 20562 7900 20572 8080
rect 20628 7900 20638 8080
rect 20672 8066 20718 8078
rect 20384 7678 20430 7690
rect 20466 7676 20476 7856
rect 20532 7676 20542 7856
rect 20576 7690 20582 7900
rect 20616 7690 20622 7900
rect 20672 7856 20678 8066
rect 20712 7856 20718 8066
rect 20754 7900 20764 8080
rect 20820 7900 20830 8080
rect 20864 8066 20910 8078
rect 20576 7678 20622 7690
rect 20658 7676 20668 7856
rect 20724 7676 20734 7856
rect 20768 7690 20774 7900
rect 20808 7690 20814 7900
rect 20864 7856 20870 8066
rect 20904 7856 20910 8066
rect 20946 7900 20956 8080
rect 21012 7900 21022 8080
rect 21056 8066 21102 8078
rect 20768 7678 20814 7690
rect 20850 7676 20860 7856
rect 20916 7676 20926 7856
rect 20960 7690 20966 7900
rect 21000 7690 21006 7900
rect 21056 7856 21062 8066
rect 21096 7856 21102 8066
rect 21138 7900 21148 8080
rect 21204 7900 21214 8080
rect 21248 8066 21294 8078
rect 20960 7678 21006 7690
rect 21042 7676 21052 7856
rect 21108 7676 21118 7856
rect 21152 7690 21158 7900
rect 21192 7690 21198 7900
rect 21248 7856 21254 8066
rect 21288 7856 21294 8066
rect 21330 7900 21340 8080
rect 21396 7900 21406 8080
rect 21440 8066 21486 8078
rect 21152 7678 21198 7690
rect 21234 7676 21244 7856
rect 21300 7676 21310 7856
rect 21344 7690 21350 7900
rect 21384 7690 21390 7900
rect 21440 7856 21446 8066
rect 21480 7856 21486 8066
rect 21344 7678 21390 7690
rect 21426 7676 21436 7856
rect 21492 7676 21500 7856
rect 21528 7648 21696 8108
rect 19556 7640 21696 7648
rect 19556 7606 19574 7640
rect 19608 7606 19766 7640
rect 19800 7606 19958 7640
rect 19992 7606 20150 7640
rect 20184 7606 20342 7640
rect 20376 7606 20534 7640
rect 20568 7606 20726 7640
rect 20760 7606 20918 7640
rect 20952 7606 21110 7640
rect 21144 7606 21302 7640
rect 21336 7606 21696 7640
rect 19556 7572 21696 7606
rect 19792 7552 21696 7572
rect 16120 7472 18612 7480
rect 16120 7438 16138 7472
rect 16172 7438 16330 7472
rect 16364 7438 16522 7472
rect 16556 7438 16714 7472
rect 16748 7438 16906 7472
rect 16940 7438 17098 7472
rect 17132 7438 17290 7472
rect 17324 7438 17482 7472
rect 17516 7438 17674 7472
rect 17708 7438 17866 7472
rect 17900 7438 18612 7472
rect 16120 7372 18612 7438
rect 20772 7512 20968 7552
rect 21320 7512 21696 7552
rect 20772 7384 20784 7512
rect 15920 7328 16468 7336
rect 16928 7328 17244 7334
rect 15920 7268 16072 7328
rect 16456 7268 16468 7328
rect 16926 7268 16936 7328
rect 17232 7268 17244 7328
rect 15920 7260 16468 7268
rect 16928 7262 17244 7268
rect 17864 7328 18180 7334
rect 17864 7268 17876 7328
rect 18168 7268 18180 7328
rect 17864 7262 18180 7268
rect 15920 7004 16004 7260
rect 18328 7228 18612 7372
rect 16216 7162 18612 7228
rect 16216 7128 16234 7162
rect 16268 7128 16426 7162
rect 16460 7128 16618 7162
rect 16652 7128 16810 7162
rect 16844 7128 17002 7162
rect 17036 7128 17194 7162
rect 17228 7128 17386 7162
rect 17420 7128 17578 7162
rect 17612 7128 17770 7162
rect 17804 7128 17962 7162
rect 17996 7128 18612 7162
rect 16216 7120 18612 7128
rect 15920 6748 15936 7004
rect 15996 6748 16004 7004
rect 16084 7078 16130 7090
rect 16084 6868 16090 7078
rect 16124 6868 16130 7078
rect 16166 6912 16176 7092
rect 16228 6912 16238 7092
rect 16276 7078 16322 7090
rect 15920 6520 16004 6748
rect 16070 6688 16080 6868
rect 16132 6688 16142 6868
rect 16180 6702 16186 6912
rect 16220 6702 16226 6912
rect 16276 6868 16282 7078
rect 16316 6868 16322 7078
rect 16358 6912 16368 7092
rect 16420 6912 16430 7092
rect 16468 7078 16514 7090
rect 16180 6690 16226 6702
rect 16262 6688 16272 6868
rect 16324 6688 16334 6868
rect 16372 6702 16378 6912
rect 16412 6702 16418 6912
rect 16468 6868 16474 7078
rect 16508 6868 16514 7078
rect 16550 6912 16560 7092
rect 16612 6912 16622 7092
rect 16660 7078 16706 7090
rect 16372 6690 16418 6702
rect 16454 6688 16464 6868
rect 16516 6688 16526 6868
rect 16564 6702 16570 6912
rect 16604 6702 16610 6912
rect 16660 6868 16666 7078
rect 16700 6868 16706 7078
rect 16742 6912 16752 7092
rect 16804 6912 16814 7092
rect 16852 7078 16898 7090
rect 16564 6690 16610 6702
rect 16646 6688 16656 6868
rect 16708 6688 16718 6868
rect 16756 6702 16762 6912
rect 16796 6702 16802 6912
rect 16852 6868 16858 7078
rect 16892 6868 16898 7078
rect 16934 6912 16944 7092
rect 16996 6912 17006 7092
rect 17044 7078 17090 7090
rect 16756 6690 16802 6702
rect 16838 6688 16848 6868
rect 16900 6688 16910 6868
rect 16948 6702 16954 6912
rect 16988 6702 16994 6912
rect 17044 6868 17050 7078
rect 17084 6868 17090 7078
rect 17126 6912 17136 7092
rect 17188 6912 17198 7092
rect 17236 7078 17282 7090
rect 16948 6690 16994 6702
rect 17030 6688 17040 6868
rect 17092 6688 17102 6868
rect 17140 6702 17146 6912
rect 17180 6702 17186 6912
rect 17236 6868 17242 7078
rect 17276 6868 17282 7078
rect 17318 6912 17328 7092
rect 17380 6912 17390 7092
rect 17428 7078 17474 7090
rect 17140 6690 17186 6702
rect 17222 6688 17232 6868
rect 17284 6688 17294 6868
rect 17332 6702 17338 6912
rect 17372 6702 17378 6912
rect 17428 6868 17434 7078
rect 17468 6868 17474 7078
rect 17510 6912 17520 7092
rect 17572 6912 17582 7092
rect 17620 7078 17666 7090
rect 17332 6690 17378 6702
rect 17414 6688 17424 6868
rect 17476 6688 17486 6868
rect 17524 6702 17530 6912
rect 17564 6702 17570 6912
rect 17620 6868 17626 7078
rect 17660 6868 17666 7078
rect 17702 6912 17712 7092
rect 17764 6912 17774 7092
rect 17812 7078 17858 7090
rect 17524 6690 17570 6702
rect 17606 6688 17616 6868
rect 17668 6688 17678 6868
rect 17716 6702 17722 6912
rect 17756 6702 17762 6912
rect 17812 6868 17818 7078
rect 17852 6868 17858 7078
rect 17894 6912 17904 7092
rect 17956 6912 17966 7092
rect 18004 7078 18050 7090
rect 17716 6690 17762 6702
rect 17798 6688 17808 6868
rect 17860 6688 17870 6868
rect 17908 6702 17914 6912
rect 17948 6702 17954 6912
rect 18004 6868 18010 7078
rect 18044 6868 18050 7078
rect 18134 7012 18206 7024
rect 17908 6690 17954 6702
rect 17990 6688 18000 6868
rect 18052 6688 18062 6868
rect 18130 6756 18140 7012
rect 18200 6756 18210 7012
rect 18134 6744 18206 6756
rect 18328 6660 18612 7120
rect 20774 7000 20784 7384
rect 21476 7392 21696 7512
rect 21724 8596 21976 8980
rect 22020 9014 22066 9026
rect 22020 8808 22026 9014
rect 22060 8808 22066 9014
rect 22102 8844 22112 9028
rect 22168 8844 22178 9028
rect 22212 9014 22258 9026
rect 22006 8624 22016 8808
rect 22072 8624 22082 8808
rect 22116 8638 22122 8844
rect 22156 8638 22162 8844
rect 22212 8808 22218 9014
rect 22252 8808 22258 9014
rect 22294 8844 22304 9028
rect 22360 8844 22370 9028
rect 22404 9014 22450 9026
rect 22116 8626 22162 8638
rect 22198 8624 22208 8808
rect 22264 8624 22274 8808
rect 22308 8638 22314 8844
rect 22348 8638 22354 8844
rect 22404 8808 22410 9014
rect 22444 8808 22450 9014
rect 22486 8844 22496 9028
rect 22552 8844 22562 9028
rect 22596 9014 22642 9026
rect 22308 8626 22354 8638
rect 22390 8624 22400 8808
rect 22456 8624 22466 8808
rect 22500 8638 22506 8844
rect 22540 8638 22546 8844
rect 22596 8808 22602 9014
rect 22636 8808 22642 9014
rect 22678 8844 22688 9028
rect 22744 8844 22754 9028
rect 22788 9014 22834 9026
rect 22500 8626 22546 8638
rect 22582 8624 22592 8808
rect 22648 8624 22658 8808
rect 22692 8638 22698 8844
rect 22732 8638 22738 8844
rect 22788 8808 22794 9014
rect 22828 8808 22834 9014
rect 22870 8844 22880 9028
rect 22936 8844 22946 9028
rect 22980 9014 23026 9026
rect 22692 8626 22738 8638
rect 22774 8624 22784 8808
rect 22840 8624 22850 8808
rect 22884 8638 22890 8844
rect 22924 8638 22930 8844
rect 22980 8808 22986 9014
rect 23020 8808 23026 9014
rect 23062 8844 23072 9028
rect 23128 8844 23138 9028
rect 23172 9014 23218 9026
rect 22884 8626 22930 8638
rect 22966 8624 22976 8808
rect 23032 8624 23042 8808
rect 23076 8638 23082 8844
rect 23116 8638 23122 8844
rect 23172 8808 23178 9014
rect 23212 8808 23218 9014
rect 23254 8844 23264 9028
rect 23320 8844 23330 9028
rect 23364 9014 23410 9026
rect 23076 8626 23122 8638
rect 23158 8624 23168 8808
rect 23224 8624 23234 8808
rect 23268 8638 23274 8844
rect 23308 8638 23314 8844
rect 23364 8808 23370 9014
rect 23404 8808 23410 9014
rect 23446 8844 23456 9028
rect 23512 8844 23522 9028
rect 23556 9014 23602 9026
rect 23268 8626 23314 8638
rect 23350 8624 23360 8808
rect 23416 8624 23426 8808
rect 23460 8638 23466 8844
rect 23500 8638 23506 8844
rect 23556 8808 23562 9014
rect 23596 8808 23602 9014
rect 23638 8844 23648 9028
rect 23704 8844 23714 9028
rect 23748 9014 23794 9026
rect 23460 8626 23506 8638
rect 23542 8624 23552 8808
rect 23608 8624 23618 8808
rect 23652 8638 23658 8844
rect 23692 8638 23698 8844
rect 23748 8808 23754 9014
rect 23788 8808 23794 9014
rect 23830 8844 23840 9028
rect 23896 8844 23906 9028
rect 23940 9014 23986 9026
rect 23652 8626 23698 8638
rect 23734 8624 23744 8808
rect 23800 8624 23810 8808
rect 23844 8638 23850 8844
rect 23884 8638 23890 8844
rect 23940 8808 23946 9014
rect 23980 8808 23986 9014
rect 23844 8626 23890 8638
rect 23926 8624 23936 8808
rect 23992 8624 24002 8808
rect 21724 8588 23852 8596
rect 21724 8554 22074 8588
rect 22108 8554 22266 8588
rect 22300 8554 22458 8588
rect 22492 8554 22650 8588
rect 22684 8554 22842 8588
rect 22876 8554 23034 8588
rect 23068 8554 23226 8588
rect 23260 8554 23418 8588
rect 23452 8554 23610 8588
rect 23644 8554 23802 8588
rect 23836 8554 23852 8588
rect 21724 8480 23852 8554
rect 21724 8446 22074 8480
rect 22108 8446 22266 8480
rect 22300 8446 22458 8480
rect 22492 8446 22650 8480
rect 22684 8446 22842 8480
rect 22876 8446 23034 8480
rect 23068 8446 23226 8480
rect 23260 8446 23418 8480
rect 23452 8446 23610 8480
rect 23644 8446 23802 8480
rect 23836 8446 23852 8480
rect 21724 8440 23852 8446
rect 21724 7976 21976 8440
rect 22020 8396 22066 8408
rect 22020 8192 22026 8396
rect 22060 8192 22066 8396
rect 22102 8228 22112 8412
rect 22168 8228 22178 8412
rect 22212 8396 22258 8408
rect 22006 8008 22016 8192
rect 22072 8008 22082 8192
rect 22116 8020 22122 8228
rect 22156 8020 22162 8228
rect 22212 8192 22218 8396
rect 22252 8192 22258 8396
rect 22294 8228 22304 8412
rect 22360 8228 22370 8412
rect 22404 8396 22450 8408
rect 22116 8008 22162 8020
rect 22198 8008 22208 8192
rect 22264 8008 22274 8192
rect 22308 8020 22314 8228
rect 22348 8020 22354 8228
rect 22404 8192 22410 8396
rect 22444 8192 22450 8396
rect 22486 8228 22496 8412
rect 22552 8228 22562 8412
rect 22596 8396 22642 8408
rect 22308 8008 22354 8020
rect 22390 8008 22400 8192
rect 22456 8008 22466 8192
rect 22500 8020 22506 8228
rect 22540 8020 22546 8228
rect 22596 8192 22602 8396
rect 22636 8192 22642 8396
rect 22678 8228 22688 8412
rect 22744 8228 22754 8412
rect 22788 8396 22834 8408
rect 22500 8008 22546 8020
rect 22582 8008 22592 8192
rect 22648 8008 22658 8192
rect 22692 8020 22698 8228
rect 22732 8020 22738 8228
rect 22788 8192 22794 8396
rect 22828 8192 22834 8396
rect 22870 8228 22880 8412
rect 22936 8228 22946 8412
rect 22980 8396 23026 8408
rect 22692 8008 22738 8020
rect 22774 8008 22784 8192
rect 22840 8008 22850 8192
rect 22884 8020 22890 8228
rect 22924 8020 22930 8228
rect 22980 8192 22986 8396
rect 23020 8192 23026 8396
rect 23062 8228 23072 8412
rect 23128 8228 23138 8412
rect 23172 8396 23218 8408
rect 22884 8008 22930 8020
rect 22966 8008 22976 8192
rect 23032 8008 23042 8192
rect 23076 8020 23082 8228
rect 23116 8020 23122 8228
rect 23172 8192 23178 8396
rect 23212 8192 23218 8396
rect 23254 8228 23264 8412
rect 23320 8228 23330 8412
rect 23364 8396 23410 8408
rect 23076 8008 23122 8020
rect 23158 8008 23168 8192
rect 23224 8008 23234 8192
rect 23268 8020 23274 8228
rect 23308 8020 23314 8228
rect 23364 8192 23370 8396
rect 23404 8192 23410 8396
rect 23446 8228 23456 8412
rect 23512 8228 23522 8412
rect 23556 8396 23602 8408
rect 23268 8008 23314 8020
rect 23350 8008 23360 8192
rect 23416 8008 23426 8192
rect 23460 8020 23466 8228
rect 23500 8020 23506 8228
rect 23556 8192 23562 8396
rect 23596 8192 23602 8396
rect 23638 8228 23648 8412
rect 23704 8228 23714 8412
rect 23748 8396 23794 8408
rect 23460 8008 23506 8020
rect 23542 8008 23552 8192
rect 23608 8008 23618 8192
rect 23652 8020 23658 8228
rect 23692 8020 23698 8228
rect 23748 8192 23754 8396
rect 23788 8192 23794 8396
rect 23830 8228 23840 8412
rect 23896 8228 23906 8412
rect 23940 8396 23986 8408
rect 23652 8008 23698 8020
rect 23734 8008 23744 8192
rect 23800 8008 23810 8192
rect 23844 8020 23850 8228
rect 23884 8020 23890 8228
rect 23940 8192 23946 8396
rect 23980 8192 23986 8396
rect 23844 8008 23890 8020
rect 23926 8008 23936 8192
rect 23992 8008 24002 8192
rect 21724 7970 23948 7976
rect 21724 7936 22170 7970
rect 22204 7936 22362 7970
rect 22396 7936 22554 7970
rect 22588 7936 22746 7970
rect 22780 7936 22938 7970
rect 22972 7936 23130 7970
rect 23164 7936 23322 7970
rect 23356 7936 23514 7970
rect 23548 7936 23706 7970
rect 23740 7936 23898 7970
rect 23932 7936 23948 7970
rect 21724 7862 23948 7936
rect 21724 7828 22170 7862
rect 22204 7828 22362 7862
rect 22396 7828 22554 7862
rect 22588 7828 22746 7862
rect 22780 7828 22938 7862
rect 22972 7828 23130 7862
rect 23164 7828 23322 7862
rect 23356 7828 23514 7862
rect 23548 7828 23706 7862
rect 23740 7828 23898 7862
rect 23932 7828 23948 7862
rect 21724 7820 23948 7828
rect 21476 7000 21486 7392
rect 21724 7360 21976 7820
rect 22020 7778 22066 7790
rect 22020 7572 22026 7778
rect 22060 7572 22066 7778
rect 22102 7608 22112 7792
rect 22168 7608 22178 7792
rect 22212 7778 22258 7790
rect 22006 7388 22016 7572
rect 22072 7388 22082 7572
rect 22116 7402 22122 7608
rect 22156 7402 22162 7608
rect 22212 7572 22218 7778
rect 22252 7572 22258 7778
rect 22294 7608 22304 7792
rect 22360 7608 22370 7792
rect 22404 7778 22450 7790
rect 22116 7390 22162 7402
rect 22198 7388 22208 7572
rect 22264 7388 22274 7572
rect 22308 7402 22314 7608
rect 22348 7402 22354 7608
rect 22404 7572 22410 7778
rect 22444 7572 22450 7778
rect 22486 7608 22496 7792
rect 22552 7608 22562 7792
rect 22596 7778 22642 7790
rect 22308 7390 22354 7402
rect 22390 7388 22400 7572
rect 22456 7388 22466 7572
rect 22500 7402 22506 7608
rect 22540 7402 22546 7608
rect 22596 7572 22602 7778
rect 22636 7572 22642 7778
rect 22678 7608 22688 7792
rect 22744 7608 22754 7792
rect 22788 7778 22834 7790
rect 22500 7390 22546 7402
rect 22582 7388 22592 7572
rect 22648 7388 22658 7572
rect 22692 7402 22698 7608
rect 22732 7402 22738 7608
rect 22788 7572 22794 7778
rect 22828 7572 22834 7778
rect 22870 7608 22880 7792
rect 22936 7608 22946 7792
rect 22980 7778 23026 7790
rect 22692 7390 22738 7402
rect 22774 7388 22784 7572
rect 22840 7388 22850 7572
rect 22884 7402 22890 7608
rect 22924 7402 22930 7608
rect 22980 7572 22986 7778
rect 23020 7572 23026 7778
rect 23062 7608 23072 7792
rect 23128 7608 23138 7792
rect 23172 7778 23218 7790
rect 22884 7390 22930 7402
rect 22966 7388 22976 7572
rect 23032 7388 23042 7572
rect 23076 7402 23082 7608
rect 23116 7402 23122 7608
rect 23172 7572 23178 7778
rect 23212 7572 23218 7778
rect 23254 7608 23264 7792
rect 23320 7608 23330 7792
rect 23364 7778 23410 7790
rect 23076 7390 23122 7402
rect 23158 7388 23168 7572
rect 23224 7388 23234 7572
rect 23268 7402 23274 7608
rect 23308 7402 23314 7608
rect 23364 7572 23370 7778
rect 23404 7572 23410 7778
rect 23446 7608 23456 7792
rect 23512 7608 23522 7792
rect 23556 7778 23602 7790
rect 23268 7390 23314 7402
rect 23350 7388 23360 7572
rect 23416 7388 23426 7572
rect 23460 7402 23466 7608
rect 23500 7402 23506 7608
rect 23556 7572 23562 7778
rect 23596 7572 23602 7778
rect 23638 7608 23648 7792
rect 23704 7608 23714 7792
rect 23748 7778 23794 7790
rect 23460 7390 23506 7402
rect 23542 7388 23552 7572
rect 23608 7388 23618 7572
rect 23652 7402 23658 7608
rect 23692 7402 23698 7608
rect 23748 7572 23754 7778
rect 23788 7572 23794 7778
rect 23830 7608 23840 7792
rect 23896 7608 23906 7792
rect 23940 7778 23986 7790
rect 23652 7390 23698 7402
rect 23734 7388 23744 7572
rect 23800 7388 23810 7572
rect 23844 7402 23850 7608
rect 23884 7402 23890 7608
rect 23940 7572 23946 7778
rect 23980 7572 23986 7778
rect 23844 7390 23890 7402
rect 23926 7388 23936 7572
rect 23992 7388 24002 7572
rect 21556 7352 23852 7360
rect 21556 7318 22074 7352
rect 22108 7318 22266 7352
rect 22300 7318 22458 7352
rect 22492 7318 22650 7352
rect 22684 7318 22842 7352
rect 22876 7318 23034 7352
rect 23068 7318 23226 7352
rect 23260 7318 23418 7352
rect 23452 7318 23610 7352
rect 23644 7318 23802 7352
rect 23836 7318 23852 7352
rect 21556 7244 23852 7318
rect 21556 7210 22074 7244
rect 22108 7210 22266 7244
rect 22300 7210 22458 7244
rect 22492 7210 22650 7244
rect 22684 7210 22842 7244
rect 22876 7210 23034 7244
rect 23068 7210 23226 7244
rect 23260 7210 23418 7244
rect 23452 7210 23610 7244
rect 23644 7210 23802 7244
rect 23836 7210 23852 7244
rect 21556 7204 23852 7210
rect 21556 6928 21976 7204
rect 22020 7160 22066 7172
rect 22020 6956 22026 7160
rect 22060 6956 22066 7160
rect 22102 6992 22112 7176
rect 22168 6992 22178 7176
rect 22212 7160 22258 7172
rect 16124 6652 18612 6660
rect 16124 6618 16138 6652
rect 16172 6618 16330 6652
rect 16364 6618 16522 6652
rect 16556 6618 16714 6652
rect 16748 6618 16906 6652
rect 16940 6618 17098 6652
rect 17132 6618 17290 6652
rect 17324 6618 17482 6652
rect 17516 6618 17674 6652
rect 17708 6618 17866 6652
rect 17900 6618 18612 6652
rect 16124 6552 18612 6618
rect 21390 6600 21400 6928
rect 21928 6740 21976 6928
rect 22006 6772 22016 6956
rect 22072 6772 22082 6956
rect 22116 6784 22122 6992
rect 22156 6784 22162 6992
rect 22212 6956 22218 7160
rect 22252 6956 22258 7160
rect 22294 6992 22304 7176
rect 22360 6992 22370 7176
rect 22404 7160 22450 7172
rect 22116 6772 22162 6784
rect 22198 6772 22208 6956
rect 22264 6772 22274 6956
rect 22308 6784 22314 6992
rect 22348 6784 22354 6992
rect 22404 6956 22410 7160
rect 22444 6956 22450 7160
rect 22486 6992 22496 7176
rect 22552 6992 22562 7176
rect 22596 7160 22642 7172
rect 22308 6772 22354 6784
rect 22390 6772 22400 6956
rect 22456 6772 22466 6956
rect 22500 6784 22506 6992
rect 22540 6784 22546 6992
rect 22596 6956 22602 7160
rect 22636 6956 22642 7160
rect 22678 6992 22688 7176
rect 22744 6992 22754 7176
rect 22788 7160 22834 7172
rect 22500 6772 22546 6784
rect 22582 6772 22592 6956
rect 22648 6772 22658 6956
rect 22692 6784 22698 6992
rect 22732 6784 22738 6992
rect 22788 6956 22794 7160
rect 22828 6956 22834 7160
rect 22870 6992 22880 7176
rect 22936 6992 22946 7176
rect 22980 7160 23026 7172
rect 22692 6772 22738 6784
rect 22774 6772 22784 6956
rect 22840 6772 22850 6956
rect 22884 6784 22890 6992
rect 22924 6784 22930 6992
rect 22980 6956 22986 7160
rect 23020 6956 23026 7160
rect 23062 6992 23072 7176
rect 23128 6992 23138 7176
rect 23172 7160 23218 7172
rect 22884 6772 22930 6784
rect 22966 6772 22976 6956
rect 23032 6772 23042 6956
rect 23076 6784 23082 6992
rect 23116 6784 23122 6992
rect 23172 6956 23178 7160
rect 23212 6956 23218 7160
rect 23254 6992 23264 7176
rect 23320 6992 23330 7176
rect 23364 7160 23410 7172
rect 23076 6772 23122 6784
rect 23158 6772 23168 6956
rect 23224 6772 23234 6956
rect 23268 6784 23274 6992
rect 23308 6784 23314 6992
rect 23364 6956 23370 7160
rect 23404 6956 23410 7160
rect 23446 6992 23456 7176
rect 23512 6992 23522 7176
rect 23556 7160 23602 7172
rect 23268 6772 23314 6784
rect 23350 6772 23360 6956
rect 23416 6772 23426 6956
rect 23460 6784 23466 6992
rect 23500 6784 23506 6992
rect 23556 6956 23562 7160
rect 23596 6956 23602 7160
rect 23638 6992 23648 7176
rect 23704 6992 23714 7176
rect 23748 7160 23794 7172
rect 23460 6772 23506 6784
rect 23542 6772 23552 6956
rect 23608 6772 23618 6956
rect 23652 6784 23658 6992
rect 23692 6784 23698 6992
rect 23748 6956 23754 7160
rect 23788 6956 23794 7160
rect 23830 6992 23840 7176
rect 23896 6992 23906 7176
rect 23940 7160 23986 7172
rect 23652 6772 23698 6784
rect 23734 6772 23744 6956
rect 23800 6772 23810 6956
rect 23844 6784 23850 6992
rect 23884 6784 23890 6992
rect 23940 6956 23946 7160
rect 23980 6956 23986 7160
rect 23844 6772 23890 6784
rect 23926 6772 23936 6956
rect 23992 6772 24002 6956
rect 21928 6734 23948 6740
rect 21928 6700 22170 6734
rect 22204 6700 22362 6734
rect 22396 6700 22554 6734
rect 22588 6700 22746 6734
rect 22780 6700 22938 6734
rect 22972 6700 23130 6734
rect 23164 6700 23322 6734
rect 23356 6700 23514 6734
rect 23548 6700 23706 6734
rect 23740 6700 23898 6734
rect 23932 6700 23948 6734
rect 21928 6626 23948 6700
rect 21928 6600 22170 6626
rect 21556 6592 22170 6600
rect 22204 6592 22362 6626
rect 22396 6592 22554 6626
rect 22588 6592 22746 6626
rect 22780 6592 22938 6626
rect 22972 6592 23130 6626
rect 23164 6592 23322 6626
rect 23356 6592 23514 6626
rect 23548 6592 23706 6626
rect 23740 6592 23898 6626
rect 23932 6592 23948 6626
rect 21556 6584 23948 6592
rect 16060 6520 16376 6522
rect 15920 6516 16376 6520
rect 15920 6456 16072 6516
rect 16364 6456 16376 6516
rect 15920 6448 16376 6456
rect 16928 6516 17244 6522
rect 16928 6456 16940 6516
rect 17232 6456 17244 6516
rect 16928 6450 17244 6456
rect 17864 6512 18180 6518
rect 17864 6452 17876 6512
rect 18168 6452 18180 6512
rect 21556 6472 21976 6584
rect 17864 6446 18180 6452
rect 21350 6156 21360 6472
rect 21856 6156 21976 6472
rect 22020 6542 22066 6554
rect 22020 6336 22026 6542
rect 22060 6336 22066 6542
rect 22102 6372 22112 6556
rect 22168 6372 22178 6556
rect 22212 6542 22258 6554
rect 21556 6124 21976 6156
rect 22006 6152 22016 6336
rect 22072 6152 22082 6336
rect 22116 6166 22122 6372
rect 22156 6166 22162 6372
rect 22212 6336 22218 6542
rect 22252 6336 22258 6542
rect 22294 6372 22304 6556
rect 22360 6372 22370 6556
rect 22404 6542 22450 6554
rect 22116 6154 22162 6166
rect 22198 6152 22208 6336
rect 22264 6152 22274 6336
rect 22308 6166 22314 6372
rect 22348 6166 22354 6372
rect 22404 6336 22410 6542
rect 22444 6336 22450 6542
rect 22486 6372 22496 6556
rect 22552 6372 22562 6556
rect 22596 6542 22642 6554
rect 22308 6154 22354 6166
rect 22390 6152 22400 6336
rect 22456 6152 22466 6336
rect 22500 6166 22506 6372
rect 22540 6166 22546 6372
rect 22596 6336 22602 6542
rect 22636 6336 22642 6542
rect 22678 6372 22688 6556
rect 22744 6372 22754 6556
rect 22788 6542 22834 6554
rect 22500 6154 22546 6166
rect 22582 6152 22592 6336
rect 22648 6152 22658 6336
rect 22692 6166 22698 6372
rect 22732 6166 22738 6372
rect 22788 6336 22794 6542
rect 22828 6336 22834 6542
rect 22870 6372 22880 6556
rect 22936 6372 22946 6556
rect 22980 6542 23026 6554
rect 22692 6154 22738 6166
rect 22774 6152 22784 6336
rect 22840 6152 22850 6336
rect 22884 6166 22890 6372
rect 22924 6166 22930 6372
rect 22980 6336 22986 6542
rect 23020 6336 23026 6542
rect 23062 6372 23072 6556
rect 23128 6372 23138 6556
rect 23172 6542 23218 6554
rect 22884 6154 22930 6166
rect 22966 6152 22976 6336
rect 23032 6152 23042 6336
rect 23076 6166 23082 6372
rect 23116 6166 23122 6372
rect 23172 6336 23178 6542
rect 23212 6336 23218 6542
rect 23254 6372 23264 6556
rect 23320 6372 23330 6556
rect 23364 6542 23410 6554
rect 23076 6154 23122 6166
rect 23158 6152 23168 6336
rect 23224 6152 23234 6336
rect 23268 6166 23274 6372
rect 23308 6166 23314 6372
rect 23364 6336 23370 6542
rect 23404 6336 23410 6542
rect 23446 6372 23456 6556
rect 23512 6372 23522 6556
rect 23556 6542 23602 6554
rect 23268 6154 23314 6166
rect 23350 6152 23360 6336
rect 23416 6152 23426 6336
rect 23460 6166 23466 6372
rect 23500 6166 23506 6372
rect 23556 6336 23562 6542
rect 23596 6336 23602 6542
rect 23638 6372 23648 6556
rect 23704 6372 23714 6556
rect 23748 6542 23794 6554
rect 23460 6154 23506 6166
rect 23542 6152 23552 6336
rect 23608 6152 23618 6336
rect 23652 6166 23658 6372
rect 23692 6166 23698 6372
rect 23748 6336 23754 6542
rect 23788 6336 23794 6542
rect 23830 6372 23840 6556
rect 23896 6372 23906 6556
rect 23940 6542 23986 6554
rect 23652 6154 23698 6166
rect 23734 6152 23744 6336
rect 23800 6152 23810 6336
rect 23844 6166 23850 6372
rect 23884 6166 23890 6372
rect 23940 6336 23946 6542
rect 23980 6336 23986 6542
rect 23844 6154 23890 6166
rect 23926 6152 23936 6336
rect 23992 6152 24002 6336
rect 21556 6116 23852 6124
rect 21556 6082 22074 6116
rect 22108 6082 22266 6116
rect 22300 6082 22458 6116
rect 22492 6082 22650 6116
rect 22684 6082 22842 6116
rect 22876 6082 23034 6116
rect 23068 6082 23226 6116
rect 23260 6082 23418 6116
rect 23452 6082 23610 6116
rect 23644 6082 23802 6116
rect 23836 6082 23852 6116
rect 21556 6080 23852 6082
rect 14004 5988 21064 6052
rect 14004 5984 21168 5988
rect 14004 5946 21304 5984
rect 14004 5912 14770 5946
rect 14804 5912 14962 5946
rect 14996 5912 15154 5946
rect 15188 5912 15346 5946
rect 15380 5912 15538 5946
rect 15572 5912 16570 5946
rect 16604 5912 16762 5946
rect 16796 5912 16954 5946
rect 16988 5912 17146 5946
rect 17180 5912 17338 5946
rect 17372 5912 18370 5946
rect 18404 5912 18562 5946
rect 18596 5912 18754 5946
rect 18788 5912 18946 5946
rect 18980 5912 19138 5946
rect 19172 5912 20170 5946
rect 20204 5912 20362 5946
rect 20396 5912 20554 5946
rect 20588 5912 20746 5946
rect 20780 5912 20938 5946
rect 20972 5912 21304 5946
rect 14004 5908 21304 5912
rect 14004 5436 14484 5908
rect 14758 5906 14816 5908
rect 14950 5906 15008 5908
rect 15142 5906 15200 5908
rect 15334 5906 15392 5908
rect 15526 5906 15584 5908
rect 14620 5862 14666 5874
rect 14620 5652 14626 5862
rect 14660 5652 14666 5862
rect 14702 5696 14712 5876
rect 14764 5696 14774 5876
rect 14812 5862 14858 5874
rect 14606 5472 14616 5652
rect 14668 5472 14678 5652
rect 14716 5486 14722 5696
rect 14756 5486 14762 5696
rect 14812 5652 14818 5862
rect 14852 5652 14858 5862
rect 14894 5696 14904 5876
rect 14956 5696 14966 5876
rect 15004 5862 15050 5874
rect 14716 5474 14762 5486
rect 14798 5472 14808 5652
rect 14860 5472 14870 5652
rect 14908 5486 14914 5696
rect 14948 5486 14954 5696
rect 15004 5652 15010 5862
rect 15044 5652 15050 5862
rect 15086 5696 15096 5876
rect 15148 5696 15158 5876
rect 15196 5862 15242 5874
rect 14908 5474 14954 5486
rect 14990 5472 15000 5652
rect 15052 5472 15062 5652
rect 15100 5486 15106 5696
rect 15140 5486 15146 5696
rect 15196 5652 15202 5862
rect 15236 5652 15242 5862
rect 15278 5696 15288 5876
rect 15340 5696 15350 5876
rect 15388 5862 15434 5874
rect 15100 5474 15146 5486
rect 15182 5472 15192 5652
rect 15244 5472 15254 5652
rect 15292 5486 15298 5696
rect 15332 5486 15338 5696
rect 15388 5652 15394 5862
rect 15428 5652 15434 5862
rect 15470 5696 15480 5876
rect 15532 5696 15542 5876
rect 15580 5862 15626 5874
rect 15292 5474 15338 5486
rect 15374 5472 15384 5652
rect 15436 5472 15446 5652
rect 15484 5486 15490 5696
rect 15524 5486 15530 5696
rect 15580 5652 15586 5862
rect 15620 5652 15626 5862
rect 15484 5474 15530 5486
rect 15566 5472 15576 5652
rect 15628 5472 15638 5652
rect 14662 5436 14720 5442
rect 14854 5436 14912 5442
rect 15046 5436 15104 5442
rect 15238 5436 15296 5442
rect 15430 5436 15488 5442
rect 15668 5436 15900 5908
rect 16558 5906 16616 5908
rect 16750 5906 16808 5908
rect 16942 5906 17000 5908
rect 17134 5906 17192 5908
rect 17326 5906 17384 5908
rect 16420 5862 16466 5874
rect 16420 5652 16426 5862
rect 16460 5652 16466 5862
rect 16502 5696 16512 5876
rect 16564 5696 16574 5876
rect 16612 5862 16658 5874
rect 16406 5472 16416 5652
rect 16468 5472 16478 5652
rect 16516 5486 16522 5696
rect 16556 5486 16562 5696
rect 16612 5652 16618 5862
rect 16652 5652 16658 5862
rect 16694 5696 16704 5876
rect 16756 5696 16766 5876
rect 16804 5862 16850 5874
rect 16516 5474 16562 5486
rect 16598 5472 16608 5652
rect 16660 5472 16670 5652
rect 16708 5486 16714 5696
rect 16748 5486 16754 5696
rect 16804 5652 16810 5862
rect 16844 5652 16850 5862
rect 16886 5696 16896 5876
rect 16948 5696 16958 5876
rect 16996 5862 17042 5874
rect 16708 5474 16754 5486
rect 16790 5472 16800 5652
rect 16852 5472 16862 5652
rect 16900 5486 16906 5696
rect 16940 5486 16946 5696
rect 16996 5652 17002 5862
rect 17036 5652 17042 5862
rect 17078 5696 17088 5876
rect 17140 5696 17150 5876
rect 17188 5862 17234 5874
rect 16900 5474 16946 5486
rect 16982 5472 16992 5652
rect 17044 5472 17054 5652
rect 17092 5486 17098 5696
rect 17132 5486 17138 5696
rect 17188 5652 17194 5862
rect 17228 5652 17234 5862
rect 17270 5696 17280 5876
rect 17332 5696 17342 5876
rect 17380 5862 17426 5874
rect 17092 5474 17138 5486
rect 17174 5472 17184 5652
rect 17236 5472 17246 5652
rect 17284 5486 17290 5696
rect 17324 5486 17330 5696
rect 17380 5652 17386 5862
rect 17420 5652 17426 5862
rect 17284 5474 17330 5486
rect 17366 5472 17376 5652
rect 17428 5472 17438 5652
rect 16462 5436 16520 5442
rect 16654 5436 16712 5442
rect 16846 5436 16904 5442
rect 17038 5436 17096 5442
rect 17230 5436 17288 5442
rect 17468 5436 17704 5908
rect 18358 5906 18416 5908
rect 18550 5906 18608 5908
rect 18742 5906 18800 5908
rect 18934 5906 18992 5908
rect 19126 5906 19184 5908
rect 18220 5862 18266 5874
rect 18220 5652 18226 5862
rect 18260 5652 18266 5862
rect 18302 5696 18312 5876
rect 18364 5696 18374 5876
rect 18412 5862 18458 5874
rect 18206 5472 18216 5652
rect 18268 5472 18278 5652
rect 18316 5486 18322 5696
rect 18356 5486 18362 5696
rect 18412 5652 18418 5862
rect 18452 5652 18458 5862
rect 18494 5696 18504 5876
rect 18556 5696 18566 5876
rect 18604 5862 18650 5874
rect 18316 5474 18362 5486
rect 18398 5472 18408 5652
rect 18460 5472 18470 5652
rect 18508 5486 18514 5696
rect 18548 5486 18554 5696
rect 18604 5652 18610 5862
rect 18644 5652 18650 5862
rect 18686 5696 18696 5876
rect 18748 5696 18758 5876
rect 18796 5862 18842 5874
rect 18508 5474 18554 5486
rect 18590 5472 18600 5652
rect 18652 5472 18662 5652
rect 18700 5486 18706 5696
rect 18740 5486 18746 5696
rect 18796 5652 18802 5862
rect 18836 5652 18842 5862
rect 18878 5696 18888 5876
rect 18940 5696 18950 5876
rect 18988 5862 19034 5874
rect 18700 5474 18746 5486
rect 18782 5472 18792 5652
rect 18844 5472 18854 5652
rect 18892 5486 18898 5696
rect 18932 5486 18938 5696
rect 18988 5652 18994 5862
rect 19028 5652 19034 5862
rect 19070 5696 19080 5876
rect 19132 5696 19142 5876
rect 19180 5862 19226 5874
rect 18892 5474 18938 5486
rect 18974 5472 18984 5652
rect 19036 5472 19046 5652
rect 19084 5486 19090 5696
rect 19124 5486 19130 5696
rect 19180 5652 19186 5862
rect 19220 5652 19226 5862
rect 19084 5474 19130 5486
rect 19166 5472 19176 5652
rect 19228 5472 19238 5652
rect 18262 5436 18320 5442
rect 18454 5436 18512 5442
rect 18646 5436 18704 5442
rect 18838 5436 18896 5442
rect 19030 5436 19088 5442
rect 19268 5436 19504 5908
rect 20158 5906 20216 5908
rect 20350 5906 20408 5908
rect 20542 5906 20600 5908
rect 20734 5906 20792 5908
rect 20926 5906 20984 5908
rect 20020 5862 20066 5874
rect 20020 5652 20026 5862
rect 20060 5652 20066 5862
rect 20102 5696 20112 5876
rect 20164 5696 20174 5876
rect 20212 5862 20258 5874
rect 20006 5472 20016 5652
rect 20068 5472 20078 5652
rect 20116 5486 20122 5696
rect 20156 5486 20162 5696
rect 20212 5652 20218 5862
rect 20252 5652 20258 5862
rect 20294 5696 20304 5876
rect 20356 5696 20366 5876
rect 20404 5862 20450 5874
rect 20116 5474 20162 5486
rect 20198 5472 20208 5652
rect 20260 5472 20270 5652
rect 20308 5486 20314 5696
rect 20348 5486 20354 5696
rect 20404 5652 20410 5862
rect 20444 5652 20450 5862
rect 20486 5696 20496 5876
rect 20548 5696 20558 5876
rect 20596 5862 20642 5874
rect 20308 5474 20354 5486
rect 20390 5472 20400 5652
rect 20452 5472 20462 5652
rect 20500 5486 20506 5696
rect 20540 5486 20546 5696
rect 20596 5652 20602 5862
rect 20636 5652 20642 5862
rect 20678 5696 20688 5876
rect 20740 5696 20750 5876
rect 20788 5862 20834 5874
rect 20500 5474 20546 5486
rect 20582 5472 20592 5652
rect 20644 5472 20654 5652
rect 20692 5486 20698 5696
rect 20732 5486 20738 5696
rect 20788 5652 20794 5862
rect 20828 5652 20834 5862
rect 20870 5696 20880 5876
rect 20932 5696 20942 5876
rect 20980 5862 21026 5874
rect 20692 5474 20738 5486
rect 20774 5472 20784 5652
rect 20836 5472 20846 5652
rect 20884 5486 20890 5696
rect 20924 5486 20930 5696
rect 20980 5652 20986 5862
rect 21020 5652 21026 5862
rect 20884 5474 20930 5486
rect 20966 5472 20976 5652
rect 21028 5472 21038 5652
rect 20062 5436 20120 5442
rect 20254 5436 20312 5442
rect 20446 5436 20504 5442
rect 20638 5436 20696 5442
rect 20830 5436 20888 5442
rect 21068 5436 21304 5908
rect 21478 5580 21488 6080
rect 21772 6008 23852 6080
rect 21772 5974 22074 6008
rect 22108 5974 22266 6008
rect 22300 5974 22458 6008
rect 22492 5974 22650 6008
rect 22684 5974 22842 6008
rect 22876 5974 23034 6008
rect 23068 5974 23226 6008
rect 23260 5974 23418 6008
rect 23452 5974 23610 6008
rect 23644 5974 23802 6008
rect 23836 5974 23852 6008
rect 21772 5968 23852 5974
rect 21772 5580 21976 5968
rect 22020 5924 22066 5936
rect 22020 5720 22026 5924
rect 22060 5720 22066 5924
rect 22102 5756 22112 5940
rect 22168 5756 22178 5940
rect 22212 5924 22258 5936
rect 14004 5402 14674 5436
rect 14708 5402 14866 5436
rect 14900 5402 15058 5436
rect 15092 5402 15250 5436
rect 15284 5402 15442 5436
rect 15476 5402 16474 5436
rect 16508 5402 16666 5436
rect 16700 5402 16858 5436
rect 16892 5402 17050 5436
rect 17084 5402 17242 5436
rect 17276 5402 18274 5436
rect 18308 5402 18466 5436
rect 18500 5402 18658 5436
rect 18692 5402 18850 5436
rect 18884 5402 19042 5436
rect 19076 5402 20074 5436
rect 20108 5402 20266 5436
rect 20300 5402 20458 5436
rect 20492 5402 20650 5436
rect 20684 5402 20842 5436
rect 20876 5402 21304 5436
rect 14004 5328 21304 5402
rect 14004 5294 14674 5328
rect 14708 5294 14866 5328
rect 14900 5294 15058 5328
rect 15092 5294 15250 5328
rect 15284 5294 15442 5328
rect 15476 5294 16474 5328
rect 16508 5294 16666 5328
rect 16700 5294 16858 5328
rect 16892 5294 17050 5328
rect 17084 5294 17242 5328
rect 17276 5294 18274 5328
rect 18308 5294 18466 5328
rect 18500 5294 18658 5328
rect 18692 5294 18850 5328
rect 18884 5294 19042 5328
rect 19076 5294 20074 5328
rect 20108 5294 20266 5328
rect 20300 5294 20458 5328
rect 20492 5294 20650 5328
rect 20684 5294 20842 5328
rect 20876 5294 21304 5328
rect 14004 5292 21304 5294
rect 14004 5092 14484 5292
rect 14662 5288 14720 5292
rect 14854 5288 14912 5292
rect 15046 5288 15104 5292
rect 15238 5288 15296 5292
rect 15430 5288 15488 5292
rect 11400 4860 11900 4920
rect 11400 4580 11480 4860
rect 11820 4580 11900 4860
rect 11400 4520 11900 4580
rect 11480 4500 11900 4520
rect 13986 4400 13996 5092
rect 14428 4820 14484 5092
rect 14620 5244 14666 5256
rect 14620 5036 14626 5244
rect 14660 5036 14666 5244
rect 14702 5080 14712 5260
rect 14764 5080 14774 5260
rect 14812 5244 14858 5256
rect 14606 4856 14616 5036
rect 14668 4856 14678 5036
rect 14716 4868 14722 5080
rect 14756 4868 14762 5080
rect 14812 5036 14818 5244
rect 14852 5036 14858 5244
rect 14894 5080 14904 5260
rect 14956 5080 14966 5260
rect 15004 5244 15050 5256
rect 14716 4856 14762 4868
rect 14798 4856 14808 5036
rect 14860 4856 14870 5036
rect 14908 4868 14914 5080
rect 14948 4868 14954 5080
rect 15004 5036 15010 5244
rect 15044 5036 15050 5244
rect 15086 5080 15096 5260
rect 15148 5080 15158 5260
rect 15196 5244 15242 5256
rect 14908 4856 14954 4868
rect 14990 4856 15000 5036
rect 15052 4856 15062 5036
rect 15100 4868 15106 5080
rect 15140 4868 15146 5080
rect 15196 5036 15202 5244
rect 15236 5036 15242 5244
rect 15278 5080 15288 5260
rect 15340 5080 15350 5260
rect 15388 5244 15434 5256
rect 15100 4856 15146 4868
rect 15182 4856 15192 5036
rect 15244 4856 15254 5036
rect 15292 4868 15298 5080
rect 15332 4868 15338 5080
rect 15388 5036 15394 5244
rect 15428 5036 15434 5244
rect 15470 5080 15480 5260
rect 15532 5080 15542 5260
rect 15580 5244 15626 5256
rect 15292 4856 15338 4868
rect 15374 4856 15384 5036
rect 15436 4856 15446 5036
rect 15484 4868 15490 5080
rect 15524 4868 15530 5080
rect 15580 5036 15586 5244
rect 15620 5036 15626 5244
rect 15484 4856 15530 4868
rect 15566 4856 15576 5036
rect 15628 4856 15638 5036
rect 14758 4820 14816 4824
rect 14950 4820 15008 4824
rect 15142 4820 15200 4824
rect 15334 4820 15392 4824
rect 15526 4820 15584 4824
rect 15668 4820 15900 5292
rect 16462 5288 16520 5292
rect 16654 5288 16712 5292
rect 16846 5288 16904 5292
rect 17038 5288 17096 5292
rect 17230 5288 17288 5292
rect 16420 5244 16466 5256
rect 16420 5036 16426 5244
rect 16460 5036 16466 5244
rect 16502 5080 16512 5260
rect 16564 5080 16574 5260
rect 16612 5244 16658 5256
rect 16406 4856 16416 5036
rect 16468 4856 16478 5036
rect 16516 4868 16522 5080
rect 16556 4868 16562 5080
rect 16612 5036 16618 5244
rect 16652 5036 16658 5244
rect 16694 5080 16704 5260
rect 16756 5080 16766 5260
rect 16804 5244 16850 5256
rect 16516 4856 16562 4868
rect 16598 4856 16608 5036
rect 16660 4856 16670 5036
rect 16708 4868 16714 5080
rect 16748 4868 16754 5080
rect 16804 5036 16810 5244
rect 16844 5036 16850 5244
rect 16886 5080 16896 5260
rect 16948 5080 16958 5260
rect 16996 5244 17042 5256
rect 16708 4856 16754 4868
rect 16790 4856 16800 5036
rect 16852 4856 16862 5036
rect 16900 4868 16906 5080
rect 16940 4868 16946 5080
rect 16996 5036 17002 5244
rect 17036 5036 17042 5244
rect 17078 5080 17088 5260
rect 17140 5080 17150 5260
rect 17188 5244 17234 5256
rect 16900 4856 16946 4868
rect 16982 4856 16992 5036
rect 17044 4856 17054 5036
rect 17092 4868 17098 5080
rect 17132 4868 17138 5080
rect 17188 5036 17194 5244
rect 17228 5036 17234 5244
rect 17270 5080 17280 5260
rect 17332 5080 17342 5260
rect 17380 5244 17426 5256
rect 17092 4856 17138 4868
rect 17174 4856 17184 5036
rect 17236 4856 17246 5036
rect 17284 4868 17290 5080
rect 17324 4868 17330 5080
rect 17380 5036 17386 5244
rect 17420 5036 17426 5244
rect 17284 4856 17330 4868
rect 17366 4856 17376 5036
rect 17428 4856 17438 5036
rect 16558 4820 16616 4824
rect 16750 4820 16808 4824
rect 16942 4820 17000 4824
rect 17134 4820 17192 4824
rect 17326 4820 17384 4824
rect 17468 4820 17704 5292
rect 18262 5288 18320 5292
rect 18454 5288 18512 5292
rect 18646 5288 18704 5292
rect 18838 5288 18896 5292
rect 19030 5288 19088 5292
rect 18220 5244 18266 5256
rect 18220 5036 18226 5244
rect 18260 5036 18266 5244
rect 18302 5080 18312 5260
rect 18364 5080 18374 5260
rect 18412 5244 18458 5256
rect 18206 4856 18216 5036
rect 18268 4856 18278 5036
rect 18316 4868 18322 5080
rect 18356 4868 18362 5080
rect 18412 5036 18418 5244
rect 18452 5036 18458 5244
rect 18494 5080 18504 5260
rect 18556 5080 18566 5260
rect 18604 5244 18650 5256
rect 18316 4856 18362 4868
rect 18398 4856 18408 5036
rect 18460 4856 18470 5036
rect 18508 4868 18514 5080
rect 18548 4868 18554 5080
rect 18604 5036 18610 5244
rect 18644 5036 18650 5244
rect 18686 5080 18696 5260
rect 18748 5080 18758 5260
rect 18796 5244 18842 5256
rect 18508 4856 18554 4868
rect 18590 4856 18600 5036
rect 18652 4856 18662 5036
rect 18700 4868 18706 5080
rect 18740 4868 18746 5080
rect 18796 5036 18802 5244
rect 18836 5036 18842 5244
rect 18878 5080 18888 5260
rect 18940 5080 18950 5260
rect 18988 5244 19034 5256
rect 18700 4856 18746 4868
rect 18782 4856 18792 5036
rect 18844 4856 18854 5036
rect 18892 4868 18898 5080
rect 18932 4868 18938 5080
rect 18988 5036 18994 5244
rect 19028 5036 19034 5244
rect 19070 5080 19080 5260
rect 19132 5080 19142 5260
rect 19180 5244 19226 5256
rect 18892 4856 18938 4868
rect 18974 4856 18984 5036
rect 19036 4856 19046 5036
rect 19084 4868 19090 5080
rect 19124 4868 19130 5080
rect 19180 5036 19186 5244
rect 19220 5036 19226 5244
rect 19084 4856 19130 4868
rect 19166 4856 19176 5036
rect 19228 4856 19238 5036
rect 18358 4820 18416 4824
rect 18550 4820 18608 4824
rect 18742 4820 18800 4824
rect 18934 4820 18992 4824
rect 19126 4820 19184 4824
rect 19268 4820 19504 5292
rect 20062 5288 20120 5292
rect 20254 5288 20312 5292
rect 20446 5288 20504 5292
rect 20638 5288 20696 5292
rect 20830 5288 20888 5292
rect 20020 5244 20066 5256
rect 20020 5036 20026 5244
rect 20060 5036 20066 5244
rect 20102 5080 20112 5260
rect 20164 5080 20174 5260
rect 20212 5244 20258 5256
rect 20006 4856 20016 5036
rect 20068 4856 20078 5036
rect 20116 4868 20122 5080
rect 20156 4868 20162 5080
rect 20212 5036 20218 5244
rect 20252 5036 20258 5244
rect 20294 5080 20304 5260
rect 20356 5080 20366 5260
rect 20404 5244 20450 5256
rect 20116 4856 20162 4868
rect 20198 4856 20208 5036
rect 20260 4856 20270 5036
rect 20308 4868 20314 5080
rect 20348 4868 20354 5080
rect 20404 5036 20410 5244
rect 20444 5036 20450 5244
rect 20486 5080 20496 5260
rect 20548 5080 20558 5260
rect 20596 5244 20642 5256
rect 20308 4856 20354 4868
rect 20390 4856 20400 5036
rect 20452 4856 20462 5036
rect 20500 4868 20506 5080
rect 20540 4868 20546 5080
rect 20596 5036 20602 5244
rect 20636 5036 20642 5244
rect 20678 5080 20688 5260
rect 20740 5080 20750 5260
rect 20788 5244 20834 5256
rect 20500 4856 20546 4868
rect 20582 4856 20592 5036
rect 20644 4856 20654 5036
rect 20692 4868 20698 5080
rect 20732 4868 20738 5080
rect 20788 5036 20794 5244
rect 20828 5036 20834 5244
rect 20870 5080 20880 5260
rect 20932 5080 20942 5260
rect 20980 5244 21026 5256
rect 20692 4856 20738 4868
rect 20774 4856 20784 5036
rect 20836 4856 20846 5036
rect 20884 4868 20890 5080
rect 20924 4868 20930 5080
rect 20980 5036 20986 5244
rect 21020 5036 21026 5244
rect 20884 4856 20930 4868
rect 20966 4856 20976 5036
rect 21028 4856 21038 5036
rect 20158 4820 20216 4824
rect 20350 4820 20408 4824
rect 20542 4820 20600 4824
rect 20734 4820 20792 4824
rect 20926 4820 20984 4824
rect 21068 4820 21304 5292
rect 14428 4818 21304 4820
rect 14428 4784 14770 4818
rect 14804 4784 14962 4818
rect 14996 4784 15154 4818
rect 15188 4784 15346 4818
rect 15380 4784 15538 4818
rect 15572 4784 16570 4818
rect 16604 4784 16762 4818
rect 16796 4784 16954 4818
rect 16988 4784 17146 4818
rect 17180 4784 17338 4818
rect 17372 4784 18370 4818
rect 18404 4784 18562 4818
rect 18596 4784 18754 4818
rect 18788 4784 18946 4818
rect 18980 4784 19138 4818
rect 19172 4784 20170 4818
rect 20204 4784 20362 4818
rect 20396 4784 20554 4818
rect 20588 4784 20746 4818
rect 20780 4784 20938 4818
rect 20972 4784 21304 4818
rect 21556 5504 21976 5580
rect 22006 5536 22016 5720
rect 22072 5536 22082 5720
rect 22116 5548 22122 5756
rect 22156 5548 22162 5756
rect 22212 5720 22218 5924
rect 22252 5720 22258 5924
rect 22294 5756 22304 5940
rect 22360 5756 22370 5940
rect 22404 5924 22450 5936
rect 22116 5536 22162 5548
rect 22198 5536 22208 5720
rect 22264 5536 22274 5720
rect 22308 5548 22314 5756
rect 22348 5548 22354 5756
rect 22404 5720 22410 5924
rect 22444 5720 22450 5924
rect 22486 5756 22496 5940
rect 22552 5756 22562 5940
rect 22596 5924 22642 5936
rect 22308 5536 22354 5548
rect 22390 5536 22400 5720
rect 22456 5536 22466 5720
rect 22500 5548 22506 5756
rect 22540 5548 22546 5756
rect 22596 5720 22602 5924
rect 22636 5720 22642 5924
rect 22678 5756 22688 5940
rect 22744 5756 22754 5940
rect 22788 5924 22834 5936
rect 22500 5536 22546 5548
rect 22582 5536 22592 5720
rect 22648 5536 22658 5720
rect 22692 5548 22698 5756
rect 22732 5548 22738 5756
rect 22788 5720 22794 5924
rect 22828 5720 22834 5924
rect 22870 5756 22880 5940
rect 22936 5756 22946 5940
rect 22980 5924 23026 5936
rect 22692 5536 22738 5548
rect 22774 5536 22784 5720
rect 22840 5536 22850 5720
rect 22884 5548 22890 5756
rect 22924 5548 22930 5756
rect 22980 5720 22986 5924
rect 23020 5720 23026 5924
rect 23062 5756 23072 5940
rect 23128 5756 23138 5940
rect 23172 5924 23218 5936
rect 22884 5536 22930 5548
rect 22966 5536 22976 5720
rect 23032 5536 23042 5720
rect 23076 5548 23082 5756
rect 23116 5548 23122 5756
rect 23172 5720 23178 5924
rect 23212 5720 23218 5924
rect 23254 5756 23264 5940
rect 23320 5756 23330 5940
rect 23364 5924 23410 5936
rect 23076 5536 23122 5548
rect 23158 5536 23168 5720
rect 23224 5536 23234 5720
rect 23268 5548 23274 5756
rect 23308 5548 23314 5756
rect 23364 5720 23370 5924
rect 23404 5720 23410 5924
rect 23446 5756 23456 5940
rect 23512 5756 23522 5940
rect 23556 5924 23602 5936
rect 23268 5536 23314 5548
rect 23350 5536 23360 5720
rect 23416 5536 23426 5720
rect 23460 5548 23466 5756
rect 23500 5548 23506 5756
rect 23556 5720 23562 5924
rect 23596 5720 23602 5924
rect 23638 5756 23648 5940
rect 23704 5756 23714 5940
rect 23748 5924 23794 5936
rect 23460 5536 23506 5548
rect 23542 5536 23552 5720
rect 23608 5536 23618 5720
rect 23652 5548 23658 5756
rect 23692 5548 23698 5756
rect 23748 5720 23754 5924
rect 23788 5720 23794 5924
rect 23830 5756 23840 5940
rect 23896 5756 23906 5940
rect 23940 5924 23986 5936
rect 23652 5536 23698 5548
rect 23734 5536 23744 5720
rect 23800 5536 23810 5720
rect 23844 5548 23850 5756
rect 23884 5548 23890 5756
rect 23940 5720 23946 5924
rect 23980 5720 23986 5924
rect 23844 5536 23890 5548
rect 23926 5536 23936 5720
rect 23992 5536 24002 5720
rect 21556 5498 23948 5504
rect 21556 5464 22170 5498
rect 22204 5464 22362 5498
rect 22396 5464 22554 5498
rect 22588 5464 22746 5498
rect 22780 5464 22938 5498
rect 22972 5464 23130 5498
rect 23164 5464 23322 5498
rect 23356 5464 23514 5498
rect 23548 5464 23706 5498
rect 23740 5464 23898 5498
rect 23932 5464 23948 5498
rect 21556 5390 23948 5464
rect 21556 5356 22170 5390
rect 22204 5356 22362 5390
rect 22396 5356 22554 5390
rect 22588 5356 22746 5390
rect 22780 5356 22938 5390
rect 22972 5356 23130 5390
rect 23164 5356 23322 5390
rect 23356 5356 23514 5390
rect 23548 5356 23706 5390
rect 23740 5356 23898 5390
rect 23932 5356 23948 5390
rect 21556 5348 23948 5356
rect 21556 4888 21976 5348
rect 22020 5306 22066 5318
rect 22020 5100 22026 5306
rect 22060 5100 22066 5306
rect 22102 5136 22112 5320
rect 22168 5136 22178 5320
rect 22212 5306 22258 5318
rect 22006 4916 22016 5100
rect 22072 4916 22082 5100
rect 22116 4930 22122 5136
rect 22156 4930 22162 5136
rect 22212 5100 22218 5306
rect 22252 5100 22258 5306
rect 22294 5136 22304 5320
rect 22360 5136 22370 5320
rect 22404 5306 22450 5318
rect 22116 4918 22162 4930
rect 22198 4916 22208 5100
rect 22264 4916 22274 5100
rect 22308 4930 22314 5136
rect 22348 4930 22354 5136
rect 22404 5100 22410 5306
rect 22444 5100 22450 5306
rect 22486 5136 22496 5320
rect 22552 5136 22562 5320
rect 22596 5306 22642 5318
rect 22308 4918 22354 4930
rect 22390 4916 22400 5100
rect 22456 4916 22466 5100
rect 22500 4930 22506 5136
rect 22540 4930 22546 5136
rect 22596 5100 22602 5306
rect 22636 5100 22642 5306
rect 22678 5136 22688 5320
rect 22744 5136 22754 5320
rect 22788 5306 22834 5318
rect 22500 4918 22546 4930
rect 22582 4916 22592 5100
rect 22648 4916 22658 5100
rect 22692 4930 22698 5136
rect 22732 4930 22738 5136
rect 22788 5100 22794 5306
rect 22828 5100 22834 5306
rect 22870 5136 22880 5320
rect 22936 5136 22946 5320
rect 22980 5306 23026 5318
rect 22692 4918 22738 4930
rect 22774 4916 22784 5100
rect 22840 4916 22850 5100
rect 22884 4930 22890 5136
rect 22924 4930 22930 5136
rect 22980 5100 22986 5306
rect 23020 5100 23026 5306
rect 23062 5136 23072 5320
rect 23128 5136 23138 5320
rect 23172 5306 23218 5318
rect 22884 4918 22930 4930
rect 22966 4916 22976 5100
rect 23032 4916 23042 5100
rect 23076 4930 23082 5136
rect 23116 4930 23122 5136
rect 23172 5100 23178 5306
rect 23212 5100 23218 5306
rect 23254 5136 23264 5320
rect 23320 5136 23330 5320
rect 23364 5306 23410 5318
rect 23076 4918 23122 4930
rect 23158 4916 23168 5100
rect 23224 4916 23234 5100
rect 23268 4930 23274 5136
rect 23308 4930 23314 5136
rect 23364 5100 23370 5306
rect 23404 5100 23410 5306
rect 23446 5136 23456 5320
rect 23512 5136 23522 5320
rect 23556 5306 23602 5318
rect 23268 4918 23314 4930
rect 23350 4916 23360 5100
rect 23416 4916 23426 5100
rect 23460 4930 23466 5136
rect 23500 4930 23506 5136
rect 23556 5100 23562 5306
rect 23596 5100 23602 5306
rect 23638 5136 23648 5320
rect 23704 5136 23714 5320
rect 23748 5306 23794 5318
rect 23460 4918 23506 4930
rect 23542 4916 23552 5100
rect 23608 4916 23618 5100
rect 23652 4930 23658 5136
rect 23692 4930 23698 5136
rect 23748 5100 23754 5306
rect 23788 5100 23794 5306
rect 23830 5136 23840 5320
rect 23896 5136 23906 5320
rect 23940 5306 23986 5318
rect 23652 4918 23698 4930
rect 23734 4916 23744 5100
rect 23800 4916 23810 5100
rect 23844 4930 23850 5136
rect 23884 4930 23890 5136
rect 23940 5100 23946 5306
rect 23980 5100 23986 5306
rect 23844 4918 23890 4930
rect 23926 4916 23936 5100
rect 23992 4916 24002 5100
rect 21556 4880 23852 4888
rect 21556 4846 22074 4880
rect 22108 4846 22266 4880
rect 22300 4846 22458 4880
rect 22492 4846 22650 4880
rect 22684 4846 22842 4880
rect 22876 4846 23034 4880
rect 23068 4846 23226 4880
rect 23260 4846 23418 4880
rect 23452 4846 23610 4880
rect 23644 4846 23802 4880
rect 23836 4846 23852 4880
rect 21556 4792 23852 4846
rect 14428 4710 21304 4784
rect 14428 4676 14770 4710
rect 14804 4676 14962 4710
rect 14996 4676 15154 4710
rect 15188 4676 15346 4710
rect 15380 4676 15538 4710
rect 15572 4676 16570 4710
rect 16604 4676 16762 4710
rect 16796 4676 16954 4710
rect 16988 4676 17146 4710
rect 17180 4676 17338 4710
rect 17372 4676 18370 4710
rect 18404 4676 18562 4710
rect 18596 4676 18754 4710
rect 18788 4676 18946 4710
rect 18980 4676 19138 4710
rect 19172 4676 20170 4710
rect 20204 4676 20362 4710
rect 20396 4676 20554 4710
rect 20588 4676 20746 4710
rect 20780 4676 20938 4710
rect 20972 4676 21304 4710
rect 24520 4700 24900 11500
rect 14428 4400 14484 4676
rect 14758 4670 14816 4676
rect 14950 4670 15008 4676
rect 15142 4670 15200 4676
rect 15334 4670 15392 4676
rect 15526 4670 15584 4676
rect 14620 4626 14666 4638
rect 14620 4416 14626 4626
rect 14660 4416 14666 4626
rect 14702 4460 14712 4640
rect 14764 4460 14774 4640
rect 14812 4626 14858 4638
rect 14004 4200 14484 4400
rect 14606 4236 14616 4416
rect 14668 4236 14678 4416
rect 14716 4250 14722 4460
rect 14756 4250 14762 4460
rect 14812 4416 14818 4626
rect 14852 4416 14858 4626
rect 14894 4460 14904 4640
rect 14956 4460 14966 4640
rect 15004 4626 15050 4638
rect 14716 4238 14762 4250
rect 14798 4236 14808 4416
rect 14860 4236 14870 4416
rect 14908 4250 14914 4460
rect 14948 4250 14954 4460
rect 15004 4416 15010 4626
rect 15044 4416 15050 4626
rect 15086 4460 15096 4640
rect 15148 4460 15158 4640
rect 15196 4626 15242 4638
rect 14908 4238 14954 4250
rect 14990 4236 15000 4416
rect 15052 4236 15062 4416
rect 15100 4250 15106 4460
rect 15140 4250 15146 4460
rect 15196 4416 15202 4626
rect 15236 4416 15242 4626
rect 15278 4460 15288 4640
rect 15340 4460 15350 4640
rect 15388 4626 15434 4638
rect 15100 4238 15146 4250
rect 15182 4236 15192 4416
rect 15244 4236 15254 4416
rect 15292 4250 15298 4460
rect 15332 4250 15338 4460
rect 15388 4416 15394 4626
rect 15428 4416 15434 4626
rect 15470 4460 15480 4640
rect 15532 4460 15542 4640
rect 15580 4626 15626 4638
rect 15292 4238 15338 4250
rect 15374 4236 15384 4416
rect 15436 4236 15446 4416
rect 15484 4250 15490 4460
rect 15524 4250 15530 4460
rect 15580 4416 15586 4626
rect 15620 4416 15626 4626
rect 15484 4238 15530 4250
rect 15566 4236 15576 4416
rect 15628 4236 15638 4416
rect 14662 4200 14720 4206
rect 14854 4200 14912 4206
rect 15046 4200 15104 4206
rect 15238 4200 15296 4206
rect 15430 4200 15488 4206
rect 15668 4200 15900 4676
rect 16558 4670 16616 4676
rect 16750 4670 16808 4676
rect 16942 4670 17000 4676
rect 17134 4670 17192 4676
rect 17326 4670 17384 4676
rect 16420 4626 16466 4638
rect 16420 4416 16426 4626
rect 16460 4416 16466 4626
rect 16502 4460 16512 4640
rect 16564 4460 16574 4640
rect 16612 4626 16658 4638
rect 16406 4236 16416 4416
rect 16468 4236 16478 4416
rect 16516 4250 16522 4460
rect 16556 4250 16562 4460
rect 16612 4416 16618 4626
rect 16652 4416 16658 4626
rect 16694 4460 16704 4640
rect 16756 4460 16766 4640
rect 16804 4626 16850 4638
rect 16516 4238 16562 4250
rect 16598 4236 16608 4416
rect 16660 4236 16670 4416
rect 16708 4250 16714 4460
rect 16748 4250 16754 4460
rect 16804 4416 16810 4626
rect 16844 4416 16850 4626
rect 16886 4460 16896 4640
rect 16948 4460 16958 4640
rect 16996 4626 17042 4638
rect 16708 4238 16754 4250
rect 16790 4236 16800 4416
rect 16852 4236 16862 4416
rect 16900 4250 16906 4460
rect 16940 4250 16946 4460
rect 16996 4416 17002 4626
rect 17036 4416 17042 4626
rect 17078 4460 17088 4640
rect 17140 4460 17150 4640
rect 17188 4626 17234 4638
rect 16900 4238 16946 4250
rect 16982 4236 16992 4416
rect 17044 4236 17054 4416
rect 17092 4250 17098 4460
rect 17132 4250 17138 4460
rect 17188 4416 17194 4626
rect 17228 4416 17234 4626
rect 17270 4460 17280 4640
rect 17332 4460 17342 4640
rect 17380 4626 17426 4638
rect 17092 4238 17138 4250
rect 17174 4236 17184 4416
rect 17236 4236 17246 4416
rect 17284 4250 17290 4460
rect 17324 4250 17330 4460
rect 17380 4416 17386 4626
rect 17420 4416 17426 4626
rect 17284 4238 17330 4250
rect 17366 4236 17376 4416
rect 17428 4236 17438 4416
rect 16462 4200 16520 4206
rect 16654 4200 16712 4206
rect 16846 4200 16904 4206
rect 17038 4200 17096 4206
rect 17230 4200 17288 4206
rect 17468 4200 17704 4676
rect 18358 4670 18416 4676
rect 18550 4670 18608 4676
rect 18742 4670 18800 4676
rect 18934 4670 18992 4676
rect 19126 4670 19184 4676
rect 18220 4626 18266 4638
rect 18220 4416 18226 4626
rect 18260 4416 18266 4626
rect 18302 4460 18312 4640
rect 18364 4460 18374 4640
rect 18412 4626 18458 4638
rect 18206 4236 18216 4416
rect 18268 4236 18278 4416
rect 18316 4250 18322 4460
rect 18356 4250 18362 4460
rect 18412 4416 18418 4626
rect 18452 4416 18458 4626
rect 18494 4460 18504 4640
rect 18556 4460 18566 4640
rect 18604 4626 18650 4638
rect 18316 4238 18362 4250
rect 18398 4236 18408 4416
rect 18460 4236 18470 4416
rect 18508 4250 18514 4460
rect 18548 4250 18554 4460
rect 18604 4416 18610 4626
rect 18644 4416 18650 4626
rect 18686 4460 18696 4640
rect 18748 4460 18758 4640
rect 18796 4626 18842 4638
rect 18508 4238 18554 4250
rect 18590 4236 18600 4416
rect 18652 4236 18662 4416
rect 18700 4250 18706 4460
rect 18740 4250 18746 4460
rect 18796 4416 18802 4626
rect 18836 4416 18842 4626
rect 18878 4460 18888 4640
rect 18940 4460 18950 4640
rect 18988 4626 19034 4638
rect 18700 4238 18746 4250
rect 18782 4236 18792 4416
rect 18844 4236 18854 4416
rect 18892 4250 18898 4460
rect 18932 4250 18938 4460
rect 18988 4416 18994 4626
rect 19028 4416 19034 4626
rect 19070 4460 19080 4640
rect 19132 4460 19142 4640
rect 19180 4626 19226 4638
rect 18892 4238 18938 4250
rect 18974 4236 18984 4416
rect 19036 4236 19046 4416
rect 19084 4250 19090 4460
rect 19124 4250 19130 4460
rect 19180 4416 19186 4626
rect 19220 4416 19226 4626
rect 19084 4238 19130 4250
rect 19166 4236 19176 4416
rect 19228 4236 19238 4416
rect 18262 4200 18320 4206
rect 18454 4200 18512 4206
rect 18646 4200 18704 4206
rect 18838 4200 18896 4206
rect 19030 4200 19088 4206
rect 19268 4200 19504 4676
rect 20158 4670 20216 4676
rect 20350 4670 20408 4676
rect 20542 4670 20600 4676
rect 20734 4670 20792 4676
rect 20926 4670 20984 4676
rect 20020 4626 20066 4638
rect 20020 4416 20026 4626
rect 20060 4416 20066 4626
rect 20102 4460 20112 4640
rect 20164 4460 20174 4640
rect 20212 4626 20258 4638
rect 20006 4236 20016 4416
rect 20068 4236 20078 4416
rect 20116 4250 20122 4460
rect 20156 4250 20162 4460
rect 20212 4416 20218 4626
rect 20252 4416 20258 4626
rect 20294 4460 20304 4640
rect 20356 4460 20366 4640
rect 20404 4626 20450 4638
rect 20116 4238 20162 4250
rect 20198 4236 20208 4416
rect 20260 4236 20270 4416
rect 20308 4250 20314 4460
rect 20348 4250 20354 4460
rect 20404 4416 20410 4626
rect 20444 4416 20450 4626
rect 20486 4460 20496 4640
rect 20548 4460 20558 4640
rect 20596 4626 20642 4638
rect 20308 4238 20354 4250
rect 20390 4236 20400 4416
rect 20452 4236 20462 4416
rect 20500 4250 20506 4460
rect 20540 4250 20546 4460
rect 20596 4416 20602 4626
rect 20636 4416 20642 4626
rect 20678 4460 20688 4640
rect 20740 4460 20750 4640
rect 20788 4626 20834 4638
rect 20500 4238 20546 4250
rect 20582 4236 20592 4416
rect 20644 4236 20654 4416
rect 20692 4250 20698 4460
rect 20732 4250 20738 4460
rect 20788 4416 20794 4626
rect 20828 4416 20834 4626
rect 20870 4460 20880 4640
rect 20932 4460 20942 4640
rect 20980 4626 21026 4638
rect 20692 4238 20738 4250
rect 20774 4236 20784 4416
rect 20836 4236 20846 4416
rect 20884 4250 20890 4460
rect 20924 4250 20930 4460
rect 20980 4416 20986 4626
rect 21020 4416 21026 4626
rect 20884 4238 20930 4250
rect 20966 4236 20976 4416
rect 21028 4236 21038 4416
rect 20062 4200 20120 4206
rect 20254 4200 20312 4206
rect 20446 4200 20504 4206
rect 20638 4200 20696 4206
rect 20830 4200 20888 4206
rect 21068 4200 21304 4676
rect 24510 4360 24520 4700
rect 24900 4360 24910 4700
rect -3192 4196 84 4200
rect 256 4196 274 4200
rect -3192 4166 274 4196
rect 308 4166 466 4200
rect 500 4166 658 4200
rect 692 4166 850 4200
rect 884 4166 1042 4200
rect 1076 4196 1500 4200
rect 2056 4196 2074 4200
rect 1076 4166 2074 4196
rect 2108 4166 2266 4200
rect 2300 4166 2458 4200
rect 2492 4166 2650 4200
rect 2684 4166 2842 4200
rect 2876 4196 3304 4200
rect 3856 4196 3874 4200
rect 2876 4166 3874 4196
rect 3908 4166 4066 4200
rect 4100 4166 4258 4200
rect 4292 4166 4450 4200
rect 4484 4166 4642 4200
rect 4676 4196 5104 4200
rect 5656 4196 5674 4200
rect 4676 4166 5674 4196
rect 5708 4166 5866 4200
rect 5900 4166 6058 4200
rect 6092 4166 6250 4200
rect 6284 4166 6442 4200
rect 6476 4196 6904 4200
rect 7040 4196 14484 4200
rect 14656 4196 14674 4200
rect 6476 4166 14674 4196
rect 14708 4166 14866 4200
rect 14900 4166 15058 4200
rect 15092 4166 15250 4200
rect 15284 4166 15442 4200
rect 15476 4196 15900 4200
rect 16456 4196 16474 4200
rect 15476 4166 16474 4196
rect 16508 4166 16666 4200
rect 16700 4166 16858 4200
rect 16892 4166 17050 4200
rect 17084 4166 17242 4200
rect 17276 4196 17704 4200
rect 18256 4196 18274 4200
rect 17276 4166 18274 4196
rect 18308 4166 18466 4200
rect 18500 4166 18658 4200
rect 18692 4166 18850 4200
rect 18884 4166 19042 4200
rect 19076 4196 19504 4200
rect 20056 4196 20074 4200
rect 19076 4166 20074 4196
rect 20108 4166 20266 4200
rect 20300 4166 20458 4200
rect 20492 4166 20650 4200
rect 20684 4166 20842 4200
rect 20876 4196 21304 4200
rect 20876 4166 21536 4196
rect -10012 4080 -8772 4100
rect -10012 4046 -9988 4080
rect -9820 4046 -9730 4080
rect -9562 4046 -9472 4080
rect -9304 4046 -9214 4080
rect -9046 4046 -8956 4080
rect -8788 4046 -8772 4080
rect -3192 4048 21536 4166
rect -10012 4040 -8772 4046
rect -10070 3828 -10060 4008
rect -10008 3828 -9998 4008
rect -9798 3996 -9752 4008
rect -10056 3620 -10050 3828
rect -10016 3620 -10010 3828
rect -9798 3788 -9792 3996
rect -9758 3788 -9752 3996
rect -10056 3608 -10010 3620
rect -9810 3608 -9800 3788
rect -9748 3608 -9738 3788
rect -9708 3576 -9588 4040
rect -9554 3828 -9544 4008
rect -9492 3828 -9482 4008
rect -9540 3620 -9534 3828
rect -9500 3620 -9494 3828
rect -9540 3608 -9494 3620
rect -9448 3576 -9328 4040
rect -9282 3996 -9236 4008
rect -9282 3788 -9276 3996
rect -9242 3788 -9236 3996
rect -9294 3608 -9284 3788
rect -9232 3608 -9222 3788
rect -9188 3576 -9068 4040
rect -9038 3828 -9028 4008
rect -8976 3828 -8966 4008
rect -8766 3996 -8720 4008
rect -9024 3620 -9018 3828
rect -8984 3620 -8978 3828
rect -8766 3788 -8760 3996
rect -8726 3788 -8720 3996
rect -3224 3800 21536 4048
rect -3224 3788 288 3800
rect -9024 3608 -8978 3620
rect -8778 3608 -8768 3788
rect -8716 3608 -8706 3788
rect -3224 3780 80 3788
rect 264 3766 288 3788
rect 456 3766 546 3800
rect 714 3766 804 3800
rect 972 3766 1062 3800
rect 1230 3766 1320 3800
rect 1488 3788 2088 3800
rect 1488 3766 1504 3788
rect 264 3760 1504 3766
rect 2064 3766 2088 3788
rect 2256 3766 2346 3800
rect 2514 3766 2604 3800
rect 2772 3766 2862 3800
rect 3030 3766 3120 3800
rect 3288 3788 3888 3800
rect 3288 3766 3304 3788
rect 2064 3760 3304 3766
rect 3864 3766 3888 3788
rect 4056 3766 4146 3800
rect 4314 3766 4404 3800
rect 4572 3766 4662 3800
rect 4830 3766 4920 3800
rect 5088 3788 5688 3800
rect 5088 3766 5104 3788
rect 3864 3760 5104 3766
rect 5664 3766 5688 3788
rect 5856 3766 5946 3800
rect 6114 3766 6204 3800
rect 6372 3766 6462 3800
rect 6630 3766 6720 3800
rect 6888 3788 14688 3800
rect 6888 3766 6904 3788
rect 7040 3780 14220 3788
rect 5664 3760 6904 3766
rect 14664 3766 14688 3788
rect 14856 3766 14946 3800
rect 15114 3766 15204 3800
rect 15372 3766 15462 3800
rect 15630 3766 15720 3800
rect 15888 3788 16488 3800
rect 15888 3766 15904 3788
rect 14664 3760 15904 3766
rect 16464 3766 16488 3788
rect 16656 3766 16746 3800
rect 16914 3766 17004 3800
rect 17172 3766 17262 3800
rect 17430 3766 17520 3800
rect 17688 3788 18288 3800
rect 17688 3766 17704 3788
rect 16464 3760 17704 3766
rect 18264 3766 18288 3788
rect 18456 3766 18546 3800
rect 18714 3766 18804 3800
rect 18972 3766 19062 3800
rect 19230 3766 19320 3800
rect 19488 3788 20088 3800
rect 19488 3766 19504 3788
rect 18264 3760 19504 3766
rect 20064 3766 20088 3788
rect 20256 3766 20346 3800
rect 20514 3766 20604 3800
rect 20772 3766 20862 3800
rect 21030 3766 21120 3800
rect 21288 3788 21536 3800
rect 21288 3766 21304 3788
rect 20064 3760 21304 3766
rect -10012 3572 -8772 3576
rect -10016 3570 -8772 3572
rect -10016 3536 -9988 3570
rect -9820 3536 -9730 3570
rect -9562 3536 -9472 3570
rect -9304 3536 -9214 3570
rect -9046 3536 -8956 3570
rect -8788 3536 -8772 3570
rect 206 3548 216 3728
rect 268 3548 278 3728
rect 478 3716 524 3728
rect -10016 3462 -8772 3536
rect -10016 3428 -9988 3462
rect -9820 3428 -9730 3462
rect -9562 3428 -9472 3462
rect -9304 3428 -9214 3462
rect -9046 3428 -8956 3462
rect -8788 3428 -8772 3462
rect -10016 3424 -8772 3428
rect -10000 3422 -9808 3424
rect -9742 3422 -9550 3424
rect -9484 3422 -9292 3424
rect -9226 3422 -9034 3424
rect -8968 3422 -8776 3424
rect -10070 3212 -10060 3392
rect -10008 3212 -9998 3392
rect -9798 3378 -9752 3390
rect -10056 3002 -10050 3212
rect -10016 3002 -10010 3212
rect -9798 3172 -9792 3378
rect -9758 3172 -9752 3378
rect -10056 2990 -10010 3002
rect -9810 2992 -9800 3172
rect -9748 2992 -9738 3172
rect -9798 2990 -9752 2992
rect -9708 2958 -9588 3422
rect -9554 3212 -9544 3392
rect -9492 3212 -9482 3392
rect -9540 3002 -9534 3212
rect -9500 3002 -9494 3212
rect -9540 2990 -9494 3002
rect -9448 2960 -9328 3422
rect -9282 3378 -9236 3390
rect -9282 3172 -9276 3378
rect -9242 3172 -9236 3378
rect -9294 2992 -9284 3172
rect -9232 2992 -9222 3172
rect -9282 2990 -9236 2992
rect -9460 2958 -9316 2960
rect -9188 2958 -9068 3422
rect -9038 3212 -9028 3392
rect -8976 3212 -8966 3392
rect -8766 3378 -8720 3390
rect -9024 3002 -9018 3212
rect -8984 3002 -8978 3212
rect -8766 3172 -8760 3378
rect -8726 3172 -8720 3378
rect 220 3340 226 3548
rect 260 3340 266 3548
rect 478 3508 484 3716
rect 518 3508 524 3716
rect 220 3328 266 3340
rect 466 3328 476 3508
rect 528 3328 538 3508
rect 568 3296 688 3760
rect 722 3548 732 3728
rect 784 3548 794 3728
rect 736 3340 742 3548
rect 776 3340 782 3548
rect 736 3328 782 3340
rect 828 3296 948 3760
rect 994 3716 1040 3728
rect 994 3508 1000 3716
rect 1034 3508 1040 3716
rect 982 3328 992 3508
rect 1044 3328 1054 3508
rect 1088 3296 1208 3760
rect 1238 3548 1248 3728
rect 1300 3548 1310 3728
rect 1510 3716 1556 3728
rect 1252 3340 1258 3548
rect 1292 3340 1298 3548
rect 1510 3508 1516 3716
rect 1550 3508 1556 3716
rect 2006 3548 2016 3728
rect 2068 3548 2078 3728
rect 2278 3716 2324 3728
rect 1252 3328 1298 3340
rect 1498 3328 1508 3508
rect 1560 3328 1570 3508
rect 2020 3340 2026 3548
rect 2060 3340 2066 3548
rect 2278 3508 2284 3716
rect 2318 3508 2324 3716
rect 2020 3328 2066 3340
rect 2266 3328 2276 3508
rect 2328 3328 2338 3508
rect 2368 3296 2488 3760
rect 2522 3548 2532 3728
rect 2584 3548 2594 3728
rect 2536 3340 2542 3548
rect 2576 3340 2582 3548
rect 2536 3328 2582 3340
rect 2628 3296 2748 3760
rect 2794 3716 2840 3728
rect 2794 3508 2800 3716
rect 2834 3508 2840 3716
rect 2782 3328 2792 3508
rect 2844 3328 2854 3508
rect 2888 3296 3008 3760
rect 3038 3548 3048 3728
rect 3100 3548 3110 3728
rect 3310 3716 3356 3728
rect 3052 3340 3058 3548
rect 3092 3340 3098 3548
rect 3310 3508 3316 3716
rect 3350 3508 3356 3716
rect 3806 3548 3816 3728
rect 3868 3548 3878 3728
rect 4078 3716 4124 3728
rect 3052 3328 3098 3340
rect 3298 3328 3308 3508
rect 3360 3328 3370 3508
rect 3820 3340 3826 3548
rect 3860 3340 3866 3548
rect 4078 3508 4084 3716
rect 4118 3508 4124 3716
rect 3820 3328 3866 3340
rect 4066 3328 4076 3508
rect 4128 3328 4138 3508
rect 4168 3296 4288 3760
rect 4322 3548 4332 3728
rect 4384 3548 4394 3728
rect 4336 3340 4342 3548
rect 4376 3340 4382 3548
rect 4336 3328 4382 3340
rect 4428 3296 4548 3760
rect 4594 3716 4640 3728
rect 4594 3508 4600 3716
rect 4634 3508 4640 3716
rect 4582 3328 4592 3508
rect 4644 3328 4654 3508
rect 4688 3296 4808 3760
rect 4838 3548 4848 3728
rect 4900 3548 4910 3728
rect 5110 3716 5156 3728
rect 4852 3340 4858 3548
rect 4892 3340 4898 3548
rect 5110 3508 5116 3716
rect 5150 3508 5156 3716
rect 5606 3548 5616 3728
rect 5668 3548 5678 3728
rect 5878 3716 5924 3728
rect 4852 3328 4898 3340
rect 5098 3328 5108 3508
rect 5160 3328 5170 3508
rect 5620 3340 5626 3548
rect 5660 3340 5666 3548
rect 5878 3508 5884 3716
rect 5918 3508 5924 3716
rect 5620 3328 5666 3340
rect 5866 3328 5876 3508
rect 5928 3328 5938 3508
rect 5968 3296 6088 3760
rect 6122 3548 6132 3728
rect 6184 3548 6194 3728
rect 6136 3340 6142 3548
rect 6176 3340 6182 3548
rect 6136 3328 6182 3340
rect 6228 3296 6348 3760
rect 6394 3716 6440 3728
rect 6394 3508 6400 3716
rect 6434 3508 6440 3716
rect 6382 3328 6392 3508
rect 6444 3328 6454 3508
rect 6488 3296 6608 3760
rect 6638 3548 6648 3728
rect 6700 3548 6710 3728
rect 6910 3716 6956 3728
rect 6652 3340 6658 3548
rect 6692 3340 6698 3548
rect 6910 3508 6916 3716
rect 6950 3508 6956 3716
rect 14606 3548 14616 3728
rect 14668 3548 14678 3728
rect 14878 3716 14924 3728
rect 6652 3328 6698 3340
rect 6898 3328 6908 3508
rect 6960 3328 6970 3508
rect 14620 3340 14626 3548
rect 14660 3340 14666 3548
rect 14878 3508 14884 3716
rect 14918 3508 14924 3716
rect 14620 3328 14666 3340
rect 14866 3328 14876 3508
rect 14928 3328 14938 3508
rect 14968 3296 15088 3760
rect 15122 3548 15132 3728
rect 15184 3548 15194 3728
rect 15136 3340 15142 3548
rect 15176 3340 15182 3548
rect 15136 3328 15182 3340
rect 15228 3296 15348 3760
rect 15394 3716 15440 3728
rect 15394 3508 15400 3716
rect 15434 3508 15440 3716
rect 15382 3328 15392 3508
rect 15444 3328 15454 3508
rect 15488 3296 15608 3760
rect 15638 3548 15648 3728
rect 15700 3548 15710 3728
rect 15910 3716 15956 3728
rect 15652 3340 15658 3548
rect 15692 3340 15698 3548
rect 15910 3508 15916 3716
rect 15950 3508 15956 3716
rect 16406 3548 16416 3728
rect 16468 3548 16478 3728
rect 16678 3716 16724 3728
rect 15652 3328 15698 3340
rect 15898 3328 15908 3508
rect 15960 3328 15970 3508
rect 16420 3340 16426 3548
rect 16460 3340 16466 3548
rect 16678 3508 16684 3716
rect 16718 3508 16724 3716
rect 16420 3328 16466 3340
rect 16666 3328 16676 3508
rect 16728 3328 16738 3508
rect 16768 3296 16888 3760
rect 16922 3548 16932 3728
rect 16984 3548 16994 3728
rect 16936 3340 16942 3548
rect 16976 3340 16982 3548
rect 16936 3328 16982 3340
rect 17028 3296 17148 3760
rect 17194 3716 17240 3728
rect 17194 3508 17200 3716
rect 17234 3508 17240 3716
rect 17182 3328 17192 3508
rect 17244 3328 17254 3508
rect 17288 3296 17408 3760
rect 17438 3548 17448 3728
rect 17500 3548 17510 3728
rect 17710 3716 17756 3728
rect 17452 3340 17458 3548
rect 17492 3340 17498 3548
rect 17710 3508 17716 3716
rect 17750 3508 17756 3716
rect 18206 3548 18216 3728
rect 18268 3548 18278 3728
rect 18478 3716 18524 3728
rect 17452 3328 17498 3340
rect 17698 3328 17708 3508
rect 17760 3328 17770 3508
rect 18220 3340 18226 3548
rect 18260 3340 18266 3548
rect 18478 3508 18484 3716
rect 18518 3508 18524 3716
rect 18220 3328 18266 3340
rect 18466 3328 18476 3508
rect 18528 3328 18538 3508
rect 18568 3296 18688 3760
rect 18722 3548 18732 3728
rect 18784 3548 18794 3728
rect 18736 3340 18742 3548
rect 18776 3340 18782 3548
rect 18736 3328 18782 3340
rect 18828 3296 18948 3760
rect 18994 3716 19040 3728
rect 18994 3508 19000 3716
rect 19034 3508 19040 3716
rect 18982 3328 18992 3508
rect 19044 3328 19054 3508
rect 19088 3296 19208 3760
rect 19238 3548 19248 3728
rect 19300 3548 19310 3728
rect 19510 3716 19556 3728
rect 19252 3340 19258 3548
rect 19292 3340 19298 3548
rect 19510 3508 19516 3716
rect 19550 3508 19556 3716
rect 20006 3548 20016 3728
rect 20068 3548 20078 3728
rect 20278 3716 20324 3728
rect 19252 3328 19298 3340
rect 19498 3328 19508 3508
rect 19560 3328 19570 3508
rect 20020 3340 20026 3548
rect 20060 3340 20066 3548
rect 20278 3508 20284 3716
rect 20318 3508 20324 3716
rect 20020 3328 20066 3340
rect 20266 3328 20276 3508
rect 20328 3328 20338 3508
rect 20368 3296 20488 3760
rect 20522 3548 20532 3728
rect 20584 3548 20594 3728
rect 20536 3340 20542 3548
rect 20576 3340 20582 3548
rect 20536 3328 20582 3340
rect 20628 3296 20748 3760
rect 20794 3716 20840 3728
rect 20794 3508 20800 3716
rect 20834 3508 20840 3716
rect 20782 3328 20792 3508
rect 20844 3328 20854 3508
rect 20888 3296 21008 3760
rect 21038 3548 21048 3728
rect 21100 3548 21110 3728
rect 21310 3716 21356 3728
rect 21052 3340 21058 3548
rect 21092 3340 21098 3548
rect 21310 3508 21316 3716
rect 21350 3508 21356 3716
rect 21052 3328 21098 3340
rect 21298 3328 21308 3508
rect 21360 3328 21370 3508
rect 24520 3420 24900 4360
rect 264 3292 1504 3296
rect 2064 3292 3304 3296
rect 3864 3292 5104 3296
rect 5664 3292 6904 3296
rect 14664 3292 15904 3296
rect 16464 3292 17704 3296
rect 18264 3292 19504 3296
rect 20064 3292 21304 3296
rect 260 3290 1504 3292
rect 260 3256 288 3290
rect 456 3256 546 3290
rect 714 3256 804 3290
rect 972 3256 1062 3290
rect 1230 3256 1320 3290
rect 1488 3256 1504 3290
rect 260 3182 1504 3256
rect -9024 2990 -8978 3002
rect -8778 2992 -8768 3172
rect -8716 2992 -8706 3172
rect 260 3148 288 3182
rect 456 3148 546 3182
rect 714 3148 804 3182
rect 972 3148 1062 3182
rect 1230 3148 1320 3182
rect 1488 3148 1504 3182
rect 260 3144 1504 3148
rect 2060 3290 3304 3292
rect 2060 3256 2088 3290
rect 2256 3256 2346 3290
rect 2514 3256 2604 3290
rect 2772 3256 2862 3290
rect 3030 3256 3120 3290
rect 3288 3256 3304 3290
rect 2060 3182 3304 3256
rect 2060 3148 2088 3182
rect 2256 3148 2346 3182
rect 2514 3148 2604 3182
rect 2772 3148 2862 3182
rect 3030 3148 3120 3182
rect 3288 3148 3304 3182
rect 2060 3144 3304 3148
rect 3860 3290 5104 3292
rect 3860 3256 3888 3290
rect 4056 3256 4146 3290
rect 4314 3256 4404 3290
rect 4572 3256 4662 3290
rect 4830 3256 4920 3290
rect 5088 3256 5104 3290
rect 3860 3182 5104 3256
rect 3860 3148 3888 3182
rect 4056 3148 4146 3182
rect 4314 3148 4404 3182
rect 4572 3148 4662 3182
rect 4830 3148 4920 3182
rect 5088 3148 5104 3182
rect 3860 3144 5104 3148
rect 5660 3290 6904 3292
rect 5660 3256 5688 3290
rect 5856 3256 5946 3290
rect 6114 3256 6204 3290
rect 6372 3256 6462 3290
rect 6630 3256 6720 3290
rect 6888 3256 6904 3290
rect 5660 3182 6904 3256
rect 5660 3148 5688 3182
rect 5856 3148 5946 3182
rect 6114 3148 6204 3182
rect 6372 3148 6462 3182
rect 6630 3148 6720 3182
rect 6888 3148 6904 3182
rect 5660 3144 6904 3148
rect 14660 3290 15904 3292
rect 14660 3256 14688 3290
rect 14856 3256 14946 3290
rect 15114 3256 15204 3290
rect 15372 3256 15462 3290
rect 15630 3256 15720 3290
rect 15888 3256 15904 3290
rect 14660 3182 15904 3256
rect 14660 3148 14688 3182
rect 14856 3148 14946 3182
rect 15114 3148 15204 3182
rect 15372 3148 15462 3182
rect 15630 3148 15720 3182
rect 15888 3148 15904 3182
rect 14660 3144 15904 3148
rect 16460 3290 17704 3292
rect 16460 3256 16488 3290
rect 16656 3256 16746 3290
rect 16914 3256 17004 3290
rect 17172 3256 17262 3290
rect 17430 3256 17520 3290
rect 17688 3256 17704 3290
rect 16460 3182 17704 3256
rect 16460 3148 16488 3182
rect 16656 3148 16746 3182
rect 16914 3148 17004 3182
rect 17172 3148 17262 3182
rect 17430 3148 17520 3182
rect 17688 3148 17704 3182
rect 16460 3144 17704 3148
rect 18260 3290 19504 3292
rect 18260 3256 18288 3290
rect 18456 3256 18546 3290
rect 18714 3256 18804 3290
rect 18972 3256 19062 3290
rect 19230 3256 19320 3290
rect 19488 3256 19504 3290
rect 18260 3182 19504 3256
rect 18260 3148 18288 3182
rect 18456 3148 18546 3182
rect 18714 3148 18804 3182
rect 18972 3148 19062 3182
rect 19230 3148 19320 3182
rect 19488 3148 19504 3182
rect 18260 3144 19504 3148
rect 20060 3290 21304 3292
rect 20060 3256 20088 3290
rect 20256 3256 20346 3290
rect 20514 3256 20604 3290
rect 20772 3256 20862 3290
rect 21030 3256 21120 3290
rect 21288 3256 21304 3290
rect 20060 3182 21304 3256
rect 20060 3148 20088 3182
rect 20256 3148 20346 3182
rect 20514 3148 20604 3182
rect 20772 3148 20862 3182
rect 21030 3148 21120 3182
rect 21288 3148 21304 3182
rect 20060 3144 21304 3148
rect 276 3142 468 3144
rect 534 3142 726 3144
rect 792 3142 984 3144
rect 1050 3142 1242 3144
rect 1308 3142 1500 3144
rect 2076 3142 2268 3144
rect 2334 3142 2526 3144
rect 2592 3142 2784 3144
rect 2850 3142 3042 3144
rect 3108 3142 3300 3144
rect 3876 3142 4068 3144
rect 4134 3142 4326 3144
rect 4392 3142 4584 3144
rect 4650 3142 4842 3144
rect 4908 3142 5100 3144
rect 5676 3142 5868 3144
rect 5934 3142 6126 3144
rect 6192 3142 6384 3144
rect 6450 3142 6642 3144
rect 6708 3142 6900 3144
rect 14676 3142 14868 3144
rect 14934 3142 15126 3144
rect 15192 3142 15384 3144
rect 15450 3142 15642 3144
rect 15708 3142 15900 3144
rect 16476 3142 16668 3144
rect 16734 3142 16926 3144
rect 16992 3142 17184 3144
rect 17250 3142 17442 3144
rect 17508 3142 17700 3144
rect 18276 3142 18468 3144
rect 18534 3142 18726 3144
rect 18792 3142 18984 3144
rect 19050 3142 19242 3144
rect 19308 3142 19500 3144
rect 20076 3142 20268 3144
rect 20334 3142 20526 3144
rect 20592 3142 20784 3144
rect 20850 3142 21042 3144
rect 21108 3142 21300 3144
rect -8766 2990 -8720 2992
rect -10000 2956 -9808 2958
rect -9742 2956 -9550 2958
rect -9484 2956 -9292 2958
rect -9226 2956 -9034 2958
rect -8968 2956 -8776 2958
rect -10012 2952 -8772 2956
rect -10012 2918 -9988 2952
rect -9820 2918 -9730 2952
rect -9562 2918 -9472 2952
rect -9304 2918 -9214 2952
rect -9046 2918 -8956 2952
rect -8788 2918 -8768 2952
rect 206 2932 216 3112
rect 268 2932 278 3112
rect 478 3098 524 3110
rect -10012 2844 -8768 2918
rect -10012 2810 -9988 2844
rect -9820 2810 -9730 2844
rect -9562 2810 -9472 2844
rect -9304 2810 -9214 2844
rect -9046 2810 -8956 2844
rect -8788 2810 -8768 2844
rect -10012 2804 -8768 2810
rect -10070 2592 -10060 2772
rect -10008 2592 -9998 2772
rect -9798 2760 -9752 2772
rect -10056 2384 -10050 2592
rect -10016 2384 -10010 2592
rect -9798 2552 -9792 2760
rect -9758 2552 -9752 2760
rect -10056 2372 -10010 2384
rect -9810 2372 -9800 2552
rect -9748 2372 -9738 2552
rect -9708 2340 -9588 2804
rect -9554 2592 -9544 2772
rect -9492 2592 -9482 2772
rect -9540 2384 -9534 2592
rect -9500 2384 -9494 2592
rect -9540 2372 -9494 2384
rect -9448 2340 -9328 2804
rect -9282 2760 -9236 2772
rect -9282 2552 -9276 2760
rect -9242 2552 -9236 2760
rect -9294 2372 -9284 2552
rect -9232 2372 -9222 2552
rect -9188 2340 -9068 2804
rect -9038 2592 -9028 2772
rect -8976 2592 -8966 2772
rect -8766 2760 -8720 2772
rect -9024 2384 -9018 2592
rect -8984 2384 -8978 2592
rect -8766 2552 -8760 2760
rect -8726 2552 -8720 2760
rect 220 2722 226 2932
rect 260 2722 266 2932
rect 478 2892 484 3098
rect 518 2892 524 3098
rect 220 2710 266 2722
rect 466 2712 476 2892
rect 528 2712 538 2892
rect 478 2710 524 2712
rect 568 2678 688 3142
rect 722 2932 732 3112
rect 784 2932 794 3112
rect 736 2722 742 2932
rect 776 2722 782 2932
rect 736 2710 782 2722
rect 828 2680 948 3142
rect 994 3098 1040 3110
rect 994 2892 1000 3098
rect 1034 2892 1040 3098
rect 982 2712 992 2892
rect 1044 2712 1054 2892
rect 994 2710 1040 2712
rect 816 2678 960 2680
rect 1088 2678 1208 3142
rect 1238 2932 1248 3112
rect 1300 2932 1310 3112
rect 1510 3098 1556 3110
rect 1252 2722 1258 2932
rect 1292 2722 1298 2932
rect 1510 2892 1516 3098
rect 1550 2892 1556 3098
rect 2006 2932 2016 3112
rect 2068 2932 2078 3112
rect 2278 3098 2324 3110
rect 1252 2710 1298 2722
rect 1498 2712 1508 2892
rect 1560 2712 1570 2892
rect 2020 2722 2026 2932
rect 2060 2722 2066 2932
rect 2278 2892 2284 3098
rect 2318 2892 2324 3098
rect 1510 2710 1556 2712
rect 2020 2710 2066 2722
rect 2266 2712 2276 2892
rect 2328 2712 2338 2892
rect 2278 2710 2324 2712
rect 2368 2678 2488 3142
rect 2522 2932 2532 3112
rect 2584 2932 2594 3112
rect 2536 2722 2542 2932
rect 2576 2722 2582 2932
rect 2536 2710 2582 2722
rect 2628 2680 2748 3142
rect 2794 3098 2840 3110
rect 2794 2892 2800 3098
rect 2834 2892 2840 3098
rect 2782 2712 2792 2892
rect 2844 2712 2854 2892
rect 2794 2710 2840 2712
rect 2616 2678 2760 2680
rect 2888 2678 3008 3142
rect 3038 2932 3048 3112
rect 3100 2932 3110 3112
rect 3310 3098 3356 3110
rect 3052 2722 3058 2932
rect 3092 2722 3098 2932
rect 3310 2892 3316 3098
rect 3350 2892 3356 3098
rect 3806 2932 3816 3112
rect 3868 2932 3878 3112
rect 4078 3098 4124 3110
rect 3052 2710 3098 2722
rect 3298 2712 3308 2892
rect 3360 2712 3370 2892
rect 3820 2722 3826 2932
rect 3860 2722 3866 2932
rect 4078 2892 4084 3098
rect 4118 2892 4124 3098
rect 3310 2710 3356 2712
rect 3820 2710 3866 2722
rect 4066 2712 4076 2892
rect 4128 2712 4138 2892
rect 4078 2710 4124 2712
rect 4168 2678 4288 3142
rect 4322 2932 4332 3112
rect 4384 2932 4394 3112
rect 4336 2722 4342 2932
rect 4376 2722 4382 2932
rect 4336 2710 4382 2722
rect 4428 2680 4548 3142
rect 4594 3098 4640 3110
rect 4594 2892 4600 3098
rect 4634 2892 4640 3098
rect 4582 2712 4592 2892
rect 4644 2712 4654 2892
rect 4594 2710 4640 2712
rect 4416 2678 4560 2680
rect 4688 2678 4808 3142
rect 4838 2932 4848 3112
rect 4900 2932 4910 3112
rect 5110 3098 5156 3110
rect 4852 2722 4858 2932
rect 4892 2722 4898 2932
rect 5110 2892 5116 3098
rect 5150 2892 5156 3098
rect 5606 2932 5616 3112
rect 5668 2932 5678 3112
rect 5878 3098 5924 3110
rect 4852 2710 4898 2722
rect 5098 2712 5108 2892
rect 5160 2712 5170 2892
rect 5620 2722 5626 2932
rect 5660 2722 5666 2932
rect 5878 2892 5884 3098
rect 5918 2892 5924 3098
rect 5110 2710 5156 2712
rect 5620 2710 5666 2722
rect 5866 2712 5876 2892
rect 5928 2712 5938 2892
rect 5878 2710 5924 2712
rect 5968 2678 6088 3142
rect 6122 2932 6132 3112
rect 6184 2932 6194 3112
rect 6136 2722 6142 2932
rect 6176 2722 6182 2932
rect 6136 2710 6182 2722
rect 6228 2680 6348 3142
rect 6394 3098 6440 3110
rect 6394 2892 6400 3098
rect 6434 2892 6440 3098
rect 6382 2712 6392 2892
rect 6444 2712 6454 2892
rect 6394 2710 6440 2712
rect 6216 2678 6360 2680
rect 6488 2678 6608 3142
rect 6638 2932 6648 3112
rect 6700 2932 6710 3112
rect 6910 3098 6956 3110
rect 6652 2722 6658 2932
rect 6692 2722 6698 2932
rect 6910 2892 6916 3098
rect 6950 2892 6956 3098
rect 14606 2932 14616 3112
rect 14668 2932 14678 3112
rect 14878 3098 14924 3110
rect 6652 2710 6698 2722
rect 6898 2712 6908 2892
rect 6960 2712 6970 2892
rect 14620 2722 14626 2932
rect 14660 2722 14666 2932
rect 14878 2892 14884 3098
rect 14918 2892 14924 3098
rect 6910 2710 6956 2712
rect 14620 2710 14666 2722
rect 14866 2712 14876 2892
rect 14928 2712 14938 2892
rect 14878 2710 14924 2712
rect 14968 2678 15088 3142
rect 15122 2932 15132 3112
rect 15184 2932 15194 3112
rect 15136 2722 15142 2932
rect 15176 2722 15182 2932
rect 15136 2710 15182 2722
rect 15228 2680 15348 3142
rect 15394 3098 15440 3110
rect 15394 2892 15400 3098
rect 15434 2892 15440 3098
rect 15382 2712 15392 2892
rect 15444 2712 15454 2892
rect 15394 2710 15440 2712
rect 15216 2678 15360 2680
rect 15488 2678 15608 3142
rect 15638 2932 15648 3112
rect 15700 2932 15710 3112
rect 15910 3098 15956 3110
rect 15652 2722 15658 2932
rect 15692 2722 15698 2932
rect 15910 2892 15916 3098
rect 15950 2892 15956 3098
rect 16406 2932 16416 3112
rect 16468 2932 16478 3112
rect 16678 3098 16724 3110
rect 15652 2710 15698 2722
rect 15898 2712 15908 2892
rect 15960 2712 15970 2892
rect 16420 2722 16426 2932
rect 16460 2722 16466 2932
rect 16678 2892 16684 3098
rect 16718 2892 16724 3098
rect 15910 2710 15956 2712
rect 16420 2710 16466 2722
rect 16666 2712 16676 2892
rect 16728 2712 16738 2892
rect 16678 2710 16724 2712
rect 16768 2678 16888 3142
rect 16922 2932 16932 3112
rect 16984 2932 16994 3112
rect 16936 2722 16942 2932
rect 16976 2722 16982 2932
rect 16936 2710 16982 2722
rect 17028 2680 17148 3142
rect 17194 3098 17240 3110
rect 17194 2892 17200 3098
rect 17234 2892 17240 3098
rect 17182 2712 17192 2892
rect 17244 2712 17254 2892
rect 17194 2710 17240 2712
rect 17016 2678 17160 2680
rect 17288 2678 17408 3142
rect 17438 2932 17448 3112
rect 17500 2932 17510 3112
rect 17710 3098 17756 3110
rect 17452 2722 17458 2932
rect 17492 2722 17498 2932
rect 17710 2892 17716 3098
rect 17750 2892 17756 3098
rect 18206 2932 18216 3112
rect 18268 2932 18278 3112
rect 18478 3098 18524 3110
rect 17452 2710 17498 2722
rect 17698 2712 17708 2892
rect 17760 2712 17770 2892
rect 18220 2722 18226 2932
rect 18260 2722 18266 2932
rect 18478 2892 18484 3098
rect 18518 2892 18524 3098
rect 17710 2710 17756 2712
rect 18220 2710 18266 2722
rect 18466 2712 18476 2892
rect 18528 2712 18538 2892
rect 18478 2710 18524 2712
rect 18568 2678 18688 3142
rect 18722 2932 18732 3112
rect 18784 2932 18794 3112
rect 18736 2722 18742 2932
rect 18776 2722 18782 2932
rect 18736 2710 18782 2722
rect 18828 2680 18948 3142
rect 18994 3098 19040 3110
rect 18994 2892 19000 3098
rect 19034 2892 19040 3098
rect 18982 2712 18992 2892
rect 19044 2712 19054 2892
rect 18994 2710 19040 2712
rect 18816 2678 18960 2680
rect 19088 2678 19208 3142
rect 19238 2932 19248 3112
rect 19300 2932 19310 3112
rect 19510 3098 19556 3110
rect 19252 2722 19258 2932
rect 19292 2722 19298 2932
rect 19510 2892 19516 3098
rect 19550 2892 19556 3098
rect 20006 2932 20016 3112
rect 20068 2932 20078 3112
rect 20278 3098 20324 3110
rect 19252 2710 19298 2722
rect 19498 2712 19508 2892
rect 19560 2712 19570 2892
rect 20020 2722 20026 2932
rect 20060 2722 20066 2932
rect 20278 2892 20284 3098
rect 20318 2892 20324 3098
rect 19510 2710 19556 2712
rect 20020 2710 20066 2722
rect 20266 2712 20276 2892
rect 20328 2712 20338 2892
rect 20278 2710 20324 2712
rect 20368 2678 20488 3142
rect 20522 2932 20532 3112
rect 20584 2932 20594 3112
rect 20536 2722 20542 2932
rect 20576 2722 20582 2932
rect 20536 2710 20582 2722
rect 20628 2680 20748 3142
rect 20794 3098 20840 3110
rect 20794 2892 20800 3098
rect 20834 2892 20840 3098
rect 20782 2712 20792 2892
rect 20844 2712 20854 2892
rect 20794 2710 20840 2712
rect 20616 2678 20760 2680
rect 20888 2678 21008 3142
rect 21038 2932 21048 3112
rect 21100 2932 21110 3112
rect 21310 3098 21356 3110
rect 21052 2722 21058 2932
rect 21092 2722 21098 2932
rect 21310 2892 21316 3098
rect 21350 2892 21356 3098
rect 21052 2710 21098 2722
rect 21298 2712 21308 2892
rect 21360 2712 21370 2892
rect 21310 2710 21356 2712
rect 276 2676 468 2678
rect 534 2676 726 2678
rect 792 2676 984 2678
rect 1050 2676 1242 2678
rect 1308 2676 1500 2678
rect 2076 2676 2268 2678
rect 2334 2676 2526 2678
rect 2592 2676 2784 2678
rect 2850 2676 3042 2678
rect 3108 2676 3300 2678
rect 3876 2676 4068 2678
rect 4134 2676 4326 2678
rect 4392 2676 4584 2678
rect 4650 2676 4842 2678
rect 4908 2676 5100 2678
rect 5676 2676 5868 2678
rect 5934 2676 6126 2678
rect 6192 2676 6384 2678
rect 6450 2676 6642 2678
rect 6708 2676 6900 2678
rect 14676 2676 14868 2678
rect 14934 2676 15126 2678
rect 15192 2676 15384 2678
rect 15450 2676 15642 2678
rect 15708 2676 15900 2678
rect 16476 2676 16668 2678
rect 16734 2676 16926 2678
rect 16992 2676 17184 2678
rect 17250 2676 17442 2678
rect 17508 2676 17700 2678
rect 18276 2676 18468 2678
rect 18534 2676 18726 2678
rect 18792 2676 18984 2678
rect 19050 2676 19242 2678
rect 19308 2676 19500 2678
rect 20076 2676 20268 2678
rect 20334 2676 20526 2678
rect 20592 2676 20784 2678
rect 20850 2676 21042 2678
rect 21108 2676 21300 2678
rect 264 2672 1504 2676
rect 2064 2672 3304 2676
rect 3864 2672 5104 2676
rect 5664 2672 6904 2676
rect 14664 2672 15904 2676
rect 16464 2672 17704 2676
rect 18264 2672 19504 2676
rect 20064 2672 21304 2676
rect 264 2638 288 2672
rect 456 2638 546 2672
rect 714 2638 804 2672
rect 972 2638 1062 2672
rect 1230 2638 1320 2672
rect 1488 2638 1508 2672
rect 264 2564 1508 2638
rect -9024 2372 -8978 2384
rect -8778 2372 -8768 2552
rect -8716 2372 -8706 2552
rect 264 2530 288 2564
rect 456 2530 546 2564
rect 714 2530 804 2564
rect 972 2530 1062 2564
rect 1230 2530 1320 2564
rect 1488 2530 1508 2564
rect 264 2524 1508 2530
rect 2064 2638 2088 2672
rect 2256 2638 2346 2672
rect 2514 2638 2604 2672
rect 2772 2638 2862 2672
rect 3030 2638 3120 2672
rect 3288 2638 3308 2672
rect 2064 2564 3308 2638
rect 2064 2530 2088 2564
rect 2256 2530 2346 2564
rect 2514 2530 2604 2564
rect 2772 2530 2862 2564
rect 3030 2530 3120 2564
rect 3288 2530 3308 2564
rect 2064 2524 3308 2530
rect 3864 2638 3888 2672
rect 4056 2638 4146 2672
rect 4314 2638 4404 2672
rect 4572 2638 4662 2672
rect 4830 2638 4920 2672
rect 5088 2638 5108 2672
rect 3864 2564 5108 2638
rect 3864 2530 3888 2564
rect 4056 2530 4146 2564
rect 4314 2530 4404 2564
rect 4572 2530 4662 2564
rect 4830 2530 4920 2564
rect 5088 2530 5108 2564
rect 3864 2524 5108 2530
rect 5664 2638 5688 2672
rect 5856 2638 5946 2672
rect 6114 2638 6204 2672
rect 6372 2638 6462 2672
rect 6630 2638 6720 2672
rect 6888 2638 6908 2672
rect 5664 2564 6908 2638
rect 5664 2530 5688 2564
rect 5856 2530 5946 2564
rect 6114 2530 6204 2564
rect 6372 2530 6462 2564
rect 6630 2530 6720 2564
rect 6888 2530 6908 2564
rect 5664 2524 6908 2530
rect 14664 2638 14688 2672
rect 14856 2638 14946 2672
rect 15114 2638 15204 2672
rect 15372 2638 15462 2672
rect 15630 2638 15720 2672
rect 15888 2638 15908 2672
rect 14664 2564 15908 2638
rect 14664 2530 14688 2564
rect 14856 2530 14946 2564
rect 15114 2530 15204 2564
rect 15372 2530 15462 2564
rect 15630 2530 15720 2564
rect 15888 2530 15908 2564
rect 14664 2524 15908 2530
rect 16464 2638 16488 2672
rect 16656 2638 16746 2672
rect 16914 2638 17004 2672
rect 17172 2638 17262 2672
rect 17430 2638 17520 2672
rect 17688 2638 17708 2672
rect 16464 2564 17708 2638
rect 16464 2530 16488 2564
rect 16656 2530 16746 2564
rect 16914 2530 17004 2564
rect 17172 2530 17262 2564
rect 17430 2530 17520 2564
rect 17688 2530 17708 2564
rect 16464 2524 17708 2530
rect 18264 2638 18288 2672
rect 18456 2638 18546 2672
rect 18714 2638 18804 2672
rect 18972 2638 19062 2672
rect 19230 2638 19320 2672
rect 19488 2638 19508 2672
rect 18264 2564 19508 2638
rect 18264 2530 18288 2564
rect 18456 2530 18546 2564
rect 18714 2530 18804 2564
rect 18972 2530 19062 2564
rect 19230 2530 19320 2564
rect 19488 2530 19508 2564
rect 18264 2524 19508 2530
rect 20064 2638 20088 2672
rect 20256 2638 20346 2672
rect 20514 2638 20604 2672
rect 20772 2638 20862 2672
rect 21030 2638 21120 2672
rect 21288 2638 21308 2672
rect 20064 2564 21308 2638
rect 20064 2530 20088 2564
rect 20256 2530 20346 2564
rect 20514 2530 20604 2564
rect 20772 2530 20862 2564
rect 21030 2530 21120 2564
rect 21288 2530 21308 2564
rect 20064 2524 21308 2530
rect -10012 2336 -9808 2340
rect -10016 2334 -9808 2336
rect -10016 2300 -9988 2334
rect -9820 2304 -9808 2334
rect -9742 2334 -9292 2340
rect -9742 2304 -9730 2334
rect -9820 2300 -9730 2304
rect -9562 2300 -9472 2334
rect -9304 2304 -9292 2334
rect -9226 2334 -8776 2340
rect -9226 2304 -9214 2334
rect -9304 2300 -9214 2304
rect -9046 2300 -8956 2334
rect -8788 2304 -8776 2334
rect 206 2312 216 2492
rect 268 2312 278 2492
rect 478 2480 524 2492
rect -8788 2300 -8772 2304
rect -10016 2226 -8772 2300
rect -10016 2192 -9988 2226
rect -9820 2192 -9730 2226
rect -9562 2192 -9472 2226
rect -9304 2192 -9214 2226
rect -9046 2192 -8956 2226
rect -8788 2192 -8772 2226
rect -10016 2188 -8772 2192
rect -10000 2186 -9808 2188
rect -9742 2186 -9550 2188
rect -9484 2186 -9292 2188
rect -9226 2186 -9034 2188
rect -8968 2186 -8776 2188
rect -10070 1976 -10060 2156
rect -10008 1976 -9998 2156
rect -9798 2142 -9752 2154
rect -10056 1766 -10050 1976
rect -10016 1766 -10010 1976
rect -9798 1936 -9792 2142
rect -9758 1936 -9752 2142
rect -10056 1754 -10010 1766
rect -9810 1756 -9800 1936
rect -9748 1756 -9738 1936
rect -9798 1754 -9752 1756
rect -9708 1722 -9588 2186
rect -9460 2184 -9316 2186
rect -9554 1976 -9544 2156
rect -9492 1976 -9482 2156
rect -9540 1766 -9534 1976
rect -9500 1766 -9494 1976
rect -9540 1754 -9494 1766
rect -9448 1722 -9328 2184
rect -9282 2142 -9236 2154
rect -9282 1936 -9276 2142
rect -9242 1936 -9236 2142
rect -9294 1756 -9284 1936
rect -9232 1756 -9222 1936
rect -9282 1754 -9236 1756
rect -9188 1722 -9068 2186
rect -9038 1976 -9028 2156
rect -8976 1976 -8966 2156
rect -8766 2142 -8720 2154
rect -9024 1766 -9018 1976
rect -8984 1766 -8978 1976
rect -8766 1936 -8760 2142
rect -8726 1936 -8720 2142
rect 220 2104 226 2312
rect 260 2104 266 2312
rect 478 2272 484 2480
rect 518 2272 524 2480
rect 220 2092 266 2104
rect 466 2092 476 2272
rect 528 2092 538 2272
rect 568 2060 688 2524
rect 722 2312 732 2492
rect 784 2312 794 2492
rect 736 2104 742 2312
rect 776 2104 782 2312
rect 736 2092 782 2104
rect 828 2060 948 2524
rect 994 2480 1040 2492
rect 994 2272 1000 2480
rect 1034 2272 1040 2480
rect 982 2092 992 2272
rect 1044 2092 1054 2272
rect 1088 2060 1208 2524
rect 1238 2312 1248 2492
rect 1300 2312 1310 2492
rect 1510 2480 1556 2492
rect 1252 2104 1258 2312
rect 1292 2104 1298 2312
rect 1510 2272 1516 2480
rect 1550 2272 1556 2480
rect 2006 2312 2016 2492
rect 2068 2312 2078 2492
rect 2278 2480 2324 2492
rect 1252 2092 1298 2104
rect 1498 2092 1508 2272
rect 1560 2092 1570 2272
rect 2020 2104 2026 2312
rect 2060 2104 2066 2312
rect 2278 2272 2284 2480
rect 2318 2272 2324 2480
rect 2020 2092 2066 2104
rect 2266 2092 2276 2272
rect 2328 2092 2338 2272
rect 2368 2060 2488 2524
rect 2522 2312 2532 2492
rect 2584 2312 2594 2492
rect 2536 2104 2542 2312
rect 2576 2104 2582 2312
rect 2536 2092 2582 2104
rect 2628 2060 2748 2524
rect 2794 2480 2840 2492
rect 2794 2272 2800 2480
rect 2834 2272 2840 2480
rect 2782 2092 2792 2272
rect 2844 2092 2854 2272
rect 2888 2060 3008 2524
rect 3038 2312 3048 2492
rect 3100 2312 3110 2492
rect 3310 2480 3356 2492
rect 3052 2104 3058 2312
rect 3092 2104 3098 2312
rect 3310 2272 3316 2480
rect 3350 2272 3356 2480
rect 3806 2312 3816 2492
rect 3868 2312 3878 2492
rect 4078 2480 4124 2492
rect 3052 2092 3098 2104
rect 3298 2092 3308 2272
rect 3360 2092 3370 2272
rect 3820 2104 3826 2312
rect 3860 2104 3866 2312
rect 4078 2272 4084 2480
rect 4118 2272 4124 2480
rect 3820 2092 3866 2104
rect 4066 2092 4076 2272
rect 4128 2092 4138 2272
rect 4168 2060 4288 2524
rect 4322 2312 4332 2492
rect 4384 2312 4394 2492
rect 4336 2104 4342 2312
rect 4376 2104 4382 2312
rect 4336 2092 4382 2104
rect 4428 2060 4548 2524
rect 4594 2480 4640 2492
rect 4594 2272 4600 2480
rect 4634 2272 4640 2480
rect 4582 2092 4592 2272
rect 4644 2092 4654 2272
rect 4688 2060 4808 2524
rect 4838 2312 4848 2492
rect 4900 2312 4910 2492
rect 5110 2480 5156 2492
rect 4852 2104 4858 2312
rect 4892 2104 4898 2312
rect 5110 2272 5116 2480
rect 5150 2272 5156 2480
rect 5606 2312 5616 2492
rect 5668 2312 5678 2492
rect 5878 2480 5924 2492
rect 4852 2092 4898 2104
rect 5098 2092 5108 2272
rect 5160 2092 5170 2272
rect 5620 2104 5626 2312
rect 5660 2104 5666 2312
rect 5878 2272 5884 2480
rect 5918 2272 5924 2480
rect 5620 2092 5666 2104
rect 5866 2092 5876 2272
rect 5928 2092 5938 2272
rect 5968 2060 6088 2524
rect 6122 2312 6132 2492
rect 6184 2312 6194 2492
rect 6136 2104 6142 2312
rect 6176 2104 6182 2312
rect 6136 2092 6182 2104
rect 6228 2060 6348 2524
rect 6394 2480 6440 2492
rect 6394 2272 6400 2480
rect 6434 2272 6440 2480
rect 6382 2092 6392 2272
rect 6444 2092 6454 2272
rect 6488 2060 6608 2524
rect 6638 2312 6648 2492
rect 6700 2312 6710 2492
rect 6910 2480 6956 2492
rect 6652 2104 6658 2312
rect 6692 2104 6698 2312
rect 6910 2272 6916 2480
rect 6950 2272 6956 2480
rect 14606 2312 14616 2492
rect 14668 2312 14678 2492
rect 14878 2480 14924 2492
rect 6652 2092 6698 2104
rect 6898 2092 6908 2272
rect 6960 2092 6970 2272
rect 14620 2104 14626 2312
rect 14660 2104 14666 2312
rect 14878 2272 14884 2480
rect 14918 2272 14924 2480
rect 14620 2092 14666 2104
rect 14866 2092 14876 2272
rect 14928 2092 14938 2272
rect 14968 2060 15088 2524
rect 15122 2312 15132 2492
rect 15184 2312 15194 2492
rect 15136 2104 15142 2312
rect 15176 2104 15182 2312
rect 15136 2092 15182 2104
rect 15228 2060 15348 2524
rect 15394 2480 15440 2492
rect 15394 2272 15400 2480
rect 15434 2272 15440 2480
rect 15382 2092 15392 2272
rect 15444 2092 15454 2272
rect 15488 2060 15608 2524
rect 15638 2312 15648 2492
rect 15700 2312 15710 2492
rect 15910 2480 15956 2492
rect 15652 2104 15658 2312
rect 15692 2104 15698 2312
rect 15910 2272 15916 2480
rect 15950 2272 15956 2480
rect 16406 2312 16416 2492
rect 16468 2312 16478 2492
rect 16678 2480 16724 2492
rect 15652 2092 15698 2104
rect 15898 2092 15908 2272
rect 15960 2092 15970 2272
rect 16420 2104 16426 2312
rect 16460 2104 16466 2312
rect 16678 2272 16684 2480
rect 16718 2272 16724 2480
rect 16420 2092 16466 2104
rect 16666 2092 16676 2272
rect 16728 2092 16738 2272
rect 16768 2060 16888 2524
rect 16922 2312 16932 2492
rect 16984 2312 16994 2492
rect 16936 2104 16942 2312
rect 16976 2104 16982 2312
rect 16936 2092 16982 2104
rect 17028 2060 17148 2524
rect 17194 2480 17240 2492
rect 17194 2272 17200 2480
rect 17234 2272 17240 2480
rect 17182 2092 17192 2272
rect 17244 2092 17254 2272
rect 17288 2060 17408 2524
rect 17438 2312 17448 2492
rect 17500 2312 17510 2492
rect 17710 2480 17756 2492
rect 17452 2104 17458 2312
rect 17492 2104 17498 2312
rect 17710 2272 17716 2480
rect 17750 2272 17756 2480
rect 18206 2312 18216 2492
rect 18268 2312 18278 2492
rect 18478 2480 18524 2492
rect 17452 2092 17498 2104
rect 17698 2092 17708 2272
rect 17760 2092 17770 2272
rect 18220 2104 18226 2312
rect 18260 2104 18266 2312
rect 18478 2272 18484 2480
rect 18518 2272 18524 2480
rect 18220 2092 18266 2104
rect 18466 2092 18476 2272
rect 18528 2092 18538 2272
rect 18568 2060 18688 2524
rect 18722 2312 18732 2492
rect 18784 2312 18794 2492
rect 18736 2104 18742 2312
rect 18776 2104 18782 2312
rect 18736 2092 18782 2104
rect 18828 2060 18948 2524
rect 18994 2480 19040 2492
rect 18994 2272 19000 2480
rect 19034 2272 19040 2480
rect 18982 2092 18992 2272
rect 19044 2092 19054 2272
rect 19088 2060 19208 2524
rect 19238 2312 19248 2492
rect 19300 2312 19310 2492
rect 19510 2480 19556 2492
rect 19252 2104 19258 2312
rect 19292 2104 19298 2312
rect 19510 2272 19516 2480
rect 19550 2272 19556 2480
rect 20006 2312 20016 2492
rect 20068 2312 20078 2492
rect 20278 2480 20324 2492
rect 19252 2092 19298 2104
rect 19498 2092 19508 2272
rect 19560 2092 19570 2272
rect 20020 2104 20026 2312
rect 20060 2104 20066 2312
rect 20278 2272 20284 2480
rect 20318 2272 20324 2480
rect 20020 2092 20066 2104
rect 20266 2092 20276 2272
rect 20328 2092 20338 2272
rect 20368 2060 20488 2524
rect 20522 2312 20532 2492
rect 20584 2312 20594 2492
rect 20536 2104 20542 2312
rect 20576 2104 20582 2312
rect 20536 2092 20582 2104
rect 20628 2060 20748 2524
rect 20794 2480 20840 2492
rect 20794 2272 20800 2480
rect 20834 2272 20840 2480
rect 20782 2092 20792 2272
rect 20844 2092 20854 2272
rect 20888 2060 21008 2524
rect 21038 2312 21048 2492
rect 21100 2312 21110 2492
rect 21310 2480 21356 2492
rect 21052 2104 21058 2312
rect 21092 2104 21098 2312
rect 21310 2272 21316 2480
rect 21350 2272 21356 2480
rect 21052 2092 21098 2104
rect 21298 2092 21308 2272
rect 21360 2092 21370 2272
rect 264 2056 468 2060
rect 260 2054 468 2056
rect 260 2020 288 2054
rect 456 2024 468 2054
rect 534 2054 984 2060
rect 534 2024 546 2054
rect 456 2020 546 2024
rect 714 2020 804 2054
rect 972 2024 984 2054
rect 1050 2054 1500 2060
rect 2064 2056 2268 2060
rect 1050 2024 1062 2054
rect 972 2020 1062 2024
rect 1230 2020 1320 2054
rect 1488 2024 1500 2054
rect 2060 2054 2268 2056
rect 1488 2020 1504 2024
rect 260 1946 1504 2020
rect -9024 1754 -8978 1766
rect -8778 1756 -8768 1936
rect -8716 1756 -8706 1936
rect 260 1912 288 1946
rect 456 1912 546 1946
rect 714 1912 804 1946
rect 972 1912 1062 1946
rect 1230 1912 1320 1946
rect 1488 1912 1504 1946
rect 260 1908 1504 1912
rect 2060 2020 2088 2054
rect 2256 2024 2268 2054
rect 2334 2054 2784 2060
rect 2334 2024 2346 2054
rect 2256 2020 2346 2024
rect 2514 2020 2604 2054
rect 2772 2024 2784 2054
rect 2850 2054 3300 2060
rect 3864 2056 4068 2060
rect 2850 2024 2862 2054
rect 2772 2020 2862 2024
rect 3030 2020 3120 2054
rect 3288 2024 3300 2054
rect 3860 2054 4068 2056
rect 3288 2020 3304 2024
rect 2060 1946 3304 2020
rect 2060 1912 2088 1946
rect 2256 1912 2346 1946
rect 2514 1912 2604 1946
rect 2772 1912 2862 1946
rect 3030 1912 3120 1946
rect 3288 1912 3304 1946
rect 2060 1908 3304 1912
rect 3860 2020 3888 2054
rect 4056 2024 4068 2054
rect 4134 2054 4584 2060
rect 4134 2024 4146 2054
rect 4056 2020 4146 2024
rect 4314 2020 4404 2054
rect 4572 2024 4584 2054
rect 4650 2054 5100 2060
rect 5664 2056 5868 2060
rect 4650 2024 4662 2054
rect 4572 2020 4662 2024
rect 4830 2020 4920 2054
rect 5088 2024 5100 2054
rect 5660 2054 5868 2056
rect 5088 2020 5104 2024
rect 3860 1946 5104 2020
rect 3860 1912 3888 1946
rect 4056 1912 4146 1946
rect 4314 1912 4404 1946
rect 4572 1912 4662 1946
rect 4830 1912 4920 1946
rect 5088 1912 5104 1946
rect 3860 1908 5104 1912
rect 5660 2020 5688 2054
rect 5856 2024 5868 2054
rect 5934 2054 6384 2060
rect 5934 2024 5946 2054
rect 5856 2020 5946 2024
rect 6114 2020 6204 2054
rect 6372 2024 6384 2054
rect 6450 2054 6900 2060
rect 14664 2056 14868 2060
rect 6450 2024 6462 2054
rect 6372 2020 6462 2024
rect 6630 2020 6720 2054
rect 6888 2024 6900 2054
rect 14660 2054 14868 2056
rect 6888 2020 6904 2024
rect 5660 1946 6904 2020
rect 5660 1912 5688 1946
rect 5856 1912 5946 1946
rect 6114 1912 6204 1946
rect 6372 1912 6462 1946
rect 6630 1912 6720 1946
rect 6888 1912 6904 1946
rect 5660 1908 6904 1912
rect 14660 2020 14688 2054
rect 14856 2024 14868 2054
rect 14934 2054 15384 2060
rect 14934 2024 14946 2054
rect 14856 2020 14946 2024
rect 15114 2020 15204 2054
rect 15372 2024 15384 2054
rect 15450 2054 15900 2060
rect 16464 2056 16668 2060
rect 15450 2024 15462 2054
rect 15372 2020 15462 2024
rect 15630 2020 15720 2054
rect 15888 2024 15900 2054
rect 16460 2054 16668 2056
rect 15888 2020 15904 2024
rect 14660 1946 15904 2020
rect 14660 1912 14688 1946
rect 14856 1912 14946 1946
rect 15114 1912 15204 1946
rect 15372 1912 15462 1946
rect 15630 1912 15720 1946
rect 15888 1912 15904 1946
rect 14660 1908 15904 1912
rect 16460 2020 16488 2054
rect 16656 2024 16668 2054
rect 16734 2054 17184 2060
rect 16734 2024 16746 2054
rect 16656 2020 16746 2024
rect 16914 2020 17004 2054
rect 17172 2024 17184 2054
rect 17250 2054 17700 2060
rect 18264 2056 18468 2060
rect 17250 2024 17262 2054
rect 17172 2020 17262 2024
rect 17430 2020 17520 2054
rect 17688 2024 17700 2054
rect 18260 2054 18468 2056
rect 17688 2020 17704 2024
rect 16460 1946 17704 2020
rect 16460 1912 16488 1946
rect 16656 1912 16746 1946
rect 16914 1912 17004 1946
rect 17172 1912 17262 1946
rect 17430 1912 17520 1946
rect 17688 1912 17704 1946
rect 16460 1908 17704 1912
rect 18260 2020 18288 2054
rect 18456 2024 18468 2054
rect 18534 2054 18984 2060
rect 18534 2024 18546 2054
rect 18456 2020 18546 2024
rect 18714 2020 18804 2054
rect 18972 2024 18984 2054
rect 19050 2054 19500 2060
rect 20064 2056 20268 2060
rect 19050 2024 19062 2054
rect 18972 2020 19062 2024
rect 19230 2020 19320 2054
rect 19488 2024 19500 2054
rect 20060 2054 20268 2056
rect 19488 2020 19504 2024
rect 18260 1946 19504 2020
rect 18260 1912 18288 1946
rect 18456 1912 18546 1946
rect 18714 1912 18804 1946
rect 18972 1912 19062 1946
rect 19230 1912 19320 1946
rect 19488 1912 19504 1946
rect 18260 1908 19504 1912
rect 20060 2020 20088 2054
rect 20256 2024 20268 2054
rect 20334 2054 20784 2060
rect 20334 2024 20346 2054
rect 20256 2020 20346 2024
rect 20514 2020 20604 2054
rect 20772 2024 20784 2054
rect 20850 2054 21300 2060
rect 20850 2024 20862 2054
rect 20772 2020 20862 2024
rect 21030 2020 21120 2054
rect 21288 2024 21300 2054
rect 21288 2020 21304 2024
rect 20060 1946 21304 2020
rect 20060 1912 20088 1946
rect 20256 1912 20346 1946
rect 20514 1912 20604 1946
rect 20772 1912 20862 1946
rect 21030 1912 21120 1946
rect 21288 1912 21304 1946
rect 20060 1908 21304 1912
rect 276 1906 468 1908
rect 534 1906 726 1908
rect 792 1906 984 1908
rect 1050 1906 1242 1908
rect 1308 1906 1500 1908
rect 2076 1906 2268 1908
rect 2334 1906 2526 1908
rect 2592 1906 2784 1908
rect 2850 1906 3042 1908
rect 3108 1906 3300 1908
rect 3876 1906 4068 1908
rect 4134 1906 4326 1908
rect 4392 1906 4584 1908
rect 4650 1906 4842 1908
rect 4908 1906 5100 1908
rect 5676 1906 5868 1908
rect 5934 1906 6126 1908
rect 6192 1906 6384 1908
rect 6450 1906 6642 1908
rect 6708 1906 6900 1908
rect 14676 1906 14868 1908
rect 14934 1906 15126 1908
rect 15192 1906 15384 1908
rect 15450 1906 15642 1908
rect 15708 1906 15900 1908
rect 16476 1906 16668 1908
rect 16734 1906 16926 1908
rect 16992 1906 17184 1908
rect 17250 1906 17442 1908
rect 17508 1906 17700 1908
rect 18276 1906 18468 1908
rect 18534 1906 18726 1908
rect 18792 1906 18984 1908
rect 19050 1906 19242 1908
rect 19308 1906 19500 1908
rect 20076 1906 20268 1908
rect 20334 1906 20526 1908
rect 20592 1906 20784 1908
rect 20850 1906 21042 1908
rect 21108 1906 21300 1908
rect -8766 1754 -8720 1756
rect -10000 1720 -9808 1722
rect -9742 1720 -9550 1722
rect -9484 1720 -9292 1722
rect -9226 1720 -9034 1722
rect -8968 1720 -8776 1722
rect -10012 1716 -8772 1720
rect -10012 1682 -9988 1716
rect -9820 1682 -9730 1716
rect -9562 1682 -9472 1716
rect -9304 1682 -9214 1716
rect -9046 1682 -8956 1716
rect -8788 1682 -8768 1716
rect 206 1696 216 1876
rect 268 1696 278 1876
rect 478 1862 524 1874
rect -10012 1608 -8768 1682
rect -10012 1574 -9988 1608
rect -9820 1574 -9730 1608
rect -9562 1574 -9472 1608
rect -9304 1574 -9214 1608
rect -9046 1574 -8956 1608
rect -8788 1574 -8768 1608
rect -10012 1568 -8768 1574
rect -10070 1356 -10060 1536
rect -10008 1356 -9998 1536
rect -9798 1524 -9752 1536
rect -10056 1148 -10050 1356
rect -10016 1148 -10010 1356
rect -9798 1316 -9792 1524
rect -9758 1316 -9752 1524
rect -10056 1136 -10010 1148
rect -9810 1136 -9800 1316
rect -9748 1136 -9738 1316
rect -9708 1104 -9588 1568
rect -9554 1356 -9544 1536
rect -9492 1356 -9482 1536
rect -9540 1148 -9534 1356
rect -9500 1148 -9494 1356
rect -9540 1136 -9494 1148
rect -9448 1104 -9328 1568
rect -9282 1524 -9236 1536
rect -9282 1316 -9276 1524
rect -9242 1316 -9236 1524
rect -9294 1136 -9284 1316
rect -9232 1136 -9222 1316
rect -9188 1104 -9068 1568
rect -9038 1356 -9028 1536
rect -8976 1356 -8966 1536
rect -8766 1524 -8720 1536
rect -9024 1148 -9018 1356
rect -8984 1148 -8978 1356
rect -8766 1316 -8760 1524
rect -8726 1316 -8720 1524
rect 220 1486 226 1696
rect 260 1486 266 1696
rect 478 1656 484 1862
rect 518 1656 524 1862
rect 220 1474 266 1486
rect 466 1476 476 1656
rect 528 1476 538 1656
rect 478 1474 524 1476
rect 568 1442 688 1906
rect 816 1904 960 1906
rect 722 1696 732 1876
rect 784 1696 794 1876
rect 736 1486 742 1696
rect 776 1486 782 1696
rect 736 1474 782 1486
rect 828 1442 948 1904
rect 994 1862 1040 1874
rect 994 1656 1000 1862
rect 1034 1656 1040 1862
rect 982 1476 992 1656
rect 1044 1476 1054 1656
rect 994 1474 1040 1476
rect 1088 1442 1208 1906
rect 1238 1696 1248 1876
rect 1300 1696 1310 1876
rect 1510 1862 1556 1874
rect 1252 1486 1258 1696
rect 1292 1486 1298 1696
rect 1510 1656 1516 1862
rect 1550 1656 1556 1862
rect 2006 1696 2016 1876
rect 2068 1696 2078 1876
rect 2278 1862 2324 1874
rect 1252 1474 1298 1486
rect 1498 1476 1508 1656
rect 1560 1476 1570 1656
rect 2020 1486 2026 1696
rect 2060 1486 2066 1696
rect 2278 1656 2284 1862
rect 2318 1656 2324 1862
rect 1510 1474 1556 1476
rect 2020 1474 2066 1486
rect 2266 1476 2276 1656
rect 2328 1476 2338 1656
rect 2278 1474 2324 1476
rect 2368 1442 2488 1906
rect 2616 1904 2760 1906
rect 2522 1696 2532 1876
rect 2584 1696 2594 1876
rect 2536 1486 2542 1696
rect 2576 1486 2582 1696
rect 2536 1474 2582 1486
rect 2628 1442 2748 1904
rect 2794 1862 2840 1874
rect 2794 1656 2800 1862
rect 2834 1656 2840 1862
rect 2782 1476 2792 1656
rect 2844 1476 2854 1656
rect 2794 1474 2840 1476
rect 2888 1442 3008 1906
rect 3038 1696 3048 1876
rect 3100 1696 3110 1876
rect 3310 1862 3356 1874
rect 3052 1486 3058 1696
rect 3092 1486 3098 1696
rect 3310 1656 3316 1862
rect 3350 1656 3356 1862
rect 3806 1696 3816 1876
rect 3868 1696 3878 1876
rect 4078 1862 4124 1874
rect 3052 1474 3098 1486
rect 3298 1476 3308 1656
rect 3360 1476 3370 1656
rect 3820 1486 3826 1696
rect 3860 1486 3866 1696
rect 4078 1656 4084 1862
rect 4118 1656 4124 1862
rect 3310 1474 3356 1476
rect 3820 1474 3866 1486
rect 4066 1476 4076 1656
rect 4128 1476 4138 1656
rect 4078 1474 4124 1476
rect 4168 1442 4288 1906
rect 4416 1904 4560 1906
rect 4322 1696 4332 1876
rect 4384 1696 4394 1876
rect 4336 1486 4342 1696
rect 4376 1486 4382 1696
rect 4336 1474 4382 1486
rect 4428 1442 4548 1904
rect 4594 1862 4640 1874
rect 4594 1656 4600 1862
rect 4634 1656 4640 1862
rect 4582 1476 4592 1656
rect 4644 1476 4654 1656
rect 4594 1474 4640 1476
rect 4688 1442 4808 1906
rect 4838 1696 4848 1876
rect 4900 1696 4910 1876
rect 5110 1862 5156 1874
rect 4852 1486 4858 1696
rect 4892 1486 4898 1696
rect 5110 1656 5116 1862
rect 5150 1656 5156 1862
rect 5606 1696 5616 1876
rect 5668 1696 5678 1876
rect 5878 1862 5924 1874
rect 4852 1474 4898 1486
rect 5098 1476 5108 1656
rect 5160 1476 5170 1656
rect 5620 1486 5626 1696
rect 5660 1486 5666 1696
rect 5878 1656 5884 1862
rect 5918 1656 5924 1862
rect 5110 1474 5156 1476
rect 5620 1474 5666 1486
rect 5866 1476 5876 1656
rect 5928 1476 5938 1656
rect 5878 1474 5924 1476
rect 5968 1442 6088 1906
rect 6216 1904 6360 1906
rect 6122 1696 6132 1876
rect 6184 1696 6194 1876
rect 6136 1486 6142 1696
rect 6176 1486 6182 1696
rect 6136 1474 6182 1486
rect 6228 1442 6348 1904
rect 6394 1862 6440 1874
rect 6394 1656 6400 1862
rect 6434 1656 6440 1862
rect 6382 1476 6392 1656
rect 6444 1476 6454 1656
rect 6394 1474 6440 1476
rect 6488 1442 6608 1906
rect 6638 1696 6648 1876
rect 6700 1696 6710 1876
rect 6910 1862 6956 1874
rect 6652 1486 6658 1696
rect 6692 1486 6698 1696
rect 6910 1656 6916 1862
rect 6950 1656 6956 1862
rect 14606 1696 14616 1876
rect 14668 1696 14678 1876
rect 14878 1862 14924 1874
rect 6652 1474 6698 1486
rect 6898 1476 6908 1656
rect 6960 1476 6970 1656
rect 14620 1486 14626 1696
rect 14660 1486 14666 1696
rect 14878 1656 14884 1862
rect 14918 1656 14924 1862
rect 6910 1474 6956 1476
rect 14620 1474 14666 1486
rect 14866 1476 14876 1656
rect 14928 1476 14938 1656
rect 14878 1474 14924 1476
rect 14968 1442 15088 1906
rect 15216 1904 15360 1906
rect 15122 1696 15132 1876
rect 15184 1696 15194 1876
rect 15136 1486 15142 1696
rect 15176 1486 15182 1696
rect 15136 1474 15182 1486
rect 15228 1442 15348 1904
rect 15394 1862 15440 1874
rect 15394 1656 15400 1862
rect 15434 1656 15440 1862
rect 15382 1476 15392 1656
rect 15444 1476 15454 1656
rect 15394 1474 15440 1476
rect 15488 1442 15608 1906
rect 15638 1696 15648 1876
rect 15700 1696 15710 1876
rect 15910 1862 15956 1874
rect 15652 1486 15658 1696
rect 15692 1486 15698 1696
rect 15910 1656 15916 1862
rect 15950 1656 15956 1862
rect 16406 1696 16416 1876
rect 16468 1696 16478 1876
rect 16678 1862 16724 1874
rect 15652 1474 15698 1486
rect 15898 1476 15908 1656
rect 15960 1476 15970 1656
rect 16420 1486 16426 1696
rect 16460 1486 16466 1696
rect 16678 1656 16684 1862
rect 16718 1656 16724 1862
rect 15910 1474 15956 1476
rect 16420 1474 16466 1486
rect 16666 1476 16676 1656
rect 16728 1476 16738 1656
rect 16678 1474 16724 1476
rect 16768 1442 16888 1906
rect 17016 1904 17160 1906
rect 16922 1696 16932 1876
rect 16984 1696 16994 1876
rect 16936 1486 16942 1696
rect 16976 1486 16982 1696
rect 16936 1474 16982 1486
rect 17028 1442 17148 1904
rect 17194 1862 17240 1874
rect 17194 1656 17200 1862
rect 17234 1656 17240 1862
rect 17182 1476 17192 1656
rect 17244 1476 17254 1656
rect 17194 1474 17240 1476
rect 17288 1442 17408 1906
rect 17438 1696 17448 1876
rect 17500 1696 17510 1876
rect 17710 1862 17756 1874
rect 17452 1486 17458 1696
rect 17492 1486 17498 1696
rect 17710 1656 17716 1862
rect 17750 1656 17756 1862
rect 18206 1696 18216 1876
rect 18268 1696 18278 1876
rect 18478 1862 18524 1874
rect 17452 1474 17498 1486
rect 17698 1476 17708 1656
rect 17760 1476 17770 1656
rect 18220 1486 18226 1696
rect 18260 1486 18266 1696
rect 18478 1656 18484 1862
rect 18518 1656 18524 1862
rect 17710 1474 17756 1476
rect 18220 1474 18266 1486
rect 18466 1476 18476 1656
rect 18528 1476 18538 1656
rect 18478 1474 18524 1476
rect 18568 1442 18688 1906
rect 18816 1904 18960 1906
rect 18722 1696 18732 1876
rect 18784 1696 18794 1876
rect 18736 1486 18742 1696
rect 18776 1486 18782 1696
rect 18736 1474 18782 1486
rect 18828 1442 18948 1904
rect 18994 1862 19040 1874
rect 18994 1656 19000 1862
rect 19034 1656 19040 1862
rect 18982 1476 18992 1656
rect 19044 1476 19054 1656
rect 18994 1474 19040 1476
rect 19088 1442 19208 1906
rect 19238 1696 19248 1876
rect 19300 1696 19310 1876
rect 19510 1862 19556 1874
rect 19252 1486 19258 1696
rect 19292 1486 19298 1696
rect 19510 1656 19516 1862
rect 19550 1656 19556 1862
rect 20006 1696 20016 1876
rect 20068 1696 20078 1876
rect 20278 1862 20324 1874
rect 19252 1474 19298 1486
rect 19498 1476 19508 1656
rect 19560 1476 19570 1656
rect 20020 1486 20026 1696
rect 20060 1486 20066 1696
rect 20278 1656 20284 1862
rect 20318 1656 20324 1862
rect 19510 1474 19556 1476
rect 20020 1474 20066 1486
rect 20266 1476 20276 1656
rect 20328 1476 20338 1656
rect 20278 1474 20324 1476
rect 20368 1442 20488 1906
rect 20616 1904 20760 1906
rect 20522 1696 20532 1876
rect 20584 1696 20594 1876
rect 20536 1486 20542 1696
rect 20576 1486 20582 1696
rect 20536 1474 20582 1486
rect 20628 1442 20748 1904
rect 20794 1862 20840 1874
rect 20794 1656 20800 1862
rect 20834 1656 20840 1862
rect 20782 1476 20792 1656
rect 20844 1476 20854 1656
rect 20794 1474 20840 1476
rect 20888 1442 21008 1906
rect 21038 1696 21048 1876
rect 21100 1696 21110 1876
rect 21310 1862 21356 1874
rect 21052 1486 21058 1696
rect 21092 1486 21098 1696
rect 21310 1656 21316 1862
rect 21350 1656 21356 1862
rect 21052 1474 21098 1486
rect 21298 1476 21308 1656
rect 21360 1476 21370 1656
rect 21310 1474 21356 1476
rect 276 1440 468 1442
rect 534 1440 726 1442
rect 792 1440 984 1442
rect 1050 1440 1242 1442
rect 1308 1440 1500 1442
rect 2076 1440 2268 1442
rect 2334 1440 2526 1442
rect 2592 1440 2784 1442
rect 2850 1440 3042 1442
rect 3108 1440 3300 1442
rect 3876 1440 4068 1442
rect 4134 1440 4326 1442
rect 4392 1440 4584 1442
rect 4650 1440 4842 1442
rect 4908 1440 5100 1442
rect 5676 1440 5868 1442
rect 5934 1440 6126 1442
rect 6192 1440 6384 1442
rect 6450 1440 6642 1442
rect 6708 1440 6900 1442
rect 14676 1440 14868 1442
rect 14934 1440 15126 1442
rect 15192 1440 15384 1442
rect 15450 1440 15642 1442
rect 15708 1440 15900 1442
rect 16476 1440 16668 1442
rect 16734 1440 16926 1442
rect 16992 1440 17184 1442
rect 17250 1440 17442 1442
rect 17508 1440 17700 1442
rect 18276 1440 18468 1442
rect 18534 1440 18726 1442
rect 18792 1440 18984 1442
rect 19050 1440 19242 1442
rect 19308 1440 19500 1442
rect 20076 1440 20268 1442
rect 20334 1440 20526 1442
rect 20592 1440 20784 1442
rect 20850 1440 21042 1442
rect 21108 1440 21300 1442
rect 264 1436 1504 1440
rect 2064 1436 3304 1440
rect 3864 1436 5104 1440
rect 5664 1436 6904 1440
rect 14664 1436 15904 1440
rect 16464 1436 17704 1440
rect 18264 1436 19504 1440
rect 20064 1436 21304 1440
rect 264 1402 288 1436
rect 456 1402 546 1436
rect 714 1402 804 1436
rect 972 1402 1062 1436
rect 1230 1402 1320 1436
rect 1488 1402 1508 1436
rect 264 1328 1508 1402
rect -9024 1136 -8978 1148
rect -8778 1136 -8768 1316
rect -8716 1136 -8706 1316
rect 264 1294 288 1328
rect 456 1294 546 1328
rect 714 1294 804 1328
rect 972 1294 1062 1328
rect 1230 1294 1320 1328
rect 1488 1294 1508 1328
rect 264 1288 1508 1294
rect 2064 1402 2088 1436
rect 2256 1402 2346 1436
rect 2514 1402 2604 1436
rect 2772 1402 2862 1436
rect 3030 1402 3120 1436
rect 3288 1402 3308 1436
rect 2064 1328 3308 1402
rect 2064 1294 2088 1328
rect 2256 1294 2346 1328
rect 2514 1294 2604 1328
rect 2772 1294 2862 1328
rect 3030 1294 3120 1328
rect 3288 1294 3308 1328
rect 2064 1288 3308 1294
rect 3864 1402 3888 1436
rect 4056 1402 4146 1436
rect 4314 1402 4404 1436
rect 4572 1402 4662 1436
rect 4830 1402 4920 1436
rect 5088 1402 5108 1436
rect 3864 1328 5108 1402
rect 3864 1294 3888 1328
rect 4056 1294 4146 1328
rect 4314 1294 4404 1328
rect 4572 1294 4662 1328
rect 4830 1294 4920 1328
rect 5088 1294 5108 1328
rect 3864 1288 5108 1294
rect 5664 1402 5688 1436
rect 5856 1402 5946 1436
rect 6114 1402 6204 1436
rect 6372 1402 6462 1436
rect 6630 1402 6720 1436
rect 6888 1402 6908 1436
rect 5664 1328 6908 1402
rect 5664 1294 5688 1328
rect 5856 1294 5946 1328
rect 6114 1294 6204 1328
rect 6372 1294 6462 1328
rect 6630 1294 6720 1328
rect 6888 1294 6908 1328
rect 5664 1288 6908 1294
rect 14664 1402 14688 1436
rect 14856 1402 14946 1436
rect 15114 1402 15204 1436
rect 15372 1402 15462 1436
rect 15630 1402 15720 1436
rect 15888 1402 15908 1436
rect 14664 1328 15908 1402
rect 14664 1294 14688 1328
rect 14856 1294 14946 1328
rect 15114 1294 15204 1328
rect 15372 1294 15462 1328
rect 15630 1294 15720 1328
rect 15888 1294 15908 1328
rect 14664 1288 15908 1294
rect 16464 1402 16488 1436
rect 16656 1402 16746 1436
rect 16914 1402 17004 1436
rect 17172 1402 17262 1436
rect 17430 1402 17520 1436
rect 17688 1402 17708 1436
rect 16464 1328 17708 1402
rect 16464 1294 16488 1328
rect 16656 1294 16746 1328
rect 16914 1294 17004 1328
rect 17172 1294 17262 1328
rect 17430 1294 17520 1328
rect 17688 1294 17708 1328
rect 16464 1288 17708 1294
rect 18264 1402 18288 1436
rect 18456 1402 18546 1436
rect 18714 1402 18804 1436
rect 18972 1402 19062 1436
rect 19230 1402 19320 1436
rect 19488 1402 19508 1436
rect 18264 1328 19508 1402
rect 18264 1294 18288 1328
rect 18456 1294 18546 1328
rect 18714 1294 18804 1328
rect 18972 1294 19062 1328
rect 19230 1294 19320 1328
rect 19488 1294 19508 1328
rect 18264 1288 19508 1294
rect 20064 1402 20088 1436
rect 20256 1402 20346 1436
rect 20514 1402 20604 1436
rect 20772 1402 20862 1436
rect 21030 1402 21120 1436
rect 21288 1402 21308 1436
rect 20064 1328 21308 1402
rect 20064 1294 20088 1328
rect 20256 1294 20346 1328
rect 20514 1294 20604 1328
rect 20772 1294 20862 1328
rect 21030 1294 21120 1328
rect 21288 1294 21308 1328
rect 20064 1288 21308 1294
rect -10012 1098 -9808 1104
rect -10012 1064 -9988 1098
rect -9820 1088 -9808 1098
rect -9742 1098 -9292 1104
rect -9742 1088 -9730 1098
rect -9820 1064 -9730 1088
rect -9562 1064 -9472 1098
rect -9304 1088 -9292 1098
rect -9226 1098 -8776 1104
rect -9226 1088 -9214 1098
rect -9304 1064 -9214 1088
rect -9046 1064 -8956 1098
rect -8788 1088 -8776 1098
rect -8788 1064 -8768 1088
rect 206 1076 216 1256
rect 268 1076 278 1256
rect 478 1244 524 1256
rect -10012 990 -8768 1064
rect -10012 956 -9988 990
rect -9820 956 -9730 990
rect -9562 956 -9472 990
rect -9304 956 -9214 990
rect -9046 956 -8956 990
rect -8788 956 -8768 990
rect -10012 952 -8768 956
rect -10000 950 -9808 952
rect -9742 950 -9550 952
rect -9484 950 -9292 952
rect -9226 950 -9034 952
rect -8968 950 -8776 952
rect -10070 740 -10060 920
rect -10008 740 -9998 920
rect -9798 906 -9752 918
rect -10056 530 -10050 740
rect -10016 530 -10010 740
rect -9798 700 -9792 906
rect -9758 700 -9752 906
rect -10056 518 -10010 530
rect -9810 520 -9800 700
rect -9748 520 -9738 700
rect -9798 518 -9752 520
rect -9708 488 -9588 950
rect -9554 740 -9544 920
rect -9492 740 -9482 920
rect -9540 530 -9534 740
rect -9500 530 -9494 740
rect -9540 518 -9494 530
rect -9448 488 -9328 950
rect -9282 906 -9236 918
rect -9282 700 -9276 906
rect -9242 700 -9236 906
rect -9294 520 -9284 700
rect -9232 520 -9222 700
rect -9282 518 -9236 520
rect -9188 488 -9068 950
rect -9038 740 -9028 920
rect -8976 740 -8966 920
rect -8766 906 -8720 918
rect -9024 530 -9018 740
rect -8984 530 -8978 740
rect -8766 700 -8760 906
rect -8726 700 -8720 906
rect 220 868 226 1076
rect 260 868 266 1076
rect 478 1036 484 1244
rect 518 1036 524 1244
rect 220 856 266 868
rect 466 856 476 1036
rect 528 856 538 1036
rect 568 824 688 1288
rect 722 1076 732 1256
rect 784 1076 794 1256
rect 736 868 742 1076
rect 776 868 782 1076
rect 736 856 782 868
rect 828 824 948 1288
rect 994 1244 1040 1256
rect 994 1036 1000 1244
rect 1034 1036 1040 1244
rect 982 856 992 1036
rect 1044 856 1054 1036
rect 1088 824 1208 1288
rect 1238 1076 1248 1256
rect 1300 1076 1310 1256
rect 1510 1244 1556 1256
rect 1252 868 1258 1076
rect 1292 868 1298 1076
rect 1510 1036 1516 1244
rect 1550 1036 1556 1244
rect 2006 1076 2016 1256
rect 2068 1076 2078 1256
rect 2278 1244 2324 1256
rect 1252 856 1298 868
rect 1498 856 1508 1036
rect 1560 856 1570 1036
rect 2020 868 2026 1076
rect 2060 868 2066 1076
rect 2278 1036 2284 1244
rect 2318 1036 2324 1244
rect 2020 856 2066 868
rect 2266 856 2276 1036
rect 2328 856 2338 1036
rect 2368 824 2488 1288
rect 2522 1076 2532 1256
rect 2584 1076 2594 1256
rect 2536 868 2542 1076
rect 2576 868 2582 1076
rect 2536 856 2582 868
rect 2628 824 2748 1288
rect 2794 1244 2840 1256
rect 2794 1036 2800 1244
rect 2834 1036 2840 1244
rect 2782 856 2792 1036
rect 2844 856 2854 1036
rect 2888 824 3008 1288
rect 3038 1076 3048 1256
rect 3100 1076 3110 1256
rect 3310 1244 3356 1256
rect 3052 868 3058 1076
rect 3092 868 3098 1076
rect 3310 1036 3316 1244
rect 3350 1036 3356 1244
rect 3806 1076 3816 1256
rect 3868 1076 3878 1256
rect 4078 1244 4124 1256
rect 3052 856 3098 868
rect 3298 856 3308 1036
rect 3360 856 3370 1036
rect 3820 868 3826 1076
rect 3860 868 3866 1076
rect 4078 1036 4084 1244
rect 4118 1036 4124 1244
rect 3820 856 3866 868
rect 4066 856 4076 1036
rect 4128 856 4138 1036
rect 4168 824 4288 1288
rect 4322 1076 4332 1256
rect 4384 1076 4394 1256
rect 4336 868 4342 1076
rect 4376 868 4382 1076
rect 4336 856 4382 868
rect 4428 824 4548 1288
rect 4594 1244 4640 1256
rect 4594 1036 4600 1244
rect 4634 1036 4640 1244
rect 4582 856 4592 1036
rect 4644 856 4654 1036
rect 4688 824 4808 1288
rect 4838 1076 4848 1256
rect 4900 1076 4910 1256
rect 5110 1244 5156 1256
rect 4852 868 4858 1076
rect 4892 868 4898 1076
rect 5110 1036 5116 1244
rect 5150 1036 5156 1244
rect 5606 1076 5616 1256
rect 5668 1076 5678 1256
rect 5878 1244 5924 1256
rect 4852 856 4898 868
rect 5098 856 5108 1036
rect 5160 856 5170 1036
rect 5620 868 5626 1076
rect 5660 868 5666 1076
rect 5878 1036 5884 1244
rect 5918 1036 5924 1244
rect 5620 856 5666 868
rect 5866 856 5876 1036
rect 5928 856 5938 1036
rect 5968 824 6088 1288
rect 6122 1076 6132 1256
rect 6184 1076 6194 1256
rect 6136 868 6142 1076
rect 6176 868 6182 1076
rect 6136 856 6182 868
rect 6228 824 6348 1288
rect 6394 1244 6440 1256
rect 6394 1036 6400 1244
rect 6434 1036 6440 1244
rect 6382 856 6392 1036
rect 6444 856 6454 1036
rect 6488 824 6608 1288
rect 6638 1076 6648 1256
rect 6700 1076 6710 1256
rect 6910 1244 6956 1256
rect 6652 868 6658 1076
rect 6692 868 6698 1076
rect 6910 1036 6916 1244
rect 6950 1036 6956 1244
rect 14606 1076 14616 1256
rect 14668 1076 14678 1256
rect 14878 1244 14924 1256
rect 6652 856 6698 868
rect 6898 856 6908 1036
rect 6960 856 6970 1036
rect 14620 868 14626 1076
rect 14660 868 14666 1076
rect 14878 1036 14884 1244
rect 14918 1036 14924 1244
rect 14620 856 14666 868
rect 14866 856 14876 1036
rect 14928 856 14938 1036
rect 14968 824 15088 1288
rect 15122 1076 15132 1256
rect 15184 1076 15194 1256
rect 15136 868 15142 1076
rect 15176 868 15182 1076
rect 15136 856 15182 868
rect 15228 824 15348 1288
rect 15394 1244 15440 1256
rect 15394 1036 15400 1244
rect 15434 1036 15440 1244
rect 15382 856 15392 1036
rect 15444 856 15454 1036
rect 15488 824 15608 1288
rect 15638 1076 15648 1256
rect 15700 1076 15710 1256
rect 15910 1244 15956 1256
rect 15652 868 15658 1076
rect 15692 868 15698 1076
rect 15910 1036 15916 1244
rect 15950 1036 15956 1244
rect 16406 1076 16416 1256
rect 16468 1076 16478 1256
rect 16678 1244 16724 1256
rect 15652 856 15698 868
rect 15898 856 15908 1036
rect 15960 856 15970 1036
rect 16420 868 16426 1076
rect 16460 868 16466 1076
rect 16678 1036 16684 1244
rect 16718 1036 16724 1244
rect 16420 856 16466 868
rect 16666 856 16676 1036
rect 16728 856 16738 1036
rect 16768 824 16888 1288
rect 16922 1076 16932 1256
rect 16984 1076 16994 1256
rect 16936 868 16942 1076
rect 16976 868 16982 1076
rect 16936 856 16982 868
rect 17028 824 17148 1288
rect 17194 1244 17240 1256
rect 17194 1036 17200 1244
rect 17234 1036 17240 1244
rect 17182 856 17192 1036
rect 17244 856 17254 1036
rect 17288 824 17408 1288
rect 17438 1076 17448 1256
rect 17500 1076 17510 1256
rect 17710 1244 17756 1256
rect 17452 868 17458 1076
rect 17492 868 17498 1076
rect 17710 1036 17716 1244
rect 17750 1036 17756 1244
rect 18206 1076 18216 1256
rect 18268 1076 18278 1256
rect 18478 1244 18524 1256
rect 17452 856 17498 868
rect 17698 856 17708 1036
rect 17760 856 17770 1036
rect 18220 868 18226 1076
rect 18260 868 18266 1076
rect 18478 1036 18484 1244
rect 18518 1036 18524 1244
rect 18220 856 18266 868
rect 18466 856 18476 1036
rect 18528 856 18538 1036
rect 18568 824 18688 1288
rect 18722 1076 18732 1256
rect 18784 1076 18794 1256
rect 18736 868 18742 1076
rect 18776 868 18782 1076
rect 18736 856 18782 868
rect 18828 824 18948 1288
rect 18994 1244 19040 1256
rect 18994 1036 19000 1244
rect 19034 1036 19040 1244
rect 18982 856 18992 1036
rect 19044 856 19054 1036
rect 19088 824 19208 1288
rect 19238 1076 19248 1256
rect 19300 1076 19310 1256
rect 19510 1244 19556 1256
rect 19252 868 19258 1076
rect 19292 868 19298 1076
rect 19510 1036 19516 1244
rect 19550 1036 19556 1244
rect 20006 1076 20016 1256
rect 20068 1076 20078 1256
rect 20278 1244 20324 1256
rect 19252 856 19298 868
rect 19498 856 19508 1036
rect 19560 856 19570 1036
rect 20020 868 20026 1076
rect 20060 868 20066 1076
rect 20278 1036 20284 1244
rect 20318 1036 20324 1244
rect 20020 856 20066 868
rect 20266 856 20276 1036
rect 20328 856 20338 1036
rect 20368 824 20488 1288
rect 20522 1076 20532 1256
rect 20584 1076 20594 1256
rect 20536 868 20542 1076
rect 20576 868 20582 1076
rect 20536 856 20582 868
rect 20628 824 20748 1288
rect 20794 1244 20840 1256
rect 20794 1036 20800 1244
rect 20834 1036 20840 1244
rect 20782 856 20792 1036
rect 20844 856 20854 1036
rect 20888 824 21008 1288
rect 21038 1076 21048 1256
rect 21100 1076 21110 1256
rect 21310 1244 21356 1256
rect 21052 868 21058 1076
rect 21092 868 21098 1076
rect 21310 1036 21316 1244
rect 21350 1036 21356 1244
rect 21052 856 21098 868
rect 21298 856 21308 1036
rect 21360 856 21370 1036
rect 264 818 468 824
rect 264 784 288 818
rect 456 808 468 818
rect 534 818 984 824
rect 534 808 546 818
rect 456 784 546 808
rect 714 784 804 818
rect 972 808 984 818
rect 1050 818 1500 824
rect 1050 808 1062 818
rect 972 784 1062 808
rect 1230 784 1320 818
rect 1488 808 1500 818
rect 2064 818 2268 824
rect 1488 784 1508 808
rect 264 710 1508 784
rect -9024 518 -8978 530
rect -8778 520 -8768 700
rect -8716 520 -8706 700
rect 264 676 288 710
rect 456 676 546 710
rect 714 676 804 710
rect 972 676 1062 710
rect 1230 676 1320 710
rect 1488 676 1508 710
rect 264 672 1508 676
rect 2064 784 2088 818
rect 2256 808 2268 818
rect 2334 818 2784 824
rect 2334 808 2346 818
rect 2256 784 2346 808
rect 2514 784 2604 818
rect 2772 808 2784 818
rect 2850 818 3300 824
rect 2850 808 2862 818
rect 2772 784 2862 808
rect 3030 784 3120 818
rect 3288 808 3300 818
rect 3864 818 4068 824
rect 3288 784 3308 808
rect 2064 710 3308 784
rect 2064 676 2088 710
rect 2256 676 2346 710
rect 2514 676 2604 710
rect 2772 676 2862 710
rect 3030 676 3120 710
rect 3288 676 3308 710
rect 2064 672 3308 676
rect 3864 784 3888 818
rect 4056 808 4068 818
rect 4134 818 4584 824
rect 4134 808 4146 818
rect 4056 784 4146 808
rect 4314 784 4404 818
rect 4572 808 4584 818
rect 4650 818 5100 824
rect 4650 808 4662 818
rect 4572 784 4662 808
rect 4830 784 4920 818
rect 5088 808 5100 818
rect 5664 818 5868 824
rect 5088 784 5108 808
rect 3864 710 5108 784
rect 3864 676 3888 710
rect 4056 676 4146 710
rect 4314 676 4404 710
rect 4572 676 4662 710
rect 4830 676 4920 710
rect 5088 676 5108 710
rect 3864 672 5108 676
rect 5664 784 5688 818
rect 5856 808 5868 818
rect 5934 818 6384 824
rect 5934 808 5946 818
rect 5856 784 5946 808
rect 6114 784 6204 818
rect 6372 808 6384 818
rect 6450 818 6900 824
rect 6450 808 6462 818
rect 6372 784 6462 808
rect 6630 784 6720 818
rect 6888 808 6900 818
rect 14664 818 14868 824
rect 6888 784 6908 808
rect 5664 710 6908 784
rect 5664 676 5688 710
rect 5856 676 5946 710
rect 6114 676 6204 710
rect 6372 676 6462 710
rect 6630 676 6720 710
rect 6888 676 6908 710
rect 5664 672 6908 676
rect 14664 784 14688 818
rect 14856 808 14868 818
rect 14934 818 15384 824
rect 14934 808 14946 818
rect 14856 784 14946 808
rect 15114 784 15204 818
rect 15372 808 15384 818
rect 15450 818 15900 824
rect 15450 808 15462 818
rect 15372 784 15462 808
rect 15630 784 15720 818
rect 15888 808 15900 818
rect 16464 818 16668 824
rect 15888 784 15908 808
rect 14664 710 15908 784
rect 14664 676 14688 710
rect 14856 676 14946 710
rect 15114 676 15204 710
rect 15372 676 15462 710
rect 15630 676 15720 710
rect 15888 676 15908 710
rect 14664 672 15908 676
rect 16464 784 16488 818
rect 16656 808 16668 818
rect 16734 818 17184 824
rect 16734 808 16746 818
rect 16656 784 16746 808
rect 16914 784 17004 818
rect 17172 808 17184 818
rect 17250 818 17700 824
rect 17250 808 17262 818
rect 17172 784 17262 808
rect 17430 784 17520 818
rect 17688 808 17700 818
rect 18264 818 18468 824
rect 17688 784 17708 808
rect 16464 710 17708 784
rect 16464 676 16488 710
rect 16656 676 16746 710
rect 16914 676 17004 710
rect 17172 676 17262 710
rect 17430 676 17520 710
rect 17688 676 17708 710
rect 16464 672 17708 676
rect 18264 784 18288 818
rect 18456 808 18468 818
rect 18534 818 18984 824
rect 18534 808 18546 818
rect 18456 784 18546 808
rect 18714 784 18804 818
rect 18972 808 18984 818
rect 19050 818 19500 824
rect 19050 808 19062 818
rect 18972 784 19062 808
rect 19230 784 19320 818
rect 19488 808 19500 818
rect 20064 818 20268 824
rect 19488 784 19508 808
rect 18264 710 19508 784
rect 18264 676 18288 710
rect 18456 676 18546 710
rect 18714 676 18804 710
rect 18972 676 19062 710
rect 19230 676 19320 710
rect 19488 676 19508 710
rect 18264 672 19508 676
rect 20064 784 20088 818
rect 20256 808 20268 818
rect 20334 818 20784 824
rect 20334 808 20346 818
rect 20256 784 20346 808
rect 20514 784 20604 818
rect 20772 808 20784 818
rect 20850 818 21300 824
rect 20850 808 20862 818
rect 20772 784 20862 808
rect 21030 784 21120 818
rect 21288 808 21300 818
rect 21288 784 21308 808
rect 20064 710 21308 784
rect 20064 676 20088 710
rect 20256 676 20346 710
rect 20514 676 20604 710
rect 20772 676 20862 710
rect 21030 676 21120 710
rect 21288 676 21308 710
rect 20064 672 21308 676
rect 276 670 468 672
rect 534 670 726 672
rect 792 670 984 672
rect 1050 670 1242 672
rect 1308 670 1500 672
rect 2076 670 2268 672
rect 2334 670 2526 672
rect 2592 670 2784 672
rect 2850 670 3042 672
rect 3108 670 3300 672
rect 3876 670 4068 672
rect 4134 670 4326 672
rect 4392 670 4584 672
rect 4650 670 4842 672
rect 4908 670 5100 672
rect 5676 670 5868 672
rect 5934 670 6126 672
rect 6192 670 6384 672
rect 6450 670 6642 672
rect 6708 670 6900 672
rect 14676 670 14868 672
rect 14934 670 15126 672
rect 15192 670 15384 672
rect 15450 670 15642 672
rect 15708 670 15900 672
rect 16476 670 16668 672
rect 16734 670 16926 672
rect 16992 670 17184 672
rect 17250 670 17442 672
rect 17508 670 17700 672
rect 18276 670 18468 672
rect 18534 670 18726 672
rect 18792 670 18984 672
rect 19050 670 19242 672
rect 19308 670 19500 672
rect 20076 670 20268 672
rect 20334 670 20526 672
rect 20592 670 20784 672
rect 20850 670 21042 672
rect 21108 670 21300 672
rect -8766 518 -8720 520
rect -8506 508 -8354 520
rect -10012 480 -8772 488
rect -10012 446 -9988 480
rect -9820 446 -9730 480
rect -9562 446 -9472 480
rect -9304 446 -9214 480
rect -9046 446 -8956 480
rect -8788 446 -8772 480
rect -10012 428 -8772 446
rect -8510 348 -8500 508
rect -8360 348 -8350 508
rect 206 460 216 640
rect 268 460 278 640
rect 478 626 524 638
rect -8506 336 -8354 348
rect 220 250 226 460
rect 260 250 266 460
rect 478 420 484 626
rect 518 420 524 626
rect 220 238 266 250
rect 466 240 476 420
rect 528 240 538 420
rect 478 238 524 240
rect 568 208 688 670
rect 722 460 732 640
rect 784 460 794 640
rect 736 250 742 460
rect 776 250 782 460
rect 736 238 782 250
rect 828 208 948 670
rect 994 626 1040 638
rect 994 420 1000 626
rect 1034 420 1040 626
rect 982 240 992 420
rect 1044 240 1054 420
rect 994 238 1040 240
rect 1088 208 1208 670
rect 1238 460 1248 640
rect 1300 460 1310 640
rect 1510 626 1556 638
rect 1252 250 1258 460
rect 1292 250 1298 460
rect 1510 420 1516 626
rect 1550 420 1556 626
rect 2006 460 2016 640
rect 2068 460 2078 640
rect 2278 626 2324 638
rect 1252 238 1298 250
rect 1498 240 1508 420
rect 1560 240 1570 420
rect 1690 268 1882 280
rect 1510 238 1556 240
rect 264 200 1504 208
rect 264 166 288 200
rect 456 166 546 200
rect 714 166 804 200
rect 972 166 1062 200
rect 1230 166 1320 200
rect 1488 166 1504 200
rect 264 148 1504 166
rect 1686 68 1696 268
rect 1876 68 1886 268
rect 2020 250 2026 460
rect 2060 250 2066 460
rect 2278 420 2284 626
rect 2318 420 2324 626
rect 2020 238 2066 250
rect 2266 240 2276 420
rect 2328 240 2338 420
rect 2278 238 2324 240
rect 2368 208 2488 670
rect 2522 460 2532 640
rect 2584 460 2594 640
rect 2536 250 2542 460
rect 2576 250 2582 460
rect 2536 238 2582 250
rect 2628 208 2748 670
rect 2794 626 2840 638
rect 2794 420 2800 626
rect 2834 420 2840 626
rect 2782 240 2792 420
rect 2844 240 2854 420
rect 2794 238 2840 240
rect 2888 208 3008 670
rect 3038 460 3048 640
rect 3100 460 3110 640
rect 3310 626 3356 638
rect 3052 250 3058 460
rect 3092 250 3098 460
rect 3310 420 3316 626
rect 3350 420 3356 626
rect 3806 460 3816 640
rect 3868 460 3878 640
rect 4078 626 4124 638
rect 3052 238 3098 250
rect 3298 240 3308 420
rect 3360 240 3370 420
rect 3506 276 3698 288
rect 3310 238 3356 240
rect 2064 200 3304 208
rect 2064 166 2088 200
rect 2256 166 2346 200
rect 2514 166 2604 200
rect 2772 166 2862 200
rect 3030 166 3120 200
rect 3288 166 3304 200
rect 2064 148 3304 166
rect 1690 56 1882 68
rect 3502 64 3512 276
rect 3692 64 3702 276
rect 3820 250 3826 460
rect 3860 250 3866 460
rect 4078 420 4084 626
rect 4118 420 4124 626
rect 3820 238 3866 250
rect 4066 240 4076 420
rect 4128 240 4138 420
rect 4078 238 4124 240
rect 4168 208 4288 670
rect 4322 460 4332 640
rect 4384 460 4394 640
rect 4336 250 4342 460
rect 4376 250 4382 460
rect 4336 238 4382 250
rect 4428 208 4548 670
rect 4594 626 4640 638
rect 4594 420 4600 626
rect 4634 420 4640 626
rect 4582 240 4592 420
rect 4644 240 4654 420
rect 4594 238 4640 240
rect 4688 208 4808 670
rect 4838 460 4848 640
rect 4900 460 4910 640
rect 5110 626 5156 638
rect 4852 250 4858 460
rect 4892 250 4898 460
rect 5110 420 5116 626
rect 5150 420 5156 626
rect 5606 460 5616 640
rect 5668 460 5678 640
rect 5878 626 5924 638
rect 4852 238 4898 250
rect 5098 240 5108 420
rect 5160 240 5170 420
rect 5282 276 5474 288
rect 5110 238 5156 240
rect 3864 200 5104 208
rect 3864 166 3888 200
rect 4056 166 4146 200
rect 4314 166 4404 200
rect 4572 166 4662 200
rect 4830 166 4920 200
rect 5088 166 5104 200
rect 3864 148 5104 166
rect 5278 64 5288 276
rect 5468 64 5478 276
rect 5620 250 5626 460
rect 5660 250 5666 460
rect 5878 420 5884 626
rect 5918 420 5924 626
rect 5620 238 5666 250
rect 5866 240 5876 420
rect 5928 240 5938 420
rect 5878 238 5924 240
rect 5968 208 6088 670
rect 6122 460 6132 640
rect 6184 460 6194 640
rect 6136 250 6142 460
rect 6176 250 6182 460
rect 6136 238 6182 250
rect 6228 208 6348 670
rect 6394 626 6440 638
rect 6394 420 6400 626
rect 6434 420 6440 626
rect 6382 240 6392 420
rect 6444 240 6454 420
rect 6394 238 6440 240
rect 6488 208 6608 670
rect 6638 460 6648 640
rect 6700 460 6710 640
rect 6910 626 6956 638
rect 6652 250 6658 460
rect 6692 250 6698 460
rect 6910 420 6916 626
rect 6950 420 6956 626
rect 14606 460 14616 640
rect 14668 460 14678 640
rect 14878 626 14924 638
rect 6652 238 6698 250
rect 6898 240 6908 420
rect 6960 240 6970 420
rect 14620 250 14626 460
rect 14660 250 14666 460
rect 14878 420 14884 626
rect 14918 420 14924 626
rect 6910 238 6956 240
rect 14620 238 14666 250
rect 14866 240 14876 420
rect 14928 240 14938 420
rect 14878 238 14924 240
rect 14968 208 15088 670
rect 15122 460 15132 640
rect 15184 460 15194 640
rect 15136 250 15142 460
rect 15176 250 15182 460
rect 15136 238 15182 250
rect 15228 208 15348 670
rect 15394 626 15440 638
rect 15394 420 15400 626
rect 15434 420 15440 626
rect 15382 240 15392 420
rect 15444 240 15454 420
rect 15394 238 15440 240
rect 15488 208 15608 670
rect 15638 460 15648 640
rect 15700 460 15710 640
rect 15910 626 15956 638
rect 15652 250 15658 460
rect 15692 250 15698 460
rect 15910 420 15916 626
rect 15950 420 15956 626
rect 16406 460 16416 640
rect 16468 460 16478 640
rect 16678 626 16724 638
rect 15652 238 15698 250
rect 15898 240 15908 420
rect 15960 240 15970 420
rect 16090 268 16282 280
rect 15910 238 15956 240
rect 5664 200 6904 208
rect 5664 166 5688 200
rect 5856 166 5946 200
rect 6114 166 6204 200
rect 6372 166 6462 200
rect 6630 166 6720 200
rect 6888 166 6904 200
rect 5664 148 6904 166
rect 14664 200 15904 208
rect 14664 166 14688 200
rect 14856 166 14946 200
rect 15114 166 15204 200
rect 15372 166 15462 200
rect 15630 166 15720 200
rect 15888 166 15904 200
rect 14664 148 15904 166
rect 16086 68 16096 268
rect 16276 68 16286 268
rect 16420 250 16426 460
rect 16460 250 16466 460
rect 16678 420 16684 626
rect 16718 420 16724 626
rect 16420 238 16466 250
rect 16666 240 16676 420
rect 16728 240 16738 420
rect 16678 238 16724 240
rect 16768 208 16888 670
rect 16922 460 16932 640
rect 16984 460 16994 640
rect 16936 250 16942 460
rect 16976 250 16982 460
rect 16936 238 16982 250
rect 17028 208 17148 670
rect 17194 626 17240 638
rect 17194 420 17200 626
rect 17234 420 17240 626
rect 17182 240 17192 420
rect 17244 240 17254 420
rect 17194 238 17240 240
rect 17288 208 17408 670
rect 17438 460 17448 640
rect 17500 460 17510 640
rect 17710 626 17756 638
rect 17452 250 17458 460
rect 17492 250 17498 460
rect 17710 420 17716 626
rect 17750 420 17756 626
rect 18206 460 18216 640
rect 18268 460 18278 640
rect 18478 626 18524 638
rect 17452 238 17498 250
rect 17698 240 17708 420
rect 17760 240 17770 420
rect 17906 276 18098 288
rect 17710 238 17756 240
rect 16464 200 17704 208
rect 16464 166 16488 200
rect 16656 166 16746 200
rect 16914 166 17004 200
rect 17172 166 17262 200
rect 17430 166 17520 200
rect 17688 166 17704 200
rect 16464 148 17704 166
rect 3506 52 3698 64
rect 5282 52 5474 64
rect 16090 56 16282 68
rect 17902 64 17912 276
rect 18092 64 18102 276
rect 18220 250 18226 460
rect 18260 250 18266 460
rect 18478 420 18484 626
rect 18518 420 18524 626
rect 18220 238 18266 250
rect 18466 240 18476 420
rect 18528 240 18538 420
rect 18478 238 18524 240
rect 18568 208 18688 670
rect 18722 460 18732 640
rect 18784 460 18794 640
rect 18736 250 18742 460
rect 18776 250 18782 460
rect 18736 238 18782 250
rect 18828 208 18948 670
rect 18994 626 19040 638
rect 18994 420 19000 626
rect 19034 420 19040 626
rect 18982 240 18992 420
rect 19044 240 19054 420
rect 18994 238 19040 240
rect 19088 208 19208 670
rect 19238 460 19248 640
rect 19300 460 19310 640
rect 19510 626 19556 638
rect 19252 250 19258 460
rect 19292 250 19298 460
rect 19510 420 19516 626
rect 19550 420 19556 626
rect 20006 460 20016 640
rect 20068 460 20078 640
rect 20278 626 20324 638
rect 19252 238 19298 250
rect 19498 240 19508 420
rect 19560 240 19570 420
rect 19682 276 19874 288
rect 19510 238 19556 240
rect 18264 200 19504 208
rect 18264 166 18288 200
rect 18456 166 18546 200
rect 18714 166 18804 200
rect 18972 166 19062 200
rect 19230 166 19320 200
rect 19488 166 19504 200
rect 18264 148 19504 166
rect 19678 64 19688 276
rect 19868 64 19878 276
rect 20020 250 20026 460
rect 20060 250 20066 460
rect 20278 420 20284 626
rect 20318 420 20324 626
rect 20020 238 20066 250
rect 20266 240 20276 420
rect 20328 240 20338 420
rect 20278 238 20324 240
rect 20368 208 20488 670
rect 20522 460 20532 640
rect 20584 460 20594 640
rect 20536 250 20542 460
rect 20576 250 20582 460
rect 20536 238 20582 250
rect 20628 208 20748 670
rect 20794 626 20840 638
rect 20794 420 20800 626
rect 20834 420 20840 626
rect 20782 240 20792 420
rect 20844 240 20854 420
rect 20794 238 20840 240
rect 20888 208 21008 670
rect 21038 460 21048 640
rect 21100 460 21110 640
rect 21310 626 21356 638
rect 21052 250 21058 460
rect 21092 250 21098 460
rect 21310 420 21316 626
rect 21350 420 21356 626
rect 21052 238 21098 250
rect 21298 240 21308 420
rect 21360 240 21370 420
rect 21310 238 21356 240
rect 20064 200 21304 208
rect 20064 166 20088 200
rect 20256 166 20346 200
rect 20514 166 20604 200
rect 20772 166 20862 200
rect 21030 166 21120 200
rect 21288 166 21304 200
rect 20064 148 21304 166
rect 17906 52 18098 64
rect 19682 52 19874 64
rect -2778 -1188 -2768 -382
rect -1960 -1188 -1950 -382
rect 11622 -1188 11632 -382
rect 12440 -1188 12450 -382
<< via1 >>
rect 7440 27336 7540 27436
rect 6632 27075 6696 27092
rect 6632 26912 6648 27075
rect 6648 26912 6682 27075
rect 6682 26912 6696 27075
rect 6476 26699 6490 26868
rect 6490 26699 6524 26868
rect 6524 26699 6540 26868
rect 6476 26688 6540 26699
rect 6948 27075 7012 27092
rect 6948 26912 6964 27075
rect 6964 26912 6998 27075
rect 6998 26912 7012 27075
rect 6792 26699 6806 26868
rect 6806 26699 6840 26868
rect 6840 26699 6856 26868
rect 6792 26688 6856 26699
rect 7264 27075 7328 27092
rect 7264 26912 7280 27075
rect 7280 26912 7314 27075
rect 7314 26912 7328 27075
rect 7108 26699 7122 26868
rect 7122 26699 7156 26868
rect 7156 26699 7172 26868
rect 7108 26688 7172 26699
rect 7580 27075 7644 27092
rect 7580 26912 7596 27075
rect 7596 26912 7630 27075
rect 7630 26912 7644 27075
rect 7424 26699 7438 26868
rect 7438 26699 7472 26868
rect 7472 26699 7488 26868
rect 7424 26688 7488 26699
rect 7896 27075 7960 27092
rect 7896 26912 7912 27075
rect 7912 26912 7946 27075
rect 7946 26912 7960 27075
rect 7740 26699 7754 26868
rect 7754 26699 7788 26868
rect 7788 26699 7804 26868
rect 7740 26688 7804 26699
rect 8056 26699 8070 26868
rect 8070 26699 8104 26868
rect 8104 26699 8120 26868
rect 8056 26688 8120 26699
rect 8852 27075 8916 27092
rect 8852 26912 8868 27075
rect 8868 26912 8902 27075
rect 8902 26912 8916 27075
rect 8696 26699 8710 26868
rect 8710 26699 8744 26868
rect 8744 26699 8760 26868
rect 8696 26688 8760 26699
rect 9168 27075 9232 27092
rect 9168 26912 9184 27075
rect 9184 26912 9218 27075
rect 9218 26912 9232 27075
rect 9012 26699 9026 26868
rect 9026 26699 9060 26868
rect 9060 26699 9076 26868
rect 9012 26688 9076 26699
rect 9484 27075 9548 27092
rect 9484 26912 9500 27075
rect 9500 26912 9534 27075
rect 9534 26912 9548 27075
rect 9328 26699 9342 26868
rect 9342 26699 9376 26868
rect 9376 26699 9392 26868
rect 9328 26688 9392 26699
rect 9800 27075 9864 27092
rect 9800 26912 9816 27075
rect 9816 26912 9850 27075
rect 9850 26912 9864 27075
rect 9644 26699 9658 26868
rect 9658 26699 9692 26868
rect 9692 26699 9708 26868
rect 9644 26688 9708 26699
rect 10116 27075 10180 27092
rect 10116 26912 10132 27075
rect 10132 26912 10166 27075
rect 10166 26912 10180 27075
rect 9960 26699 9974 26868
rect 9974 26699 10008 26868
rect 10008 26699 10024 26868
rect 9960 26688 10024 26699
rect 10276 26699 10290 26868
rect 10290 26699 10324 26868
rect 10324 26699 10340 26868
rect 10276 26688 10340 26699
rect 11032 27075 11096 27092
rect 11032 26912 11048 27075
rect 11048 26912 11082 27075
rect 11082 26912 11096 27075
rect 10876 26699 10890 26868
rect 10890 26699 10924 26868
rect 10924 26699 10940 26868
rect 10876 26688 10940 26699
rect 11348 27075 11412 27092
rect 11348 26912 11364 27075
rect 11364 26912 11398 27075
rect 11398 26912 11412 27075
rect 11192 26699 11206 26868
rect 11206 26699 11240 26868
rect 11240 26699 11256 26868
rect 11192 26688 11256 26699
rect 11664 27075 11728 27092
rect 11664 26912 11680 27075
rect 11680 26912 11714 27075
rect 11714 26912 11728 27075
rect 11508 26699 11522 26868
rect 11522 26699 11556 26868
rect 11556 26699 11572 26868
rect 11508 26688 11572 26699
rect 11980 27075 12044 27092
rect 11980 26912 11996 27075
rect 11996 26912 12030 27075
rect 12030 26912 12044 27075
rect 11824 26699 11838 26868
rect 11838 26699 11872 26868
rect 11872 26699 11888 26868
rect 11824 26688 11888 26699
rect 12296 27075 12360 27092
rect 12296 26912 12312 27075
rect 12312 26912 12346 27075
rect 12346 26912 12360 27075
rect 12140 26699 12154 26868
rect 12154 26699 12188 26868
rect 12188 26699 12204 26868
rect 12140 26688 12204 26699
rect 12456 26699 12470 26868
rect 12470 26699 12504 26868
rect 12504 26699 12520 26868
rect 12456 26688 12520 26699
rect 13212 27075 13276 27092
rect 13212 26912 13228 27075
rect 13228 26912 13262 27075
rect 13262 26912 13276 27075
rect 13056 26699 13070 26868
rect 13070 26699 13104 26868
rect 13104 26699 13120 26868
rect 13056 26688 13120 26699
rect 13528 27075 13592 27092
rect 13528 26912 13544 27075
rect 13544 26912 13578 27075
rect 13578 26912 13592 27075
rect 13372 26699 13386 26868
rect 13386 26699 13420 26868
rect 13420 26699 13436 26868
rect 13372 26688 13436 26699
rect 13844 27075 13908 27092
rect 13844 26912 13860 27075
rect 13860 26912 13894 27075
rect 13894 26912 13908 27075
rect 13688 26699 13702 26868
rect 13702 26699 13736 26868
rect 13736 26699 13752 26868
rect 13688 26688 13752 26699
rect 14160 27075 14224 27092
rect 14160 26912 14176 27075
rect 14176 26912 14210 27075
rect 14210 26912 14224 27075
rect 14004 26699 14018 26868
rect 14018 26699 14052 26868
rect 14052 26699 14068 26868
rect 14004 26688 14068 26699
rect 14476 27075 14540 27092
rect 14476 26912 14492 27075
rect 14492 26912 14526 27075
rect 14526 26912 14540 27075
rect 14320 26699 14334 26868
rect 14334 26699 14368 26868
rect 14368 26699 14384 26868
rect 14320 26688 14384 26699
rect 14636 26699 14650 26868
rect 14650 26699 14684 26868
rect 14684 26699 14700 26868
rect 14636 26688 14700 26699
rect 15412 27075 15476 27092
rect 15412 26912 15428 27075
rect 15428 26912 15462 27075
rect 15462 26912 15476 27075
rect 15256 26699 15270 26868
rect 15270 26699 15304 26868
rect 15304 26699 15320 26868
rect 15256 26688 15320 26699
rect 15728 27075 15792 27092
rect 15728 26912 15744 27075
rect 15744 26912 15778 27075
rect 15778 26912 15792 27075
rect 15572 26699 15586 26868
rect 15586 26699 15620 26868
rect 15620 26699 15636 26868
rect 15572 26688 15636 26699
rect 16044 27075 16108 27092
rect 16044 26912 16060 27075
rect 16060 26912 16094 27075
rect 16094 26912 16108 27075
rect 15888 26699 15902 26868
rect 15902 26699 15936 26868
rect 15936 26699 15952 26868
rect 15888 26688 15952 26699
rect 16360 27075 16424 27092
rect 16360 26912 16376 27075
rect 16376 26912 16410 27075
rect 16410 26912 16424 27075
rect 16204 26699 16218 26868
rect 16218 26699 16252 26868
rect 16252 26699 16268 26868
rect 16204 26688 16268 26699
rect 16676 27075 16740 27092
rect 16676 26912 16692 27075
rect 16692 26912 16726 27075
rect 16726 26912 16740 27075
rect 16520 26699 16534 26868
rect 16534 26699 16568 26868
rect 16568 26699 16584 26868
rect 16520 26688 16584 26699
rect 16836 26699 16850 26868
rect 16850 26699 16884 26868
rect 16884 26699 16900 26868
rect 16836 26688 16900 26699
rect 6632 26439 6696 26456
rect 6632 26276 6648 26439
rect 6648 26276 6682 26439
rect 6682 26276 6696 26439
rect 6476 26063 6490 26232
rect 6490 26063 6524 26232
rect 6524 26063 6540 26232
rect 6476 26052 6540 26063
rect 6948 26439 7012 26456
rect 6948 26276 6964 26439
rect 6964 26276 6998 26439
rect 6998 26276 7012 26439
rect 6792 26063 6806 26232
rect 6806 26063 6840 26232
rect 6840 26063 6856 26232
rect 6792 26052 6856 26063
rect 7264 26439 7328 26456
rect 7264 26276 7280 26439
rect 7280 26276 7314 26439
rect 7314 26276 7328 26439
rect 7108 26063 7122 26232
rect 7122 26063 7156 26232
rect 7156 26063 7172 26232
rect 7108 26052 7172 26063
rect 7580 26439 7644 26456
rect 7580 26276 7596 26439
rect 7596 26276 7630 26439
rect 7630 26276 7644 26439
rect 7424 26063 7438 26232
rect 7438 26063 7472 26232
rect 7472 26063 7488 26232
rect 7424 26052 7488 26063
rect 7896 26439 7960 26456
rect 7896 26276 7912 26439
rect 7912 26276 7946 26439
rect 7946 26276 7960 26439
rect 7740 26063 7754 26232
rect 7754 26063 7788 26232
rect 7788 26063 7804 26232
rect 7740 26052 7804 26063
rect 8056 26063 8070 26232
rect 8070 26063 8104 26232
rect 8104 26063 8120 26232
rect 8056 26052 8120 26063
rect 8852 26439 8916 26456
rect 8852 26276 8868 26439
rect 8868 26276 8902 26439
rect 8902 26276 8916 26439
rect 8696 26063 8710 26232
rect 8710 26063 8744 26232
rect 8744 26063 8760 26232
rect 8696 26052 8760 26063
rect 9168 26439 9232 26456
rect 9168 26276 9184 26439
rect 9184 26276 9218 26439
rect 9218 26276 9232 26439
rect 9012 26063 9026 26232
rect 9026 26063 9060 26232
rect 9060 26063 9076 26232
rect 9012 26052 9076 26063
rect 9484 26439 9548 26456
rect 9484 26276 9500 26439
rect 9500 26276 9534 26439
rect 9534 26276 9548 26439
rect 9328 26063 9342 26232
rect 9342 26063 9376 26232
rect 9376 26063 9392 26232
rect 9328 26052 9392 26063
rect 9800 26439 9864 26456
rect 9800 26276 9816 26439
rect 9816 26276 9850 26439
rect 9850 26276 9864 26439
rect 9644 26063 9658 26232
rect 9658 26063 9692 26232
rect 9692 26063 9708 26232
rect 9644 26052 9708 26063
rect 10116 26439 10180 26456
rect 10116 26276 10132 26439
rect 10132 26276 10166 26439
rect 10166 26276 10180 26439
rect 9960 26063 9974 26232
rect 9974 26063 10008 26232
rect 10008 26063 10024 26232
rect 9960 26052 10024 26063
rect 10276 26063 10290 26232
rect 10290 26063 10324 26232
rect 10324 26063 10340 26232
rect 10276 26052 10340 26063
rect 11032 26439 11096 26456
rect 11032 26276 11048 26439
rect 11048 26276 11082 26439
rect 11082 26276 11096 26439
rect 10876 26063 10890 26232
rect 10890 26063 10924 26232
rect 10924 26063 10940 26232
rect 10876 26052 10940 26063
rect 11348 26439 11412 26456
rect 11348 26276 11364 26439
rect 11364 26276 11398 26439
rect 11398 26276 11412 26439
rect 11192 26063 11206 26232
rect 11206 26063 11240 26232
rect 11240 26063 11256 26232
rect 11192 26052 11256 26063
rect 11664 26439 11728 26456
rect 11664 26276 11680 26439
rect 11680 26276 11714 26439
rect 11714 26276 11728 26439
rect 11508 26063 11522 26232
rect 11522 26063 11556 26232
rect 11556 26063 11572 26232
rect 11508 26052 11572 26063
rect 11980 26439 12044 26456
rect 11980 26276 11996 26439
rect 11996 26276 12030 26439
rect 12030 26276 12044 26439
rect 11824 26063 11838 26232
rect 11838 26063 11872 26232
rect 11872 26063 11888 26232
rect 11824 26052 11888 26063
rect 12296 26439 12360 26456
rect 12296 26276 12312 26439
rect 12312 26276 12346 26439
rect 12346 26276 12360 26439
rect 12140 26063 12154 26232
rect 12154 26063 12188 26232
rect 12188 26063 12204 26232
rect 12140 26052 12204 26063
rect 12456 26063 12470 26232
rect 12470 26063 12504 26232
rect 12504 26063 12520 26232
rect 12456 26052 12520 26063
rect 13212 26439 13276 26456
rect 13212 26276 13228 26439
rect 13228 26276 13262 26439
rect 13262 26276 13276 26439
rect 13056 26063 13070 26232
rect 13070 26063 13104 26232
rect 13104 26063 13120 26232
rect 13056 26052 13120 26063
rect 13528 26439 13592 26456
rect 13528 26276 13544 26439
rect 13544 26276 13578 26439
rect 13578 26276 13592 26439
rect 13372 26063 13386 26232
rect 13386 26063 13420 26232
rect 13420 26063 13436 26232
rect 13372 26052 13436 26063
rect 13844 26439 13908 26456
rect 13844 26276 13860 26439
rect 13860 26276 13894 26439
rect 13894 26276 13908 26439
rect 13688 26063 13702 26232
rect 13702 26063 13736 26232
rect 13736 26063 13752 26232
rect 13688 26052 13752 26063
rect 14160 26439 14224 26456
rect 14160 26276 14176 26439
rect 14176 26276 14210 26439
rect 14210 26276 14224 26439
rect 14004 26063 14018 26232
rect 14018 26063 14052 26232
rect 14052 26063 14068 26232
rect 14004 26052 14068 26063
rect 14476 26439 14540 26456
rect 14476 26276 14492 26439
rect 14492 26276 14526 26439
rect 14526 26276 14540 26439
rect 14320 26063 14334 26232
rect 14334 26063 14368 26232
rect 14368 26063 14384 26232
rect 14320 26052 14384 26063
rect 14636 26063 14650 26232
rect 14650 26063 14684 26232
rect 14684 26063 14700 26232
rect 14636 26052 14700 26063
rect 15412 26439 15476 26456
rect 15412 26276 15428 26439
rect 15428 26276 15462 26439
rect 15462 26276 15476 26439
rect 15256 26063 15270 26232
rect 15270 26063 15304 26232
rect 15304 26063 15320 26232
rect 15256 26052 15320 26063
rect 15728 26439 15792 26456
rect 15728 26276 15744 26439
rect 15744 26276 15778 26439
rect 15778 26276 15792 26439
rect 15572 26063 15586 26232
rect 15586 26063 15620 26232
rect 15620 26063 15636 26232
rect 15572 26052 15636 26063
rect 16044 26439 16108 26456
rect 16044 26276 16060 26439
rect 16060 26276 16094 26439
rect 16094 26276 16108 26439
rect 15888 26063 15902 26232
rect 15902 26063 15936 26232
rect 15936 26063 15952 26232
rect 15888 26052 15952 26063
rect 16360 26439 16424 26456
rect 16360 26276 16376 26439
rect 16376 26276 16410 26439
rect 16410 26276 16424 26439
rect 16204 26063 16218 26232
rect 16218 26063 16252 26232
rect 16252 26063 16268 26232
rect 16204 26052 16268 26063
rect 16676 26439 16740 26456
rect 16676 26276 16692 26439
rect 16692 26276 16726 26439
rect 16726 26276 16740 26439
rect 16520 26063 16534 26232
rect 16534 26063 16568 26232
rect 16568 26063 16584 26232
rect 16520 26052 16584 26063
rect 16836 26063 16850 26232
rect 16850 26063 16884 26232
rect 16884 26063 16900 26232
rect 16836 26052 16900 26063
rect 6632 25803 6696 25816
rect 6632 25636 6648 25803
rect 6648 25636 6682 25803
rect 6682 25636 6696 25803
rect 6476 25427 6490 25592
rect 6490 25427 6524 25592
rect 6524 25427 6540 25592
rect 6476 25412 6540 25427
rect 6948 25803 7012 25816
rect 6948 25636 6964 25803
rect 6964 25636 6998 25803
rect 6998 25636 7012 25803
rect 6792 25427 6806 25592
rect 6806 25427 6840 25592
rect 6840 25427 6856 25592
rect 6792 25412 6856 25427
rect 7264 25803 7328 25816
rect 7264 25636 7280 25803
rect 7280 25636 7314 25803
rect 7314 25636 7328 25803
rect 7108 25427 7122 25592
rect 7122 25427 7156 25592
rect 7156 25427 7172 25592
rect 7108 25412 7172 25427
rect 7580 25803 7644 25816
rect 7580 25636 7596 25803
rect 7596 25636 7630 25803
rect 7630 25636 7644 25803
rect 7424 25427 7438 25592
rect 7438 25427 7472 25592
rect 7472 25427 7488 25592
rect 7424 25412 7488 25427
rect 7896 25803 7960 25816
rect 7896 25636 7912 25803
rect 7912 25636 7946 25803
rect 7946 25636 7960 25803
rect 7740 25427 7754 25592
rect 7754 25427 7788 25592
rect 7788 25427 7804 25592
rect 7740 25412 7804 25427
rect 8056 25427 8070 25592
rect 8070 25427 8104 25592
rect 8104 25427 8120 25592
rect 8056 25412 8120 25427
rect 8852 25803 8916 25816
rect 8852 25636 8868 25803
rect 8868 25636 8902 25803
rect 8902 25636 8916 25803
rect 8696 25427 8710 25592
rect 8710 25427 8744 25592
rect 8744 25427 8760 25592
rect 8696 25412 8760 25427
rect 9168 25803 9232 25816
rect 9168 25636 9184 25803
rect 9184 25636 9218 25803
rect 9218 25636 9232 25803
rect 9012 25427 9026 25592
rect 9026 25427 9060 25592
rect 9060 25427 9076 25592
rect 9012 25412 9076 25427
rect 9484 25803 9548 25816
rect 9484 25636 9500 25803
rect 9500 25636 9534 25803
rect 9534 25636 9548 25803
rect 9328 25427 9342 25592
rect 9342 25427 9376 25592
rect 9376 25427 9392 25592
rect 9328 25412 9392 25427
rect 9800 25803 9864 25816
rect 9800 25636 9816 25803
rect 9816 25636 9850 25803
rect 9850 25636 9864 25803
rect 9644 25427 9658 25592
rect 9658 25427 9692 25592
rect 9692 25427 9708 25592
rect 9644 25412 9708 25427
rect 10116 25803 10180 25816
rect 10116 25636 10132 25803
rect 10132 25636 10166 25803
rect 10166 25636 10180 25803
rect 9960 25427 9974 25592
rect 9974 25427 10008 25592
rect 10008 25427 10024 25592
rect 9960 25412 10024 25427
rect 10276 25427 10290 25592
rect 10290 25427 10324 25592
rect 10324 25427 10340 25592
rect 10276 25412 10340 25427
rect 11032 25803 11096 25816
rect 11032 25636 11048 25803
rect 11048 25636 11082 25803
rect 11082 25636 11096 25803
rect 10876 25427 10890 25592
rect 10890 25427 10924 25592
rect 10924 25427 10940 25592
rect 10876 25412 10940 25427
rect 11348 25803 11412 25816
rect 11348 25636 11364 25803
rect 11364 25636 11398 25803
rect 11398 25636 11412 25803
rect 11192 25427 11206 25592
rect 11206 25427 11240 25592
rect 11240 25427 11256 25592
rect 11192 25412 11256 25427
rect 11664 25803 11728 25816
rect 11664 25636 11680 25803
rect 11680 25636 11714 25803
rect 11714 25636 11728 25803
rect 11508 25427 11522 25592
rect 11522 25427 11556 25592
rect 11556 25427 11572 25592
rect 11508 25412 11572 25427
rect 11980 25803 12044 25816
rect 11980 25636 11996 25803
rect 11996 25636 12030 25803
rect 12030 25636 12044 25803
rect 11824 25427 11838 25592
rect 11838 25427 11872 25592
rect 11872 25427 11888 25592
rect 11824 25412 11888 25427
rect 12296 25803 12360 25816
rect 12296 25636 12312 25803
rect 12312 25636 12346 25803
rect 12346 25636 12360 25803
rect 12140 25427 12154 25592
rect 12154 25427 12188 25592
rect 12188 25427 12204 25592
rect 12140 25412 12204 25427
rect 12456 25427 12470 25592
rect 12470 25427 12504 25592
rect 12504 25427 12520 25592
rect 12456 25412 12520 25427
rect 13212 25803 13276 25816
rect 13212 25636 13228 25803
rect 13228 25636 13262 25803
rect 13262 25636 13276 25803
rect 13056 25427 13070 25592
rect 13070 25427 13104 25592
rect 13104 25427 13120 25592
rect 13056 25412 13120 25427
rect 13528 25803 13592 25816
rect 13528 25636 13544 25803
rect 13544 25636 13578 25803
rect 13578 25636 13592 25803
rect 13372 25427 13386 25592
rect 13386 25427 13420 25592
rect 13420 25427 13436 25592
rect 13372 25412 13436 25427
rect 13844 25803 13908 25816
rect 13844 25636 13860 25803
rect 13860 25636 13894 25803
rect 13894 25636 13908 25803
rect 13688 25427 13702 25592
rect 13702 25427 13736 25592
rect 13736 25427 13752 25592
rect 13688 25412 13752 25427
rect 14160 25803 14224 25816
rect 14160 25636 14176 25803
rect 14176 25636 14210 25803
rect 14210 25636 14224 25803
rect 14004 25427 14018 25592
rect 14018 25427 14052 25592
rect 14052 25427 14068 25592
rect 14004 25412 14068 25427
rect 14476 25803 14540 25816
rect 14476 25636 14492 25803
rect 14492 25636 14526 25803
rect 14526 25636 14540 25803
rect 14320 25427 14334 25592
rect 14334 25427 14368 25592
rect 14368 25427 14384 25592
rect 14320 25412 14384 25427
rect 14636 25427 14650 25592
rect 14650 25427 14684 25592
rect 14684 25427 14700 25592
rect 14636 25412 14700 25427
rect 15412 25803 15476 25816
rect 15412 25636 15428 25803
rect 15428 25636 15462 25803
rect 15462 25636 15476 25803
rect 15256 25427 15270 25592
rect 15270 25427 15304 25592
rect 15304 25427 15320 25592
rect 15256 25412 15320 25427
rect 15728 25803 15792 25816
rect 15728 25636 15744 25803
rect 15744 25636 15778 25803
rect 15778 25636 15792 25803
rect 15572 25427 15586 25592
rect 15586 25427 15620 25592
rect 15620 25427 15636 25592
rect 15572 25412 15636 25427
rect 16044 25803 16108 25816
rect 16044 25636 16060 25803
rect 16060 25636 16094 25803
rect 16094 25636 16108 25803
rect 15888 25427 15902 25592
rect 15902 25427 15936 25592
rect 15936 25427 15952 25592
rect 15888 25412 15952 25427
rect 16360 25803 16424 25816
rect 16360 25636 16376 25803
rect 16376 25636 16410 25803
rect 16410 25636 16424 25803
rect 16204 25427 16218 25592
rect 16218 25427 16252 25592
rect 16252 25427 16268 25592
rect 16204 25412 16268 25427
rect 16676 25803 16740 25816
rect 16676 25636 16692 25803
rect 16692 25636 16726 25803
rect 16726 25636 16740 25803
rect 16520 25427 16534 25592
rect 16534 25427 16568 25592
rect 16568 25427 16584 25592
rect 16520 25412 16584 25427
rect 16836 25427 16850 25592
rect 16850 25427 16884 25592
rect 16884 25427 16900 25592
rect 16836 25412 16900 25427
rect 6572 24979 6636 24992
rect 6572 24812 6586 24979
rect 6586 24812 6620 24979
rect 6620 24812 6636 24979
rect 6476 24603 6490 24768
rect 6490 24603 6524 24768
rect 6524 24603 6540 24768
rect 6476 24588 6540 24603
rect 6764 24979 6828 24992
rect 6764 24812 6778 24979
rect 6778 24812 6812 24979
rect 6812 24812 6828 24979
rect 6664 24603 6682 24768
rect 6682 24603 6716 24768
rect 6716 24603 6728 24768
rect 6664 24588 6728 24603
rect 6956 24979 7020 24992
rect 6956 24812 6970 24979
rect 6970 24812 7004 24979
rect 7004 24812 7020 24979
rect 6856 24603 6874 24768
rect 6874 24603 6908 24768
rect 6908 24603 6920 24768
rect 6856 24588 6920 24603
rect 7148 24979 7212 24992
rect 7148 24812 7162 24979
rect 7162 24812 7196 24979
rect 7196 24812 7212 24979
rect 7052 24603 7066 24768
rect 7066 24603 7100 24768
rect 7100 24603 7116 24768
rect 7052 24588 7116 24603
rect 7340 24979 7404 24992
rect 7340 24812 7354 24979
rect 7354 24812 7388 24979
rect 7388 24812 7404 24979
rect 7244 24603 7258 24768
rect 7258 24603 7292 24768
rect 7292 24603 7308 24768
rect 7244 24588 7308 24603
rect 7532 24979 7596 24992
rect 7532 24812 7546 24979
rect 7546 24812 7580 24979
rect 7580 24812 7596 24979
rect 7436 24603 7450 24768
rect 7450 24603 7484 24768
rect 7484 24603 7500 24768
rect 7436 24588 7500 24603
rect 7724 24979 7788 24992
rect 7724 24812 7738 24979
rect 7738 24812 7772 24979
rect 7772 24812 7788 24979
rect 7628 24603 7642 24768
rect 7642 24603 7676 24768
rect 7676 24603 7692 24768
rect 7628 24588 7692 24603
rect 7916 24979 7980 24992
rect 7916 24812 7930 24979
rect 7930 24812 7964 24979
rect 7964 24812 7980 24979
rect 7820 24603 7834 24768
rect 7834 24603 7868 24768
rect 7868 24603 7884 24768
rect 7820 24588 7884 24603
rect 8792 24979 8856 24992
rect 8792 24812 8806 24979
rect 8806 24812 8840 24979
rect 8840 24812 8856 24979
rect 8696 24603 8710 24768
rect 8710 24603 8744 24768
rect 8744 24603 8760 24768
rect 8696 24588 8760 24603
rect 8984 24979 9048 24992
rect 8984 24812 8998 24979
rect 8998 24812 9032 24979
rect 9032 24812 9048 24979
rect 8884 24603 8902 24768
rect 8902 24603 8936 24768
rect 8936 24603 8948 24768
rect 8884 24588 8948 24603
rect 9176 24979 9240 24992
rect 9176 24812 9190 24979
rect 9190 24812 9224 24979
rect 9224 24812 9240 24979
rect 9076 24603 9094 24768
rect 9094 24603 9128 24768
rect 9128 24603 9140 24768
rect 9076 24588 9140 24603
rect 9368 24979 9432 24992
rect 9368 24812 9382 24979
rect 9382 24812 9416 24979
rect 9416 24812 9432 24979
rect 9272 24603 9286 24768
rect 9286 24603 9320 24768
rect 9320 24603 9336 24768
rect 9272 24588 9336 24603
rect 9560 24979 9624 24992
rect 9560 24812 9574 24979
rect 9574 24812 9608 24979
rect 9608 24812 9624 24979
rect 9464 24603 9478 24768
rect 9478 24603 9512 24768
rect 9512 24603 9528 24768
rect 9464 24588 9528 24603
rect 9752 24979 9816 24992
rect 9752 24812 9766 24979
rect 9766 24812 9800 24979
rect 9800 24812 9816 24979
rect 9656 24603 9670 24768
rect 9670 24603 9704 24768
rect 9704 24603 9720 24768
rect 9656 24588 9720 24603
rect 9944 24979 10008 24992
rect 9944 24812 9958 24979
rect 9958 24812 9992 24979
rect 9992 24812 10008 24979
rect 9848 24603 9862 24768
rect 9862 24603 9896 24768
rect 9896 24603 9912 24768
rect 9848 24588 9912 24603
rect 10136 24979 10200 24992
rect 10136 24812 10150 24979
rect 10150 24812 10184 24979
rect 10184 24812 10200 24979
rect 10040 24603 10054 24768
rect 10054 24603 10088 24768
rect 10088 24603 10104 24768
rect 10040 24588 10104 24603
rect 10972 24979 11036 24992
rect 10972 24812 10986 24979
rect 10986 24812 11020 24979
rect 11020 24812 11036 24979
rect 10876 24603 10890 24768
rect 10890 24603 10924 24768
rect 10924 24603 10940 24768
rect 10876 24588 10940 24603
rect 11164 24979 11228 24992
rect 11164 24812 11178 24979
rect 11178 24812 11212 24979
rect 11212 24812 11228 24979
rect 11064 24603 11082 24768
rect 11082 24603 11116 24768
rect 11116 24603 11128 24768
rect 11064 24588 11128 24603
rect 11356 24979 11420 24992
rect 11356 24812 11370 24979
rect 11370 24812 11404 24979
rect 11404 24812 11420 24979
rect 11256 24603 11274 24768
rect 11274 24603 11308 24768
rect 11308 24603 11320 24768
rect 11256 24588 11320 24603
rect 11548 24979 11612 24992
rect 11548 24812 11562 24979
rect 11562 24812 11596 24979
rect 11596 24812 11612 24979
rect 11452 24603 11466 24768
rect 11466 24603 11500 24768
rect 11500 24603 11516 24768
rect 11452 24588 11516 24603
rect 11740 24979 11804 24992
rect 11740 24812 11754 24979
rect 11754 24812 11788 24979
rect 11788 24812 11804 24979
rect 11644 24603 11658 24768
rect 11658 24603 11692 24768
rect 11692 24603 11708 24768
rect 11644 24588 11708 24603
rect 11932 24979 11996 24992
rect 11932 24812 11946 24979
rect 11946 24812 11980 24979
rect 11980 24812 11996 24979
rect 11836 24603 11850 24768
rect 11850 24603 11884 24768
rect 11884 24603 11900 24768
rect 11836 24588 11900 24603
rect 12124 24979 12188 24992
rect 12124 24812 12138 24979
rect 12138 24812 12172 24979
rect 12172 24812 12188 24979
rect 12028 24603 12042 24768
rect 12042 24603 12076 24768
rect 12076 24603 12092 24768
rect 12028 24588 12092 24603
rect 12316 24979 12380 24992
rect 12316 24812 12330 24979
rect 12330 24812 12364 24979
rect 12364 24812 12380 24979
rect 12220 24603 12234 24768
rect 12234 24603 12268 24768
rect 12268 24603 12284 24768
rect 12220 24588 12284 24603
rect 13152 24979 13216 24992
rect 13152 24812 13166 24979
rect 13166 24812 13200 24979
rect 13200 24812 13216 24979
rect 13056 24603 13070 24768
rect 13070 24603 13104 24768
rect 13104 24603 13120 24768
rect 13056 24588 13120 24603
rect 13344 24979 13408 24992
rect 13344 24812 13358 24979
rect 13358 24812 13392 24979
rect 13392 24812 13408 24979
rect 13244 24603 13262 24768
rect 13262 24603 13296 24768
rect 13296 24603 13308 24768
rect 13244 24588 13308 24603
rect 13536 24979 13600 24992
rect 13536 24812 13550 24979
rect 13550 24812 13584 24979
rect 13584 24812 13600 24979
rect 13436 24603 13454 24768
rect 13454 24603 13488 24768
rect 13488 24603 13500 24768
rect 13436 24588 13500 24603
rect 13728 24979 13792 24992
rect 13728 24812 13742 24979
rect 13742 24812 13776 24979
rect 13776 24812 13792 24979
rect 13632 24603 13646 24768
rect 13646 24603 13680 24768
rect 13680 24603 13696 24768
rect 13632 24588 13696 24603
rect 13920 24979 13984 24992
rect 13920 24812 13934 24979
rect 13934 24812 13968 24979
rect 13968 24812 13984 24979
rect 13824 24603 13838 24768
rect 13838 24603 13872 24768
rect 13872 24603 13888 24768
rect 13824 24588 13888 24603
rect 14112 24979 14176 24992
rect 14112 24812 14126 24979
rect 14126 24812 14160 24979
rect 14160 24812 14176 24979
rect 14016 24603 14030 24768
rect 14030 24603 14064 24768
rect 14064 24603 14080 24768
rect 14016 24588 14080 24603
rect 14304 24979 14368 24992
rect 14304 24812 14318 24979
rect 14318 24812 14352 24979
rect 14352 24812 14368 24979
rect 14208 24603 14222 24768
rect 14222 24603 14256 24768
rect 14256 24603 14272 24768
rect 14208 24588 14272 24603
rect 14496 24979 14560 24992
rect 14496 24812 14510 24979
rect 14510 24812 14544 24979
rect 14544 24812 14560 24979
rect 14400 24603 14414 24768
rect 14414 24603 14448 24768
rect 14448 24603 14464 24768
rect 14400 24588 14464 24603
rect 15352 24979 15416 24992
rect 15352 24812 15366 24979
rect 15366 24812 15400 24979
rect 15400 24812 15416 24979
rect 15256 24603 15270 24768
rect 15270 24603 15304 24768
rect 15304 24603 15320 24768
rect 15256 24588 15320 24603
rect 15544 24979 15608 24992
rect 15544 24812 15558 24979
rect 15558 24812 15592 24979
rect 15592 24812 15608 24979
rect 15444 24603 15462 24768
rect 15462 24603 15496 24768
rect 15496 24603 15508 24768
rect 15444 24588 15508 24603
rect 15736 24979 15800 24992
rect 15736 24812 15750 24979
rect 15750 24812 15784 24979
rect 15784 24812 15800 24979
rect 15636 24603 15654 24768
rect 15654 24603 15688 24768
rect 15688 24603 15700 24768
rect 15636 24588 15700 24603
rect 15928 24979 15992 24992
rect 15928 24812 15942 24979
rect 15942 24812 15976 24979
rect 15976 24812 15992 24979
rect 15832 24603 15846 24768
rect 15846 24603 15880 24768
rect 15880 24603 15896 24768
rect 15832 24588 15896 24603
rect 16120 24979 16184 24992
rect 16120 24812 16134 24979
rect 16134 24812 16168 24979
rect 16168 24812 16184 24979
rect 16024 24603 16038 24768
rect 16038 24603 16072 24768
rect 16072 24603 16088 24768
rect 16024 24588 16088 24603
rect 16312 24979 16376 24992
rect 16312 24812 16326 24979
rect 16326 24812 16360 24979
rect 16360 24812 16376 24979
rect 16216 24603 16230 24768
rect 16230 24603 16264 24768
rect 16264 24603 16280 24768
rect 16216 24588 16280 24603
rect 16504 24979 16568 24992
rect 16504 24812 16518 24979
rect 16518 24812 16552 24979
rect 16552 24812 16568 24979
rect 16408 24603 16422 24768
rect 16422 24603 16456 24768
rect 16456 24603 16472 24768
rect 16408 24588 16472 24603
rect 16696 24979 16760 24992
rect 16696 24812 16710 24979
rect 16710 24812 16744 24979
rect 16744 24812 16760 24979
rect 16600 24603 16614 24768
rect 16614 24603 16648 24768
rect 16648 24603 16664 24768
rect 16600 24588 16664 24603
rect 18280 25068 18640 25120
rect 18280 24671 18342 25068
rect 18342 24671 18592 25068
rect 18592 24671 18640 25068
rect 18280 24600 18640 24671
rect 19040 25082 19240 25260
rect 19040 25048 19051 25082
rect 19051 25048 19227 25082
rect 19227 25048 19240 25082
rect 19040 25040 19240 25048
rect 6572 24343 6636 24356
rect 6572 24176 6586 24343
rect 6586 24176 6620 24343
rect 6620 24176 6636 24343
rect 6476 23967 6490 24132
rect 6490 23967 6524 24132
rect 6524 23967 6540 24132
rect 6476 23952 6540 23967
rect 6764 24343 6828 24356
rect 6764 24176 6778 24343
rect 6778 24176 6812 24343
rect 6812 24176 6828 24343
rect 6664 23967 6682 24132
rect 6682 23967 6716 24132
rect 6716 23967 6728 24132
rect 6664 23952 6728 23967
rect 6956 24343 7020 24356
rect 6956 24176 6970 24343
rect 6970 24176 7004 24343
rect 7004 24176 7020 24343
rect 6856 23967 6874 24132
rect 6874 23967 6908 24132
rect 6908 23967 6920 24132
rect 6856 23952 6920 23967
rect 7148 24343 7212 24356
rect 7148 24176 7162 24343
rect 7162 24176 7196 24343
rect 7196 24176 7212 24343
rect 7052 23967 7066 24132
rect 7066 23967 7100 24132
rect 7100 23967 7116 24132
rect 7052 23952 7116 23967
rect 7340 24343 7404 24356
rect 7340 24176 7354 24343
rect 7354 24176 7388 24343
rect 7388 24176 7404 24343
rect 7244 23967 7258 24132
rect 7258 23967 7292 24132
rect 7292 23967 7308 24132
rect 7244 23952 7308 23967
rect 7532 24343 7596 24356
rect 7532 24176 7546 24343
rect 7546 24176 7580 24343
rect 7580 24176 7596 24343
rect 7436 23967 7450 24132
rect 7450 23967 7484 24132
rect 7484 23967 7500 24132
rect 7436 23952 7500 23967
rect 7724 24343 7788 24356
rect 7724 24176 7738 24343
rect 7738 24176 7772 24343
rect 7772 24176 7788 24343
rect 7628 23967 7642 24132
rect 7642 23967 7676 24132
rect 7676 23967 7692 24132
rect 7628 23952 7692 23967
rect 7916 24343 7980 24356
rect 7916 24176 7930 24343
rect 7930 24176 7964 24343
rect 7964 24176 7980 24343
rect 8156 24212 8328 24436
rect 7820 23967 7834 24132
rect 7834 23967 7868 24132
rect 7868 23967 7884 24132
rect 7820 23952 7884 23967
rect 8792 24343 8856 24356
rect 8792 24176 8806 24343
rect 8806 24176 8840 24343
rect 8840 24176 8856 24343
rect 8696 23967 8710 24132
rect 8710 23967 8744 24132
rect 8744 23967 8760 24132
rect 8696 23952 8760 23967
rect 8984 24343 9048 24356
rect 8984 24176 8998 24343
rect 8998 24176 9032 24343
rect 9032 24176 9048 24343
rect 8884 23967 8902 24132
rect 8902 23967 8936 24132
rect 8936 23967 8948 24132
rect 8884 23952 8948 23967
rect 9176 24343 9240 24356
rect 9176 24176 9190 24343
rect 9190 24176 9224 24343
rect 9224 24176 9240 24343
rect 9076 23967 9094 24132
rect 9094 23967 9128 24132
rect 9128 23967 9140 24132
rect 9076 23952 9140 23967
rect 9368 24343 9432 24356
rect 9368 24176 9382 24343
rect 9382 24176 9416 24343
rect 9416 24176 9432 24343
rect 9272 23967 9286 24132
rect 9286 23967 9320 24132
rect 9320 23967 9336 24132
rect 9272 23952 9336 23967
rect 9560 24343 9624 24356
rect 9560 24176 9574 24343
rect 9574 24176 9608 24343
rect 9608 24176 9624 24343
rect 9464 23967 9478 24132
rect 9478 23967 9512 24132
rect 9512 23967 9528 24132
rect 9464 23952 9528 23967
rect 9752 24343 9816 24356
rect 9752 24176 9766 24343
rect 9766 24176 9800 24343
rect 9800 24176 9816 24343
rect 9656 23967 9670 24132
rect 9670 23967 9704 24132
rect 9704 23967 9720 24132
rect 9656 23952 9720 23967
rect 9944 24343 10008 24356
rect 9944 24176 9958 24343
rect 9958 24176 9992 24343
rect 9992 24176 10008 24343
rect 9848 23967 9862 24132
rect 9862 23967 9896 24132
rect 9896 23967 9912 24132
rect 9848 23952 9912 23967
rect 10136 24343 10200 24356
rect 10136 24176 10150 24343
rect 10150 24176 10184 24343
rect 10184 24176 10200 24343
rect 10040 23967 10054 24132
rect 10054 23967 10088 24132
rect 10088 23967 10104 24132
rect 10040 23952 10104 23967
rect 10972 24343 11036 24356
rect 10972 24176 10986 24343
rect 10986 24176 11020 24343
rect 11020 24176 11036 24343
rect 10876 23967 10890 24132
rect 10890 23967 10924 24132
rect 10924 23967 10940 24132
rect 10876 23952 10940 23967
rect 11164 24343 11228 24356
rect 11164 24176 11178 24343
rect 11178 24176 11212 24343
rect 11212 24176 11228 24343
rect 11064 23967 11082 24132
rect 11082 23967 11116 24132
rect 11116 23967 11128 24132
rect 11064 23952 11128 23967
rect 11356 24343 11420 24356
rect 11356 24176 11370 24343
rect 11370 24176 11404 24343
rect 11404 24176 11420 24343
rect 11256 23967 11274 24132
rect 11274 23967 11308 24132
rect 11308 23967 11320 24132
rect 11256 23952 11320 23967
rect 11548 24343 11612 24356
rect 11548 24176 11562 24343
rect 11562 24176 11596 24343
rect 11596 24176 11612 24343
rect 11452 23967 11466 24132
rect 11466 23967 11500 24132
rect 11500 23967 11516 24132
rect 11452 23952 11516 23967
rect 11740 24343 11804 24356
rect 11740 24176 11754 24343
rect 11754 24176 11788 24343
rect 11788 24176 11804 24343
rect 11644 23967 11658 24132
rect 11658 23967 11692 24132
rect 11692 23967 11708 24132
rect 11644 23952 11708 23967
rect 11932 24343 11996 24356
rect 11932 24176 11946 24343
rect 11946 24176 11980 24343
rect 11980 24176 11996 24343
rect 11836 23967 11850 24132
rect 11850 23967 11884 24132
rect 11884 23967 11900 24132
rect 11836 23952 11900 23967
rect 12124 24343 12188 24356
rect 12124 24176 12138 24343
rect 12138 24176 12172 24343
rect 12172 24176 12188 24343
rect 12028 23967 12042 24132
rect 12042 23967 12076 24132
rect 12076 23967 12092 24132
rect 12028 23952 12092 23967
rect 12316 24343 12380 24356
rect 12316 24176 12330 24343
rect 12330 24176 12364 24343
rect 12364 24176 12380 24343
rect 12220 23967 12234 24132
rect 12234 23967 12268 24132
rect 12268 23967 12284 24132
rect 12220 23952 12284 23967
rect 13152 24343 13216 24356
rect 13152 24176 13166 24343
rect 13166 24176 13200 24343
rect 13200 24176 13216 24343
rect 13056 23967 13070 24132
rect 13070 23967 13104 24132
rect 13104 23967 13120 24132
rect 13056 23952 13120 23967
rect 13344 24343 13408 24356
rect 13344 24176 13358 24343
rect 13358 24176 13392 24343
rect 13392 24176 13408 24343
rect 13244 23967 13262 24132
rect 13262 23967 13296 24132
rect 13296 23967 13308 24132
rect 13244 23952 13308 23967
rect 13536 24343 13600 24356
rect 13536 24176 13550 24343
rect 13550 24176 13584 24343
rect 13584 24176 13600 24343
rect 13436 23967 13454 24132
rect 13454 23967 13488 24132
rect 13488 23967 13500 24132
rect 13436 23952 13500 23967
rect 13728 24343 13792 24356
rect 13728 24176 13742 24343
rect 13742 24176 13776 24343
rect 13776 24176 13792 24343
rect 13632 23967 13646 24132
rect 13646 23967 13680 24132
rect 13680 23967 13696 24132
rect 13632 23952 13696 23967
rect 13920 24343 13984 24356
rect 13920 24176 13934 24343
rect 13934 24176 13968 24343
rect 13968 24176 13984 24343
rect 13824 23967 13838 24132
rect 13838 23967 13872 24132
rect 13872 23967 13888 24132
rect 13824 23952 13888 23967
rect 14112 24343 14176 24356
rect 14112 24176 14126 24343
rect 14126 24176 14160 24343
rect 14160 24176 14176 24343
rect 14016 23967 14030 24132
rect 14030 23967 14064 24132
rect 14064 23967 14080 24132
rect 14016 23952 14080 23967
rect 14304 24343 14368 24356
rect 14304 24176 14318 24343
rect 14318 24176 14352 24343
rect 14352 24176 14368 24343
rect 14208 23967 14222 24132
rect 14222 23967 14256 24132
rect 14256 23967 14272 24132
rect 14208 23952 14272 23967
rect 14496 24343 14560 24356
rect 14496 24176 14510 24343
rect 14510 24176 14544 24343
rect 14544 24176 14560 24343
rect 14400 23967 14414 24132
rect 14414 23967 14448 24132
rect 14448 23967 14464 24132
rect 14400 23952 14464 23967
rect 15352 24343 15416 24356
rect 15352 24176 15366 24343
rect 15366 24176 15400 24343
rect 15400 24176 15416 24343
rect 15256 23967 15270 24132
rect 15270 23967 15304 24132
rect 15304 23967 15320 24132
rect 15256 23952 15320 23967
rect 15544 24343 15608 24356
rect 15544 24176 15558 24343
rect 15558 24176 15592 24343
rect 15592 24176 15608 24343
rect 15444 23967 15462 24132
rect 15462 23967 15496 24132
rect 15496 23967 15508 24132
rect 15444 23952 15508 23967
rect 15736 24343 15800 24356
rect 15736 24176 15750 24343
rect 15750 24176 15784 24343
rect 15784 24176 15800 24343
rect 15636 23967 15654 24132
rect 15654 23967 15688 24132
rect 15688 23967 15700 24132
rect 15636 23952 15700 23967
rect 15928 24343 15992 24356
rect 15928 24176 15942 24343
rect 15942 24176 15976 24343
rect 15976 24176 15992 24343
rect 15832 23967 15846 24132
rect 15846 23967 15880 24132
rect 15880 23967 15896 24132
rect 15832 23952 15896 23967
rect 16120 24343 16184 24356
rect 16120 24176 16134 24343
rect 16134 24176 16168 24343
rect 16168 24176 16184 24343
rect 16024 23967 16038 24132
rect 16038 23967 16072 24132
rect 16072 23967 16088 24132
rect 16024 23952 16088 23967
rect 16312 24343 16376 24356
rect 16312 24176 16326 24343
rect 16326 24176 16360 24343
rect 16360 24176 16376 24343
rect 16216 23967 16230 24132
rect 16230 23967 16264 24132
rect 16264 23967 16280 24132
rect 16216 23952 16280 23967
rect 16504 24343 16568 24356
rect 16504 24176 16518 24343
rect 16518 24176 16552 24343
rect 16552 24176 16568 24343
rect 16408 23967 16422 24132
rect 16422 23967 16456 24132
rect 16456 23967 16472 24132
rect 16408 23952 16472 23967
rect 16696 24343 16760 24356
rect 16696 24176 16710 24343
rect 16710 24176 16744 24343
rect 16744 24176 16760 24343
rect 16600 23967 16614 24132
rect 16614 23967 16648 24132
rect 16648 23967 16664 24132
rect 16600 23952 16664 23967
rect 6696 23410 6748 23424
rect 6696 23244 6706 23410
rect 6706 23244 6740 23410
rect 6740 23244 6748 23410
rect 6600 23034 6610 23200
rect 6610 23034 6644 23200
rect 6644 23034 6652 23200
rect 6600 23020 6652 23034
rect 6888 23410 6940 23424
rect 6888 23244 6898 23410
rect 6898 23244 6932 23410
rect 6932 23244 6940 23410
rect 6792 23034 6802 23200
rect 6802 23034 6836 23200
rect 6836 23034 6844 23200
rect 6792 23020 6844 23034
rect 7080 23410 7132 23424
rect 7080 23244 7090 23410
rect 7090 23244 7124 23410
rect 7124 23244 7132 23410
rect 6984 23034 6994 23200
rect 6994 23034 7028 23200
rect 7028 23034 7036 23200
rect 6984 23020 7036 23034
rect 7272 23410 7324 23424
rect 7272 23244 7282 23410
rect 7282 23244 7316 23410
rect 7316 23244 7324 23410
rect 7176 23034 7186 23200
rect 7186 23034 7220 23200
rect 7220 23034 7228 23200
rect 7176 23020 7228 23034
rect 7464 23410 7516 23424
rect 7464 23244 7474 23410
rect 7474 23244 7508 23410
rect 7508 23244 7516 23410
rect 7368 23034 7378 23200
rect 7378 23034 7412 23200
rect 7412 23034 7420 23200
rect 7368 23020 7420 23034
rect 7560 23034 7570 23200
rect 7570 23034 7604 23200
rect 7604 23034 7612 23200
rect 7560 23020 7612 23034
rect 8416 23410 8468 23424
rect 8416 23244 8426 23410
rect 8426 23244 8460 23410
rect 8460 23244 8468 23410
rect 8320 23034 8330 23200
rect 8330 23034 8364 23200
rect 8364 23034 8372 23200
rect 8320 23020 8372 23034
rect 8608 23410 8660 23424
rect 8608 23244 8618 23410
rect 8618 23244 8652 23410
rect 8652 23244 8660 23410
rect 8512 23034 8522 23200
rect 8522 23034 8556 23200
rect 8556 23034 8564 23200
rect 8512 23020 8564 23034
rect 8800 23410 8852 23424
rect 8800 23244 8810 23410
rect 8810 23244 8844 23410
rect 8844 23244 8852 23410
rect 8704 23034 8714 23200
rect 8714 23034 8748 23200
rect 8748 23034 8756 23200
rect 8704 23020 8756 23034
rect 8992 23410 9044 23424
rect 8992 23244 9002 23410
rect 9002 23244 9036 23410
rect 9036 23244 9044 23410
rect 8896 23034 8906 23200
rect 8906 23034 8940 23200
rect 8940 23034 8948 23200
rect 8896 23020 8948 23034
rect 9184 23410 9236 23424
rect 9184 23244 9194 23410
rect 9194 23244 9228 23410
rect 9228 23244 9236 23410
rect 9088 23034 9098 23200
rect 9098 23034 9132 23200
rect 9132 23034 9140 23200
rect 9088 23020 9140 23034
rect 9280 23034 9290 23200
rect 9290 23034 9324 23200
rect 9324 23034 9332 23200
rect 9280 23020 9332 23034
rect 18328 23837 18688 23852
rect 18328 23440 18342 23837
rect 18342 23440 18592 23837
rect 18592 23440 18688 23837
rect 18328 23420 18688 23440
rect 19044 23424 19232 23448
rect 19044 23390 19051 23424
rect 19051 23390 19227 23424
rect 19227 23390 19232 23424
rect 19044 23364 19232 23390
rect 6696 22792 6748 22808
rect 6696 22628 6706 22792
rect 6706 22628 6740 22792
rect 6740 22628 6748 22792
rect 6600 22416 6610 22584
rect 6610 22416 6644 22584
rect 6644 22416 6652 22584
rect 6600 22404 6652 22416
rect 6888 22792 6940 22808
rect 6888 22628 6898 22792
rect 6898 22628 6932 22792
rect 6932 22628 6940 22792
rect 6792 22416 6802 22584
rect 6802 22416 6836 22584
rect 6836 22416 6844 22584
rect 6792 22404 6844 22416
rect 7080 22792 7132 22808
rect 7080 22628 7090 22792
rect 7090 22628 7124 22792
rect 7124 22628 7132 22792
rect 6984 22416 6994 22584
rect 6994 22416 7028 22584
rect 7028 22416 7036 22584
rect 6984 22404 7036 22416
rect 7272 22792 7324 22808
rect 7272 22628 7282 22792
rect 7282 22628 7316 22792
rect 7316 22628 7324 22792
rect 7176 22416 7186 22584
rect 7186 22416 7220 22584
rect 7220 22416 7228 22584
rect 7176 22404 7228 22416
rect 7464 22792 7516 22808
rect 7464 22628 7474 22792
rect 7474 22628 7508 22792
rect 7508 22628 7516 22792
rect 7368 22416 7378 22584
rect 7378 22416 7412 22584
rect 7412 22416 7420 22584
rect 7368 22404 7420 22416
rect 7560 22416 7570 22584
rect 7570 22416 7604 22584
rect 7604 22416 7612 22584
rect 7560 22404 7612 22416
rect 8416 22792 8468 22808
rect 8416 22628 8426 22792
rect 8426 22628 8460 22792
rect 8460 22628 8468 22792
rect 8320 22416 8330 22584
rect 8330 22416 8364 22584
rect 8364 22416 8372 22584
rect 8320 22404 8372 22416
rect 8608 22792 8660 22808
rect 8608 22628 8618 22792
rect 8618 22628 8652 22792
rect 8652 22628 8660 22792
rect 8512 22416 8522 22584
rect 8522 22416 8556 22584
rect 8556 22416 8564 22584
rect 8512 22404 8564 22416
rect 8800 22792 8852 22808
rect 8800 22628 8810 22792
rect 8810 22628 8844 22792
rect 8844 22628 8852 22792
rect 8704 22416 8714 22584
rect 8714 22416 8748 22584
rect 8748 22416 8756 22584
rect 8704 22404 8756 22416
rect 8992 22792 9044 22808
rect 8992 22628 9002 22792
rect 9002 22628 9036 22792
rect 9036 22628 9044 22792
rect 8896 22416 8906 22584
rect 8906 22416 8940 22584
rect 8940 22416 8948 22584
rect 8896 22404 8948 22416
rect 9184 22792 9236 22808
rect 9184 22628 9194 22792
rect 9194 22628 9228 22792
rect 9228 22628 9236 22792
rect 9088 22416 9098 22584
rect 9098 22416 9132 22584
rect 9132 22416 9140 22584
rect 9088 22404 9140 22416
rect 9280 22416 9290 22584
rect 9290 22416 9324 22584
rect 9324 22416 9332 22584
rect 9280 22404 9332 22416
rect 18396 23011 18448 23024
rect 18396 22844 18406 23011
rect 18406 22844 18440 23011
rect 18440 22844 18448 23011
rect 18300 22635 18310 22800
rect 18310 22635 18344 22800
rect 18344 22635 18352 22800
rect 18300 22620 18352 22635
rect 18588 23011 18640 23024
rect 18588 22844 18598 23011
rect 18598 22844 18632 23011
rect 18632 22844 18640 23011
rect 18492 22635 18502 22800
rect 18502 22635 18536 22800
rect 18536 22635 18544 22800
rect 18492 22620 18544 22635
rect 18780 23011 18832 23024
rect 18780 22844 18790 23011
rect 18790 22844 18824 23011
rect 18824 22844 18832 23011
rect 18684 22635 18694 22800
rect 18694 22635 18728 22800
rect 18728 22635 18736 22800
rect 18684 22620 18736 22635
rect 18972 23011 19024 23024
rect 18972 22844 18982 23011
rect 18982 22844 19016 23011
rect 19016 22844 19024 23011
rect 18876 22635 18886 22800
rect 18886 22635 18920 22800
rect 18920 22635 18928 22800
rect 18876 22620 18928 22635
rect 19164 23011 19216 23024
rect 19164 22844 19174 23011
rect 19174 22844 19208 23011
rect 19208 22844 19216 23011
rect 19068 22635 19078 22800
rect 19078 22635 19112 22800
rect 19112 22635 19120 22800
rect 19068 22620 19120 22635
rect 19260 22635 19270 22800
rect 19270 22635 19304 22800
rect 19304 22635 19312 22800
rect 19260 22620 19312 22635
rect 18272 22542 18358 22572
rect 18358 22542 18392 22572
rect 18392 22542 18550 22572
rect 18550 22542 18584 22572
rect 18584 22542 18742 22572
rect 18742 22542 18776 22572
rect 18776 22542 18860 22572
rect 18272 22472 18860 22542
rect 6696 22174 6748 22188
rect 6696 22008 6706 22174
rect 6706 22008 6740 22174
rect 6740 22008 6748 22174
rect 6600 21798 6610 21964
rect 6610 21798 6644 21964
rect 6644 21798 6652 21964
rect 6600 21784 6652 21798
rect 6888 22174 6940 22188
rect 6888 22008 6898 22174
rect 6898 22008 6932 22174
rect 6932 22008 6940 22174
rect 6792 21798 6802 21964
rect 6802 21798 6836 21964
rect 6836 21798 6844 21964
rect 6792 21784 6844 21798
rect 7080 22174 7132 22188
rect 7080 22008 7090 22174
rect 7090 22008 7124 22174
rect 7124 22008 7132 22174
rect 6984 21798 6994 21964
rect 6994 21798 7028 21964
rect 7028 21798 7036 21964
rect 6984 21784 7036 21798
rect 7272 22174 7324 22188
rect 7272 22008 7282 22174
rect 7282 22008 7316 22174
rect 7316 22008 7324 22174
rect 7176 21798 7186 21964
rect 7186 21798 7220 21964
rect 7220 21798 7228 21964
rect 7176 21784 7228 21798
rect 7464 22174 7516 22188
rect 7464 22008 7474 22174
rect 7474 22008 7508 22174
rect 7508 22008 7516 22174
rect 7368 21798 7378 21964
rect 7378 21798 7412 21964
rect 7412 21798 7420 21964
rect 7368 21784 7420 21798
rect 7560 21798 7570 21964
rect 7570 21798 7604 21964
rect 7604 21798 7612 21964
rect 7560 21784 7612 21798
rect 8416 22174 8468 22188
rect 8416 22008 8426 22174
rect 8426 22008 8460 22174
rect 8460 22008 8468 22174
rect 8320 21798 8330 21964
rect 8330 21798 8364 21964
rect 8364 21798 8372 21964
rect 8320 21784 8372 21798
rect 8608 22174 8660 22188
rect 8608 22008 8618 22174
rect 8618 22008 8652 22174
rect 8652 22008 8660 22174
rect 8512 21798 8522 21964
rect 8522 21798 8556 21964
rect 8556 21798 8564 21964
rect 8512 21784 8564 21798
rect 8800 22174 8852 22188
rect 8800 22008 8810 22174
rect 8810 22008 8844 22174
rect 8844 22008 8852 22174
rect 8704 21798 8714 21964
rect 8714 21798 8748 21964
rect 8748 21798 8756 21964
rect 8704 21784 8756 21798
rect 8992 22174 9044 22188
rect 8992 22008 9002 22174
rect 9002 22008 9036 22174
rect 9036 22008 9044 22174
rect 8896 21798 8906 21964
rect 8906 21798 8940 21964
rect 8940 21798 8948 21964
rect 8896 21784 8948 21798
rect 9184 22174 9236 22188
rect 9184 22008 9194 22174
rect 9194 22008 9228 22174
rect 9228 22008 9236 22174
rect 9088 21798 9098 21964
rect 9098 21798 9132 21964
rect 9132 21798 9140 21964
rect 9088 21784 9140 21798
rect 9280 21798 9290 21964
rect 9290 21798 9324 21964
rect 9324 21798 9332 21964
rect 9280 21784 9332 21798
rect 18392 22152 18444 22168
rect 18392 21988 18406 22152
rect 18406 21988 18440 22152
rect 18440 21988 18444 22152
rect 18300 21776 18310 21944
rect 18310 21776 18344 21944
rect 18344 21776 18352 21944
rect 18300 21764 18352 21776
rect 18584 22152 18636 22168
rect 18584 21988 18598 22152
rect 18598 21988 18632 22152
rect 18632 21988 18636 22152
rect 18488 21776 18502 21944
rect 18502 21776 18536 21944
rect 18536 21776 18540 21944
rect 18488 21764 18540 21776
rect 18776 22152 18828 22168
rect 18776 21988 18790 22152
rect 18790 21988 18824 22152
rect 18824 21988 18828 22152
rect 18680 21776 18694 21944
rect 18694 21776 18728 21944
rect 18728 21776 18732 21944
rect 18680 21764 18732 21776
rect 18968 22152 19020 22168
rect 18968 21988 18982 22152
rect 18982 21988 19016 22152
rect 19016 21988 19020 22152
rect 18872 21776 18886 21944
rect 18886 21776 18920 21944
rect 18920 21776 18924 21944
rect 18872 21764 18924 21776
rect 19160 22152 19212 22168
rect 19160 21988 19174 22152
rect 19174 21988 19208 22152
rect 19208 21988 19212 22152
rect 19064 21776 19078 21944
rect 19078 21776 19112 21944
rect 19112 21776 19116 21944
rect 19064 21764 19116 21776
rect 19256 21776 19270 21944
rect 19270 21776 19304 21944
rect 19304 21776 19308 21944
rect 19256 21764 19308 21776
rect 6600 21264 6652 21276
rect 6600 21096 6610 21264
rect 6610 21096 6644 21264
rect 6644 21096 6652 21264
rect 6860 20888 6868 21056
rect 6868 20888 6902 21056
rect 6902 20888 6912 21056
rect 6860 20876 6912 20888
rect 7116 21264 7168 21276
rect 7116 21096 7126 21264
rect 7126 21096 7160 21264
rect 7160 21096 7168 21264
rect 7376 20888 7384 21056
rect 7384 20888 7418 21056
rect 7418 20888 7428 21056
rect 7376 20876 7428 20888
rect 7632 21264 7684 21276
rect 7632 21096 7642 21264
rect 7642 21096 7676 21264
rect 7676 21096 7684 21264
rect 8320 21264 8372 21276
rect 8320 21096 8330 21264
rect 8330 21096 8364 21264
rect 8364 21096 8372 21264
rect 7892 20888 7900 21056
rect 7900 20888 7934 21056
rect 7934 20888 7944 21056
rect 7892 20876 7944 20888
rect 8580 20888 8588 21056
rect 8588 20888 8622 21056
rect 8622 20888 8632 21056
rect 8580 20876 8632 20888
rect 8836 21264 8888 21276
rect 8836 21096 8846 21264
rect 8846 21096 8880 21264
rect 8880 21096 8888 21264
rect 9096 20888 9104 21056
rect 9104 20888 9138 21056
rect 9138 20888 9148 21056
rect 9096 20876 9148 20888
rect 9352 21264 9404 21276
rect 9352 21096 9362 21264
rect 9362 21096 9396 21264
rect 9396 21096 9404 21264
rect 9612 20888 9620 21056
rect 9620 20888 9654 21056
rect 9654 20888 9664 21056
rect 9612 20876 9664 20888
rect 10380 20860 10840 21220
rect 6600 20646 6652 20660
rect 6600 20480 6610 20646
rect 6610 20480 6644 20646
rect 6644 20480 6652 20646
rect 6860 20270 6868 20440
rect 6868 20270 6902 20440
rect 6902 20270 6912 20440
rect 6860 20260 6912 20270
rect 7116 20646 7168 20660
rect 7116 20480 7126 20646
rect 7126 20480 7160 20646
rect 7160 20480 7168 20646
rect 7376 20270 7384 20440
rect 7384 20270 7418 20440
rect 7418 20270 7428 20440
rect 7376 20260 7428 20270
rect 7632 20646 7684 20660
rect 7632 20480 7642 20646
rect 7642 20480 7676 20646
rect 7676 20480 7684 20646
rect 8320 20646 8372 20660
rect 8320 20480 8330 20646
rect 8330 20480 8364 20646
rect 8364 20480 8372 20646
rect 7892 20270 7900 20440
rect 7900 20270 7934 20440
rect 7934 20270 7944 20440
rect 7892 20260 7944 20270
rect 8580 20270 8588 20440
rect 8588 20270 8622 20440
rect 8622 20270 8632 20440
rect 8580 20260 8632 20270
rect 8836 20646 8888 20660
rect 8836 20480 8846 20646
rect 8846 20480 8880 20646
rect 8880 20480 8888 20646
rect 9096 20270 9104 20440
rect 9104 20270 9138 20440
rect 9138 20270 9148 20440
rect 9096 20260 9148 20270
rect 9352 20646 9404 20660
rect 9352 20480 9362 20646
rect 9362 20480 9396 20646
rect 9396 20480 9404 20646
rect 9612 20270 9620 20440
rect 9620 20270 9654 20440
rect 9654 20270 9664 20440
rect 9612 20260 9664 20270
rect 6600 20028 6652 20040
rect 6600 19860 6610 20028
rect 6610 19860 6644 20028
rect 6644 19860 6652 20028
rect 6860 19652 6868 19820
rect 6868 19652 6902 19820
rect 6902 19652 6912 19820
rect 6860 19640 6912 19652
rect 7116 20028 7168 20040
rect 7116 19860 7126 20028
rect 7126 19860 7160 20028
rect 7160 19860 7168 20028
rect 7376 19652 7384 19820
rect 7384 19652 7418 19820
rect 7418 19652 7428 19820
rect 7376 19640 7428 19652
rect 7632 20028 7684 20040
rect 7632 19860 7642 20028
rect 7642 19860 7676 20028
rect 7676 19860 7684 20028
rect 8320 20028 8372 20040
rect 8320 19860 8330 20028
rect 8330 19860 8364 20028
rect 8364 19860 8372 20028
rect 7892 19652 7900 19820
rect 7900 19652 7934 19820
rect 7934 19652 7944 19820
rect 7892 19640 7944 19652
rect 8580 19652 8588 19820
rect 8588 19652 8622 19820
rect 8622 19652 8632 19820
rect 8580 19640 8632 19652
rect 8836 20028 8888 20040
rect 8836 19860 8846 20028
rect 8846 19860 8880 20028
rect 8880 19860 8888 20028
rect 9096 19652 9104 19820
rect 9104 19652 9138 19820
rect 9138 19652 9148 19820
rect 9096 19640 9148 19652
rect 9352 20028 9404 20040
rect 9352 19860 9362 20028
rect 9362 19860 9396 20028
rect 9396 19860 9404 20028
rect 9612 19652 9620 19820
rect 9620 19652 9654 19820
rect 9654 19652 9664 19820
rect 9612 19640 9664 19652
rect 10188 19768 10260 19836
rect 6600 19410 6652 19424
rect 6600 19244 6610 19410
rect 6610 19244 6644 19410
rect 6644 19244 6652 19410
rect 6860 19034 6868 19204
rect 6868 19034 6902 19204
rect 6902 19034 6912 19204
rect 6860 19024 6912 19034
rect 7116 19410 7168 19424
rect 7116 19244 7126 19410
rect 7126 19244 7160 19410
rect 7160 19244 7168 19410
rect 7376 19034 7384 19204
rect 7384 19034 7418 19204
rect 7418 19034 7428 19204
rect 7376 19024 7428 19034
rect 7632 19410 7684 19424
rect 7632 19244 7642 19410
rect 7642 19244 7676 19410
rect 7676 19244 7684 19410
rect 8320 19410 8372 19424
rect 8320 19244 8330 19410
rect 8330 19244 8364 19410
rect 8364 19244 8372 19410
rect 7892 19034 7900 19204
rect 7900 19034 7934 19204
rect 7934 19034 7944 19204
rect 7892 19024 7944 19034
rect 8580 19034 8588 19204
rect 8588 19034 8622 19204
rect 8622 19034 8632 19204
rect 8580 19024 8632 19034
rect 8836 19410 8888 19424
rect 8836 19244 8846 19410
rect 8846 19244 8880 19410
rect 8880 19244 8888 19410
rect 9096 19034 9104 19204
rect 9104 19034 9138 19204
rect 9138 19034 9148 19204
rect 9096 19024 9148 19034
rect 9352 19410 9404 19424
rect 9352 19244 9362 19410
rect 9362 19244 9396 19410
rect 9396 19244 9404 19410
rect 10252 19714 10312 19728
rect 10252 19548 10266 19714
rect 10266 19548 10300 19714
rect 10300 19548 10312 19714
rect 10160 19338 10170 19504
rect 10170 19338 10204 19504
rect 10204 19338 10220 19504
rect 10160 19324 10220 19338
rect 10444 19714 10504 19728
rect 10444 19548 10458 19714
rect 10458 19548 10492 19714
rect 10492 19548 10504 19714
rect 10348 19338 10362 19504
rect 10362 19338 10396 19504
rect 10396 19338 10408 19504
rect 10348 19324 10408 19338
rect 10636 19714 10696 19728
rect 10636 19548 10650 19714
rect 10650 19548 10684 19714
rect 10684 19548 10696 19714
rect 10540 19338 10554 19504
rect 10554 19338 10588 19504
rect 10588 19338 10600 19504
rect 10540 19324 10600 19338
rect 10828 19714 10888 19728
rect 10828 19548 10842 19714
rect 10842 19548 10876 19714
rect 10876 19548 10888 19714
rect 10732 19338 10746 19504
rect 10746 19338 10780 19504
rect 10780 19338 10792 19504
rect 10732 19324 10792 19338
rect 9612 19034 9620 19204
rect 9620 19034 9654 19204
rect 9654 19034 9664 19204
rect 9612 19024 9664 19034
rect 6600 18792 6652 18804
rect 6600 18624 6610 18792
rect 6610 18624 6644 18792
rect 6644 18624 6652 18792
rect 6860 18416 6868 18584
rect 6868 18416 6902 18584
rect 6902 18416 6912 18584
rect 6860 18404 6912 18416
rect 7116 18792 7168 18804
rect 7116 18624 7126 18792
rect 7126 18624 7160 18792
rect 7160 18624 7168 18792
rect 7376 18416 7384 18584
rect 7384 18416 7418 18584
rect 7418 18416 7428 18584
rect 7376 18404 7428 18416
rect 7632 18792 7684 18804
rect 7632 18624 7642 18792
rect 7642 18624 7676 18792
rect 7676 18624 7684 18792
rect 8320 18792 8372 18804
rect 8320 18624 8330 18792
rect 8330 18624 8364 18792
rect 8364 18624 8372 18792
rect 7892 18416 7900 18584
rect 7900 18416 7934 18584
rect 7934 18416 7944 18584
rect 7892 18404 7944 18416
rect 8580 18416 8588 18584
rect 8588 18416 8622 18584
rect 8622 18416 8632 18584
rect 8580 18404 8632 18416
rect 8836 18792 8888 18804
rect 8836 18624 8846 18792
rect 8846 18624 8880 18792
rect 8880 18624 8888 18792
rect 9096 18416 9104 18584
rect 9104 18416 9138 18584
rect 9138 18416 9148 18584
rect 9096 18404 9148 18416
rect 9352 18792 9404 18804
rect 9352 18624 9362 18792
rect 9362 18624 9396 18792
rect 9396 18624 9404 18792
rect 9612 18416 9620 18584
rect 9620 18416 9654 18584
rect 9654 18416 9664 18584
rect 9612 18404 9664 18416
rect 10252 18792 10312 18804
rect 10252 18624 10266 18792
rect 10266 18624 10300 18792
rect 10300 18624 10312 18792
rect 10160 18416 10170 18584
rect 10170 18416 10204 18584
rect 10204 18416 10220 18584
rect 10160 18404 10220 18416
rect 10444 18792 10504 18804
rect 10444 18624 10458 18792
rect 10458 18624 10492 18792
rect 10492 18624 10504 18792
rect 10348 18416 10362 18584
rect 10362 18416 10396 18584
rect 10396 18416 10408 18584
rect 10348 18404 10408 18416
rect 10636 18792 10696 18804
rect 10636 18624 10650 18792
rect 10650 18624 10684 18792
rect 10684 18624 10696 18792
rect 10540 18416 10554 18584
rect 10554 18416 10588 18584
rect 10588 18416 10600 18584
rect 10540 18404 10600 18416
rect 10828 18792 10888 18804
rect 10828 18624 10842 18792
rect 10842 18624 10876 18792
rect 10876 18624 10888 18792
rect 10732 18416 10746 18584
rect 10746 18416 10780 18584
rect 10780 18416 10792 18584
rect 10732 18404 10792 18416
rect 11020 18792 11080 18804
rect 11020 18624 11034 18792
rect 11034 18624 11068 18792
rect 11068 18624 11080 18792
rect 10924 18416 10938 18584
rect 10938 18416 10972 18584
rect 10972 18416 10984 18584
rect 10924 18404 10984 18416
rect 11116 18416 11130 18584
rect 11130 18416 11164 18584
rect 11164 18416 11176 18584
rect 11116 18404 11176 18416
rect 6600 18174 6652 18188
rect 6600 18008 6610 18174
rect 6610 18008 6644 18174
rect 6644 18008 6652 18174
rect 6860 17798 6868 17968
rect 6868 17798 6902 17968
rect 6902 17798 6912 17968
rect 6860 17788 6912 17798
rect 7116 18174 7168 18188
rect 7116 18008 7126 18174
rect 7126 18008 7160 18174
rect 7160 18008 7168 18174
rect 7376 17798 7384 17968
rect 7384 17798 7418 17968
rect 7418 17798 7428 17968
rect 7376 17788 7428 17798
rect 7632 18174 7684 18188
rect 7632 18008 7642 18174
rect 7642 18008 7676 18174
rect 7676 18008 7684 18174
rect 8320 18174 8372 18188
rect 8320 18008 8330 18174
rect 8330 18008 8364 18174
rect 8364 18008 8372 18174
rect 7892 17798 7900 17968
rect 7900 17798 7934 17968
rect 7934 17798 7944 17968
rect 7892 17788 7944 17798
rect 8580 17798 8588 17968
rect 8588 17798 8622 17968
rect 8622 17798 8632 17968
rect 8580 17788 8632 17798
rect 8040 17616 8220 17776
rect 8836 18174 8888 18188
rect 8836 18008 8846 18174
rect 8846 18008 8880 18174
rect 8880 18008 8888 18174
rect 9096 17798 9104 17968
rect 9104 17798 9138 17968
rect 9138 17798 9148 17968
rect 9096 17788 9148 17798
rect 9352 18174 9404 18188
rect 9352 18008 9362 18174
rect 9362 18008 9396 18174
rect 9396 18008 9404 18174
rect 9612 17798 9620 17968
rect 9620 17798 9654 17968
rect 9654 17798 9664 17968
rect 9612 17788 9664 17798
rect 10252 18174 10312 18188
rect 10252 18008 10266 18174
rect 10266 18008 10300 18174
rect 10300 18008 10312 18174
rect 10160 17798 10170 17964
rect 10170 17798 10204 17964
rect 10204 17798 10220 17964
rect 10160 17784 10220 17798
rect 10444 18174 10504 18188
rect 10444 18008 10458 18174
rect 10458 18008 10492 18174
rect 10492 18008 10504 18174
rect 10348 17798 10362 17964
rect 10362 17798 10396 17964
rect 10396 17798 10408 17964
rect 10348 17784 10408 17798
rect 10636 18174 10696 18188
rect 10636 18008 10650 18174
rect 10650 18008 10684 18174
rect 10684 18008 10696 18174
rect 10540 17798 10554 17964
rect 10554 17798 10588 17964
rect 10588 17798 10600 17964
rect 10540 17784 10600 17798
rect 10828 18174 10888 18188
rect 10828 18008 10842 18174
rect 10842 18008 10876 18174
rect 10876 18008 10888 18174
rect 10732 17798 10746 17964
rect 10746 17798 10780 17964
rect 10780 17798 10792 17964
rect 10732 17784 10792 17798
rect 11020 18174 11080 18188
rect 11020 18008 11034 18174
rect 11034 18008 11068 18174
rect 11068 18008 11080 18174
rect 10924 17798 10938 17964
rect 10938 17798 10972 17964
rect 10972 17798 10984 17964
rect 10924 17784 10984 17798
rect 11116 17798 11130 17964
rect 11130 17798 11164 17964
rect 11164 17798 11176 17964
rect 11116 17784 11176 17798
rect 1300 10532 1568 10768
rect 2588 11100 4792 11148
rect 2588 10703 2618 11100
rect 2618 10703 2868 11100
rect 2868 10703 2996 11100
rect 2996 10703 3246 11100
rect 3246 10703 3374 11100
rect 3374 10703 3624 11100
rect 3624 10703 3752 11100
rect 3752 10703 4002 11100
rect 4002 10703 4130 11100
rect 4130 10703 4380 11100
rect 4380 10703 4508 11100
rect 4508 10703 4758 11100
rect 4758 10703 4792 11100
rect 2588 10660 4792 10703
rect 6096 10608 6276 10808
rect 5212 10271 5268 10284
rect 5212 10104 5222 10271
rect 5222 10104 5256 10271
rect 5256 10104 5268 10271
rect 2588 9869 4780 9908
rect 2588 9472 2618 9869
rect 2618 9472 2868 9869
rect 2868 9472 2996 9869
rect 2996 9472 3246 9869
rect 3246 9472 3374 9869
rect 3374 9472 3624 9869
rect 3624 9472 3752 9869
rect 3752 9472 4002 9869
rect 4002 9472 4130 9869
rect 4130 9472 4380 9869
rect 4380 9472 4508 9869
rect 4508 9472 4758 9869
rect 4758 9472 4780 9869
rect 2588 9440 4780 9472
rect 5116 9895 5126 10060
rect 5126 9895 5160 10060
rect 5160 9895 5172 10060
rect 5116 9880 5172 9895
rect 5404 10271 5460 10284
rect 5404 10104 5414 10271
rect 5414 10104 5448 10271
rect 5448 10104 5460 10271
rect 5308 9895 5318 10060
rect 5318 9895 5352 10060
rect 5352 9895 5364 10060
rect 5308 9880 5364 9895
rect 5596 10271 5652 10284
rect 5596 10104 5606 10271
rect 5606 10104 5640 10271
rect 5640 10104 5652 10271
rect 5500 9895 5510 10060
rect 5510 9895 5544 10060
rect 5544 9895 5556 10060
rect 5500 9880 5556 9895
rect 5788 10271 5844 10284
rect 5788 10104 5798 10271
rect 5798 10104 5832 10271
rect 5832 10104 5844 10271
rect 5692 9895 5702 10060
rect 5702 9895 5736 10060
rect 5736 9895 5748 10060
rect 5692 9880 5748 9895
rect 5980 10271 6036 10284
rect 5980 10104 5990 10271
rect 5990 10104 6024 10271
rect 6024 10104 6036 10271
rect 5884 9895 5894 10060
rect 5894 9895 5928 10060
rect 5928 9895 5940 10060
rect 5884 9880 5940 9895
rect 6172 10271 6228 10284
rect 6172 10104 6182 10271
rect 6182 10104 6216 10271
rect 6216 10104 6228 10271
rect 6076 9895 6086 10060
rect 6086 9895 6120 10060
rect 6120 9895 6132 10060
rect 6076 9880 6132 9895
rect 6364 10271 6420 10284
rect 6364 10104 6374 10271
rect 6374 10104 6408 10271
rect 6408 10104 6420 10271
rect 6268 9895 6278 10060
rect 6278 9895 6312 10060
rect 6312 9895 6324 10060
rect 6268 9880 6324 9895
rect 6556 10271 6612 10284
rect 6556 10104 6566 10271
rect 6566 10104 6600 10271
rect 6600 10104 6612 10271
rect 6460 9895 6470 10060
rect 6470 9895 6504 10060
rect 6504 9895 6516 10060
rect 6460 9880 6516 9895
rect 6748 10271 6804 10284
rect 6748 10104 6758 10271
rect 6758 10104 6792 10271
rect 6792 10104 6804 10271
rect 6652 9895 6662 10060
rect 6662 9895 6696 10060
rect 6696 9895 6708 10060
rect 6652 9880 6708 9895
rect 6940 10271 6996 10284
rect 6940 10104 6950 10271
rect 6950 10104 6984 10271
rect 6984 10104 6996 10271
rect 6844 9895 6854 10060
rect 6854 9895 6888 10060
rect 6888 9895 6900 10060
rect 6844 9880 6900 9895
rect 7036 9895 7046 10060
rect 7046 9895 7080 10060
rect 7080 9895 7092 10060
rect 7036 9880 7092 9895
rect 7712 10250 7768 10264
rect 7712 10080 7722 10250
rect 7722 10080 7756 10250
rect 7756 10080 7768 10250
rect 7616 9874 7626 10044
rect 7626 9874 7660 10044
rect 7660 9874 7672 10044
rect 7616 9860 7672 9874
rect 7904 10250 7960 10264
rect 7904 10080 7914 10250
rect 7914 10080 7948 10250
rect 7948 10080 7960 10250
rect 7808 9874 7818 10044
rect 7818 9874 7852 10044
rect 7852 9874 7864 10044
rect 7808 9860 7864 9874
rect 8096 10250 8152 10264
rect 8096 10080 8106 10250
rect 8106 10080 8140 10250
rect 8140 10080 8152 10250
rect 8000 9874 8010 10044
rect 8010 9874 8044 10044
rect 8044 9874 8056 10044
rect 8000 9860 8056 9874
rect 8288 10250 8344 10264
rect 8288 10080 8298 10250
rect 8298 10080 8332 10250
rect 8332 10080 8344 10250
rect 8192 9874 8202 10044
rect 8202 9874 8236 10044
rect 8236 9874 8248 10044
rect 8192 9860 8248 9874
rect 8480 10250 8536 10264
rect 8480 10080 8490 10250
rect 8490 10080 8524 10250
rect 8524 10080 8536 10250
rect 8384 9874 8394 10044
rect 8394 9874 8428 10044
rect 8428 9874 8440 10044
rect 8384 9860 8440 9874
rect 8672 10250 8728 10264
rect 8672 10080 8682 10250
rect 8682 10080 8716 10250
rect 8716 10080 8728 10250
rect 8576 9874 8586 10044
rect 8586 9874 8620 10044
rect 8620 9874 8632 10044
rect 8576 9860 8632 9874
rect 8864 10250 8920 10264
rect 8864 10080 8874 10250
rect 8874 10080 8908 10250
rect 8908 10080 8920 10250
rect 8768 9874 8778 10044
rect 8778 9874 8812 10044
rect 8812 9874 8824 10044
rect 8768 9860 8824 9874
rect 9056 10250 9112 10264
rect 9056 10080 9066 10250
rect 9066 10080 9100 10250
rect 9100 10080 9112 10250
rect 8960 9874 8970 10044
rect 8970 9874 9004 10044
rect 9004 9874 9016 10044
rect 8960 9860 9016 9874
rect 9248 10250 9304 10264
rect 9248 10080 9258 10250
rect 9258 10080 9292 10250
rect 9292 10080 9304 10250
rect 9152 9874 9162 10044
rect 9162 9874 9196 10044
rect 9196 9874 9208 10044
rect 9152 9860 9208 9874
rect 9440 10250 9496 10264
rect 9440 10080 9450 10250
rect 9450 10080 9484 10250
rect 9484 10080 9496 10250
rect 9344 9874 9354 10044
rect 9354 9874 9388 10044
rect 9388 9874 9400 10044
rect 9344 9860 9400 9874
rect 9536 9874 9546 10044
rect 9546 9874 9580 10044
rect 9580 9874 9592 10044
rect 9536 9860 9592 9874
rect 5212 9635 5268 9652
rect 5212 9472 5222 9635
rect 5222 9472 5256 9635
rect 5256 9472 5268 9635
rect 5116 9259 5126 9428
rect 5126 9259 5160 9428
rect 5160 9259 5172 9428
rect 5116 9248 5172 9259
rect 5404 9635 5460 9652
rect 5404 9472 5414 9635
rect 5414 9472 5448 9635
rect 5448 9472 5460 9635
rect 5308 9259 5318 9428
rect 5318 9259 5352 9428
rect 5352 9259 5364 9428
rect 5308 9248 5364 9259
rect 5596 9635 5652 9652
rect 5596 9472 5606 9635
rect 5606 9472 5640 9635
rect 5640 9472 5652 9635
rect 5500 9259 5510 9428
rect 5510 9259 5544 9428
rect 5544 9259 5556 9428
rect 5500 9248 5556 9259
rect 5788 9635 5844 9652
rect 5788 9472 5798 9635
rect 5798 9472 5832 9635
rect 5832 9472 5844 9635
rect 5692 9259 5702 9428
rect 5702 9259 5736 9428
rect 5736 9259 5748 9428
rect 5692 9248 5748 9259
rect 5980 9635 6036 9652
rect 5980 9472 5990 9635
rect 5990 9472 6024 9635
rect 6024 9472 6036 9635
rect 5884 9259 5894 9428
rect 5894 9259 5928 9428
rect 5928 9259 5940 9428
rect 5884 9248 5940 9259
rect 6172 9635 6228 9652
rect 6172 9472 6182 9635
rect 6182 9472 6216 9635
rect 6216 9472 6228 9635
rect 6076 9259 6086 9428
rect 6086 9259 6120 9428
rect 6120 9259 6132 9428
rect 6076 9248 6132 9259
rect 6364 9635 6420 9652
rect 6364 9472 6374 9635
rect 6374 9472 6408 9635
rect 6408 9472 6420 9635
rect 6268 9259 6278 9428
rect 6278 9259 6312 9428
rect 6312 9259 6324 9428
rect 6268 9248 6324 9259
rect 6556 9635 6612 9652
rect 6556 9472 6566 9635
rect 6566 9472 6600 9635
rect 6600 9472 6612 9635
rect 6460 9259 6470 9428
rect 6470 9259 6504 9428
rect 6504 9259 6516 9428
rect 6460 9248 6516 9259
rect 6748 9635 6804 9652
rect 6748 9472 6758 9635
rect 6758 9472 6792 9635
rect 6792 9472 6804 9635
rect 6652 9259 6662 9428
rect 6662 9259 6696 9428
rect 6696 9259 6708 9428
rect 6652 9248 6708 9259
rect 6940 9635 6996 9652
rect 6940 9472 6950 9635
rect 6950 9472 6984 9635
rect 6984 9472 6996 9635
rect 6844 9259 6854 9428
rect 6854 9259 6888 9428
rect 6888 9259 6900 9428
rect 6844 9248 6900 9259
rect 7036 9259 7046 9428
rect 7046 9259 7080 9428
rect 7080 9259 7092 9428
rect 7036 9248 7092 9259
rect 7712 9632 7768 9648
rect 7712 9464 7722 9632
rect 7722 9464 7756 9632
rect 7756 9464 7768 9632
rect 7616 9256 7626 9428
rect 7626 9256 7660 9428
rect 7660 9256 7672 9428
rect 7616 9244 7672 9256
rect 7904 9632 7960 9648
rect 7904 9464 7914 9632
rect 7914 9464 7948 9632
rect 7948 9464 7960 9632
rect 7808 9256 7818 9428
rect 7818 9256 7852 9428
rect 7852 9256 7864 9428
rect 7808 9244 7864 9256
rect 8096 9632 8152 9648
rect 8096 9464 8106 9632
rect 8106 9464 8140 9632
rect 8140 9464 8152 9632
rect 8000 9256 8010 9428
rect 8010 9256 8044 9428
rect 8044 9256 8056 9428
rect 8000 9244 8056 9256
rect 8288 9632 8344 9648
rect 8288 9464 8298 9632
rect 8298 9464 8332 9632
rect 8332 9464 8344 9632
rect 8192 9256 8202 9428
rect 8202 9256 8236 9428
rect 8236 9256 8248 9428
rect 8192 9244 8248 9256
rect 8480 9632 8536 9648
rect 8480 9464 8490 9632
rect 8490 9464 8524 9632
rect 8524 9464 8536 9632
rect 8384 9256 8394 9428
rect 8394 9256 8428 9428
rect 8428 9256 8440 9428
rect 8384 9244 8440 9256
rect 8672 9632 8728 9648
rect 8672 9464 8682 9632
rect 8682 9464 8716 9632
rect 8716 9464 8728 9632
rect 8576 9256 8586 9428
rect 8586 9256 8620 9428
rect 8620 9256 8632 9428
rect 8576 9244 8632 9256
rect 8864 9632 8920 9648
rect 8864 9464 8874 9632
rect 8874 9464 8908 9632
rect 8908 9464 8920 9632
rect 8768 9256 8778 9428
rect 8778 9256 8812 9428
rect 8812 9256 8824 9428
rect 8768 9244 8824 9256
rect 9056 9632 9112 9648
rect 9056 9464 9066 9632
rect 9066 9464 9100 9632
rect 9100 9464 9112 9632
rect 8960 9256 8970 9428
rect 8970 9256 9004 9428
rect 9004 9256 9016 9428
rect 8960 9244 9016 9256
rect 9248 9632 9304 9648
rect 9248 9464 9258 9632
rect 9258 9464 9292 9632
rect 9292 9464 9304 9632
rect 9152 9256 9162 9428
rect 9162 9256 9196 9428
rect 9196 9256 9208 9428
rect 9152 9244 9208 9256
rect 9440 9632 9496 9648
rect 9440 9464 9450 9632
rect 9450 9464 9484 9632
rect 9484 9464 9496 9632
rect 9344 9256 9354 9428
rect 9354 9256 9388 9428
rect 9388 9256 9400 9428
rect 9344 9244 9400 9256
rect 9536 9256 9546 9428
rect 9546 9256 9580 9428
rect 9580 9256 9592 9428
rect 9536 9244 9592 9256
rect 1764 8904 1964 8964
rect 1964 8904 2056 8964
rect 2540 8904 2832 8964
rect 3476 8904 3768 8964
rect -9044 8280 -8904 8356
rect 1776 8718 1828 8732
rect 1776 8552 1786 8718
rect 1786 8552 1820 8718
rect 1820 8552 1828 8718
rect -9964 8222 -9912 8236
rect -9964 8056 -9954 8222
rect -9954 8056 -9920 8222
rect -9920 8056 -9912 8222
rect -10060 7846 -10050 8012
rect -10050 7846 -10016 8012
rect -10016 7846 -10008 8012
rect -10060 7832 -10008 7846
rect -9772 8222 -9720 8236
rect -9772 8056 -9762 8222
rect -9762 8056 -9728 8222
rect -9728 8056 -9720 8222
rect -9868 7846 -9858 8012
rect -9858 7846 -9824 8012
rect -9824 7846 -9816 8012
rect -9868 7832 -9816 7846
rect -9580 8222 -9528 8236
rect -9580 8056 -9570 8222
rect -9570 8056 -9536 8222
rect -9536 8056 -9528 8222
rect -9676 7846 -9666 8012
rect -9666 7846 -9632 8012
rect -9632 7846 -9624 8012
rect -9676 7832 -9624 7846
rect -9388 8222 -9336 8236
rect -9388 8056 -9378 8222
rect -9378 8056 -9344 8222
rect -9344 8056 -9336 8222
rect -9484 7846 -9474 8012
rect -9474 7846 -9440 8012
rect -9440 7846 -9432 8012
rect -9484 7832 -9432 7846
rect -9196 8222 -9144 8236
rect -9196 8056 -9186 8222
rect -9186 8056 -9152 8222
rect -9152 8056 -9144 8222
rect -9292 7846 -9282 8012
rect -9282 7846 -9248 8012
rect -9248 7846 -9240 8012
rect -9292 7832 -9240 7846
rect -9100 7846 -9090 8012
rect -9090 7846 -9056 8012
rect -9056 7846 -9048 8012
rect -9100 7832 -9048 7846
rect -8660 8230 -8480 8296
rect -8660 8196 -8658 8230
rect -8658 8196 -8482 8230
rect -8482 8196 -8480 8230
rect -9964 7604 -9912 7620
rect -9964 7440 -9954 7604
rect -9954 7440 -9920 7604
rect -9920 7440 -9912 7604
rect -10060 7228 -10050 7396
rect -10050 7228 -10016 7396
rect -10016 7228 -10008 7396
rect -10060 7216 -10008 7228
rect -9772 7604 -9720 7620
rect -9772 7440 -9762 7604
rect -9762 7440 -9728 7604
rect -9728 7440 -9720 7604
rect -9868 7228 -9858 7396
rect -9858 7228 -9824 7396
rect -9824 7228 -9816 7396
rect -9868 7216 -9816 7228
rect -9580 7604 -9528 7620
rect -9580 7440 -9570 7604
rect -9570 7440 -9536 7604
rect -9536 7440 -9528 7604
rect -9676 7228 -9666 7396
rect -9666 7228 -9632 7396
rect -9632 7228 -9624 7396
rect -9676 7216 -9624 7228
rect -9388 7604 -9336 7620
rect -9388 7440 -9378 7604
rect -9378 7440 -9344 7604
rect -9344 7440 -9336 7604
rect -9484 7228 -9474 7396
rect -9474 7228 -9440 7396
rect -9440 7228 -9432 7396
rect -9484 7216 -9432 7228
rect -9196 7604 -9144 7620
rect -9196 7440 -9186 7604
rect -9186 7440 -9152 7604
rect -9152 7440 -9144 7604
rect -9292 7228 -9282 7396
rect -9282 7228 -9248 7396
rect -9248 7228 -9240 7396
rect -9292 7216 -9240 7228
rect -9100 7228 -9090 7396
rect -9090 7228 -9056 7396
rect -9056 7228 -9048 7396
rect -9100 7216 -9048 7228
rect 1680 8342 1690 8508
rect 1690 8342 1724 8508
rect 1724 8342 1732 8508
rect 1680 8328 1732 8342
rect 1968 8718 2020 8732
rect 1968 8552 1978 8718
rect 1978 8552 2012 8718
rect 2012 8552 2020 8718
rect 1872 8342 1882 8508
rect 1882 8342 1916 8508
rect 1916 8342 1924 8508
rect 1872 8328 1924 8342
rect 2160 8718 2212 8732
rect 2160 8552 2170 8718
rect 2170 8552 2204 8718
rect 2204 8552 2212 8718
rect 2064 8342 2074 8508
rect 2074 8342 2108 8508
rect 2108 8342 2116 8508
rect 2064 8328 2116 8342
rect 2352 8718 2404 8732
rect 2352 8552 2362 8718
rect 2362 8552 2396 8718
rect 2396 8552 2404 8718
rect 2256 8342 2266 8508
rect 2266 8342 2300 8508
rect 2300 8342 2308 8508
rect 2256 8328 2308 8342
rect 2544 8718 2596 8732
rect 2544 8552 2554 8718
rect 2554 8552 2588 8718
rect 2588 8552 2596 8718
rect 2448 8342 2458 8508
rect 2458 8342 2492 8508
rect 2492 8342 2500 8508
rect 2448 8328 2500 8342
rect 2736 8718 2788 8732
rect 2736 8552 2746 8718
rect 2746 8552 2780 8718
rect 2780 8552 2788 8718
rect 2640 8342 2650 8508
rect 2650 8342 2684 8508
rect 2684 8342 2692 8508
rect 2640 8328 2692 8342
rect 2928 8718 2980 8732
rect 2928 8552 2938 8718
rect 2938 8552 2972 8718
rect 2972 8552 2980 8718
rect 2832 8342 2842 8508
rect 2842 8342 2876 8508
rect 2876 8342 2884 8508
rect 2832 8328 2884 8342
rect 3120 8718 3172 8732
rect 3120 8552 3130 8718
rect 3130 8552 3164 8718
rect 3164 8552 3172 8718
rect 3024 8342 3034 8508
rect 3034 8342 3068 8508
rect 3068 8342 3076 8508
rect 3024 8328 3076 8342
rect 3312 8718 3364 8732
rect 3312 8552 3322 8718
rect 3322 8552 3356 8718
rect 3356 8552 3364 8718
rect 3216 8342 3226 8508
rect 3226 8342 3260 8508
rect 3260 8342 3268 8508
rect 3216 8328 3268 8342
rect 3504 8718 3556 8732
rect 3504 8552 3514 8718
rect 3514 8552 3548 8718
rect 3548 8552 3556 8718
rect 3408 8342 3418 8508
rect 3418 8342 3452 8508
rect 3452 8342 3460 8508
rect 3408 8328 3460 8342
rect 3600 8342 3610 8508
rect 3610 8342 3644 8508
rect 3644 8342 3652 8508
rect 3600 8328 3652 8342
rect 3740 8416 3800 8672
rect 4588 8432 5008 8984
rect 5212 8684 5268 8700
rect 5212 8520 5222 8684
rect 5222 8520 5256 8684
rect 5256 8520 5268 8684
rect 5116 8308 5126 8476
rect 5126 8308 5160 8476
rect 5160 8308 5172 8476
rect 5116 8296 5172 8308
rect 5404 8684 5460 8700
rect 5404 8520 5414 8684
rect 5414 8520 5448 8684
rect 5448 8520 5460 8684
rect 5308 8308 5318 8476
rect 5318 8308 5352 8476
rect 5352 8308 5364 8476
rect 5308 8296 5364 8308
rect 5596 8684 5652 8700
rect 5596 8520 5606 8684
rect 5606 8520 5640 8684
rect 5640 8520 5652 8684
rect 5500 8308 5510 8476
rect 5510 8308 5544 8476
rect 5544 8308 5556 8476
rect 5500 8296 5556 8308
rect 5788 8684 5844 8700
rect 5788 8520 5798 8684
rect 5798 8520 5832 8684
rect 5832 8520 5844 8684
rect 5692 8308 5702 8476
rect 5702 8308 5736 8476
rect 5736 8308 5748 8476
rect 5692 8296 5748 8308
rect 5980 8684 6036 8700
rect 5980 8520 5990 8684
rect 5990 8520 6024 8684
rect 6024 8520 6036 8684
rect 5884 8308 5894 8476
rect 5894 8308 5928 8476
rect 5928 8308 5940 8476
rect 5884 8296 5940 8308
rect 6172 8684 6228 8700
rect 6172 8520 6182 8684
rect 6182 8520 6216 8684
rect 6216 8520 6228 8684
rect 6076 8308 6086 8476
rect 6086 8308 6120 8476
rect 6120 8308 6132 8476
rect 6076 8296 6132 8308
rect 6364 8684 6420 8700
rect 6364 8520 6374 8684
rect 6374 8520 6408 8684
rect 6408 8520 6420 8684
rect 6268 8308 6278 8476
rect 6278 8308 6312 8476
rect 6312 8308 6324 8476
rect 6268 8296 6324 8308
rect 6556 8684 6612 8700
rect 6556 8520 6566 8684
rect 6566 8520 6600 8684
rect 6600 8520 6612 8684
rect 6460 8308 6470 8476
rect 6470 8308 6504 8476
rect 6504 8308 6516 8476
rect 6460 8296 6516 8308
rect 6748 8684 6804 8700
rect 6748 8520 6758 8684
rect 6758 8520 6792 8684
rect 6792 8520 6804 8684
rect 6652 8308 6662 8476
rect 6662 8308 6696 8476
rect 6696 8308 6708 8476
rect 6652 8296 6708 8308
rect 6940 8684 6996 8700
rect 6940 8520 6950 8684
rect 6950 8520 6984 8684
rect 6984 8520 6996 8684
rect 6844 8308 6854 8476
rect 6854 8308 6888 8476
rect 6888 8308 6900 8476
rect 6844 8296 6900 8308
rect 7036 8308 7046 8476
rect 7046 8308 7080 8476
rect 7080 8308 7092 8476
rect 7036 8296 7092 8308
rect 1764 8148 2056 8152
rect 1764 8088 1964 8148
rect 1964 8088 2056 8148
rect 2540 8148 2860 8152
rect 2540 8088 2860 8148
rect 3476 8092 3768 8152
rect 1776 7898 1828 7912
rect 1776 7732 1786 7898
rect 1786 7732 1820 7898
rect 1820 7732 1828 7898
rect 1680 7522 1690 7688
rect 1690 7522 1724 7688
rect 1724 7522 1732 7688
rect 1680 7508 1732 7522
rect 1968 7898 2020 7912
rect 1968 7732 1978 7898
rect 1978 7732 2012 7898
rect 2012 7732 2020 7898
rect 1872 7522 1882 7688
rect 1882 7522 1916 7688
rect 1916 7522 1924 7688
rect 1872 7508 1924 7522
rect 2160 7898 2212 7912
rect 2160 7732 2170 7898
rect 2170 7732 2204 7898
rect 2204 7732 2212 7898
rect 2064 7522 2074 7688
rect 2074 7522 2108 7688
rect 2108 7522 2116 7688
rect 2064 7508 2116 7522
rect 2352 7898 2404 7912
rect 2352 7732 2362 7898
rect 2362 7732 2396 7898
rect 2396 7732 2404 7898
rect 2256 7522 2266 7688
rect 2266 7522 2300 7688
rect 2300 7522 2308 7688
rect 2256 7508 2308 7522
rect 2544 7898 2596 7912
rect 2544 7732 2554 7898
rect 2554 7732 2588 7898
rect 2588 7732 2596 7898
rect 2448 7522 2458 7688
rect 2458 7522 2492 7688
rect 2492 7522 2500 7688
rect 2448 7508 2500 7522
rect 2736 7898 2788 7912
rect 2736 7732 2746 7898
rect 2746 7732 2780 7898
rect 2780 7732 2788 7898
rect 2640 7522 2650 7688
rect 2650 7522 2684 7688
rect 2684 7522 2692 7688
rect 2640 7508 2692 7522
rect 2928 7898 2980 7912
rect 2928 7732 2938 7898
rect 2938 7732 2972 7898
rect 2972 7732 2980 7898
rect 2832 7522 2842 7688
rect 2842 7522 2876 7688
rect 2876 7522 2884 7688
rect 2832 7508 2884 7522
rect 3120 7898 3172 7912
rect 3120 7732 3130 7898
rect 3130 7732 3164 7898
rect 3164 7732 3172 7898
rect 3024 7522 3034 7688
rect 3034 7522 3068 7688
rect 3068 7522 3076 7688
rect 3024 7508 3076 7522
rect 3312 7898 3364 7912
rect 3312 7732 3322 7898
rect 3322 7732 3356 7898
rect 3356 7732 3364 7898
rect 3216 7522 3226 7688
rect 3226 7522 3260 7688
rect 3260 7522 3268 7688
rect 3216 7508 3268 7522
rect 3504 7898 3556 7912
rect 3504 7732 3514 7898
rect 3514 7732 3548 7898
rect 3548 7732 3556 7898
rect 3408 7522 3418 7688
rect 3418 7522 3452 7688
rect 3452 7522 3460 7688
rect 3408 7508 3460 7522
rect 3600 7522 3610 7688
rect 3610 7522 3644 7688
rect 3644 7522 3652 7688
rect 3600 7508 3652 7522
rect 3740 7568 3800 7824
rect 5212 8066 5268 8080
rect 5212 7900 5222 8066
rect 5222 7900 5256 8066
rect 5256 7900 5268 8066
rect 5116 7690 5126 7856
rect 5126 7690 5160 7856
rect 5160 7690 5172 7856
rect 5116 7676 5172 7690
rect 5404 8066 5460 8080
rect 5404 7900 5414 8066
rect 5414 7900 5448 8066
rect 5448 7900 5460 8066
rect 5308 7690 5318 7856
rect 5318 7690 5352 7856
rect 5352 7690 5364 7856
rect 5308 7676 5364 7690
rect 5596 8066 5652 8080
rect 5596 7900 5606 8066
rect 5606 7900 5640 8066
rect 5640 7900 5652 8066
rect 5500 7690 5510 7856
rect 5510 7690 5544 7856
rect 5544 7690 5556 7856
rect 5500 7676 5556 7690
rect 5788 8066 5844 8080
rect 5788 7900 5798 8066
rect 5798 7900 5832 8066
rect 5832 7900 5844 8066
rect 5692 7690 5702 7856
rect 5702 7690 5736 7856
rect 5736 7690 5748 7856
rect 5692 7676 5748 7690
rect 5980 8066 6036 8080
rect 5980 7900 5990 8066
rect 5990 7900 6024 8066
rect 6024 7900 6036 8066
rect 5884 7690 5894 7856
rect 5894 7690 5928 7856
rect 5928 7690 5940 7856
rect 5884 7676 5940 7690
rect 6172 8066 6228 8080
rect 6172 7900 6182 8066
rect 6182 7900 6216 8066
rect 6216 7900 6228 8066
rect 6076 7690 6086 7856
rect 6086 7690 6120 7856
rect 6120 7690 6132 7856
rect 6076 7676 6132 7690
rect 6364 8066 6420 8080
rect 6364 7900 6374 8066
rect 6374 7900 6408 8066
rect 6408 7900 6420 8066
rect 6268 7690 6278 7856
rect 6278 7690 6312 7856
rect 6312 7690 6324 7856
rect 6268 7676 6324 7690
rect 6556 8066 6612 8080
rect 6556 7900 6566 8066
rect 6566 7900 6600 8066
rect 6600 7900 6612 8066
rect 6460 7690 6470 7856
rect 6470 7690 6504 7856
rect 6504 7690 6516 7856
rect 6460 7676 6516 7690
rect 6748 8066 6804 8080
rect 6748 7900 6758 8066
rect 6758 7900 6792 8066
rect 6792 7900 6804 8066
rect 6652 7690 6662 7856
rect 6662 7690 6696 7856
rect 6696 7690 6708 7856
rect 6652 7676 6708 7690
rect 6940 8066 6996 8080
rect 6940 7900 6950 8066
rect 6950 7900 6984 8066
rect 6984 7900 6996 8066
rect 6844 7690 6854 7856
rect 6854 7690 6888 7856
rect 6888 7690 6900 7856
rect 6844 7676 6900 7690
rect 7036 7690 7046 7856
rect 7046 7690 7080 7856
rect 7080 7690 7092 7856
rect 7036 7676 7092 7690
rect 1764 7268 1964 7328
rect 1964 7268 2056 7328
rect 2536 7268 2540 7328
rect 2540 7268 2828 7328
rect 3476 7268 3768 7328
rect -9964 6986 -9912 7000
rect -9964 6820 -9954 6986
rect -9954 6820 -9920 6986
rect -9920 6820 -9912 6986
rect -10060 6610 -10050 6776
rect -10050 6610 -10016 6776
rect -10016 6610 -10008 6776
rect -10060 6596 -10008 6610
rect -9772 6986 -9720 7000
rect -9772 6820 -9762 6986
rect -9762 6820 -9728 6986
rect -9728 6820 -9720 6986
rect -9868 6610 -9858 6776
rect -9858 6610 -9824 6776
rect -9824 6610 -9816 6776
rect -9868 6596 -9816 6610
rect -9580 6986 -9528 7000
rect -9580 6820 -9570 6986
rect -9570 6820 -9536 6986
rect -9536 6820 -9528 6986
rect -9676 6610 -9666 6776
rect -9666 6610 -9632 6776
rect -9632 6610 -9624 6776
rect -9676 6596 -9624 6610
rect -9388 6986 -9336 7000
rect -9388 6820 -9378 6986
rect -9378 6820 -9344 6986
rect -9344 6820 -9336 6986
rect -9484 6610 -9474 6776
rect -9474 6610 -9440 6776
rect -9440 6610 -9432 6776
rect -9484 6596 -9432 6610
rect -9196 6986 -9144 7000
rect -9196 6820 -9186 6986
rect -9186 6820 -9152 6986
rect -9152 6820 -9144 6986
rect -9292 6610 -9282 6776
rect -9282 6610 -9248 6776
rect -9248 6610 -9240 6776
rect -9292 6596 -9240 6610
rect -9100 6610 -9090 6776
rect -9090 6610 -9056 6776
rect -9056 6610 -9048 6776
rect -9100 6596 -9048 6610
rect -8756 6828 -8742 7040
rect -8742 6828 -8708 7040
rect -8708 6828 -8680 7040
rect -8456 6832 -8432 7044
rect -8432 6832 -8398 7044
rect -8398 6832 -8380 7044
rect 1776 7078 1828 7092
rect 1776 6912 1786 7078
rect 1786 6912 1820 7078
rect 1820 6912 1828 7078
rect -8660 6538 -8658 6572
rect -8658 6538 -8482 6572
rect -8482 6538 -8480 6572
rect -8660 6492 -8480 6538
rect 1680 6702 1690 6868
rect 1690 6702 1724 6868
rect 1724 6702 1732 6868
rect 1680 6688 1732 6702
rect 1968 7078 2020 7092
rect 1968 6912 1978 7078
rect 1978 6912 2012 7078
rect 2012 6912 2020 7078
rect 1872 6702 1882 6868
rect 1882 6702 1916 6868
rect 1916 6702 1924 6868
rect 1872 6688 1924 6702
rect 2160 7078 2212 7092
rect 2160 6912 2170 7078
rect 2170 6912 2204 7078
rect 2204 6912 2212 7078
rect 2064 6702 2074 6868
rect 2074 6702 2108 6868
rect 2108 6702 2116 6868
rect 2064 6688 2116 6702
rect 2352 7078 2404 7092
rect 2352 6912 2362 7078
rect 2362 6912 2396 7078
rect 2396 6912 2404 7078
rect 2256 6702 2266 6868
rect 2266 6702 2300 6868
rect 2300 6702 2308 6868
rect 2256 6688 2308 6702
rect 2544 7078 2596 7092
rect 2544 6912 2554 7078
rect 2554 6912 2588 7078
rect 2588 6912 2596 7078
rect 2448 6702 2458 6868
rect 2458 6702 2492 6868
rect 2492 6702 2500 6868
rect 2448 6688 2500 6702
rect 2736 7078 2788 7092
rect 2736 6912 2746 7078
rect 2746 6912 2780 7078
rect 2780 6912 2788 7078
rect 2640 6702 2650 6868
rect 2650 6702 2684 6868
rect 2684 6702 2692 6868
rect 2640 6688 2692 6702
rect 2928 7078 2980 7092
rect 2928 6912 2938 7078
rect 2938 6912 2972 7078
rect 2972 6912 2980 7078
rect 2832 6702 2842 6868
rect 2842 6702 2876 6868
rect 2876 6702 2884 6868
rect 2832 6688 2884 6702
rect 3120 7078 3172 7092
rect 3120 6912 3130 7078
rect 3130 6912 3164 7078
rect 3164 6912 3172 7078
rect 3024 6702 3034 6868
rect 3034 6702 3068 6868
rect 3068 6702 3076 6868
rect 3024 6688 3076 6702
rect 3312 7078 3364 7092
rect 3312 6912 3322 7078
rect 3322 6912 3356 7078
rect 3356 6912 3364 7078
rect 3216 6702 3226 6868
rect 3226 6702 3260 6868
rect 3260 6702 3268 6868
rect 3216 6688 3268 6702
rect 3504 7078 3556 7092
rect 3504 6912 3514 7078
rect 3514 6912 3548 7078
rect 3548 6912 3556 7078
rect 3408 6702 3418 6868
rect 3418 6702 3452 6868
rect 3452 6702 3460 6868
rect 3408 6688 3460 6702
rect 3600 6702 3610 6868
rect 3610 6702 3644 6868
rect 3644 6702 3652 6868
rect 3600 6688 3652 6702
rect 3740 6756 3800 7012
rect 6384 7000 7076 7512
rect 7712 9014 7768 9028
rect 7712 8844 7722 9014
rect 7722 8844 7756 9014
rect 7756 8844 7768 9014
rect 7616 8638 7626 8808
rect 7626 8638 7660 8808
rect 7660 8638 7672 8808
rect 7616 8624 7672 8638
rect 7904 9014 7960 9028
rect 7904 8844 7914 9014
rect 7914 8844 7948 9014
rect 7948 8844 7960 9014
rect 7808 8638 7818 8808
rect 7818 8638 7852 8808
rect 7852 8638 7864 8808
rect 7808 8624 7864 8638
rect 8096 9014 8152 9028
rect 8096 8844 8106 9014
rect 8106 8844 8140 9014
rect 8140 8844 8152 9014
rect 8000 8638 8010 8808
rect 8010 8638 8044 8808
rect 8044 8638 8056 8808
rect 8000 8624 8056 8638
rect 8288 9014 8344 9028
rect 8288 8844 8298 9014
rect 8298 8844 8332 9014
rect 8332 8844 8344 9014
rect 8192 8638 8202 8808
rect 8202 8638 8236 8808
rect 8236 8638 8248 8808
rect 8192 8624 8248 8638
rect 8480 9014 8536 9028
rect 8480 8844 8490 9014
rect 8490 8844 8524 9014
rect 8524 8844 8536 9014
rect 8384 8638 8394 8808
rect 8394 8638 8428 8808
rect 8428 8638 8440 8808
rect 8384 8624 8440 8638
rect 8672 9014 8728 9028
rect 8672 8844 8682 9014
rect 8682 8844 8716 9014
rect 8716 8844 8728 9014
rect 8576 8638 8586 8808
rect 8586 8638 8620 8808
rect 8620 8638 8632 8808
rect 8576 8624 8632 8638
rect 8864 9014 8920 9028
rect 8864 8844 8874 9014
rect 8874 8844 8908 9014
rect 8908 8844 8920 9014
rect 8768 8638 8778 8808
rect 8778 8638 8812 8808
rect 8812 8638 8824 8808
rect 8768 8624 8824 8638
rect 9056 9014 9112 9028
rect 9056 8844 9066 9014
rect 9066 8844 9100 9014
rect 9100 8844 9112 9014
rect 8960 8638 8970 8808
rect 8970 8638 9004 8808
rect 9004 8638 9016 8808
rect 8960 8624 9016 8638
rect 9248 9014 9304 9028
rect 9248 8844 9258 9014
rect 9258 8844 9292 9014
rect 9292 8844 9304 9014
rect 9152 8638 9162 8808
rect 9162 8638 9196 8808
rect 9196 8638 9208 8808
rect 9152 8624 9208 8638
rect 9440 9014 9496 9028
rect 9440 8844 9450 9014
rect 9450 8844 9484 9014
rect 9484 8844 9496 9014
rect 9344 8638 9354 8808
rect 9354 8638 9388 8808
rect 9388 8638 9400 8808
rect 9344 8624 9400 8638
rect 9536 8638 9546 8808
rect 9546 8638 9580 8808
rect 9580 8638 9592 8808
rect 9536 8624 9592 8638
rect 7712 8396 7768 8412
rect 7712 8228 7722 8396
rect 7722 8228 7756 8396
rect 7756 8228 7768 8396
rect 7616 8020 7626 8192
rect 7626 8020 7660 8192
rect 7660 8020 7672 8192
rect 7616 8008 7672 8020
rect 7904 8396 7960 8412
rect 7904 8228 7914 8396
rect 7914 8228 7948 8396
rect 7948 8228 7960 8396
rect 7808 8020 7818 8192
rect 7818 8020 7852 8192
rect 7852 8020 7864 8192
rect 7808 8008 7864 8020
rect 8096 8396 8152 8412
rect 8096 8228 8106 8396
rect 8106 8228 8140 8396
rect 8140 8228 8152 8396
rect 8000 8020 8010 8192
rect 8010 8020 8044 8192
rect 8044 8020 8056 8192
rect 8000 8008 8056 8020
rect 8288 8396 8344 8412
rect 8288 8228 8298 8396
rect 8298 8228 8332 8396
rect 8332 8228 8344 8396
rect 8192 8020 8202 8192
rect 8202 8020 8236 8192
rect 8236 8020 8248 8192
rect 8192 8008 8248 8020
rect 8480 8396 8536 8412
rect 8480 8228 8490 8396
rect 8490 8228 8524 8396
rect 8524 8228 8536 8396
rect 8384 8020 8394 8192
rect 8394 8020 8428 8192
rect 8428 8020 8440 8192
rect 8384 8008 8440 8020
rect 8672 8396 8728 8412
rect 8672 8228 8682 8396
rect 8682 8228 8716 8396
rect 8716 8228 8728 8396
rect 8576 8020 8586 8192
rect 8586 8020 8620 8192
rect 8620 8020 8632 8192
rect 8576 8008 8632 8020
rect 8864 8396 8920 8412
rect 8864 8228 8874 8396
rect 8874 8228 8908 8396
rect 8908 8228 8920 8396
rect 8768 8020 8778 8192
rect 8778 8020 8812 8192
rect 8812 8020 8824 8192
rect 8768 8008 8824 8020
rect 9056 8396 9112 8412
rect 9056 8228 9066 8396
rect 9066 8228 9100 8396
rect 9100 8228 9112 8396
rect 8960 8020 8970 8192
rect 8970 8020 9004 8192
rect 9004 8020 9016 8192
rect 8960 8008 9016 8020
rect 9248 8396 9304 8412
rect 9248 8228 9258 8396
rect 9258 8228 9292 8396
rect 9292 8228 9304 8396
rect 9152 8020 9162 8192
rect 9162 8020 9196 8192
rect 9196 8020 9208 8192
rect 9152 8008 9208 8020
rect 9440 8396 9496 8412
rect 9440 8228 9450 8396
rect 9450 8228 9484 8396
rect 9484 8228 9496 8396
rect 9344 8020 9354 8192
rect 9354 8020 9388 8192
rect 9388 8020 9400 8192
rect 9344 8008 9400 8020
rect 9536 8020 9546 8192
rect 9546 8020 9580 8192
rect 9580 8020 9592 8192
rect 9536 8008 9592 8020
rect 7712 7778 7768 7792
rect 7712 7608 7722 7778
rect 7722 7608 7756 7778
rect 7756 7608 7768 7778
rect 7616 7402 7626 7572
rect 7626 7402 7660 7572
rect 7660 7402 7672 7572
rect 7616 7388 7672 7402
rect 7904 7778 7960 7792
rect 7904 7608 7914 7778
rect 7914 7608 7948 7778
rect 7948 7608 7960 7778
rect 7808 7402 7818 7572
rect 7818 7402 7852 7572
rect 7852 7402 7864 7572
rect 7808 7388 7864 7402
rect 8096 7778 8152 7792
rect 8096 7608 8106 7778
rect 8106 7608 8140 7778
rect 8140 7608 8152 7778
rect 8000 7402 8010 7572
rect 8010 7402 8044 7572
rect 8044 7402 8056 7572
rect 8000 7388 8056 7402
rect 8288 7778 8344 7792
rect 8288 7608 8298 7778
rect 8298 7608 8332 7778
rect 8332 7608 8344 7778
rect 8192 7402 8202 7572
rect 8202 7402 8236 7572
rect 8236 7402 8248 7572
rect 8192 7388 8248 7402
rect 8480 7778 8536 7792
rect 8480 7608 8490 7778
rect 8490 7608 8524 7778
rect 8524 7608 8536 7778
rect 8384 7402 8394 7572
rect 8394 7402 8428 7572
rect 8428 7402 8440 7572
rect 8384 7388 8440 7402
rect 8672 7778 8728 7792
rect 8672 7608 8682 7778
rect 8682 7608 8716 7778
rect 8716 7608 8728 7778
rect 8576 7402 8586 7572
rect 8586 7402 8620 7572
rect 8620 7402 8632 7572
rect 8576 7388 8632 7402
rect 8864 7778 8920 7792
rect 8864 7608 8874 7778
rect 8874 7608 8908 7778
rect 8908 7608 8920 7778
rect 8768 7402 8778 7572
rect 8778 7402 8812 7572
rect 8812 7402 8824 7572
rect 8768 7388 8824 7402
rect 9056 7778 9112 7792
rect 9056 7608 9066 7778
rect 9066 7608 9100 7778
rect 9100 7608 9112 7778
rect 8960 7402 8970 7572
rect 8970 7402 9004 7572
rect 9004 7402 9016 7572
rect 8960 7388 9016 7402
rect 9248 7778 9304 7792
rect 9248 7608 9258 7778
rect 9258 7608 9292 7778
rect 9292 7608 9304 7778
rect 9152 7402 9162 7572
rect 9162 7402 9196 7572
rect 9196 7402 9208 7572
rect 9152 7388 9208 7402
rect 9440 7778 9496 7792
rect 9440 7608 9450 7778
rect 9450 7608 9484 7778
rect 9484 7608 9496 7778
rect 9344 7402 9354 7572
rect 9354 7402 9388 7572
rect 9388 7402 9400 7572
rect 9344 7388 9400 7402
rect 9536 7402 9546 7572
rect 9546 7402 9580 7572
rect 9580 7402 9592 7572
rect 9536 7388 9592 7402
rect 7712 7160 7768 7176
rect 7712 6992 7722 7160
rect 7722 6992 7756 7160
rect 7756 6992 7768 7160
rect 7000 6600 7528 6928
rect 7616 6784 7626 6956
rect 7626 6784 7660 6956
rect 7660 6784 7672 6956
rect 7616 6772 7672 6784
rect 7904 7160 7960 7176
rect 7904 6992 7914 7160
rect 7914 6992 7948 7160
rect 7948 6992 7960 7160
rect 7808 6784 7818 6956
rect 7818 6784 7852 6956
rect 7852 6784 7864 6956
rect 7808 6772 7864 6784
rect 8096 7160 8152 7176
rect 8096 6992 8106 7160
rect 8106 6992 8140 7160
rect 8140 6992 8152 7160
rect 8000 6784 8010 6956
rect 8010 6784 8044 6956
rect 8044 6784 8056 6956
rect 8000 6772 8056 6784
rect 8288 7160 8344 7176
rect 8288 6992 8298 7160
rect 8298 6992 8332 7160
rect 8332 6992 8344 7160
rect 8192 6784 8202 6956
rect 8202 6784 8236 6956
rect 8236 6784 8248 6956
rect 8192 6772 8248 6784
rect 8480 7160 8536 7176
rect 8480 6992 8490 7160
rect 8490 6992 8524 7160
rect 8524 6992 8536 7160
rect 8384 6784 8394 6956
rect 8394 6784 8428 6956
rect 8428 6784 8440 6956
rect 8384 6772 8440 6784
rect 8672 7160 8728 7176
rect 8672 6992 8682 7160
rect 8682 6992 8716 7160
rect 8716 6992 8728 7160
rect 8576 6784 8586 6956
rect 8586 6784 8620 6956
rect 8620 6784 8632 6956
rect 8576 6772 8632 6784
rect 8864 7160 8920 7176
rect 8864 6992 8874 7160
rect 8874 6992 8908 7160
rect 8908 6992 8920 7160
rect 8768 6784 8778 6956
rect 8778 6784 8812 6956
rect 8812 6784 8824 6956
rect 8768 6772 8824 6784
rect 9056 7160 9112 7176
rect 9056 6992 9066 7160
rect 9066 6992 9100 7160
rect 9100 6992 9112 7160
rect 8960 6784 8970 6956
rect 8970 6784 9004 6956
rect 9004 6784 9016 6956
rect 8960 6772 9016 6784
rect 9248 7160 9304 7176
rect 9248 6992 9258 7160
rect 9258 6992 9292 7160
rect 9292 6992 9304 7160
rect 9152 6784 9162 6956
rect 9162 6784 9196 6956
rect 9196 6784 9208 6956
rect 9152 6772 9208 6784
rect 9440 7160 9496 7176
rect 9440 6992 9450 7160
rect 9450 6992 9484 7160
rect 9484 6992 9496 7160
rect 9344 6784 9354 6956
rect 9354 6784 9388 6956
rect 9388 6784 9400 6956
rect 9344 6772 9400 6784
rect 9536 6784 9546 6956
rect 9546 6784 9580 6956
rect 9580 6784 9592 6956
rect 9536 6772 9592 6784
rect 1672 6456 1964 6516
rect 2540 6456 2832 6516
rect 3476 6452 3768 6512
rect -9964 6142 -9912 6156
rect -9964 5976 -9954 6142
rect -9954 5976 -9920 6142
rect -9920 5976 -9912 6142
rect -10060 5766 -10050 5932
rect -10050 5766 -10016 5932
rect -10016 5766 -10008 5932
rect -10060 5752 -10008 5766
rect -9772 6142 -9720 6156
rect -9772 5976 -9762 6142
rect -9762 5976 -9728 6142
rect -9728 5976 -9720 6142
rect -9868 5766 -9858 5932
rect -9858 5766 -9824 5932
rect -9824 5766 -9816 5932
rect -9868 5752 -9816 5766
rect -9580 6142 -9528 6156
rect -9580 5976 -9570 6142
rect -9570 5976 -9536 6142
rect -9536 5976 -9528 6142
rect -9676 5766 -9666 5932
rect -9666 5766 -9632 5932
rect -9632 5766 -9624 5932
rect -9676 5752 -9624 5766
rect -9388 6142 -9336 6156
rect -9388 5976 -9378 6142
rect -9378 5976 -9344 6142
rect -9344 5976 -9336 6142
rect -9484 5766 -9474 5932
rect -9474 5766 -9440 5932
rect -9440 5766 -9432 5932
rect -9484 5752 -9432 5766
rect -9196 6142 -9144 6156
rect -9196 5976 -9186 6142
rect -9186 5976 -9152 6142
rect -9152 5976 -9144 6142
rect -9292 5766 -9282 5932
rect -9282 5766 -9248 5932
rect -9248 5766 -9240 5932
rect -9292 5752 -9240 5766
rect -8992 5988 -8824 6164
rect 6960 6156 7456 6472
rect 7712 6542 7768 6556
rect 7712 6372 7722 6542
rect 7722 6372 7756 6542
rect 7756 6372 7768 6542
rect 7616 6166 7626 6336
rect 7626 6166 7660 6336
rect 7660 6166 7672 6336
rect 7616 6152 7672 6166
rect 7904 6542 7960 6556
rect 7904 6372 7914 6542
rect 7914 6372 7948 6542
rect 7948 6372 7960 6542
rect 7808 6166 7818 6336
rect 7818 6166 7852 6336
rect 7852 6166 7864 6336
rect 7808 6152 7864 6166
rect 8096 6542 8152 6556
rect 8096 6372 8106 6542
rect 8106 6372 8140 6542
rect 8140 6372 8152 6542
rect 8000 6166 8010 6336
rect 8010 6166 8044 6336
rect 8044 6166 8056 6336
rect 8000 6152 8056 6166
rect 8288 6542 8344 6556
rect 8288 6372 8298 6542
rect 8298 6372 8332 6542
rect 8332 6372 8344 6542
rect 8192 6166 8202 6336
rect 8202 6166 8236 6336
rect 8236 6166 8248 6336
rect 8192 6152 8248 6166
rect 8480 6542 8536 6556
rect 8480 6372 8490 6542
rect 8490 6372 8524 6542
rect 8524 6372 8536 6542
rect 8384 6166 8394 6336
rect 8394 6166 8428 6336
rect 8428 6166 8440 6336
rect 8384 6152 8440 6166
rect 8672 6542 8728 6556
rect 8672 6372 8682 6542
rect 8682 6372 8716 6542
rect 8716 6372 8728 6542
rect 8576 6166 8586 6336
rect 8586 6166 8620 6336
rect 8620 6166 8632 6336
rect 8576 6152 8632 6166
rect 8864 6542 8920 6556
rect 8864 6372 8874 6542
rect 8874 6372 8908 6542
rect 8908 6372 8920 6542
rect 8768 6166 8778 6336
rect 8778 6166 8812 6336
rect 8812 6166 8824 6336
rect 8768 6152 8824 6166
rect 9056 6542 9112 6556
rect 9056 6372 9066 6542
rect 9066 6372 9100 6542
rect 9100 6372 9112 6542
rect 8960 6166 8970 6336
rect 8970 6166 9004 6336
rect 9004 6166 9016 6336
rect 8960 6152 9016 6166
rect 9248 6542 9304 6556
rect 9248 6372 9258 6542
rect 9258 6372 9292 6542
rect 9292 6372 9304 6542
rect 9152 6166 9162 6336
rect 9162 6166 9196 6336
rect 9196 6166 9208 6336
rect 9152 6152 9208 6166
rect 9440 6542 9496 6556
rect 9440 6372 9450 6542
rect 9450 6372 9484 6542
rect 9484 6372 9496 6542
rect 9344 6166 9354 6336
rect 9354 6166 9388 6336
rect 9388 6166 9400 6336
rect 9344 6152 9400 6166
rect 9536 6166 9546 6336
rect 9546 6166 9580 6336
rect 9580 6166 9592 6336
rect 9536 6152 9592 6166
rect -9100 5766 -9090 5932
rect -9090 5766 -9056 5932
rect -9056 5766 -9048 5932
rect -9100 5752 -9048 5766
rect -9964 5524 -9912 5540
rect -9964 5360 -9954 5524
rect -9954 5360 -9920 5524
rect -9920 5360 -9912 5524
rect -10060 5148 -10050 5316
rect -10050 5148 -10016 5316
rect -10016 5148 -10008 5316
rect -10060 5136 -10008 5148
rect -9772 5524 -9720 5540
rect -9772 5360 -9762 5524
rect -9762 5360 -9728 5524
rect -9728 5360 -9720 5524
rect -9868 5148 -9858 5316
rect -9858 5148 -9824 5316
rect -9824 5148 -9816 5316
rect -9868 5136 -9816 5148
rect -9580 5524 -9528 5540
rect -9580 5360 -9570 5524
rect -9570 5360 -9536 5524
rect -9536 5360 -9528 5524
rect -9676 5148 -9666 5316
rect -9666 5148 -9632 5316
rect -9632 5148 -9624 5316
rect -9676 5136 -9624 5148
rect -9388 5524 -9336 5540
rect -9388 5360 -9378 5524
rect -9378 5360 -9344 5524
rect -9344 5360 -9336 5524
rect -9484 5148 -9474 5316
rect -9474 5148 -9440 5316
rect -9440 5148 -9432 5316
rect -9484 5136 -9432 5148
rect -9196 5524 -9144 5540
rect -9196 5360 -9186 5524
rect -9186 5360 -9152 5524
rect -9152 5360 -9144 5524
rect -9292 5148 -9282 5316
rect -9282 5148 -9248 5316
rect -9248 5148 -9240 5316
rect -9292 5136 -9240 5148
rect -9100 5148 -9090 5316
rect -9090 5148 -9056 5316
rect -9056 5148 -9048 5316
rect -9100 5136 -9048 5148
rect 312 5862 364 5876
rect 312 5696 322 5862
rect 322 5696 356 5862
rect 356 5696 364 5862
rect 216 5486 226 5652
rect 226 5486 260 5652
rect 260 5486 268 5652
rect 216 5472 268 5486
rect 504 5862 556 5876
rect 504 5696 514 5862
rect 514 5696 548 5862
rect 548 5696 556 5862
rect 408 5486 418 5652
rect 418 5486 452 5652
rect 452 5486 460 5652
rect 408 5472 460 5486
rect 696 5862 748 5876
rect 696 5696 706 5862
rect 706 5696 740 5862
rect 740 5696 748 5862
rect 600 5486 610 5652
rect 610 5486 644 5652
rect 644 5486 652 5652
rect 600 5472 652 5486
rect 888 5862 940 5876
rect 888 5696 898 5862
rect 898 5696 932 5862
rect 932 5696 940 5862
rect 792 5486 802 5652
rect 802 5486 836 5652
rect 836 5486 844 5652
rect 792 5472 844 5486
rect 1080 5862 1132 5876
rect 1080 5696 1090 5862
rect 1090 5696 1124 5862
rect 1124 5696 1132 5862
rect 984 5486 994 5652
rect 994 5486 1028 5652
rect 1028 5486 1036 5652
rect 984 5472 1036 5486
rect 1176 5486 1186 5652
rect 1186 5486 1220 5652
rect 1220 5486 1228 5652
rect 1176 5472 1228 5486
rect 2112 5862 2164 5876
rect 2112 5696 2122 5862
rect 2122 5696 2156 5862
rect 2156 5696 2164 5862
rect 2016 5486 2026 5652
rect 2026 5486 2060 5652
rect 2060 5486 2068 5652
rect 2016 5472 2068 5486
rect 2304 5862 2356 5876
rect 2304 5696 2314 5862
rect 2314 5696 2348 5862
rect 2348 5696 2356 5862
rect 2208 5486 2218 5652
rect 2218 5486 2252 5652
rect 2252 5486 2260 5652
rect 2208 5472 2260 5486
rect 2496 5862 2548 5876
rect 2496 5696 2506 5862
rect 2506 5696 2540 5862
rect 2540 5696 2548 5862
rect 2400 5486 2410 5652
rect 2410 5486 2444 5652
rect 2444 5486 2452 5652
rect 2400 5472 2452 5486
rect 2688 5862 2740 5876
rect 2688 5696 2698 5862
rect 2698 5696 2732 5862
rect 2732 5696 2740 5862
rect 2592 5486 2602 5652
rect 2602 5486 2636 5652
rect 2636 5486 2644 5652
rect 2592 5472 2644 5486
rect 2880 5862 2932 5876
rect 2880 5696 2890 5862
rect 2890 5696 2924 5862
rect 2924 5696 2932 5862
rect 2784 5486 2794 5652
rect 2794 5486 2828 5652
rect 2828 5486 2836 5652
rect 2784 5472 2836 5486
rect 2976 5486 2986 5652
rect 2986 5486 3020 5652
rect 3020 5486 3028 5652
rect 2976 5472 3028 5486
rect 3912 5862 3964 5876
rect 3912 5696 3922 5862
rect 3922 5696 3956 5862
rect 3956 5696 3964 5862
rect 3816 5486 3826 5652
rect 3826 5486 3860 5652
rect 3860 5486 3868 5652
rect 3816 5472 3868 5486
rect 4104 5862 4156 5876
rect 4104 5696 4114 5862
rect 4114 5696 4148 5862
rect 4148 5696 4156 5862
rect 4008 5486 4018 5652
rect 4018 5486 4052 5652
rect 4052 5486 4060 5652
rect 4008 5472 4060 5486
rect 4296 5862 4348 5876
rect 4296 5696 4306 5862
rect 4306 5696 4340 5862
rect 4340 5696 4348 5862
rect 4200 5486 4210 5652
rect 4210 5486 4244 5652
rect 4244 5486 4252 5652
rect 4200 5472 4252 5486
rect 4488 5862 4540 5876
rect 4488 5696 4498 5862
rect 4498 5696 4532 5862
rect 4532 5696 4540 5862
rect 4392 5486 4402 5652
rect 4402 5486 4436 5652
rect 4436 5486 4444 5652
rect 4392 5472 4444 5486
rect 4680 5862 4732 5876
rect 4680 5696 4690 5862
rect 4690 5696 4724 5862
rect 4724 5696 4732 5862
rect 4584 5486 4594 5652
rect 4594 5486 4628 5652
rect 4628 5486 4636 5652
rect 4584 5472 4636 5486
rect 4776 5486 4786 5652
rect 4786 5486 4820 5652
rect 4820 5486 4828 5652
rect 4776 5472 4828 5486
rect 5712 5862 5764 5876
rect 5712 5696 5722 5862
rect 5722 5696 5756 5862
rect 5756 5696 5764 5862
rect 5616 5486 5626 5652
rect 5626 5486 5660 5652
rect 5660 5486 5668 5652
rect 5616 5472 5668 5486
rect 5904 5862 5956 5876
rect 5904 5696 5914 5862
rect 5914 5696 5948 5862
rect 5948 5696 5956 5862
rect 5808 5486 5818 5652
rect 5818 5486 5852 5652
rect 5852 5486 5860 5652
rect 5808 5472 5860 5486
rect 6096 5862 6148 5876
rect 6096 5696 6106 5862
rect 6106 5696 6140 5862
rect 6140 5696 6148 5862
rect 6000 5486 6010 5652
rect 6010 5486 6044 5652
rect 6044 5486 6052 5652
rect 6000 5472 6052 5486
rect 6288 5862 6340 5876
rect 6288 5696 6298 5862
rect 6298 5696 6332 5862
rect 6332 5696 6340 5862
rect 6192 5486 6202 5652
rect 6202 5486 6236 5652
rect 6236 5486 6244 5652
rect 6192 5472 6244 5486
rect 6480 5862 6532 5876
rect 6480 5696 6490 5862
rect 6490 5696 6524 5862
rect 6524 5696 6532 5862
rect 6384 5486 6394 5652
rect 6394 5486 6428 5652
rect 6428 5486 6436 5652
rect 6384 5472 6436 5486
rect 6576 5486 6586 5652
rect 6586 5486 6620 5652
rect 6620 5486 6628 5652
rect 6576 5472 6628 5486
rect 7088 5580 7372 6080
rect 7712 5924 7768 5940
rect 7712 5756 7722 5924
rect 7722 5756 7756 5924
rect 7756 5756 7768 5924
rect -9964 4906 -9912 4920
rect -9964 4740 -9954 4906
rect -9954 4740 -9920 4906
rect -9920 4740 -9912 4906
rect -10060 4530 -10050 4696
rect -10050 4530 -10016 4696
rect -10016 4530 -10008 4696
rect -10060 4516 -10008 4530
rect -9772 4906 -9720 4920
rect -9772 4740 -9762 4906
rect -9762 4740 -9728 4906
rect -9728 4740 -9720 4906
rect -9868 4530 -9858 4696
rect -9858 4530 -9824 4696
rect -9824 4530 -9816 4696
rect -9868 4516 -9816 4530
rect -9580 4906 -9528 4920
rect -9580 4740 -9570 4906
rect -9570 4740 -9536 4906
rect -9536 4740 -9528 4906
rect -9676 4530 -9666 4696
rect -9666 4530 -9632 4696
rect -9632 4530 -9624 4696
rect -9676 4516 -9624 4530
rect -9388 4906 -9336 4920
rect -9388 4740 -9378 4906
rect -9378 4740 -9344 4906
rect -9344 4740 -9336 4906
rect -9484 4530 -9474 4696
rect -9474 4530 -9440 4696
rect -9440 4530 -9432 4696
rect -9484 4516 -9432 4530
rect -9196 4906 -9144 4920
rect -9196 4740 -9186 4906
rect -9186 4740 -9152 4906
rect -9152 4740 -9144 4906
rect -9292 4530 -9282 4696
rect -9282 4530 -9248 4696
rect -9248 4530 -9240 4696
rect -9292 4516 -9240 4530
rect -9100 4530 -9090 4696
rect -9090 4530 -9056 4696
rect -9056 4530 -9048 4696
rect -9100 4516 -9048 4530
rect -3172 4420 -3028 4532
rect -404 4400 28 5092
rect 312 5244 364 5260
rect 312 5080 322 5244
rect 322 5080 356 5244
rect 356 5080 364 5244
rect 216 4868 226 5036
rect 226 4868 260 5036
rect 260 4868 268 5036
rect 216 4856 268 4868
rect 504 5244 556 5260
rect 504 5080 514 5244
rect 514 5080 548 5244
rect 548 5080 556 5244
rect 408 4868 418 5036
rect 418 4868 452 5036
rect 452 4868 460 5036
rect 408 4856 460 4868
rect 696 5244 748 5260
rect 696 5080 706 5244
rect 706 5080 740 5244
rect 740 5080 748 5244
rect 600 4868 610 5036
rect 610 4868 644 5036
rect 644 4868 652 5036
rect 600 4856 652 4868
rect 888 5244 940 5260
rect 888 5080 898 5244
rect 898 5080 932 5244
rect 932 5080 940 5244
rect 792 4868 802 5036
rect 802 4868 836 5036
rect 836 4868 844 5036
rect 792 4856 844 4868
rect 1080 5244 1132 5260
rect 1080 5080 1090 5244
rect 1090 5080 1124 5244
rect 1124 5080 1132 5244
rect 984 4868 994 5036
rect 994 4868 1028 5036
rect 1028 4868 1036 5036
rect 984 4856 1036 4868
rect 1176 4868 1186 5036
rect 1186 4868 1220 5036
rect 1220 4868 1228 5036
rect 1176 4856 1228 4868
rect 2112 5244 2164 5260
rect 2112 5080 2122 5244
rect 2122 5080 2156 5244
rect 2156 5080 2164 5244
rect 2016 4868 2026 5036
rect 2026 4868 2060 5036
rect 2060 4868 2068 5036
rect 2016 4856 2068 4868
rect 2304 5244 2356 5260
rect 2304 5080 2314 5244
rect 2314 5080 2348 5244
rect 2348 5080 2356 5244
rect 2208 4868 2218 5036
rect 2218 4868 2252 5036
rect 2252 4868 2260 5036
rect 2208 4856 2260 4868
rect 2496 5244 2548 5260
rect 2496 5080 2506 5244
rect 2506 5080 2540 5244
rect 2540 5080 2548 5244
rect 2400 4868 2410 5036
rect 2410 4868 2444 5036
rect 2444 4868 2452 5036
rect 2400 4856 2452 4868
rect 2688 5244 2740 5260
rect 2688 5080 2698 5244
rect 2698 5080 2732 5244
rect 2732 5080 2740 5244
rect 2592 4868 2602 5036
rect 2602 4868 2636 5036
rect 2636 4868 2644 5036
rect 2592 4856 2644 4868
rect 2880 5244 2932 5260
rect 2880 5080 2890 5244
rect 2890 5080 2924 5244
rect 2924 5080 2932 5244
rect 2784 4868 2794 5036
rect 2794 4868 2828 5036
rect 2828 4868 2836 5036
rect 2784 4856 2836 4868
rect 2976 4868 2986 5036
rect 2986 4868 3020 5036
rect 3020 4868 3028 5036
rect 2976 4856 3028 4868
rect 3912 5244 3964 5260
rect 3912 5080 3922 5244
rect 3922 5080 3956 5244
rect 3956 5080 3964 5244
rect 3816 4868 3826 5036
rect 3826 4868 3860 5036
rect 3860 4868 3868 5036
rect 3816 4856 3868 4868
rect 4104 5244 4156 5260
rect 4104 5080 4114 5244
rect 4114 5080 4148 5244
rect 4148 5080 4156 5244
rect 4008 4868 4018 5036
rect 4018 4868 4052 5036
rect 4052 4868 4060 5036
rect 4008 4856 4060 4868
rect 4296 5244 4348 5260
rect 4296 5080 4306 5244
rect 4306 5080 4340 5244
rect 4340 5080 4348 5244
rect 4200 4868 4210 5036
rect 4210 4868 4244 5036
rect 4244 4868 4252 5036
rect 4200 4856 4252 4868
rect 4488 5244 4540 5260
rect 4488 5080 4498 5244
rect 4498 5080 4532 5244
rect 4532 5080 4540 5244
rect 4392 4868 4402 5036
rect 4402 4868 4436 5036
rect 4436 4868 4444 5036
rect 4392 4856 4444 4868
rect 4680 5244 4732 5260
rect 4680 5080 4690 5244
rect 4690 5080 4724 5244
rect 4724 5080 4732 5244
rect 4584 4868 4594 5036
rect 4594 4868 4628 5036
rect 4628 4868 4636 5036
rect 4584 4856 4636 4868
rect 4776 4868 4786 5036
rect 4786 4868 4820 5036
rect 4820 4868 4828 5036
rect 4776 4856 4828 4868
rect 5712 5244 5764 5260
rect 5712 5080 5722 5244
rect 5722 5080 5756 5244
rect 5756 5080 5764 5244
rect 5616 4868 5626 5036
rect 5626 4868 5660 5036
rect 5660 4868 5668 5036
rect 5616 4856 5668 4868
rect 5904 5244 5956 5260
rect 5904 5080 5914 5244
rect 5914 5080 5948 5244
rect 5948 5080 5956 5244
rect 5808 4868 5818 5036
rect 5818 4868 5852 5036
rect 5852 4868 5860 5036
rect 5808 4856 5860 4868
rect 6096 5244 6148 5260
rect 6096 5080 6106 5244
rect 6106 5080 6140 5244
rect 6140 5080 6148 5244
rect 6000 4868 6010 5036
rect 6010 4868 6044 5036
rect 6044 4868 6052 5036
rect 6000 4856 6052 4868
rect 6288 5244 6340 5260
rect 6288 5080 6298 5244
rect 6298 5080 6332 5244
rect 6332 5080 6340 5244
rect 6192 4868 6202 5036
rect 6202 4868 6236 5036
rect 6236 4868 6244 5036
rect 6192 4856 6244 4868
rect 6480 5244 6532 5260
rect 6480 5080 6490 5244
rect 6490 5080 6524 5244
rect 6524 5080 6532 5244
rect 6384 4868 6394 5036
rect 6394 4868 6428 5036
rect 6428 4868 6436 5036
rect 6384 4856 6436 4868
rect 6576 4868 6586 5036
rect 6586 4868 6620 5036
rect 6620 4868 6628 5036
rect 6576 4856 6628 4868
rect 7616 5548 7626 5720
rect 7626 5548 7660 5720
rect 7660 5548 7672 5720
rect 7616 5536 7672 5548
rect 7904 5924 7960 5940
rect 7904 5756 7914 5924
rect 7914 5756 7948 5924
rect 7948 5756 7960 5924
rect 7808 5548 7818 5720
rect 7818 5548 7852 5720
rect 7852 5548 7864 5720
rect 7808 5536 7864 5548
rect 8096 5924 8152 5940
rect 8096 5756 8106 5924
rect 8106 5756 8140 5924
rect 8140 5756 8152 5924
rect 8000 5548 8010 5720
rect 8010 5548 8044 5720
rect 8044 5548 8056 5720
rect 8000 5536 8056 5548
rect 8288 5924 8344 5940
rect 8288 5756 8298 5924
rect 8298 5756 8332 5924
rect 8332 5756 8344 5924
rect 8192 5548 8202 5720
rect 8202 5548 8236 5720
rect 8236 5548 8248 5720
rect 8192 5536 8248 5548
rect 8480 5924 8536 5940
rect 8480 5756 8490 5924
rect 8490 5756 8524 5924
rect 8524 5756 8536 5924
rect 8384 5548 8394 5720
rect 8394 5548 8428 5720
rect 8428 5548 8440 5720
rect 8384 5536 8440 5548
rect 8672 5924 8728 5940
rect 8672 5756 8682 5924
rect 8682 5756 8716 5924
rect 8716 5756 8728 5924
rect 8576 5548 8586 5720
rect 8586 5548 8620 5720
rect 8620 5548 8632 5720
rect 8576 5536 8632 5548
rect 8864 5924 8920 5940
rect 8864 5756 8874 5924
rect 8874 5756 8908 5924
rect 8908 5756 8920 5924
rect 8768 5548 8778 5720
rect 8778 5548 8812 5720
rect 8812 5548 8824 5720
rect 8768 5536 8824 5548
rect 9056 5924 9112 5940
rect 9056 5756 9066 5924
rect 9066 5756 9100 5924
rect 9100 5756 9112 5924
rect 8960 5548 8970 5720
rect 8970 5548 9004 5720
rect 9004 5548 9016 5720
rect 8960 5536 9016 5548
rect 9248 5924 9304 5940
rect 9248 5756 9258 5924
rect 9258 5756 9292 5924
rect 9292 5756 9304 5924
rect 9152 5548 9162 5720
rect 9162 5548 9196 5720
rect 9196 5548 9208 5720
rect 9152 5536 9208 5548
rect 9440 5924 9496 5940
rect 9440 5756 9450 5924
rect 9450 5756 9484 5924
rect 9484 5756 9496 5924
rect 9344 5548 9354 5720
rect 9354 5548 9388 5720
rect 9388 5548 9400 5720
rect 9344 5536 9400 5548
rect 9536 5548 9546 5720
rect 9546 5548 9580 5720
rect 9580 5548 9592 5720
rect 9536 5536 9592 5548
rect 7712 5306 7768 5320
rect 7712 5136 7722 5306
rect 7722 5136 7756 5306
rect 7756 5136 7768 5306
rect 7616 4930 7626 5100
rect 7626 4930 7660 5100
rect 7660 4930 7672 5100
rect 7616 4916 7672 4930
rect 7904 5306 7960 5320
rect 7904 5136 7914 5306
rect 7914 5136 7948 5306
rect 7948 5136 7960 5306
rect 7808 4930 7818 5100
rect 7818 4930 7852 5100
rect 7852 4930 7864 5100
rect 7808 4916 7864 4930
rect 8096 5306 8152 5320
rect 8096 5136 8106 5306
rect 8106 5136 8140 5306
rect 8140 5136 8152 5306
rect 8000 4930 8010 5100
rect 8010 4930 8044 5100
rect 8044 4930 8056 5100
rect 8000 4916 8056 4930
rect 8288 5306 8344 5320
rect 8288 5136 8298 5306
rect 8298 5136 8332 5306
rect 8332 5136 8344 5306
rect 8192 4930 8202 5100
rect 8202 4930 8236 5100
rect 8236 4930 8248 5100
rect 8192 4916 8248 4930
rect 8480 5306 8536 5320
rect 8480 5136 8490 5306
rect 8490 5136 8524 5306
rect 8524 5136 8536 5306
rect 8384 4930 8394 5100
rect 8394 4930 8428 5100
rect 8428 4930 8440 5100
rect 8384 4916 8440 4930
rect 8672 5306 8728 5320
rect 8672 5136 8682 5306
rect 8682 5136 8716 5306
rect 8716 5136 8728 5306
rect 8576 4930 8586 5100
rect 8586 4930 8620 5100
rect 8620 4930 8632 5100
rect 8576 4916 8632 4930
rect 8864 5306 8920 5320
rect 8864 5136 8874 5306
rect 8874 5136 8908 5306
rect 8908 5136 8920 5306
rect 8768 4930 8778 5100
rect 8778 4930 8812 5100
rect 8812 4930 8824 5100
rect 8768 4916 8824 4930
rect 9056 5306 9112 5320
rect 9056 5136 9066 5306
rect 9066 5136 9100 5306
rect 9100 5136 9112 5306
rect 8960 4930 8970 5100
rect 8970 4930 9004 5100
rect 9004 4930 9016 5100
rect 8960 4916 9016 4930
rect 9248 5306 9304 5320
rect 9248 5136 9258 5306
rect 9258 5136 9292 5306
rect 9292 5136 9304 5306
rect 9152 4930 9162 5100
rect 9162 4930 9196 5100
rect 9196 4930 9208 5100
rect 9152 4916 9208 4930
rect 9440 5306 9496 5320
rect 9440 5136 9450 5306
rect 9450 5136 9484 5306
rect 9484 5136 9496 5306
rect 9344 4930 9354 5100
rect 9354 4930 9388 5100
rect 9388 4930 9400 5100
rect 9344 4916 9400 4930
rect 9536 4930 9546 5100
rect 9546 4930 9580 5100
rect 9580 4930 9592 5100
rect 9536 4916 9592 4930
rect 312 4626 364 4640
rect 312 4460 322 4626
rect 322 4460 356 4626
rect 356 4460 364 4626
rect 216 4250 226 4416
rect 226 4250 260 4416
rect 260 4250 268 4416
rect 216 4236 268 4250
rect 504 4626 556 4640
rect 504 4460 514 4626
rect 514 4460 548 4626
rect 548 4460 556 4626
rect 408 4250 418 4416
rect 418 4250 452 4416
rect 452 4250 460 4416
rect 408 4236 460 4250
rect 696 4626 748 4640
rect 696 4460 706 4626
rect 706 4460 740 4626
rect 740 4460 748 4626
rect 600 4250 610 4416
rect 610 4250 644 4416
rect 644 4250 652 4416
rect 600 4236 652 4250
rect 888 4626 940 4640
rect 888 4460 898 4626
rect 898 4460 932 4626
rect 932 4460 940 4626
rect 792 4250 802 4416
rect 802 4250 836 4416
rect 836 4250 844 4416
rect 792 4236 844 4250
rect 1080 4626 1132 4640
rect 1080 4460 1090 4626
rect 1090 4460 1124 4626
rect 1124 4460 1132 4626
rect 984 4250 994 4416
rect 994 4250 1028 4416
rect 1028 4250 1036 4416
rect 984 4236 1036 4250
rect 1176 4250 1186 4416
rect 1186 4250 1220 4416
rect 1220 4250 1228 4416
rect 1176 4236 1228 4250
rect 2112 4626 2164 4640
rect 2112 4460 2122 4626
rect 2122 4460 2156 4626
rect 2156 4460 2164 4626
rect 2016 4250 2026 4416
rect 2026 4250 2060 4416
rect 2060 4250 2068 4416
rect 2016 4236 2068 4250
rect 2304 4626 2356 4640
rect 2304 4460 2314 4626
rect 2314 4460 2348 4626
rect 2348 4460 2356 4626
rect 2208 4250 2218 4416
rect 2218 4250 2252 4416
rect 2252 4250 2260 4416
rect 2208 4236 2260 4250
rect 2496 4626 2548 4640
rect 2496 4460 2506 4626
rect 2506 4460 2540 4626
rect 2540 4460 2548 4626
rect 2400 4250 2410 4416
rect 2410 4250 2444 4416
rect 2444 4250 2452 4416
rect 2400 4236 2452 4250
rect 2688 4626 2740 4640
rect 2688 4460 2698 4626
rect 2698 4460 2732 4626
rect 2732 4460 2740 4626
rect 2592 4250 2602 4416
rect 2602 4250 2636 4416
rect 2636 4250 2644 4416
rect 2592 4236 2644 4250
rect 2880 4626 2932 4640
rect 2880 4460 2890 4626
rect 2890 4460 2924 4626
rect 2924 4460 2932 4626
rect 2784 4250 2794 4416
rect 2794 4250 2828 4416
rect 2828 4250 2836 4416
rect 2784 4236 2836 4250
rect 2976 4250 2986 4416
rect 2986 4250 3020 4416
rect 3020 4250 3028 4416
rect 2976 4236 3028 4250
rect 3912 4626 3964 4640
rect 3912 4460 3922 4626
rect 3922 4460 3956 4626
rect 3956 4460 3964 4626
rect 3816 4250 3826 4416
rect 3826 4250 3860 4416
rect 3860 4250 3868 4416
rect 3816 4236 3868 4250
rect 4104 4626 4156 4640
rect 4104 4460 4114 4626
rect 4114 4460 4148 4626
rect 4148 4460 4156 4626
rect 4008 4250 4018 4416
rect 4018 4250 4052 4416
rect 4052 4250 4060 4416
rect 4008 4236 4060 4250
rect 4296 4626 4348 4640
rect 4296 4460 4306 4626
rect 4306 4460 4340 4626
rect 4340 4460 4348 4626
rect 4200 4250 4210 4416
rect 4210 4250 4244 4416
rect 4244 4250 4252 4416
rect 4200 4236 4252 4250
rect 4488 4626 4540 4640
rect 4488 4460 4498 4626
rect 4498 4460 4532 4626
rect 4532 4460 4540 4626
rect 4392 4250 4402 4416
rect 4402 4250 4436 4416
rect 4436 4250 4444 4416
rect 4392 4236 4444 4250
rect 4680 4626 4732 4640
rect 4680 4460 4690 4626
rect 4690 4460 4724 4626
rect 4724 4460 4732 4626
rect 4584 4250 4594 4416
rect 4594 4250 4628 4416
rect 4628 4250 4636 4416
rect 4584 4236 4636 4250
rect 4776 4250 4786 4416
rect 4786 4250 4820 4416
rect 4820 4250 4828 4416
rect 4776 4236 4828 4250
rect 5712 4626 5764 4640
rect 5712 4460 5722 4626
rect 5722 4460 5756 4626
rect 5756 4460 5764 4626
rect 5616 4250 5626 4416
rect 5626 4250 5660 4416
rect 5660 4250 5668 4416
rect 5616 4236 5668 4250
rect 5904 4626 5956 4640
rect 5904 4460 5914 4626
rect 5914 4460 5948 4626
rect 5948 4460 5956 4626
rect 5808 4250 5818 4416
rect 5818 4250 5852 4416
rect 5852 4250 5860 4416
rect 5808 4236 5860 4250
rect 6096 4626 6148 4640
rect 6096 4460 6106 4626
rect 6106 4460 6140 4626
rect 6140 4460 6148 4626
rect 6000 4250 6010 4416
rect 6010 4250 6044 4416
rect 6044 4250 6052 4416
rect 6000 4236 6052 4250
rect 6288 4626 6340 4640
rect 6288 4460 6298 4626
rect 6298 4460 6332 4626
rect 6332 4460 6340 4626
rect 6192 4250 6202 4416
rect 6202 4250 6236 4416
rect 6236 4250 6244 4416
rect 6192 4236 6244 4250
rect 6480 4626 6532 4640
rect 6480 4460 6490 4626
rect 6490 4460 6524 4626
rect 6524 4460 6532 4626
rect 6384 4250 6394 4416
rect 6394 4250 6428 4416
rect 6428 4250 6436 4416
rect 6384 4236 6436 4250
rect 6576 4250 6586 4416
rect 6586 4250 6620 4416
rect 6620 4250 6628 4416
rect 6576 4236 6628 4250
rect 18396 21534 18448 21548
rect 18396 21368 18406 21534
rect 18406 21368 18440 21534
rect 18440 21368 18448 21534
rect 18304 21158 18310 21324
rect 18310 21158 18344 21324
rect 18344 21158 18356 21324
rect 18304 21144 18356 21158
rect 18588 21534 18640 21548
rect 18588 21368 18598 21534
rect 18598 21368 18632 21534
rect 18632 21368 18640 21534
rect 18492 21158 18502 21324
rect 18502 21158 18536 21324
rect 18536 21158 18544 21324
rect 18492 21144 18544 21158
rect 18780 21534 18832 21548
rect 18780 21368 18790 21534
rect 18790 21368 18824 21534
rect 18824 21368 18832 21534
rect 18684 21158 18694 21324
rect 18694 21158 18728 21324
rect 18728 21158 18736 21324
rect 18684 21144 18736 21158
rect 18972 21534 19024 21548
rect 18972 21368 18982 21534
rect 18982 21368 19016 21534
rect 19016 21368 19024 21534
rect 18876 21158 18886 21324
rect 18886 21158 18920 21324
rect 18920 21158 18928 21324
rect 18876 21144 18928 21158
rect 19164 21534 19216 21548
rect 19164 21368 19174 21534
rect 19174 21368 19208 21534
rect 19208 21368 19216 21534
rect 19068 21158 19078 21324
rect 19078 21158 19112 21324
rect 19112 21158 19120 21324
rect 19068 21144 19120 21158
rect 19260 21158 19270 21324
rect 19270 21158 19304 21324
rect 19304 21158 19312 21324
rect 19260 21144 19312 21158
rect 18560 20668 18612 20684
rect 18560 20504 18568 20668
rect 18568 20504 18602 20668
rect 18602 20504 18612 20668
rect 18300 20292 18310 20460
rect 18310 20292 18344 20460
rect 18344 20292 18352 20460
rect 18300 20280 18352 20292
rect 19076 20668 19128 20684
rect 19076 20504 19084 20668
rect 19084 20504 19118 20668
rect 19118 20504 19128 20668
rect 18816 20292 18826 20460
rect 18826 20292 18860 20460
rect 18860 20292 18868 20460
rect 18816 20280 18868 20292
rect 19592 20668 19644 20684
rect 19592 20504 19600 20668
rect 19600 20504 19634 20668
rect 19634 20504 19644 20668
rect 19332 20292 19342 20460
rect 19342 20292 19376 20460
rect 19376 20292 19384 20460
rect 19332 20280 19384 20292
rect 18560 20050 18612 20064
rect 18560 19884 18568 20050
rect 18568 19884 18602 20050
rect 18602 19884 18612 20050
rect 18300 19674 18310 19840
rect 18310 19674 18344 19840
rect 18344 19674 18352 19840
rect 18300 19660 18352 19674
rect 19076 20050 19128 20064
rect 19076 19884 19084 20050
rect 19084 19884 19118 20050
rect 19118 19884 19128 20050
rect 18816 19674 18826 19840
rect 18826 19674 18860 19840
rect 18860 19674 18868 19840
rect 18816 19660 18868 19674
rect 19592 20050 19644 20064
rect 19592 19884 19600 20050
rect 19600 19884 19634 20050
rect 19634 19884 19644 20050
rect 19332 19674 19342 19840
rect 19342 19674 19376 19840
rect 19376 19674 19384 19840
rect 19332 19660 19384 19674
rect 18560 19432 18612 19448
rect 18560 19268 18568 19432
rect 18568 19268 18602 19432
rect 18602 19268 18612 19432
rect 18300 19056 18310 19224
rect 18310 19056 18344 19224
rect 18344 19056 18352 19224
rect 18300 19044 18352 19056
rect 19076 19432 19128 19448
rect 19076 19268 19084 19432
rect 19084 19268 19118 19432
rect 19118 19268 19128 19432
rect 18816 19056 18826 19224
rect 18826 19056 18860 19224
rect 18860 19056 18868 19224
rect 18816 19044 18868 19056
rect 19592 19432 19644 19448
rect 19592 19268 19600 19432
rect 19600 19268 19634 19432
rect 19634 19268 19644 19432
rect 19332 19056 19342 19224
rect 19342 19056 19376 19224
rect 19376 19056 19384 19224
rect 19332 19044 19384 19056
rect 18560 18814 18612 18828
rect 18560 18648 18568 18814
rect 18568 18648 18602 18814
rect 18602 18648 18612 18814
rect 18300 18438 18310 18604
rect 18310 18438 18344 18604
rect 18344 18438 18352 18604
rect 18300 18424 18352 18438
rect 19076 18814 19128 18828
rect 19076 18648 19084 18814
rect 19084 18648 19118 18814
rect 19118 18648 19128 18814
rect 18816 18438 18826 18604
rect 18826 18438 18860 18604
rect 18860 18438 18868 18604
rect 18816 18424 18868 18438
rect 19592 18814 19644 18828
rect 19592 18648 19600 18814
rect 19600 18648 19634 18814
rect 19634 18648 19644 18814
rect 19332 18438 19342 18604
rect 19342 18438 19376 18604
rect 19376 18438 19384 18604
rect 19332 18424 19384 18438
rect 18480 18056 18680 18156
rect 10800 7472 11300 7928
rect 15700 10532 15968 10768
rect 16988 11100 19192 11148
rect 16988 10703 17018 11100
rect 17018 10703 17268 11100
rect 17268 10703 17396 11100
rect 17396 10703 17646 11100
rect 17646 10703 17774 11100
rect 17774 10703 18024 11100
rect 18024 10703 18152 11100
rect 18152 10703 18402 11100
rect 18402 10703 18530 11100
rect 18530 10703 18780 11100
rect 18780 10703 18908 11100
rect 18908 10703 19158 11100
rect 19158 10703 19192 11100
rect 16988 10660 19192 10703
rect 20496 10608 20676 10808
rect 19612 10271 19668 10284
rect 19612 10104 19622 10271
rect 19622 10104 19656 10271
rect 19656 10104 19668 10271
rect 16988 9869 19180 9908
rect 16988 9472 17018 9869
rect 17018 9472 17268 9869
rect 17268 9472 17396 9869
rect 17396 9472 17646 9869
rect 17646 9472 17774 9869
rect 17774 9472 18024 9869
rect 18024 9472 18152 9869
rect 18152 9472 18402 9869
rect 18402 9472 18530 9869
rect 18530 9472 18780 9869
rect 18780 9472 18908 9869
rect 18908 9472 19158 9869
rect 19158 9472 19180 9869
rect 16988 9440 19180 9472
rect 19516 9895 19526 10060
rect 19526 9895 19560 10060
rect 19560 9895 19572 10060
rect 19516 9880 19572 9895
rect 19804 10271 19860 10284
rect 19804 10104 19814 10271
rect 19814 10104 19848 10271
rect 19848 10104 19860 10271
rect 19708 9895 19718 10060
rect 19718 9895 19752 10060
rect 19752 9895 19764 10060
rect 19708 9880 19764 9895
rect 19996 10271 20052 10284
rect 19996 10104 20006 10271
rect 20006 10104 20040 10271
rect 20040 10104 20052 10271
rect 19900 9895 19910 10060
rect 19910 9895 19944 10060
rect 19944 9895 19956 10060
rect 19900 9880 19956 9895
rect 20188 10271 20244 10284
rect 20188 10104 20198 10271
rect 20198 10104 20232 10271
rect 20232 10104 20244 10271
rect 20092 9895 20102 10060
rect 20102 9895 20136 10060
rect 20136 9895 20148 10060
rect 20092 9880 20148 9895
rect 20380 10271 20436 10284
rect 20380 10104 20390 10271
rect 20390 10104 20424 10271
rect 20424 10104 20436 10271
rect 20284 9895 20294 10060
rect 20294 9895 20328 10060
rect 20328 9895 20340 10060
rect 20284 9880 20340 9895
rect 20572 10271 20628 10284
rect 20572 10104 20582 10271
rect 20582 10104 20616 10271
rect 20616 10104 20628 10271
rect 20476 9895 20486 10060
rect 20486 9895 20520 10060
rect 20520 9895 20532 10060
rect 20476 9880 20532 9895
rect 20764 10271 20820 10284
rect 20764 10104 20774 10271
rect 20774 10104 20808 10271
rect 20808 10104 20820 10271
rect 20668 9895 20678 10060
rect 20678 9895 20712 10060
rect 20712 9895 20724 10060
rect 20668 9880 20724 9895
rect 20956 10271 21012 10284
rect 20956 10104 20966 10271
rect 20966 10104 21000 10271
rect 21000 10104 21012 10271
rect 20860 9895 20870 10060
rect 20870 9895 20904 10060
rect 20904 9895 20916 10060
rect 20860 9880 20916 9895
rect 21148 10271 21204 10284
rect 21148 10104 21158 10271
rect 21158 10104 21192 10271
rect 21192 10104 21204 10271
rect 21052 9895 21062 10060
rect 21062 9895 21096 10060
rect 21096 9895 21108 10060
rect 21052 9880 21108 9895
rect 21340 10271 21396 10284
rect 21340 10104 21350 10271
rect 21350 10104 21384 10271
rect 21384 10104 21396 10271
rect 21244 9895 21254 10060
rect 21254 9895 21288 10060
rect 21288 9895 21300 10060
rect 21244 9880 21300 9895
rect 21436 9895 21446 10060
rect 21446 9895 21480 10060
rect 21480 9895 21492 10060
rect 21436 9880 21492 9895
rect 22112 10250 22168 10264
rect 22112 10080 22122 10250
rect 22122 10080 22156 10250
rect 22156 10080 22168 10250
rect 22016 9874 22026 10044
rect 22026 9874 22060 10044
rect 22060 9874 22072 10044
rect 22016 9860 22072 9874
rect 22304 10250 22360 10264
rect 22304 10080 22314 10250
rect 22314 10080 22348 10250
rect 22348 10080 22360 10250
rect 22208 9874 22218 10044
rect 22218 9874 22252 10044
rect 22252 9874 22264 10044
rect 22208 9860 22264 9874
rect 22496 10250 22552 10264
rect 22496 10080 22506 10250
rect 22506 10080 22540 10250
rect 22540 10080 22552 10250
rect 22400 9874 22410 10044
rect 22410 9874 22444 10044
rect 22444 9874 22456 10044
rect 22400 9860 22456 9874
rect 22688 10250 22744 10264
rect 22688 10080 22698 10250
rect 22698 10080 22732 10250
rect 22732 10080 22744 10250
rect 22592 9874 22602 10044
rect 22602 9874 22636 10044
rect 22636 9874 22648 10044
rect 22592 9860 22648 9874
rect 22880 10250 22936 10264
rect 22880 10080 22890 10250
rect 22890 10080 22924 10250
rect 22924 10080 22936 10250
rect 22784 9874 22794 10044
rect 22794 9874 22828 10044
rect 22828 9874 22840 10044
rect 22784 9860 22840 9874
rect 23072 10250 23128 10264
rect 23072 10080 23082 10250
rect 23082 10080 23116 10250
rect 23116 10080 23128 10250
rect 22976 9874 22986 10044
rect 22986 9874 23020 10044
rect 23020 9874 23032 10044
rect 22976 9860 23032 9874
rect 23264 10250 23320 10264
rect 23264 10080 23274 10250
rect 23274 10080 23308 10250
rect 23308 10080 23320 10250
rect 23168 9874 23178 10044
rect 23178 9874 23212 10044
rect 23212 9874 23224 10044
rect 23168 9860 23224 9874
rect 23456 10250 23512 10264
rect 23456 10080 23466 10250
rect 23466 10080 23500 10250
rect 23500 10080 23512 10250
rect 23360 9874 23370 10044
rect 23370 9874 23404 10044
rect 23404 9874 23416 10044
rect 23360 9860 23416 9874
rect 23648 10250 23704 10264
rect 23648 10080 23658 10250
rect 23658 10080 23692 10250
rect 23692 10080 23704 10250
rect 23552 9874 23562 10044
rect 23562 9874 23596 10044
rect 23596 9874 23608 10044
rect 23552 9860 23608 9874
rect 23840 10250 23896 10264
rect 23840 10080 23850 10250
rect 23850 10080 23884 10250
rect 23884 10080 23896 10250
rect 23744 9874 23754 10044
rect 23754 9874 23788 10044
rect 23788 9874 23800 10044
rect 23744 9860 23800 9874
rect 23936 9874 23946 10044
rect 23946 9874 23980 10044
rect 23980 9874 23992 10044
rect 23936 9860 23992 9874
rect 19612 9635 19668 9652
rect 19612 9472 19622 9635
rect 19622 9472 19656 9635
rect 19656 9472 19668 9635
rect 19516 9259 19526 9428
rect 19526 9259 19560 9428
rect 19560 9259 19572 9428
rect 19516 9248 19572 9259
rect 19804 9635 19860 9652
rect 19804 9472 19814 9635
rect 19814 9472 19848 9635
rect 19848 9472 19860 9635
rect 19708 9259 19718 9428
rect 19718 9259 19752 9428
rect 19752 9259 19764 9428
rect 19708 9248 19764 9259
rect 19996 9635 20052 9652
rect 19996 9472 20006 9635
rect 20006 9472 20040 9635
rect 20040 9472 20052 9635
rect 19900 9259 19910 9428
rect 19910 9259 19944 9428
rect 19944 9259 19956 9428
rect 19900 9248 19956 9259
rect 20188 9635 20244 9652
rect 20188 9472 20198 9635
rect 20198 9472 20232 9635
rect 20232 9472 20244 9635
rect 20092 9259 20102 9428
rect 20102 9259 20136 9428
rect 20136 9259 20148 9428
rect 20092 9248 20148 9259
rect 20380 9635 20436 9652
rect 20380 9472 20390 9635
rect 20390 9472 20424 9635
rect 20424 9472 20436 9635
rect 20284 9259 20294 9428
rect 20294 9259 20328 9428
rect 20328 9259 20340 9428
rect 20284 9248 20340 9259
rect 20572 9635 20628 9652
rect 20572 9472 20582 9635
rect 20582 9472 20616 9635
rect 20616 9472 20628 9635
rect 20476 9259 20486 9428
rect 20486 9259 20520 9428
rect 20520 9259 20532 9428
rect 20476 9248 20532 9259
rect 20764 9635 20820 9652
rect 20764 9472 20774 9635
rect 20774 9472 20808 9635
rect 20808 9472 20820 9635
rect 20668 9259 20678 9428
rect 20678 9259 20712 9428
rect 20712 9259 20724 9428
rect 20668 9248 20724 9259
rect 20956 9635 21012 9652
rect 20956 9472 20966 9635
rect 20966 9472 21000 9635
rect 21000 9472 21012 9635
rect 20860 9259 20870 9428
rect 20870 9259 20904 9428
rect 20904 9259 20916 9428
rect 20860 9248 20916 9259
rect 21148 9635 21204 9652
rect 21148 9472 21158 9635
rect 21158 9472 21192 9635
rect 21192 9472 21204 9635
rect 21052 9259 21062 9428
rect 21062 9259 21096 9428
rect 21096 9259 21108 9428
rect 21052 9248 21108 9259
rect 21340 9635 21396 9652
rect 21340 9472 21350 9635
rect 21350 9472 21384 9635
rect 21384 9472 21396 9635
rect 21244 9259 21254 9428
rect 21254 9259 21288 9428
rect 21288 9259 21300 9428
rect 21244 9248 21300 9259
rect 21436 9259 21446 9428
rect 21446 9259 21480 9428
rect 21480 9259 21492 9428
rect 21436 9248 21492 9259
rect 22112 9632 22168 9648
rect 22112 9464 22122 9632
rect 22122 9464 22156 9632
rect 22156 9464 22168 9632
rect 22016 9256 22026 9428
rect 22026 9256 22060 9428
rect 22060 9256 22072 9428
rect 22016 9244 22072 9256
rect 22304 9632 22360 9648
rect 22304 9464 22314 9632
rect 22314 9464 22348 9632
rect 22348 9464 22360 9632
rect 22208 9256 22218 9428
rect 22218 9256 22252 9428
rect 22252 9256 22264 9428
rect 22208 9244 22264 9256
rect 22496 9632 22552 9648
rect 22496 9464 22506 9632
rect 22506 9464 22540 9632
rect 22540 9464 22552 9632
rect 22400 9256 22410 9428
rect 22410 9256 22444 9428
rect 22444 9256 22456 9428
rect 22400 9244 22456 9256
rect 22688 9632 22744 9648
rect 22688 9464 22698 9632
rect 22698 9464 22732 9632
rect 22732 9464 22744 9632
rect 22592 9256 22602 9428
rect 22602 9256 22636 9428
rect 22636 9256 22648 9428
rect 22592 9244 22648 9256
rect 22880 9632 22936 9648
rect 22880 9464 22890 9632
rect 22890 9464 22924 9632
rect 22924 9464 22936 9632
rect 22784 9256 22794 9428
rect 22794 9256 22828 9428
rect 22828 9256 22840 9428
rect 22784 9244 22840 9256
rect 23072 9632 23128 9648
rect 23072 9464 23082 9632
rect 23082 9464 23116 9632
rect 23116 9464 23128 9632
rect 22976 9256 22986 9428
rect 22986 9256 23020 9428
rect 23020 9256 23032 9428
rect 22976 9244 23032 9256
rect 23264 9632 23320 9648
rect 23264 9464 23274 9632
rect 23274 9464 23308 9632
rect 23308 9464 23320 9632
rect 23168 9256 23178 9428
rect 23178 9256 23212 9428
rect 23212 9256 23224 9428
rect 23168 9244 23224 9256
rect 23456 9632 23512 9648
rect 23456 9464 23466 9632
rect 23466 9464 23500 9632
rect 23500 9464 23512 9632
rect 23360 9256 23370 9428
rect 23370 9256 23404 9428
rect 23404 9256 23416 9428
rect 23360 9244 23416 9256
rect 23648 9632 23704 9648
rect 23648 9464 23658 9632
rect 23658 9464 23692 9632
rect 23692 9464 23704 9632
rect 23552 9256 23562 9428
rect 23562 9256 23596 9428
rect 23596 9256 23608 9428
rect 23552 9244 23608 9256
rect 23840 9632 23896 9648
rect 23840 9464 23850 9632
rect 23850 9464 23884 9632
rect 23884 9464 23896 9632
rect 23744 9256 23754 9428
rect 23754 9256 23788 9428
rect 23788 9256 23800 9428
rect 23744 9244 23800 9256
rect 23936 9256 23946 9428
rect 23946 9256 23980 9428
rect 23980 9256 23992 9428
rect 23936 9244 23992 9256
rect 16164 8904 16364 8964
rect 16364 8904 16456 8964
rect 16940 8904 17232 8964
rect 17876 8904 18168 8964
rect 16176 8718 16228 8732
rect 16176 8552 16186 8718
rect 16186 8552 16220 8718
rect 16220 8552 16228 8718
rect 16080 8342 16090 8508
rect 16090 8342 16124 8508
rect 16124 8342 16132 8508
rect 16080 8328 16132 8342
rect 16368 8718 16420 8732
rect 16368 8552 16378 8718
rect 16378 8552 16412 8718
rect 16412 8552 16420 8718
rect 16272 8342 16282 8508
rect 16282 8342 16316 8508
rect 16316 8342 16324 8508
rect 16272 8328 16324 8342
rect 16560 8718 16612 8732
rect 16560 8552 16570 8718
rect 16570 8552 16604 8718
rect 16604 8552 16612 8718
rect 16464 8342 16474 8508
rect 16474 8342 16508 8508
rect 16508 8342 16516 8508
rect 16464 8328 16516 8342
rect 16752 8718 16804 8732
rect 16752 8552 16762 8718
rect 16762 8552 16796 8718
rect 16796 8552 16804 8718
rect 16656 8342 16666 8508
rect 16666 8342 16700 8508
rect 16700 8342 16708 8508
rect 16656 8328 16708 8342
rect 16944 8718 16996 8732
rect 16944 8552 16954 8718
rect 16954 8552 16988 8718
rect 16988 8552 16996 8718
rect 16848 8342 16858 8508
rect 16858 8342 16892 8508
rect 16892 8342 16900 8508
rect 16848 8328 16900 8342
rect 17136 8718 17188 8732
rect 17136 8552 17146 8718
rect 17146 8552 17180 8718
rect 17180 8552 17188 8718
rect 17040 8342 17050 8508
rect 17050 8342 17084 8508
rect 17084 8342 17092 8508
rect 17040 8328 17092 8342
rect 17328 8718 17380 8732
rect 17328 8552 17338 8718
rect 17338 8552 17372 8718
rect 17372 8552 17380 8718
rect 17232 8342 17242 8508
rect 17242 8342 17276 8508
rect 17276 8342 17284 8508
rect 17232 8328 17284 8342
rect 17520 8718 17572 8732
rect 17520 8552 17530 8718
rect 17530 8552 17564 8718
rect 17564 8552 17572 8718
rect 17424 8342 17434 8508
rect 17434 8342 17468 8508
rect 17468 8342 17476 8508
rect 17424 8328 17476 8342
rect 17712 8718 17764 8732
rect 17712 8552 17722 8718
rect 17722 8552 17756 8718
rect 17756 8552 17764 8718
rect 17616 8342 17626 8508
rect 17626 8342 17660 8508
rect 17660 8342 17668 8508
rect 17616 8328 17668 8342
rect 17904 8718 17956 8732
rect 17904 8552 17914 8718
rect 17914 8552 17948 8718
rect 17948 8552 17956 8718
rect 17808 8342 17818 8508
rect 17818 8342 17852 8508
rect 17852 8342 17860 8508
rect 17808 8328 17860 8342
rect 18000 8342 18010 8508
rect 18010 8342 18044 8508
rect 18044 8342 18052 8508
rect 18000 8328 18052 8342
rect 18140 8416 18200 8672
rect 18988 8432 19408 8984
rect 19612 8684 19668 8700
rect 19612 8520 19622 8684
rect 19622 8520 19656 8684
rect 19656 8520 19668 8684
rect 19516 8308 19526 8476
rect 19526 8308 19560 8476
rect 19560 8308 19572 8476
rect 19516 8296 19572 8308
rect 19804 8684 19860 8700
rect 19804 8520 19814 8684
rect 19814 8520 19848 8684
rect 19848 8520 19860 8684
rect 19708 8308 19718 8476
rect 19718 8308 19752 8476
rect 19752 8308 19764 8476
rect 19708 8296 19764 8308
rect 19996 8684 20052 8700
rect 19996 8520 20006 8684
rect 20006 8520 20040 8684
rect 20040 8520 20052 8684
rect 19900 8308 19910 8476
rect 19910 8308 19944 8476
rect 19944 8308 19956 8476
rect 19900 8296 19956 8308
rect 20188 8684 20244 8700
rect 20188 8520 20198 8684
rect 20198 8520 20232 8684
rect 20232 8520 20244 8684
rect 20092 8308 20102 8476
rect 20102 8308 20136 8476
rect 20136 8308 20148 8476
rect 20092 8296 20148 8308
rect 20380 8684 20436 8700
rect 20380 8520 20390 8684
rect 20390 8520 20424 8684
rect 20424 8520 20436 8684
rect 20284 8308 20294 8476
rect 20294 8308 20328 8476
rect 20328 8308 20340 8476
rect 20284 8296 20340 8308
rect 20572 8684 20628 8700
rect 20572 8520 20582 8684
rect 20582 8520 20616 8684
rect 20616 8520 20628 8684
rect 20476 8308 20486 8476
rect 20486 8308 20520 8476
rect 20520 8308 20532 8476
rect 20476 8296 20532 8308
rect 20764 8684 20820 8700
rect 20764 8520 20774 8684
rect 20774 8520 20808 8684
rect 20808 8520 20820 8684
rect 20668 8308 20678 8476
rect 20678 8308 20712 8476
rect 20712 8308 20724 8476
rect 20668 8296 20724 8308
rect 20956 8684 21012 8700
rect 20956 8520 20966 8684
rect 20966 8520 21000 8684
rect 21000 8520 21012 8684
rect 20860 8308 20870 8476
rect 20870 8308 20904 8476
rect 20904 8308 20916 8476
rect 20860 8296 20916 8308
rect 21148 8684 21204 8700
rect 21148 8520 21158 8684
rect 21158 8520 21192 8684
rect 21192 8520 21204 8684
rect 21052 8308 21062 8476
rect 21062 8308 21096 8476
rect 21096 8308 21108 8476
rect 21052 8296 21108 8308
rect 21340 8684 21396 8700
rect 21340 8520 21350 8684
rect 21350 8520 21384 8684
rect 21384 8520 21396 8684
rect 21244 8308 21254 8476
rect 21254 8308 21288 8476
rect 21288 8308 21300 8476
rect 21244 8296 21300 8308
rect 21436 8308 21446 8476
rect 21446 8308 21480 8476
rect 21480 8308 21492 8476
rect 21436 8296 21492 8308
rect 16164 8148 16456 8152
rect 16164 8088 16364 8148
rect 16364 8088 16456 8148
rect 16940 8148 17260 8152
rect 16940 8088 17260 8148
rect 17876 8092 18168 8152
rect 16176 7898 16228 7912
rect 16176 7732 16186 7898
rect 16186 7732 16220 7898
rect 16220 7732 16228 7898
rect 16080 7522 16090 7688
rect 16090 7522 16124 7688
rect 16124 7522 16132 7688
rect 16080 7508 16132 7522
rect 16368 7898 16420 7912
rect 16368 7732 16378 7898
rect 16378 7732 16412 7898
rect 16412 7732 16420 7898
rect 16272 7522 16282 7688
rect 16282 7522 16316 7688
rect 16316 7522 16324 7688
rect 16272 7508 16324 7522
rect 16560 7898 16612 7912
rect 16560 7732 16570 7898
rect 16570 7732 16604 7898
rect 16604 7732 16612 7898
rect 16464 7522 16474 7688
rect 16474 7522 16508 7688
rect 16508 7522 16516 7688
rect 16464 7508 16516 7522
rect 16752 7898 16804 7912
rect 16752 7732 16762 7898
rect 16762 7732 16796 7898
rect 16796 7732 16804 7898
rect 16656 7522 16666 7688
rect 16666 7522 16700 7688
rect 16700 7522 16708 7688
rect 16656 7508 16708 7522
rect 16944 7898 16996 7912
rect 16944 7732 16954 7898
rect 16954 7732 16988 7898
rect 16988 7732 16996 7898
rect 16848 7522 16858 7688
rect 16858 7522 16892 7688
rect 16892 7522 16900 7688
rect 16848 7508 16900 7522
rect 17136 7898 17188 7912
rect 17136 7732 17146 7898
rect 17146 7732 17180 7898
rect 17180 7732 17188 7898
rect 17040 7522 17050 7688
rect 17050 7522 17084 7688
rect 17084 7522 17092 7688
rect 17040 7508 17092 7522
rect 17328 7898 17380 7912
rect 17328 7732 17338 7898
rect 17338 7732 17372 7898
rect 17372 7732 17380 7898
rect 17232 7522 17242 7688
rect 17242 7522 17276 7688
rect 17276 7522 17284 7688
rect 17232 7508 17284 7522
rect 17520 7898 17572 7912
rect 17520 7732 17530 7898
rect 17530 7732 17564 7898
rect 17564 7732 17572 7898
rect 17424 7522 17434 7688
rect 17434 7522 17468 7688
rect 17468 7522 17476 7688
rect 17424 7508 17476 7522
rect 17712 7898 17764 7912
rect 17712 7732 17722 7898
rect 17722 7732 17756 7898
rect 17756 7732 17764 7898
rect 17616 7522 17626 7688
rect 17626 7522 17660 7688
rect 17660 7522 17668 7688
rect 17616 7508 17668 7522
rect 17904 7898 17956 7912
rect 17904 7732 17914 7898
rect 17914 7732 17948 7898
rect 17948 7732 17956 7898
rect 17808 7522 17818 7688
rect 17818 7522 17852 7688
rect 17852 7522 17860 7688
rect 17808 7508 17860 7522
rect 18000 7522 18010 7688
rect 18010 7522 18044 7688
rect 18044 7522 18052 7688
rect 18000 7508 18052 7522
rect 18140 7568 18200 7824
rect 19612 8066 19668 8080
rect 19612 7900 19622 8066
rect 19622 7900 19656 8066
rect 19656 7900 19668 8066
rect 19516 7690 19526 7856
rect 19526 7690 19560 7856
rect 19560 7690 19572 7856
rect 19516 7676 19572 7690
rect 19804 8066 19860 8080
rect 19804 7900 19814 8066
rect 19814 7900 19848 8066
rect 19848 7900 19860 8066
rect 19708 7690 19718 7856
rect 19718 7690 19752 7856
rect 19752 7690 19764 7856
rect 19708 7676 19764 7690
rect 19996 8066 20052 8080
rect 19996 7900 20006 8066
rect 20006 7900 20040 8066
rect 20040 7900 20052 8066
rect 19900 7690 19910 7856
rect 19910 7690 19944 7856
rect 19944 7690 19956 7856
rect 19900 7676 19956 7690
rect 20188 8066 20244 8080
rect 20188 7900 20198 8066
rect 20198 7900 20232 8066
rect 20232 7900 20244 8066
rect 20092 7690 20102 7856
rect 20102 7690 20136 7856
rect 20136 7690 20148 7856
rect 20092 7676 20148 7690
rect 20380 8066 20436 8080
rect 20380 7900 20390 8066
rect 20390 7900 20424 8066
rect 20424 7900 20436 8066
rect 20284 7690 20294 7856
rect 20294 7690 20328 7856
rect 20328 7690 20340 7856
rect 20284 7676 20340 7690
rect 20572 8066 20628 8080
rect 20572 7900 20582 8066
rect 20582 7900 20616 8066
rect 20616 7900 20628 8066
rect 20476 7690 20486 7856
rect 20486 7690 20520 7856
rect 20520 7690 20532 7856
rect 20476 7676 20532 7690
rect 20764 8066 20820 8080
rect 20764 7900 20774 8066
rect 20774 7900 20808 8066
rect 20808 7900 20820 8066
rect 20668 7690 20678 7856
rect 20678 7690 20712 7856
rect 20712 7690 20724 7856
rect 20668 7676 20724 7690
rect 20956 8066 21012 8080
rect 20956 7900 20966 8066
rect 20966 7900 21000 8066
rect 21000 7900 21012 8066
rect 20860 7690 20870 7856
rect 20870 7690 20904 7856
rect 20904 7690 20916 7856
rect 20860 7676 20916 7690
rect 21148 8066 21204 8080
rect 21148 7900 21158 8066
rect 21158 7900 21192 8066
rect 21192 7900 21204 8066
rect 21052 7690 21062 7856
rect 21062 7690 21096 7856
rect 21096 7690 21108 7856
rect 21052 7676 21108 7690
rect 21340 8066 21396 8080
rect 21340 7900 21350 8066
rect 21350 7900 21384 8066
rect 21384 7900 21396 8066
rect 21244 7690 21254 7856
rect 21254 7690 21288 7856
rect 21288 7690 21300 7856
rect 21244 7676 21300 7690
rect 21436 7690 21446 7856
rect 21446 7690 21480 7856
rect 21480 7690 21492 7856
rect 21436 7676 21492 7690
rect 16164 7268 16364 7328
rect 16364 7268 16456 7328
rect 16936 7268 16940 7328
rect 16940 7268 17228 7328
rect 17876 7268 18168 7328
rect 16176 7078 16228 7092
rect 16176 6912 16186 7078
rect 16186 6912 16220 7078
rect 16220 6912 16228 7078
rect 16080 6702 16090 6868
rect 16090 6702 16124 6868
rect 16124 6702 16132 6868
rect 16080 6688 16132 6702
rect 16368 7078 16420 7092
rect 16368 6912 16378 7078
rect 16378 6912 16412 7078
rect 16412 6912 16420 7078
rect 16272 6702 16282 6868
rect 16282 6702 16316 6868
rect 16316 6702 16324 6868
rect 16272 6688 16324 6702
rect 16560 7078 16612 7092
rect 16560 6912 16570 7078
rect 16570 6912 16604 7078
rect 16604 6912 16612 7078
rect 16464 6702 16474 6868
rect 16474 6702 16508 6868
rect 16508 6702 16516 6868
rect 16464 6688 16516 6702
rect 16752 7078 16804 7092
rect 16752 6912 16762 7078
rect 16762 6912 16796 7078
rect 16796 6912 16804 7078
rect 16656 6702 16666 6868
rect 16666 6702 16700 6868
rect 16700 6702 16708 6868
rect 16656 6688 16708 6702
rect 16944 7078 16996 7092
rect 16944 6912 16954 7078
rect 16954 6912 16988 7078
rect 16988 6912 16996 7078
rect 16848 6702 16858 6868
rect 16858 6702 16892 6868
rect 16892 6702 16900 6868
rect 16848 6688 16900 6702
rect 17136 7078 17188 7092
rect 17136 6912 17146 7078
rect 17146 6912 17180 7078
rect 17180 6912 17188 7078
rect 17040 6702 17050 6868
rect 17050 6702 17084 6868
rect 17084 6702 17092 6868
rect 17040 6688 17092 6702
rect 17328 7078 17380 7092
rect 17328 6912 17338 7078
rect 17338 6912 17372 7078
rect 17372 6912 17380 7078
rect 17232 6702 17242 6868
rect 17242 6702 17276 6868
rect 17276 6702 17284 6868
rect 17232 6688 17284 6702
rect 17520 7078 17572 7092
rect 17520 6912 17530 7078
rect 17530 6912 17564 7078
rect 17564 6912 17572 7078
rect 17424 6702 17434 6868
rect 17434 6702 17468 6868
rect 17468 6702 17476 6868
rect 17424 6688 17476 6702
rect 17712 7078 17764 7092
rect 17712 6912 17722 7078
rect 17722 6912 17756 7078
rect 17756 6912 17764 7078
rect 17616 6702 17626 6868
rect 17626 6702 17660 6868
rect 17660 6702 17668 6868
rect 17616 6688 17668 6702
rect 17904 7078 17956 7092
rect 17904 6912 17914 7078
rect 17914 6912 17948 7078
rect 17948 6912 17956 7078
rect 17808 6702 17818 6868
rect 17818 6702 17852 6868
rect 17852 6702 17860 6868
rect 17808 6688 17860 6702
rect 18000 6702 18010 6868
rect 18010 6702 18044 6868
rect 18044 6702 18052 6868
rect 18000 6688 18052 6702
rect 18140 6756 18200 7012
rect 20784 7000 21476 7512
rect 22112 9014 22168 9028
rect 22112 8844 22122 9014
rect 22122 8844 22156 9014
rect 22156 8844 22168 9014
rect 22016 8638 22026 8808
rect 22026 8638 22060 8808
rect 22060 8638 22072 8808
rect 22016 8624 22072 8638
rect 22304 9014 22360 9028
rect 22304 8844 22314 9014
rect 22314 8844 22348 9014
rect 22348 8844 22360 9014
rect 22208 8638 22218 8808
rect 22218 8638 22252 8808
rect 22252 8638 22264 8808
rect 22208 8624 22264 8638
rect 22496 9014 22552 9028
rect 22496 8844 22506 9014
rect 22506 8844 22540 9014
rect 22540 8844 22552 9014
rect 22400 8638 22410 8808
rect 22410 8638 22444 8808
rect 22444 8638 22456 8808
rect 22400 8624 22456 8638
rect 22688 9014 22744 9028
rect 22688 8844 22698 9014
rect 22698 8844 22732 9014
rect 22732 8844 22744 9014
rect 22592 8638 22602 8808
rect 22602 8638 22636 8808
rect 22636 8638 22648 8808
rect 22592 8624 22648 8638
rect 22880 9014 22936 9028
rect 22880 8844 22890 9014
rect 22890 8844 22924 9014
rect 22924 8844 22936 9014
rect 22784 8638 22794 8808
rect 22794 8638 22828 8808
rect 22828 8638 22840 8808
rect 22784 8624 22840 8638
rect 23072 9014 23128 9028
rect 23072 8844 23082 9014
rect 23082 8844 23116 9014
rect 23116 8844 23128 9014
rect 22976 8638 22986 8808
rect 22986 8638 23020 8808
rect 23020 8638 23032 8808
rect 22976 8624 23032 8638
rect 23264 9014 23320 9028
rect 23264 8844 23274 9014
rect 23274 8844 23308 9014
rect 23308 8844 23320 9014
rect 23168 8638 23178 8808
rect 23178 8638 23212 8808
rect 23212 8638 23224 8808
rect 23168 8624 23224 8638
rect 23456 9014 23512 9028
rect 23456 8844 23466 9014
rect 23466 8844 23500 9014
rect 23500 8844 23512 9014
rect 23360 8638 23370 8808
rect 23370 8638 23404 8808
rect 23404 8638 23416 8808
rect 23360 8624 23416 8638
rect 23648 9014 23704 9028
rect 23648 8844 23658 9014
rect 23658 8844 23692 9014
rect 23692 8844 23704 9014
rect 23552 8638 23562 8808
rect 23562 8638 23596 8808
rect 23596 8638 23608 8808
rect 23552 8624 23608 8638
rect 23840 9014 23896 9028
rect 23840 8844 23850 9014
rect 23850 8844 23884 9014
rect 23884 8844 23896 9014
rect 23744 8638 23754 8808
rect 23754 8638 23788 8808
rect 23788 8638 23800 8808
rect 23744 8624 23800 8638
rect 23936 8638 23946 8808
rect 23946 8638 23980 8808
rect 23980 8638 23992 8808
rect 23936 8624 23992 8638
rect 22112 8396 22168 8412
rect 22112 8228 22122 8396
rect 22122 8228 22156 8396
rect 22156 8228 22168 8396
rect 22016 8020 22026 8192
rect 22026 8020 22060 8192
rect 22060 8020 22072 8192
rect 22016 8008 22072 8020
rect 22304 8396 22360 8412
rect 22304 8228 22314 8396
rect 22314 8228 22348 8396
rect 22348 8228 22360 8396
rect 22208 8020 22218 8192
rect 22218 8020 22252 8192
rect 22252 8020 22264 8192
rect 22208 8008 22264 8020
rect 22496 8396 22552 8412
rect 22496 8228 22506 8396
rect 22506 8228 22540 8396
rect 22540 8228 22552 8396
rect 22400 8020 22410 8192
rect 22410 8020 22444 8192
rect 22444 8020 22456 8192
rect 22400 8008 22456 8020
rect 22688 8396 22744 8412
rect 22688 8228 22698 8396
rect 22698 8228 22732 8396
rect 22732 8228 22744 8396
rect 22592 8020 22602 8192
rect 22602 8020 22636 8192
rect 22636 8020 22648 8192
rect 22592 8008 22648 8020
rect 22880 8396 22936 8412
rect 22880 8228 22890 8396
rect 22890 8228 22924 8396
rect 22924 8228 22936 8396
rect 22784 8020 22794 8192
rect 22794 8020 22828 8192
rect 22828 8020 22840 8192
rect 22784 8008 22840 8020
rect 23072 8396 23128 8412
rect 23072 8228 23082 8396
rect 23082 8228 23116 8396
rect 23116 8228 23128 8396
rect 22976 8020 22986 8192
rect 22986 8020 23020 8192
rect 23020 8020 23032 8192
rect 22976 8008 23032 8020
rect 23264 8396 23320 8412
rect 23264 8228 23274 8396
rect 23274 8228 23308 8396
rect 23308 8228 23320 8396
rect 23168 8020 23178 8192
rect 23178 8020 23212 8192
rect 23212 8020 23224 8192
rect 23168 8008 23224 8020
rect 23456 8396 23512 8412
rect 23456 8228 23466 8396
rect 23466 8228 23500 8396
rect 23500 8228 23512 8396
rect 23360 8020 23370 8192
rect 23370 8020 23404 8192
rect 23404 8020 23416 8192
rect 23360 8008 23416 8020
rect 23648 8396 23704 8412
rect 23648 8228 23658 8396
rect 23658 8228 23692 8396
rect 23692 8228 23704 8396
rect 23552 8020 23562 8192
rect 23562 8020 23596 8192
rect 23596 8020 23608 8192
rect 23552 8008 23608 8020
rect 23840 8396 23896 8412
rect 23840 8228 23850 8396
rect 23850 8228 23884 8396
rect 23884 8228 23896 8396
rect 23744 8020 23754 8192
rect 23754 8020 23788 8192
rect 23788 8020 23800 8192
rect 23744 8008 23800 8020
rect 23936 8020 23946 8192
rect 23946 8020 23980 8192
rect 23980 8020 23992 8192
rect 23936 8008 23992 8020
rect 22112 7778 22168 7792
rect 22112 7608 22122 7778
rect 22122 7608 22156 7778
rect 22156 7608 22168 7778
rect 22016 7402 22026 7572
rect 22026 7402 22060 7572
rect 22060 7402 22072 7572
rect 22016 7388 22072 7402
rect 22304 7778 22360 7792
rect 22304 7608 22314 7778
rect 22314 7608 22348 7778
rect 22348 7608 22360 7778
rect 22208 7402 22218 7572
rect 22218 7402 22252 7572
rect 22252 7402 22264 7572
rect 22208 7388 22264 7402
rect 22496 7778 22552 7792
rect 22496 7608 22506 7778
rect 22506 7608 22540 7778
rect 22540 7608 22552 7778
rect 22400 7402 22410 7572
rect 22410 7402 22444 7572
rect 22444 7402 22456 7572
rect 22400 7388 22456 7402
rect 22688 7778 22744 7792
rect 22688 7608 22698 7778
rect 22698 7608 22732 7778
rect 22732 7608 22744 7778
rect 22592 7402 22602 7572
rect 22602 7402 22636 7572
rect 22636 7402 22648 7572
rect 22592 7388 22648 7402
rect 22880 7778 22936 7792
rect 22880 7608 22890 7778
rect 22890 7608 22924 7778
rect 22924 7608 22936 7778
rect 22784 7402 22794 7572
rect 22794 7402 22828 7572
rect 22828 7402 22840 7572
rect 22784 7388 22840 7402
rect 23072 7778 23128 7792
rect 23072 7608 23082 7778
rect 23082 7608 23116 7778
rect 23116 7608 23128 7778
rect 22976 7402 22986 7572
rect 22986 7402 23020 7572
rect 23020 7402 23032 7572
rect 22976 7388 23032 7402
rect 23264 7778 23320 7792
rect 23264 7608 23274 7778
rect 23274 7608 23308 7778
rect 23308 7608 23320 7778
rect 23168 7402 23178 7572
rect 23178 7402 23212 7572
rect 23212 7402 23224 7572
rect 23168 7388 23224 7402
rect 23456 7778 23512 7792
rect 23456 7608 23466 7778
rect 23466 7608 23500 7778
rect 23500 7608 23512 7778
rect 23360 7402 23370 7572
rect 23370 7402 23404 7572
rect 23404 7402 23416 7572
rect 23360 7388 23416 7402
rect 23648 7778 23704 7792
rect 23648 7608 23658 7778
rect 23658 7608 23692 7778
rect 23692 7608 23704 7778
rect 23552 7402 23562 7572
rect 23562 7402 23596 7572
rect 23596 7402 23608 7572
rect 23552 7388 23608 7402
rect 23840 7778 23896 7792
rect 23840 7608 23850 7778
rect 23850 7608 23884 7778
rect 23884 7608 23896 7778
rect 23744 7402 23754 7572
rect 23754 7402 23788 7572
rect 23788 7402 23800 7572
rect 23744 7388 23800 7402
rect 23936 7402 23946 7572
rect 23946 7402 23980 7572
rect 23980 7402 23992 7572
rect 23936 7388 23992 7402
rect 22112 7160 22168 7176
rect 22112 6992 22122 7160
rect 22122 6992 22156 7160
rect 22156 6992 22168 7160
rect 21400 6600 21928 6928
rect 22016 6784 22026 6956
rect 22026 6784 22060 6956
rect 22060 6784 22072 6956
rect 22016 6772 22072 6784
rect 22304 7160 22360 7176
rect 22304 6992 22314 7160
rect 22314 6992 22348 7160
rect 22348 6992 22360 7160
rect 22208 6784 22218 6956
rect 22218 6784 22252 6956
rect 22252 6784 22264 6956
rect 22208 6772 22264 6784
rect 22496 7160 22552 7176
rect 22496 6992 22506 7160
rect 22506 6992 22540 7160
rect 22540 6992 22552 7160
rect 22400 6784 22410 6956
rect 22410 6784 22444 6956
rect 22444 6784 22456 6956
rect 22400 6772 22456 6784
rect 22688 7160 22744 7176
rect 22688 6992 22698 7160
rect 22698 6992 22732 7160
rect 22732 6992 22744 7160
rect 22592 6784 22602 6956
rect 22602 6784 22636 6956
rect 22636 6784 22648 6956
rect 22592 6772 22648 6784
rect 22880 7160 22936 7176
rect 22880 6992 22890 7160
rect 22890 6992 22924 7160
rect 22924 6992 22936 7160
rect 22784 6784 22794 6956
rect 22794 6784 22828 6956
rect 22828 6784 22840 6956
rect 22784 6772 22840 6784
rect 23072 7160 23128 7176
rect 23072 6992 23082 7160
rect 23082 6992 23116 7160
rect 23116 6992 23128 7160
rect 22976 6784 22986 6956
rect 22986 6784 23020 6956
rect 23020 6784 23032 6956
rect 22976 6772 23032 6784
rect 23264 7160 23320 7176
rect 23264 6992 23274 7160
rect 23274 6992 23308 7160
rect 23308 6992 23320 7160
rect 23168 6784 23178 6956
rect 23178 6784 23212 6956
rect 23212 6784 23224 6956
rect 23168 6772 23224 6784
rect 23456 7160 23512 7176
rect 23456 6992 23466 7160
rect 23466 6992 23500 7160
rect 23500 6992 23512 7160
rect 23360 6784 23370 6956
rect 23370 6784 23404 6956
rect 23404 6784 23416 6956
rect 23360 6772 23416 6784
rect 23648 7160 23704 7176
rect 23648 6992 23658 7160
rect 23658 6992 23692 7160
rect 23692 6992 23704 7160
rect 23552 6784 23562 6956
rect 23562 6784 23596 6956
rect 23596 6784 23608 6956
rect 23552 6772 23608 6784
rect 23840 7160 23896 7176
rect 23840 6992 23850 7160
rect 23850 6992 23884 7160
rect 23884 6992 23896 7160
rect 23744 6784 23754 6956
rect 23754 6784 23788 6956
rect 23788 6784 23800 6956
rect 23744 6772 23800 6784
rect 23936 6784 23946 6956
rect 23946 6784 23980 6956
rect 23980 6784 23992 6956
rect 23936 6772 23992 6784
rect 16072 6456 16364 6516
rect 16940 6456 17232 6516
rect 17876 6452 18168 6512
rect 21360 6156 21856 6472
rect 22112 6542 22168 6556
rect 22112 6372 22122 6542
rect 22122 6372 22156 6542
rect 22156 6372 22168 6542
rect 22016 6166 22026 6336
rect 22026 6166 22060 6336
rect 22060 6166 22072 6336
rect 22016 6152 22072 6166
rect 22304 6542 22360 6556
rect 22304 6372 22314 6542
rect 22314 6372 22348 6542
rect 22348 6372 22360 6542
rect 22208 6166 22218 6336
rect 22218 6166 22252 6336
rect 22252 6166 22264 6336
rect 22208 6152 22264 6166
rect 22496 6542 22552 6556
rect 22496 6372 22506 6542
rect 22506 6372 22540 6542
rect 22540 6372 22552 6542
rect 22400 6166 22410 6336
rect 22410 6166 22444 6336
rect 22444 6166 22456 6336
rect 22400 6152 22456 6166
rect 22688 6542 22744 6556
rect 22688 6372 22698 6542
rect 22698 6372 22732 6542
rect 22732 6372 22744 6542
rect 22592 6166 22602 6336
rect 22602 6166 22636 6336
rect 22636 6166 22648 6336
rect 22592 6152 22648 6166
rect 22880 6542 22936 6556
rect 22880 6372 22890 6542
rect 22890 6372 22924 6542
rect 22924 6372 22936 6542
rect 22784 6166 22794 6336
rect 22794 6166 22828 6336
rect 22828 6166 22840 6336
rect 22784 6152 22840 6166
rect 23072 6542 23128 6556
rect 23072 6372 23082 6542
rect 23082 6372 23116 6542
rect 23116 6372 23128 6542
rect 22976 6166 22986 6336
rect 22986 6166 23020 6336
rect 23020 6166 23032 6336
rect 22976 6152 23032 6166
rect 23264 6542 23320 6556
rect 23264 6372 23274 6542
rect 23274 6372 23308 6542
rect 23308 6372 23320 6542
rect 23168 6166 23178 6336
rect 23178 6166 23212 6336
rect 23212 6166 23224 6336
rect 23168 6152 23224 6166
rect 23456 6542 23512 6556
rect 23456 6372 23466 6542
rect 23466 6372 23500 6542
rect 23500 6372 23512 6542
rect 23360 6166 23370 6336
rect 23370 6166 23404 6336
rect 23404 6166 23416 6336
rect 23360 6152 23416 6166
rect 23648 6542 23704 6556
rect 23648 6372 23658 6542
rect 23658 6372 23692 6542
rect 23692 6372 23704 6542
rect 23552 6166 23562 6336
rect 23562 6166 23596 6336
rect 23596 6166 23608 6336
rect 23552 6152 23608 6166
rect 23840 6542 23896 6556
rect 23840 6372 23850 6542
rect 23850 6372 23884 6542
rect 23884 6372 23896 6542
rect 23744 6166 23754 6336
rect 23754 6166 23788 6336
rect 23788 6166 23800 6336
rect 23744 6152 23800 6166
rect 23936 6166 23946 6336
rect 23946 6166 23980 6336
rect 23980 6166 23992 6336
rect 23936 6152 23992 6166
rect 14712 5862 14764 5876
rect 14712 5696 14722 5862
rect 14722 5696 14756 5862
rect 14756 5696 14764 5862
rect 14616 5486 14626 5652
rect 14626 5486 14660 5652
rect 14660 5486 14668 5652
rect 14616 5472 14668 5486
rect 14904 5862 14956 5876
rect 14904 5696 14914 5862
rect 14914 5696 14948 5862
rect 14948 5696 14956 5862
rect 14808 5486 14818 5652
rect 14818 5486 14852 5652
rect 14852 5486 14860 5652
rect 14808 5472 14860 5486
rect 15096 5862 15148 5876
rect 15096 5696 15106 5862
rect 15106 5696 15140 5862
rect 15140 5696 15148 5862
rect 15000 5486 15010 5652
rect 15010 5486 15044 5652
rect 15044 5486 15052 5652
rect 15000 5472 15052 5486
rect 15288 5862 15340 5876
rect 15288 5696 15298 5862
rect 15298 5696 15332 5862
rect 15332 5696 15340 5862
rect 15192 5486 15202 5652
rect 15202 5486 15236 5652
rect 15236 5486 15244 5652
rect 15192 5472 15244 5486
rect 15480 5862 15532 5876
rect 15480 5696 15490 5862
rect 15490 5696 15524 5862
rect 15524 5696 15532 5862
rect 15384 5486 15394 5652
rect 15394 5486 15428 5652
rect 15428 5486 15436 5652
rect 15384 5472 15436 5486
rect 15576 5486 15586 5652
rect 15586 5486 15620 5652
rect 15620 5486 15628 5652
rect 15576 5472 15628 5486
rect 16512 5862 16564 5876
rect 16512 5696 16522 5862
rect 16522 5696 16556 5862
rect 16556 5696 16564 5862
rect 16416 5486 16426 5652
rect 16426 5486 16460 5652
rect 16460 5486 16468 5652
rect 16416 5472 16468 5486
rect 16704 5862 16756 5876
rect 16704 5696 16714 5862
rect 16714 5696 16748 5862
rect 16748 5696 16756 5862
rect 16608 5486 16618 5652
rect 16618 5486 16652 5652
rect 16652 5486 16660 5652
rect 16608 5472 16660 5486
rect 16896 5862 16948 5876
rect 16896 5696 16906 5862
rect 16906 5696 16940 5862
rect 16940 5696 16948 5862
rect 16800 5486 16810 5652
rect 16810 5486 16844 5652
rect 16844 5486 16852 5652
rect 16800 5472 16852 5486
rect 17088 5862 17140 5876
rect 17088 5696 17098 5862
rect 17098 5696 17132 5862
rect 17132 5696 17140 5862
rect 16992 5486 17002 5652
rect 17002 5486 17036 5652
rect 17036 5486 17044 5652
rect 16992 5472 17044 5486
rect 17280 5862 17332 5876
rect 17280 5696 17290 5862
rect 17290 5696 17324 5862
rect 17324 5696 17332 5862
rect 17184 5486 17194 5652
rect 17194 5486 17228 5652
rect 17228 5486 17236 5652
rect 17184 5472 17236 5486
rect 17376 5486 17386 5652
rect 17386 5486 17420 5652
rect 17420 5486 17428 5652
rect 17376 5472 17428 5486
rect 18312 5862 18364 5876
rect 18312 5696 18322 5862
rect 18322 5696 18356 5862
rect 18356 5696 18364 5862
rect 18216 5486 18226 5652
rect 18226 5486 18260 5652
rect 18260 5486 18268 5652
rect 18216 5472 18268 5486
rect 18504 5862 18556 5876
rect 18504 5696 18514 5862
rect 18514 5696 18548 5862
rect 18548 5696 18556 5862
rect 18408 5486 18418 5652
rect 18418 5486 18452 5652
rect 18452 5486 18460 5652
rect 18408 5472 18460 5486
rect 18696 5862 18748 5876
rect 18696 5696 18706 5862
rect 18706 5696 18740 5862
rect 18740 5696 18748 5862
rect 18600 5486 18610 5652
rect 18610 5486 18644 5652
rect 18644 5486 18652 5652
rect 18600 5472 18652 5486
rect 18888 5862 18940 5876
rect 18888 5696 18898 5862
rect 18898 5696 18932 5862
rect 18932 5696 18940 5862
rect 18792 5486 18802 5652
rect 18802 5486 18836 5652
rect 18836 5486 18844 5652
rect 18792 5472 18844 5486
rect 19080 5862 19132 5876
rect 19080 5696 19090 5862
rect 19090 5696 19124 5862
rect 19124 5696 19132 5862
rect 18984 5486 18994 5652
rect 18994 5486 19028 5652
rect 19028 5486 19036 5652
rect 18984 5472 19036 5486
rect 19176 5486 19186 5652
rect 19186 5486 19220 5652
rect 19220 5486 19228 5652
rect 19176 5472 19228 5486
rect 20112 5862 20164 5876
rect 20112 5696 20122 5862
rect 20122 5696 20156 5862
rect 20156 5696 20164 5862
rect 20016 5486 20026 5652
rect 20026 5486 20060 5652
rect 20060 5486 20068 5652
rect 20016 5472 20068 5486
rect 20304 5862 20356 5876
rect 20304 5696 20314 5862
rect 20314 5696 20348 5862
rect 20348 5696 20356 5862
rect 20208 5486 20218 5652
rect 20218 5486 20252 5652
rect 20252 5486 20260 5652
rect 20208 5472 20260 5486
rect 20496 5862 20548 5876
rect 20496 5696 20506 5862
rect 20506 5696 20540 5862
rect 20540 5696 20548 5862
rect 20400 5486 20410 5652
rect 20410 5486 20444 5652
rect 20444 5486 20452 5652
rect 20400 5472 20452 5486
rect 20688 5862 20740 5876
rect 20688 5696 20698 5862
rect 20698 5696 20732 5862
rect 20732 5696 20740 5862
rect 20592 5486 20602 5652
rect 20602 5486 20636 5652
rect 20636 5486 20644 5652
rect 20592 5472 20644 5486
rect 20880 5862 20932 5876
rect 20880 5696 20890 5862
rect 20890 5696 20924 5862
rect 20924 5696 20932 5862
rect 20784 5486 20794 5652
rect 20794 5486 20828 5652
rect 20828 5486 20836 5652
rect 20784 5472 20836 5486
rect 20976 5486 20986 5652
rect 20986 5486 21020 5652
rect 21020 5486 21028 5652
rect 20976 5472 21028 5486
rect 21488 5580 21772 6080
rect 22112 5924 22168 5940
rect 22112 5756 22122 5924
rect 22122 5756 22156 5924
rect 22156 5756 22168 5924
rect 11480 4580 11820 4860
rect 13996 4400 14428 5092
rect 14712 5244 14764 5260
rect 14712 5080 14722 5244
rect 14722 5080 14756 5244
rect 14756 5080 14764 5244
rect 14616 4868 14626 5036
rect 14626 4868 14660 5036
rect 14660 4868 14668 5036
rect 14616 4856 14668 4868
rect 14904 5244 14956 5260
rect 14904 5080 14914 5244
rect 14914 5080 14948 5244
rect 14948 5080 14956 5244
rect 14808 4868 14818 5036
rect 14818 4868 14852 5036
rect 14852 4868 14860 5036
rect 14808 4856 14860 4868
rect 15096 5244 15148 5260
rect 15096 5080 15106 5244
rect 15106 5080 15140 5244
rect 15140 5080 15148 5244
rect 15000 4868 15010 5036
rect 15010 4868 15044 5036
rect 15044 4868 15052 5036
rect 15000 4856 15052 4868
rect 15288 5244 15340 5260
rect 15288 5080 15298 5244
rect 15298 5080 15332 5244
rect 15332 5080 15340 5244
rect 15192 4868 15202 5036
rect 15202 4868 15236 5036
rect 15236 4868 15244 5036
rect 15192 4856 15244 4868
rect 15480 5244 15532 5260
rect 15480 5080 15490 5244
rect 15490 5080 15524 5244
rect 15524 5080 15532 5244
rect 15384 4868 15394 5036
rect 15394 4868 15428 5036
rect 15428 4868 15436 5036
rect 15384 4856 15436 4868
rect 15576 4868 15586 5036
rect 15586 4868 15620 5036
rect 15620 4868 15628 5036
rect 15576 4856 15628 4868
rect 16512 5244 16564 5260
rect 16512 5080 16522 5244
rect 16522 5080 16556 5244
rect 16556 5080 16564 5244
rect 16416 4868 16426 5036
rect 16426 4868 16460 5036
rect 16460 4868 16468 5036
rect 16416 4856 16468 4868
rect 16704 5244 16756 5260
rect 16704 5080 16714 5244
rect 16714 5080 16748 5244
rect 16748 5080 16756 5244
rect 16608 4868 16618 5036
rect 16618 4868 16652 5036
rect 16652 4868 16660 5036
rect 16608 4856 16660 4868
rect 16896 5244 16948 5260
rect 16896 5080 16906 5244
rect 16906 5080 16940 5244
rect 16940 5080 16948 5244
rect 16800 4868 16810 5036
rect 16810 4868 16844 5036
rect 16844 4868 16852 5036
rect 16800 4856 16852 4868
rect 17088 5244 17140 5260
rect 17088 5080 17098 5244
rect 17098 5080 17132 5244
rect 17132 5080 17140 5244
rect 16992 4868 17002 5036
rect 17002 4868 17036 5036
rect 17036 4868 17044 5036
rect 16992 4856 17044 4868
rect 17280 5244 17332 5260
rect 17280 5080 17290 5244
rect 17290 5080 17324 5244
rect 17324 5080 17332 5244
rect 17184 4868 17194 5036
rect 17194 4868 17228 5036
rect 17228 4868 17236 5036
rect 17184 4856 17236 4868
rect 17376 4868 17386 5036
rect 17386 4868 17420 5036
rect 17420 4868 17428 5036
rect 17376 4856 17428 4868
rect 18312 5244 18364 5260
rect 18312 5080 18322 5244
rect 18322 5080 18356 5244
rect 18356 5080 18364 5244
rect 18216 4868 18226 5036
rect 18226 4868 18260 5036
rect 18260 4868 18268 5036
rect 18216 4856 18268 4868
rect 18504 5244 18556 5260
rect 18504 5080 18514 5244
rect 18514 5080 18548 5244
rect 18548 5080 18556 5244
rect 18408 4868 18418 5036
rect 18418 4868 18452 5036
rect 18452 4868 18460 5036
rect 18408 4856 18460 4868
rect 18696 5244 18748 5260
rect 18696 5080 18706 5244
rect 18706 5080 18740 5244
rect 18740 5080 18748 5244
rect 18600 4868 18610 5036
rect 18610 4868 18644 5036
rect 18644 4868 18652 5036
rect 18600 4856 18652 4868
rect 18888 5244 18940 5260
rect 18888 5080 18898 5244
rect 18898 5080 18932 5244
rect 18932 5080 18940 5244
rect 18792 4868 18802 5036
rect 18802 4868 18836 5036
rect 18836 4868 18844 5036
rect 18792 4856 18844 4868
rect 19080 5244 19132 5260
rect 19080 5080 19090 5244
rect 19090 5080 19124 5244
rect 19124 5080 19132 5244
rect 18984 4868 18994 5036
rect 18994 4868 19028 5036
rect 19028 4868 19036 5036
rect 18984 4856 19036 4868
rect 19176 4868 19186 5036
rect 19186 4868 19220 5036
rect 19220 4868 19228 5036
rect 19176 4856 19228 4868
rect 20112 5244 20164 5260
rect 20112 5080 20122 5244
rect 20122 5080 20156 5244
rect 20156 5080 20164 5244
rect 20016 4868 20026 5036
rect 20026 4868 20060 5036
rect 20060 4868 20068 5036
rect 20016 4856 20068 4868
rect 20304 5244 20356 5260
rect 20304 5080 20314 5244
rect 20314 5080 20348 5244
rect 20348 5080 20356 5244
rect 20208 4868 20218 5036
rect 20218 4868 20252 5036
rect 20252 4868 20260 5036
rect 20208 4856 20260 4868
rect 20496 5244 20548 5260
rect 20496 5080 20506 5244
rect 20506 5080 20540 5244
rect 20540 5080 20548 5244
rect 20400 4868 20410 5036
rect 20410 4868 20444 5036
rect 20444 4868 20452 5036
rect 20400 4856 20452 4868
rect 20688 5244 20740 5260
rect 20688 5080 20698 5244
rect 20698 5080 20732 5244
rect 20732 5080 20740 5244
rect 20592 4868 20602 5036
rect 20602 4868 20636 5036
rect 20636 4868 20644 5036
rect 20592 4856 20644 4868
rect 20880 5244 20932 5260
rect 20880 5080 20890 5244
rect 20890 5080 20924 5244
rect 20924 5080 20932 5244
rect 20784 4868 20794 5036
rect 20794 4868 20828 5036
rect 20828 4868 20836 5036
rect 20784 4856 20836 4868
rect 20976 4868 20986 5036
rect 20986 4868 21020 5036
rect 21020 4868 21028 5036
rect 20976 4856 21028 4868
rect 22016 5548 22026 5720
rect 22026 5548 22060 5720
rect 22060 5548 22072 5720
rect 22016 5536 22072 5548
rect 22304 5924 22360 5940
rect 22304 5756 22314 5924
rect 22314 5756 22348 5924
rect 22348 5756 22360 5924
rect 22208 5548 22218 5720
rect 22218 5548 22252 5720
rect 22252 5548 22264 5720
rect 22208 5536 22264 5548
rect 22496 5924 22552 5940
rect 22496 5756 22506 5924
rect 22506 5756 22540 5924
rect 22540 5756 22552 5924
rect 22400 5548 22410 5720
rect 22410 5548 22444 5720
rect 22444 5548 22456 5720
rect 22400 5536 22456 5548
rect 22688 5924 22744 5940
rect 22688 5756 22698 5924
rect 22698 5756 22732 5924
rect 22732 5756 22744 5924
rect 22592 5548 22602 5720
rect 22602 5548 22636 5720
rect 22636 5548 22648 5720
rect 22592 5536 22648 5548
rect 22880 5924 22936 5940
rect 22880 5756 22890 5924
rect 22890 5756 22924 5924
rect 22924 5756 22936 5924
rect 22784 5548 22794 5720
rect 22794 5548 22828 5720
rect 22828 5548 22840 5720
rect 22784 5536 22840 5548
rect 23072 5924 23128 5940
rect 23072 5756 23082 5924
rect 23082 5756 23116 5924
rect 23116 5756 23128 5924
rect 22976 5548 22986 5720
rect 22986 5548 23020 5720
rect 23020 5548 23032 5720
rect 22976 5536 23032 5548
rect 23264 5924 23320 5940
rect 23264 5756 23274 5924
rect 23274 5756 23308 5924
rect 23308 5756 23320 5924
rect 23168 5548 23178 5720
rect 23178 5548 23212 5720
rect 23212 5548 23224 5720
rect 23168 5536 23224 5548
rect 23456 5924 23512 5940
rect 23456 5756 23466 5924
rect 23466 5756 23500 5924
rect 23500 5756 23512 5924
rect 23360 5548 23370 5720
rect 23370 5548 23404 5720
rect 23404 5548 23416 5720
rect 23360 5536 23416 5548
rect 23648 5924 23704 5940
rect 23648 5756 23658 5924
rect 23658 5756 23692 5924
rect 23692 5756 23704 5924
rect 23552 5548 23562 5720
rect 23562 5548 23596 5720
rect 23596 5548 23608 5720
rect 23552 5536 23608 5548
rect 23840 5924 23896 5940
rect 23840 5756 23850 5924
rect 23850 5756 23884 5924
rect 23884 5756 23896 5924
rect 23744 5548 23754 5720
rect 23754 5548 23788 5720
rect 23788 5548 23800 5720
rect 23744 5536 23800 5548
rect 23936 5548 23946 5720
rect 23946 5548 23980 5720
rect 23980 5548 23992 5720
rect 23936 5536 23992 5548
rect 22112 5306 22168 5320
rect 22112 5136 22122 5306
rect 22122 5136 22156 5306
rect 22156 5136 22168 5306
rect 22016 4930 22026 5100
rect 22026 4930 22060 5100
rect 22060 4930 22072 5100
rect 22016 4916 22072 4930
rect 22304 5306 22360 5320
rect 22304 5136 22314 5306
rect 22314 5136 22348 5306
rect 22348 5136 22360 5306
rect 22208 4930 22218 5100
rect 22218 4930 22252 5100
rect 22252 4930 22264 5100
rect 22208 4916 22264 4930
rect 22496 5306 22552 5320
rect 22496 5136 22506 5306
rect 22506 5136 22540 5306
rect 22540 5136 22552 5306
rect 22400 4930 22410 5100
rect 22410 4930 22444 5100
rect 22444 4930 22456 5100
rect 22400 4916 22456 4930
rect 22688 5306 22744 5320
rect 22688 5136 22698 5306
rect 22698 5136 22732 5306
rect 22732 5136 22744 5306
rect 22592 4930 22602 5100
rect 22602 4930 22636 5100
rect 22636 4930 22648 5100
rect 22592 4916 22648 4930
rect 22880 5306 22936 5320
rect 22880 5136 22890 5306
rect 22890 5136 22924 5306
rect 22924 5136 22936 5306
rect 22784 4930 22794 5100
rect 22794 4930 22828 5100
rect 22828 4930 22840 5100
rect 22784 4916 22840 4930
rect 23072 5306 23128 5320
rect 23072 5136 23082 5306
rect 23082 5136 23116 5306
rect 23116 5136 23128 5306
rect 22976 4930 22986 5100
rect 22986 4930 23020 5100
rect 23020 4930 23032 5100
rect 22976 4916 23032 4930
rect 23264 5306 23320 5320
rect 23264 5136 23274 5306
rect 23274 5136 23308 5306
rect 23308 5136 23320 5306
rect 23168 4930 23178 5100
rect 23178 4930 23212 5100
rect 23212 4930 23224 5100
rect 23168 4916 23224 4930
rect 23456 5306 23512 5320
rect 23456 5136 23466 5306
rect 23466 5136 23500 5306
rect 23500 5136 23512 5306
rect 23360 4930 23370 5100
rect 23370 4930 23404 5100
rect 23404 4930 23416 5100
rect 23360 4916 23416 4930
rect 23648 5306 23704 5320
rect 23648 5136 23658 5306
rect 23658 5136 23692 5306
rect 23692 5136 23704 5306
rect 23552 4930 23562 5100
rect 23562 4930 23596 5100
rect 23596 4930 23608 5100
rect 23552 4916 23608 4930
rect 23840 5306 23896 5320
rect 23840 5136 23850 5306
rect 23850 5136 23884 5306
rect 23884 5136 23896 5306
rect 23744 4930 23754 5100
rect 23754 4930 23788 5100
rect 23788 4930 23800 5100
rect 23744 4916 23800 4930
rect 23936 4930 23946 5100
rect 23946 4930 23980 5100
rect 23980 4930 23992 5100
rect 23936 4916 23992 4930
rect 14712 4626 14764 4640
rect 14712 4460 14722 4626
rect 14722 4460 14756 4626
rect 14756 4460 14764 4626
rect 14616 4250 14626 4416
rect 14626 4250 14660 4416
rect 14660 4250 14668 4416
rect 14616 4236 14668 4250
rect 14904 4626 14956 4640
rect 14904 4460 14914 4626
rect 14914 4460 14948 4626
rect 14948 4460 14956 4626
rect 14808 4250 14818 4416
rect 14818 4250 14852 4416
rect 14852 4250 14860 4416
rect 14808 4236 14860 4250
rect 15096 4626 15148 4640
rect 15096 4460 15106 4626
rect 15106 4460 15140 4626
rect 15140 4460 15148 4626
rect 15000 4250 15010 4416
rect 15010 4250 15044 4416
rect 15044 4250 15052 4416
rect 15000 4236 15052 4250
rect 15288 4626 15340 4640
rect 15288 4460 15298 4626
rect 15298 4460 15332 4626
rect 15332 4460 15340 4626
rect 15192 4250 15202 4416
rect 15202 4250 15236 4416
rect 15236 4250 15244 4416
rect 15192 4236 15244 4250
rect 15480 4626 15532 4640
rect 15480 4460 15490 4626
rect 15490 4460 15524 4626
rect 15524 4460 15532 4626
rect 15384 4250 15394 4416
rect 15394 4250 15428 4416
rect 15428 4250 15436 4416
rect 15384 4236 15436 4250
rect 15576 4250 15586 4416
rect 15586 4250 15620 4416
rect 15620 4250 15628 4416
rect 15576 4236 15628 4250
rect 16512 4626 16564 4640
rect 16512 4460 16522 4626
rect 16522 4460 16556 4626
rect 16556 4460 16564 4626
rect 16416 4250 16426 4416
rect 16426 4250 16460 4416
rect 16460 4250 16468 4416
rect 16416 4236 16468 4250
rect 16704 4626 16756 4640
rect 16704 4460 16714 4626
rect 16714 4460 16748 4626
rect 16748 4460 16756 4626
rect 16608 4250 16618 4416
rect 16618 4250 16652 4416
rect 16652 4250 16660 4416
rect 16608 4236 16660 4250
rect 16896 4626 16948 4640
rect 16896 4460 16906 4626
rect 16906 4460 16940 4626
rect 16940 4460 16948 4626
rect 16800 4250 16810 4416
rect 16810 4250 16844 4416
rect 16844 4250 16852 4416
rect 16800 4236 16852 4250
rect 17088 4626 17140 4640
rect 17088 4460 17098 4626
rect 17098 4460 17132 4626
rect 17132 4460 17140 4626
rect 16992 4250 17002 4416
rect 17002 4250 17036 4416
rect 17036 4250 17044 4416
rect 16992 4236 17044 4250
rect 17280 4626 17332 4640
rect 17280 4460 17290 4626
rect 17290 4460 17324 4626
rect 17324 4460 17332 4626
rect 17184 4250 17194 4416
rect 17194 4250 17228 4416
rect 17228 4250 17236 4416
rect 17184 4236 17236 4250
rect 17376 4250 17386 4416
rect 17386 4250 17420 4416
rect 17420 4250 17428 4416
rect 17376 4236 17428 4250
rect 18312 4626 18364 4640
rect 18312 4460 18322 4626
rect 18322 4460 18356 4626
rect 18356 4460 18364 4626
rect 18216 4250 18226 4416
rect 18226 4250 18260 4416
rect 18260 4250 18268 4416
rect 18216 4236 18268 4250
rect 18504 4626 18556 4640
rect 18504 4460 18514 4626
rect 18514 4460 18548 4626
rect 18548 4460 18556 4626
rect 18408 4250 18418 4416
rect 18418 4250 18452 4416
rect 18452 4250 18460 4416
rect 18408 4236 18460 4250
rect 18696 4626 18748 4640
rect 18696 4460 18706 4626
rect 18706 4460 18740 4626
rect 18740 4460 18748 4626
rect 18600 4250 18610 4416
rect 18610 4250 18644 4416
rect 18644 4250 18652 4416
rect 18600 4236 18652 4250
rect 18888 4626 18940 4640
rect 18888 4460 18898 4626
rect 18898 4460 18932 4626
rect 18932 4460 18940 4626
rect 18792 4250 18802 4416
rect 18802 4250 18836 4416
rect 18836 4250 18844 4416
rect 18792 4236 18844 4250
rect 19080 4626 19132 4640
rect 19080 4460 19090 4626
rect 19090 4460 19124 4626
rect 19124 4460 19132 4626
rect 18984 4250 18994 4416
rect 18994 4250 19028 4416
rect 19028 4250 19036 4416
rect 18984 4236 19036 4250
rect 19176 4250 19186 4416
rect 19186 4250 19220 4416
rect 19220 4250 19228 4416
rect 19176 4236 19228 4250
rect 20112 4626 20164 4640
rect 20112 4460 20122 4626
rect 20122 4460 20156 4626
rect 20156 4460 20164 4626
rect 20016 4250 20026 4416
rect 20026 4250 20060 4416
rect 20060 4250 20068 4416
rect 20016 4236 20068 4250
rect 20304 4626 20356 4640
rect 20304 4460 20314 4626
rect 20314 4460 20348 4626
rect 20348 4460 20356 4626
rect 20208 4250 20218 4416
rect 20218 4250 20252 4416
rect 20252 4250 20260 4416
rect 20208 4236 20260 4250
rect 20496 4626 20548 4640
rect 20496 4460 20506 4626
rect 20506 4460 20540 4626
rect 20540 4460 20548 4626
rect 20400 4250 20410 4416
rect 20410 4250 20444 4416
rect 20444 4250 20452 4416
rect 20400 4236 20452 4250
rect 20688 4626 20740 4640
rect 20688 4460 20698 4626
rect 20698 4460 20732 4626
rect 20732 4460 20740 4626
rect 20592 4250 20602 4416
rect 20602 4250 20636 4416
rect 20636 4250 20644 4416
rect 20592 4236 20644 4250
rect 20880 4626 20932 4640
rect 20880 4460 20890 4626
rect 20890 4460 20924 4626
rect 20924 4460 20932 4626
rect 20784 4250 20794 4416
rect 20794 4250 20828 4416
rect 20828 4250 20836 4416
rect 20784 4236 20836 4250
rect 20976 4250 20986 4416
rect 20986 4250 21020 4416
rect 21020 4250 21028 4416
rect 20976 4236 21028 4250
rect 24520 4360 24900 4700
rect -10060 3996 -10008 4008
rect -10060 3828 -10050 3996
rect -10050 3828 -10016 3996
rect -10016 3828 -10008 3996
rect -9800 3620 -9792 3788
rect -9792 3620 -9758 3788
rect -9758 3620 -9748 3788
rect -9800 3608 -9748 3620
rect -9544 3996 -9492 4008
rect -9544 3828 -9534 3996
rect -9534 3828 -9500 3996
rect -9500 3828 -9492 3996
rect -9284 3620 -9276 3788
rect -9276 3620 -9242 3788
rect -9242 3620 -9232 3788
rect -9284 3608 -9232 3620
rect -9028 3996 -8976 4008
rect -9028 3828 -9018 3996
rect -9018 3828 -8984 3996
rect -8984 3828 -8976 3996
rect -8768 3620 -8760 3788
rect -8760 3620 -8726 3788
rect -8726 3620 -8716 3788
rect -8768 3608 -8716 3620
rect 216 3716 268 3728
rect 216 3548 226 3716
rect 226 3548 260 3716
rect 260 3548 268 3716
rect -10060 3378 -10008 3392
rect -10060 3212 -10050 3378
rect -10050 3212 -10016 3378
rect -10016 3212 -10008 3378
rect -9800 3002 -9792 3172
rect -9792 3002 -9758 3172
rect -9758 3002 -9748 3172
rect -9800 2992 -9748 3002
rect -9544 3378 -9492 3392
rect -9544 3212 -9534 3378
rect -9534 3212 -9500 3378
rect -9500 3212 -9492 3378
rect -9284 3002 -9276 3172
rect -9276 3002 -9242 3172
rect -9242 3002 -9232 3172
rect -9284 2992 -9232 3002
rect -9028 3378 -8976 3392
rect -9028 3212 -9018 3378
rect -9018 3212 -8984 3378
rect -8984 3212 -8976 3378
rect 476 3340 484 3508
rect 484 3340 518 3508
rect 518 3340 528 3508
rect 476 3328 528 3340
rect 732 3716 784 3728
rect 732 3548 742 3716
rect 742 3548 776 3716
rect 776 3548 784 3716
rect 992 3340 1000 3508
rect 1000 3340 1034 3508
rect 1034 3340 1044 3508
rect 992 3328 1044 3340
rect 1248 3716 1300 3728
rect 1248 3548 1258 3716
rect 1258 3548 1292 3716
rect 1292 3548 1300 3716
rect 2016 3716 2068 3728
rect 2016 3548 2026 3716
rect 2026 3548 2060 3716
rect 2060 3548 2068 3716
rect 1508 3340 1516 3508
rect 1516 3340 1550 3508
rect 1550 3340 1560 3508
rect 1508 3328 1560 3340
rect 2276 3340 2284 3508
rect 2284 3340 2318 3508
rect 2318 3340 2328 3508
rect 2276 3328 2328 3340
rect 2532 3716 2584 3728
rect 2532 3548 2542 3716
rect 2542 3548 2576 3716
rect 2576 3548 2584 3716
rect 2792 3340 2800 3508
rect 2800 3340 2834 3508
rect 2834 3340 2844 3508
rect 2792 3328 2844 3340
rect 3048 3716 3100 3728
rect 3048 3548 3058 3716
rect 3058 3548 3092 3716
rect 3092 3548 3100 3716
rect 3816 3716 3868 3728
rect 3816 3548 3826 3716
rect 3826 3548 3860 3716
rect 3860 3548 3868 3716
rect 3308 3340 3316 3508
rect 3316 3340 3350 3508
rect 3350 3340 3360 3508
rect 3308 3328 3360 3340
rect 4076 3340 4084 3508
rect 4084 3340 4118 3508
rect 4118 3340 4128 3508
rect 4076 3328 4128 3340
rect 4332 3716 4384 3728
rect 4332 3548 4342 3716
rect 4342 3548 4376 3716
rect 4376 3548 4384 3716
rect 4592 3340 4600 3508
rect 4600 3340 4634 3508
rect 4634 3340 4644 3508
rect 4592 3328 4644 3340
rect 4848 3716 4900 3728
rect 4848 3548 4858 3716
rect 4858 3548 4892 3716
rect 4892 3548 4900 3716
rect 5616 3716 5668 3728
rect 5616 3548 5626 3716
rect 5626 3548 5660 3716
rect 5660 3548 5668 3716
rect 5108 3340 5116 3508
rect 5116 3340 5150 3508
rect 5150 3340 5160 3508
rect 5108 3328 5160 3340
rect 5876 3340 5884 3508
rect 5884 3340 5918 3508
rect 5918 3340 5928 3508
rect 5876 3328 5928 3340
rect 6132 3716 6184 3728
rect 6132 3548 6142 3716
rect 6142 3548 6176 3716
rect 6176 3548 6184 3716
rect 6392 3340 6400 3508
rect 6400 3340 6434 3508
rect 6434 3340 6444 3508
rect 6392 3328 6444 3340
rect 6648 3716 6700 3728
rect 6648 3548 6658 3716
rect 6658 3548 6692 3716
rect 6692 3548 6700 3716
rect 14616 3716 14668 3728
rect 14616 3548 14626 3716
rect 14626 3548 14660 3716
rect 14660 3548 14668 3716
rect 6908 3340 6916 3508
rect 6916 3340 6950 3508
rect 6950 3340 6960 3508
rect 6908 3328 6960 3340
rect 14876 3340 14884 3508
rect 14884 3340 14918 3508
rect 14918 3340 14928 3508
rect 14876 3328 14928 3340
rect 15132 3716 15184 3728
rect 15132 3548 15142 3716
rect 15142 3548 15176 3716
rect 15176 3548 15184 3716
rect 15392 3340 15400 3508
rect 15400 3340 15434 3508
rect 15434 3340 15444 3508
rect 15392 3328 15444 3340
rect 15648 3716 15700 3728
rect 15648 3548 15658 3716
rect 15658 3548 15692 3716
rect 15692 3548 15700 3716
rect 16416 3716 16468 3728
rect 16416 3548 16426 3716
rect 16426 3548 16460 3716
rect 16460 3548 16468 3716
rect 15908 3340 15916 3508
rect 15916 3340 15950 3508
rect 15950 3340 15960 3508
rect 15908 3328 15960 3340
rect 16676 3340 16684 3508
rect 16684 3340 16718 3508
rect 16718 3340 16728 3508
rect 16676 3328 16728 3340
rect 16932 3716 16984 3728
rect 16932 3548 16942 3716
rect 16942 3548 16976 3716
rect 16976 3548 16984 3716
rect 17192 3340 17200 3508
rect 17200 3340 17234 3508
rect 17234 3340 17244 3508
rect 17192 3328 17244 3340
rect 17448 3716 17500 3728
rect 17448 3548 17458 3716
rect 17458 3548 17492 3716
rect 17492 3548 17500 3716
rect 18216 3716 18268 3728
rect 18216 3548 18226 3716
rect 18226 3548 18260 3716
rect 18260 3548 18268 3716
rect 17708 3340 17716 3508
rect 17716 3340 17750 3508
rect 17750 3340 17760 3508
rect 17708 3328 17760 3340
rect 18476 3340 18484 3508
rect 18484 3340 18518 3508
rect 18518 3340 18528 3508
rect 18476 3328 18528 3340
rect 18732 3716 18784 3728
rect 18732 3548 18742 3716
rect 18742 3548 18776 3716
rect 18776 3548 18784 3716
rect 18992 3340 19000 3508
rect 19000 3340 19034 3508
rect 19034 3340 19044 3508
rect 18992 3328 19044 3340
rect 19248 3716 19300 3728
rect 19248 3548 19258 3716
rect 19258 3548 19292 3716
rect 19292 3548 19300 3716
rect 20016 3716 20068 3728
rect 20016 3548 20026 3716
rect 20026 3548 20060 3716
rect 20060 3548 20068 3716
rect 19508 3340 19516 3508
rect 19516 3340 19550 3508
rect 19550 3340 19560 3508
rect 19508 3328 19560 3340
rect 20276 3340 20284 3508
rect 20284 3340 20318 3508
rect 20318 3340 20328 3508
rect 20276 3328 20328 3340
rect 20532 3716 20584 3728
rect 20532 3548 20542 3716
rect 20542 3548 20576 3716
rect 20576 3548 20584 3716
rect 20792 3340 20800 3508
rect 20800 3340 20834 3508
rect 20834 3340 20844 3508
rect 20792 3328 20844 3340
rect 21048 3716 21100 3728
rect 21048 3548 21058 3716
rect 21058 3548 21092 3716
rect 21092 3548 21100 3716
rect 21308 3340 21316 3508
rect 21316 3340 21350 3508
rect 21350 3340 21360 3508
rect 21308 3328 21360 3340
rect -8768 3002 -8760 3172
rect -8760 3002 -8726 3172
rect -8726 3002 -8716 3172
rect -8768 2992 -8716 3002
rect 216 3098 268 3112
rect 216 2932 226 3098
rect 226 2932 260 3098
rect 260 2932 268 3098
rect -10060 2760 -10008 2772
rect -10060 2592 -10050 2760
rect -10050 2592 -10016 2760
rect -10016 2592 -10008 2760
rect -9800 2384 -9792 2552
rect -9792 2384 -9758 2552
rect -9758 2384 -9748 2552
rect -9800 2372 -9748 2384
rect -9544 2760 -9492 2772
rect -9544 2592 -9534 2760
rect -9534 2592 -9500 2760
rect -9500 2592 -9492 2760
rect -9284 2384 -9276 2552
rect -9276 2384 -9242 2552
rect -9242 2384 -9232 2552
rect -9284 2372 -9232 2384
rect -9028 2760 -8976 2772
rect -9028 2592 -9018 2760
rect -9018 2592 -8984 2760
rect -8984 2592 -8976 2760
rect 476 2722 484 2892
rect 484 2722 518 2892
rect 518 2722 528 2892
rect 476 2712 528 2722
rect 732 3098 784 3112
rect 732 2932 742 3098
rect 742 2932 776 3098
rect 776 2932 784 3098
rect 992 2722 1000 2892
rect 1000 2722 1034 2892
rect 1034 2722 1044 2892
rect 992 2712 1044 2722
rect 1248 3098 1300 3112
rect 1248 2932 1258 3098
rect 1258 2932 1292 3098
rect 1292 2932 1300 3098
rect 2016 3098 2068 3112
rect 2016 2932 2026 3098
rect 2026 2932 2060 3098
rect 2060 2932 2068 3098
rect 1508 2722 1516 2892
rect 1516 2722 1550 2892
rect 1550 2722 1560 2892
rect 1508 2712 1560 2722
rect 2276 2722 2284 2892
rect 2284 2722 2318 2892
rect 2318 2722 2328 2892
rect 2276 2712 2328 2722
rect 2532 3098 2584 3112
rect 2532 2932 2542 3098
rect 2542 2932 2576 3098
rect 2576 2932 2584 3098
rect 2792 2722 2800 2892
rect 2800 2722 2834 2892
rect 2834 2722 2844 2892
rect 2792 2712 2844 2722
rect 3048 3098 3100 3112
rect 3048 2932 3058 3098
rect 3058 2932 3092 3098
rect 3092 2932 3100 3098
rect 3816 3098 3868 3112
rect 3816 2932 3826 3098
rect 3826 2932 3860 3098
rect 3860 2932 3868 3098
rect 3308 2722 3316 2892
rect 3316 2722 3350 2892
rect 3350 2722 3360 2892
rect 3308 2712 3360 2722
rect 4076 2722 4084 2892
rect 4084 2722 4118 2892
rect 4118 2722 4128 2892
rect 4076 2712 4128 2722
rect 4332 3098 4384 3112
rect 4332 2932 4342 3098
rect 4342 2932 4376 3098
rect 4376 2932 4384 3098
rect 4592 2722 4600 2892
rect 4600 2722 4634 2892
rect 4634 2722 4644 2892
rect 4592 2712 4644 2722
rect 4848 3098 4900 3112
rect 4848 2932 4858 3098
rect 4858 2932 4892 3098
rect 4892 2932 4900 3098
rect 5616 3098 5668 3112
rect 5616 2932 5626 3098
rect 5626 2932 5660 3098
rect 5660 2932 5668 3098
rect 5108 2722 5116 2892
rect 5116 2722 5150 2892
rect 5150 2722 5160 2892
rect 5108 2712 5160 2722
rect 5876 2722 5884 2892
rect 5884 2722 5918 2892
rect 5918 2722 5928 2892
rect 5876 2712 5928 2722
rect 6132 3098 6184 3112
rect 6132 2932 6142 3098
rect 6142 2932 6176 3098
rect 6176 2932 6184 3098
rect 6392 2722 6400 2892
rect 6400 2722 6434 2892
rect 6434 2722 6444 2892
rect 6392 2712 6444 2722
rect 6648 3098 6700 3112
rect 6648 2932 6658 3098
rect 6658 2932 6692 3098
rect 6692 2932 6700 3098
rect 14616 3098 14668 3112
rect 14616 2932 14626 3098
rect 14626 2932 14660 3098
rect 14660 2932 14668 3098
rect 6908 2722 6916 2892
rect 6916 2722 6950 2892
rect 6950 2722 6960 2892
rect 6908 2712 6960 2722
rect 14876 2722 14884 2892
rect 14884 2722 14918 2892
rect 14918 2722 14928 2892
rect 14876 2712 14928 2722
rect 15132 3098 15184 3112
rect 15132 2932 15142 3098
rect 15142 2932 15176 3098
rect 15176 2932 15184 3098
rect 15392 2722 15400 2892
rect 15400 2722 15434 2892
rect 15434 2722 15444 2892
rect 15392 2712 15444 2722
rect 15648 3098 15700 3112
rect 15648 2932 15658 3098
rect 15658 2932 15692 3098
rect 15692 2932 15700 3098
rect 16416 3098 16468 3112
rect 16416 2932 16426 3098
rect 16426 2932 16460 3098
rect 16460 2932 16468 3098
rect 15908 2722 15916 2892
rect 15916 2722 15950 2892
rect 15950 2722 15960 2892
rect 15908 2712 15960 2722
rect 16676 2722 16684 2892
rect 16684 2722 16718 2892
rect 16718 2722 16728 2892
rect 16676 2712 16728 2722
rect 16932 3098 16984 3112
rect 16932 2932 16942 3098
rect 16942 2932 16976 3098
rect 16976 2932 16984 3098
rect 17192 2722 17200 2892
rect 17200 2722 17234 2892
rect 17234 2722 17244 2892
rect 17192 2712 17244 2722
rect 17448 3098 17500 3112
rect 17448 2932 17458 3098
rect 17458 2932 17492 3098
rect 17492 2932 17500 3098
rect 18216 3098 18268 3112
rect 18216 2932 18226 3098
rect 18226 2932 18260 3098
rect 18260 2932 18268 3098
rect 17708 2722 17716 2892
rect 17716 2722 17750 2892
rect 17750 2722 17760 2892
rect 17708 2712 17760 2722
rect 18476 2722 18484 2892
rect 18484 2722 18518 2892
rect 18518 2722 18528 2892
rect 18476 2712 18528 2722
rect 18732 3098 18784 3112
rect 18732 2932 18742 3098
rect 18742 2932 18776 3098
rect 18776 2932 18784 3098
rect 18992 2722 19000 2892
rect 19000 2722 19034 2892
rect 19034 2722 19044 2892
rect 18992 2712 19044 2722
rect 19248 3098 19300 3112
rect 19248 2932 19258 3098
rect 19258 2932 19292 3098
rect 19292 2932 19300 3098
rect 20016 3098 20068 3112
rect 20016 2932 20026 3098
rect 20026 2932 20060 3098
rect 20060 2932 20068 3098
rect 19508 2722 19516 2892
rect 19516 2722 19550 2892
rect 19550 2722 19560 2892
rect 19508 2712 19560 2722
rect 20276 2722 20284 2892
rect 20284 2722 20318 2892
rect 20318 2722 20328 2892
rect 20276 2712 20328 2722
rect 20532 3098 20584 3112
rect 20532 2932 20542 3098
rect 20542 2932 20576 3098
rect 20576 2932 20584 3098
rect 20792 2722 20800 2892
rect 20800 2722 20834 2892
rect 20834 2722 20844 2892
rect 20792 2712 20844 2722
rect 21048 3098 21100 3112
rect 21048 2932 21058 3098
rect 21058 2932 21092 3098
rect 21092 2932 21100 3098
rect 21308 2722 21316 2892
rect 21316 2722 21350 2892
rect 21350 2722 21360 2892
rect 21308 2712 21360 2722
rect -8768 2384 -8760 2552
rect -8760 2384 -8726 2552
rect -8726 2384 -8716 2552
rect -8768 2372 -8716 2384
rect 216 2480 268 2492
rect 216 2312 226 2480
rect 226 2312 260 2480
rect 260 2312 268 2480
rect -10060 2142 -10008 2156
rect -10060 1976 -10050 2142
rect -10050 1976 -10016 2142
rect -10016 1976 -10008 2142
rect -9800 1766 -9792 1936
rect -9792 1766 -9758 1936
rect -9758 1766 -9748 1936
rect -9800 1756 -9748 1766
rect -9544 2142 -9492 2156
rect -9544 1976 -9534 2142
rect -9534 1976 -9500 2142
rect -9500 1976 -9492 2142
rect -9284 1766 -9276 1936
rect -9276 1766 -9242 1936
rect -9242 1766 -9232 1936
rect -9284 1756 -9232 1766
rect -9028 2142 -8976 2156
rect -9028 1976 -9018 2142
rect -9018 1976 -8984 2142
rect -8984 1976 -8976 2142
rect 476 2104 484 2272
rect 484 2104 518 2272
rect 518 2104 528 2272
rect 476 2092 528 2104
rect 732 2480 784 2492
rect 732 2312 742 2480
rect 742 2312 776 2480
rect 776 2312 784 2480
rect 992 2104 1000 2272
rect 1000 2104 1034 2272
rect 1034 2104 1044 2272
rect 992 2092 1044 2104
rect 1248 2480 1300 2492
rect 1248 2312 1258 2480
rect 1258 2312 1292 2480
rect 1292 2312 1300 2480
rect 2016 2480 2068 2492
rect 2016 2312 2026 2480
rect 2026 2312 2060 2480
rect 2060 2312 2068 2480
rect 1508 2104 1516 2272
rect 1516 2104 1550 2272
rect 1550 2104 1560 2272
rect 1508 2092 1560 2104
rect 2276 2104 2284 2272
rect 2284 2104 2318 2272
rect 2318 2104 2328 2272
rect 2276 2092 2328 2104
rect 2532 2480 2584 2492
rect 2532 2312 2542 2480
rect 2542 2312 2576 2480
rect 2576 2312 2584 2480
rect 2792 2104 2800 2272
rect 2800 2104 2834 2272
rect 2834 2104 2844 2272
rect 2792 2092 2844 2104
rect 3048 2480 3100 2492
rect 3048 2312 3058 2480
rect 3058 2312 3092 2480
rect 3092 2312 3100 2480
rect 3816 2480 3868 2492
rect 3816 2312 3826 2480
rect 3826 2312 3860 2480
rect 3860 2312 3868 2480
rect 3308 2104 3316 2272
rect 3316 2104 3350 2272
rect 3350 2104 3360 2272
rect 3308 2092 3360 2104
rect 4076 2104 4084 2272
rect 4084 2104 4118 2272
rect 4118 2104 4128 2272
rect 4076 2092 4128 2104
rect 4332 2480 4384 2492
rect 4332 2312 4342 2480
rect 4342 2312 4376 2480
rect 4376 2312 4384 2480
rect 4592 2104 4600 2272
rect 4600 2104 4634 2272
rect 4634 2104 4644 2272
rect 4592 2092 4644 2104
rect 4848 2480 4900 2492
rect 4848 2312 4858 2480
rect 4858 2312 4892 2480
rect 4892 2312 4900 2480
rect 5616 2480 5668 2492
rect 5616 2312 5626 2480
rect 5626 2312 5660 2480
rect 5660 2312 5668 2480
rect 5108 2104 5116 2272
rect 5116 2104 5150 2272
rect 5150 2104 5160 2272
rect 5108 2092 5160 2104
rect 5876 2104 5884 2272
rect 5884 2104 5918 2272
rect 5918 2104 5928 2272
rect 5876 2092 5928 2104
rect 6132 2480 6184 2492
rect 6132 2312 6142 2480
rect 6142 2312 6176 2480
rect 6176 2312 6184 2480
rect 6392 2104 6400 2272
rect 6400 2104 6434 2272
rect 6434 2104 6444 2272
rect 6392 2092 6444 2104
rect 6648 2480 6700 2492
rect 6648 2312 6658 2480
rect 6658 2312 6692 2480
rect 6692 2312 6700 2480
rect 14616 2480 14668 2492
rect 14616 2312 14626 2480
rect 14626 2312 14660 2480
rect 14660 2312 14668 2480
rect 6908 2104 6916 2272
rect 6916 2104 6950 2272
rect 6950 2104 6960 2272
rect 6908 2092 6960 2104
rect 14876 2104 14884 2272
rect 14884 2104 14918 2272
rect 14918 2104 14928 2272
rect 14876 2092 14928 2104
rect 15132 2480 15184 2492
rect 15132 2312 15142 2480
rect 15142 2312 15176 2480
rect 15176 2312 15184 2480
rect 15392 2104 15400 2272
rect 15400 2104 15434 2272
rect 15434 2104 15444 2272
rect 15392 2092 15444 2104
rect 15648 2480 15700 2492
rect 15648 2312 15658 2480
rect 15658 2312 15692 2480
rect 15692 2312 15700 2480
rect 16416 2480 16468 2492
rect 16416 2312 16426 2480
rect 16426 2312 16460 2480
rect 16460 2312 16468 2480
rect 15908 2104 15916 2272
rect 15916 2104 15950 2272
rect 15950 2104 15960 2272
rect 15908 2092 15960 2104
rect 16676 2104 16684 2272
rect 16684 2104 16718 2272
rect 16718 2104 16728 2272
rect 16676 2092 16728 2104
rect 16932 2480 16984 2492
rect 16932 2312 16942 2480
rect 16942 2312 16976 2480
rect 16976 2312 16984 2480
rect 17192 2104 17200 2272
rect 17200 2104 17234 2272
rect 17234 2104 17244 2272
rect 17192 2092 17244 2104
rect 17448 2480 17500 2492
rect 17448 2312 17458 2480
rect 17458 2312 17492 2480
rect 17492 2312 17500 2480
rect 18216 2480 18268 2492
rect 18216 2312 18226 2480
rect 18226 2312 18260 2480
rect 18260 2312 18268 2480
rect 17708 2104 17716 2272
rect 17716 2104 17750 2272
rect 17750 2104 17760 2272
rect 17708 2092 17760 2104
rect 18476 2104 18484 2272
rect 18484 2104 18518 2272
rect 18518 2104 18528 2272
rect 18476 2092 18528 2104
rect 18732 2480 18784 2492
rect 18732 2312 18742 2480
rect 18742 2312 18776 2480
rect 18776 2312 18784 2480
rect 18992 2104 19000 2272
rect 19000 2104 19034 2272
rect 19034 2104 19044 2272
rect 18992 2092 19044 2104
rect 19248 2480 19300 2492
rect 19248 2312 19258 2480
rect 19258 2312 19292 2480
rect 19292 2312 19300 2480
rect 20016 2480 20068 2492
rect 20016 2312 20026 2480
rect 20026 2312 20060 2480
rect 20060 2312 20068 2480
rect 19508 2104 19516 2272
rect 19516 2104 19550 2272
rect 19550 2104 19560 2272
rect 19508 2092 19560 2104
rect 20276 2104 20284 2272
rect 20284 2104 20318 2272
rect 20318 2104 20328 2272
rect 20276 2092 20328 2104
rect 20532 2480 20584 2492
rect 20532 2312 20542 2480
rect 20542 2312 20576 2480
rect 20576 2312 20584 2480
rect 20792 2104 20800 2272
rect 20800 2104 20834 2272
rect 20834 2104 20844 2272
rect 20792 2092 20844 2104
rect 21048 2480 21100 2492
rect 21048 2312 21058 2480
rect 21058 2312 21092 2480
rect 21092 2312 21100 2480
rect 21308 2104 21316 2272
rect 21316 2104 21350 2272
rect 21350 2104 21360 2272
rect 21308 2092 21360 2104
rect -8768 1766 -8760 1936
rect -8760 1766 -8726 1936
rect -8726 1766 -8716 1936
rect -8768 1756 -8716 1766
rect 216 1862 268 1876
rect 216 1696 226 1862
rect 226 1696 260 1862
rect 260 1696 268 1862
rect -10060 1524 -10008 1536
rect -10060 1356 -10050 1524
rect -10050 1356 -10016 1524
rect -10016 1356 -10008 1524
rect -9800 1148 -9792 1316
rect -9792 1148 -9758 1316
rect -9758 1148 -9748 1316
rect -9800 1136 -9748 1148
rect -9544 1524 -9492 1536
rect -9544 1356 -9534 1524
rect -9534 1356 -9500 1524
rect -9500 1356 -9492 1524
rect -9284 1148 -9276 1316
rect -9276 1148 -9242 1316
rect -9242 1148 -9232 1316
rect -9284 1136 -9232 1148
rect -9028 1524 -8976 1536
rect -9028 1356 -9018 1524
rect -9018 1356 -8984 1524
rect -8984 1356 -8976 1524
rect 476 1486 484 1656
rect 484 1486 518 1656
rect 518 1486 528 1656
rect 476 1476 528 1486
rect 732 1862 784 1876
rect 732 1696 742 1862
rect 742 1696 776 1862
rect 776 1696 784 1862
rect 992 1486 1000 1656
rect 1000 1486 1034 1656
rect 1034 1486 1044 1656
rect 992 1476 1044 1486
rect 1248 1862 1300 1876
rect 1248 1696 1258 1862
rect 1258 1696 1292 1862
rect 1292 1696 1300 1862
rect 2016 1862 2068 1876
rect 2016 1696 2026 1862
rect 2026 1696 2060 1862
rect 2060 1696 2068 1862
rect 1508 1486 1516 1656
rect 1516 1486 1550 1656
rect 1550 1486 1560 1656
rect 1508 1476 1560 1486
rect 2276 1486 2284 1656
rect 2284 1486 2318 1656
rect 2318 1486 2328 1656
rect 2276 1476 2328 1486
rect 2532 1862 2584 1876
rect 2532 1696 2542 1862
rect 2542 1696 2576 1862
rect 2576 1696 2584 1862
rect 2792 1486 2800 1656
rect 2800 1486 2834 1656
rect 2834 1486 2844 1656
rect 2792 1476 2844 1486
rect 3048 1862 3100 1876
rect 3048 1696 3058 1862
rect 3058 1696 3092 1862
rect 3092 1696 3100 1862
rect 3816 1862 3868 1876
rect 3816 1696 3826 1862
rect 3826 1696 3860 1862
rect 3860 1696 3868 1862
rect 3308 1486 3316 1656
rect 3316 1486 3350 1656
rect 3350 1486 3360 1656
rect 3308 1476 3360 1486
rect 4076 1486 4084 1656
rect 4084 1486 4118 1656
rect 4118 1486 4128 1656
rect 4076 1476 4128 1486
rect 4332 1862 4384 1876
rect 4332 1696 4342 1862
rect 4342 1696 4376 1862
rect 4376 1696 4384 1862
rect 4592 1486 4600 1656
rect 4600 1486 4634 1656
rect 4634 1486 4644 1656
rect 4592 1476 4644 1486
rect 4848 1862 4900 1876
rect 4848 1696 4858 1862
rect 4858 1696 4892 1862
rect 4892 1696 4900 1862
rect 5616 1862 5668 1876
rect 5616 1696 5626 1862
rect 5626 1696 5660 1862
rect 5660 1696 5668 1862
rect 5108 1486 5116 1656
rect 5116 1486 5150 1656
rect 5150 1486 5160 1656
rect 5108 1476 5160 1486
rect 5876 1486 5884 1656
rect 5884 1486 5918 1656
rect 5918 1486 5928 1656
rect 5876 1476 5928 1486
rect 6132 1862 6184 1876
rect 6132 1696 6142 1862
rect 6142 1696 6176 1862
rect 6176 1696 6184 1862
rect 6392 1486 6400 1656
rect 6400 1486 6434 1656
rect 6434 1486 6444 1656
rect 6392 1476 6444 1486
rect 6648 1862 6700 1876
rect 6648 1696 6658 1862
rect 6658 1696 6692 1862
rect 6692 1696 6700 1862
rect 14616 1862 14668 1876
rect 14616 1696 14626 1862
rect 14626 1696 14660 1862
rect 14660 1696 14668 1862
rect 6908 1486 6916 1656
rect 6916 1486 6950 1656
rect 6950 1486 6960 1656
rect 6908 1476 6960 1486
rect 14876 1486 14884 1656
rect 14884 1486 14918 1656
rect 14918 1486 14928 1656
rect 14876 1476 14928 1486
rect 15132 1862 15184 1876
rect 15132 1696 15142 1862
rect 15142 1696 15176 1862
rect 15176 1696 15184 1862
rect 15392 1486 15400 1656
rect 15400 1486 15434 1656
rect 15434 1486 15444 1656
rect 15392 1476 15444 1486
rect 15648 1862 15700 1876
rect 15648 1696 15658 1862
rect 15658 1696 15692 1862
rect 15692 1696 15700 1862
rect 16416 1862 16468 1876
rect 16416 1696 16426 1862
rect 16426 1696 16460 1862
rect 16460 1696 16468 1862
rect 15908 1486 15916 1656
rect 15916 1486 15950 1656
rect 15950 1486 15960 1656
rect 15908 1476 15960 1486
rect 16676 1486 16684 1656
rect 16684 1486 16718 1656
rect 16718 1486 16728 1656
rect 16676 1476 16728 1486
rect 16932 1862 16984 1876
rect 16932 1696 16942 1862
rect 16942 1696 16976 1862
rect 16976 1696 16984 1862
rect 17192 1486 17200 1656
rect 17200 1486 17234 1656
rect 17234 1486 17244 1656
rect 17192 1476 17244 1486
rect 17448 1862 17500 1876
rect 17448 1696 17458 1862
rect 17458 1696 17492 1862
rect 17492 1696 17500 1862
rect 18216 1862 18268 1876
rect 18216 1696 18226 1862
rect 18226 1696 18260 1862
rect 18260 1696 18268 1862
rect 17708 1486 17716 1656
rect 17716 1486 17750 1656
rect 17750 1486 17760 1656
rect 17708 1476 17760 1486
rect 18476 1486 18484 1656
rect 18484 1486 18518 1656
rect 18518 1486 18528 1656
rect 18476 1476 18528 1486
rect 18732 1862 18784 1876
rect 18732 1696 18742 1862
rect 18742 1696 18776 1862
rect 18776 1696 18784 1862
rect 18992 1486 19000 1656
rect 19000 1486 19034 1656
rect 19034 1486 19044 1656
rect 18992 1476 19044 1486
rect 19248 1862 19300 1876
rect 19248 1696 19258 1862
rect 19258 1696 19292 1862
rect 19292 1696 19300 1862
rect 20016 1862 20068 1876
rect 20016 1696 20026 1862
rect 20026 1696 20060 1862
rect 20060 1696 20068 1862
rect 19508 1486 19516 1656
rect 19516 1486 19550 1656
rect 19550 1486 19560 1656
rect 19508 1476 19560 1486
rect 20276 1486 20284 1656
rect 20284 1486 20318 1656
rect 20318 1486 20328 1656
rect 20276 1476 20328 1486
rect 20532 1862 20584 1876
rect 20532 1696 20542 1862
rect 20542 1696 20576 1862
rect 20576 1696 20584 1862
rect 20792 1486 20800 1656
rect 20800 1486 20834 1656
rect 20834 1486 20844 1656
rect 20792 1476 20844 1486
rect 21048 1862 21100 1876
rect 21048 1696 21058 1862
rect 21058 1696 21092 1862
rect 21092 1696 21100 1862
rect 21308 1486 21316 1656
rect 21316 1486 21350 1656
rect 21350 1486 21360 1656
rect 21308 1476 21360 1486
rect -8768 1148 -8760 1316
rect -8760 1148 -8726 1316
rect -8726 1148 -8716 1316
rect -8768 1136 -8716 1148
rect 216 1244 268 1256
rect 216 1076 226 1244
rect 226 1076 260 1244
rect 260 1076 268 1244
rect -10060 906 -10008 920
rect -10060 740 -10050 906
rect -10050 740 -10016 906
rect -10016 740 -10008 906
rect -9800 530 -9792 700
rect -9792 530 -9758 700
rect -9758 530 -9748 700
rect -9800 520 -9748 530
rect -9544 906 -9492 920
rect -9544 740 -9534 906
rect -9534 740 -9500 906
rect -9500 740 -9492 906
rect -9284 530 -9276 700
rect -9276 530 -9242 700
rect -9242 530 -9232 700
rect -9284 520 -9232 530
rect -9028 906 -8976 920
rect -9028 740 -9018 906
rect -9018 740 -8984 906
rect -8984 740 -8976 906
rect 476 868 484 1036
rect 484 868 518 1036
rect 518 868 528 1036
rect 476 856 528 868
rect 732 1244 784 1256
rect 732 1076 742 1244
rect 742 1076 776 1244
rect 776 1076 784 1244
rect 992 868 1000 1036
rect 1000 868 1034 1036
rect 1034 868 1044 1036
rect 992 856 1044 868
rect 1248 1244 1300 1256
rect 1248 1076 1258 1244
rect 1258 1076 1292 1244
rect 1292 1076 1300 1244
rect 2016 1244 2068 1256
rect 2016 1076 2026 1244
rect 2026 1076 2060 1244
rect 2060 1076 2068 1244
rect 1508 868 1516 1036
rect 1516 868 1550 1036
rect 1550 868 1560 1036
rect 1508 856 1560 868
rect 2276 868 2284 1036
rect 2284 868 2318 1036
rect 2318 868 2328 1036
rect 2276 856 2328 868
rect 2532 1244 2584 1256
rect 2532 1076 2542 1244
rect 2542 1076 2576 1244
rect 2576 1076 2584 1244
rect 2792 868 2800 1036
rect 2800 868 2834 1036
rect 2834 868 2844 1036
rect 2792 856 2844 868
rect 3048 1244 3100 1256
rect 3048 1076 3058 1244
rect 3058 1076 3092 1244
rect 3092 1076 3100 1244
rect 3816 1244 3868 1256
rect 3816 1076 3826 1244
rect 3826 1076 3860 1244
rect 3860 1076 3868 1244
rect 3308 868 3316 1036
rect 3316 868 3350 1036
rect 3350 868 3360 1036
rect 3308 856 3360 868
rect 4076 868 4084 1036
rect 4084 868 4118 1036
rect 4118 868 4128 1036
rect 4076 856 4128 868
rect 4332 1244 4384 1256
rect 4332 1076 4342 1244
rect 4342 1076 4376 1244
rect 4376 1076 4384 1244
rect 4592 868 4600 1036
rect 4600 868 4634 1036
rect 4634 868 4644 1036
rect 4592 856 4644 868
rect 4848 1244 4900 1256
rect 4848 1076 4858 1244
rect 4858 1076 4892 1244
rect 4892 1076 4900 1244
rect 5616 1244 5668 1256
rect 5616 1076 5626 1244
rect 5626 1076 5660 1244
rect 5660 1076 5668 1244
rect 5108 868 5116 1036
rect 5116 868 5150 1036
rect 5150 868 5160 1036
rect 5108 856 5160 868
rect 5876 868 5884 1036
rect 5884 868 5918 1036
rect 5918 868 5928 1036
rect 5876 856 5928 868
rect 6132 1244 6184 1256
rect 6132 1076 6142 1244
rect 6142 1076 6176 1244
rect 6176 1076 6184 1244
rect 6392 868 6400 1036
rect 6400 868 6434 1036
rect 6434 868 6444 1036
rect 6392 856 6444 868
rect 6648 1244 6700 1256
rect 6648 1076 6658 1244
rect 6658 1076 6692 1244
rect 6692 1076 6700 1244
rect 14616 1244 14668 1256
rect 14616 1076 14626 1244
rect 14626 1076 14660 1244
rect 14660 1076 14668 1244
rect 6908 868 6916 1036
rect 6916 868 6950 1036
rect 6950 868 6960 1036
rect 6908 856 6960 868
rect 14876 868 14884 1036
rect 14884 868 14918 1036
rect 14918 868 14928 1036
rect 14876 856 14928 868
rect 15132 1244 15184 1256
rect 15132 1076 15142 1244
rect 15142 1076 15176 1244
rect 15176 1076 15184 1244
rect 15392 868 15400 1036
rect 15400 868 15434 1036
rect 15434 868 15444 1036
rect 15392 856 15444 868
rect 15648 1244 15700 1256
rect 15648 1076 15658 1244
rect 15658 1076 15692 1244
rect 15692 1076 15700 1244
rect 16416 1244 16468 1256
rect 16416 1076 16426 1244
rect 16426 1076 16460 1244
rect 16460 1076 16468 1244
rect 15908 868 15916 1036
rect 15916 868 15950 1036
rect 15950 868 15960 1036
rect 15908 856 15960 868
rect 16676 868 16684 1036
rect 16684 868 16718 1036
rect 16718 868 16728 1036
rect 16676 856 16728 868
rect 16932 1244 16984 1256
rect 16932 1076 16942 1244
rect 16942 1076 16976 1244
rect 16976 1076 16984 1244
rect 17192 868 17200 1036
rect 17200 868 17234 1036
rect 17234 868 17244 1036
rect 17192 856 17244 868
rect 17448 1244 17500 1256
rect 17448 1076 17458 1244
rect 17458 1076 17492 1244
rect 17492 1076 17500 1244
rect 18216 1244 18268 1256
rect 18216 1076 18226 1244
rect 18226 1076 18260 1244
rect 18260 1076 18268 1244
rect 17708 868 17716 1036
rect 17716 868 17750 1036
rect 17750 868 17760 1036
rect 17708 856 17760 868
rect 18476 868 18484 1036
rect 18484 868 18518 1036
rect 18518 868 18528 1036
rect 18476 856 18528 868
rect 18732 1244 18784 1256
rect 18732 1076 18742 1244
rect 18742 1076 18776 1244
rect 18776 1076 18784 1244
rect 18992 868 19000 1036
rect 19000 868 19034 1036
rect 19034 868 19044 1036
rect 18992 856 19044 868
rect 19248 1244 19300 1256
rect 19248 1076 19258 1244
rect 19258 1076 19292 1244
rect 19292 1076 19300 1244
rect 20016 1244 20068 1256
rect 20016 1076 20026 1244
rect 20026 1076 20060 1244
rect 20060 1076 20068 1244
rect 19508 868 19516 1036
rect 19516 868 19550 1036
rect 19550 868 19560 1036
rect 19508 856 19560 868
rect 20276 868 20284 1036
rect 20284 868 20318 1036
rect 20318 868 20328 1036
rect 20276 856 20328 868
rect 20532 1244 20584 1256
rect 20532 1076 20542 1244
rect 20542 1076 20576 1244
rect 20576 1076 20584 1244
rect 20792 868 20800 1036
rect 20800 868 20834 1036
rect 20834 868 20844 1036
rect 20792 856 20844 868
rect 21048 1244 21100 1256
rect 21048 1076 21058 1244
rect 21058 1076 21092 1244
rect 21092 1076 21100 1244
rect 21308 868 21316 1036
rect 21316 868 21350 1036
rect 21350 868 21360 1036
rect 21308 856 21360 868
rect -8768 530 -8760 700
rect -8760 530 -8726 700
rect -8726 530 -8716 700
rect -8768 520 -8716 530
rect -8500 348 -8360 508
rect 216 626 268 640
rect 216 460 226 626
rect 226 460 260 626
rect 260 460 268 626
rect 476 250 484 420
rect 484 250 518 420
rect 518 250 528 420
rect 476 240 528 250
rect 732 626 784 640
rect 732 460 742 626
rect 742 460 776 626
rect 776 460 784 626
rect 992 250 1000 420
rect 1000 250 1034 420
rect 1034 250 1044 420
rect 992 240 1044 250
rect 1248 626 1300 640
rect 1248 460 1258 626
rect 1258 460 1292 626
rect 1292 460 1300 626
rect 2016 626 2068 640
rect 2016 460 2026 626
rect 2026 460 2060 626
rect 2060 460 2068 626
rect 1508 250 1516 420
rect 1516 250 1550 420
rect 1550 250 1560 420
rect 1508 240 1560 250
rect 1696 68 1876 268
rect 2276 250 2284 420
rect 2284 250 2318 420
rect 2318 250 2328 420
rect 2276 240 2328 250
rect 2532 626 2584 640
rect 2532 460 2542 626
rect 2542 460 2576 626
rect 2576 460 2584 626
rect 2792 250 2800 420
rect 2800 250 2834 420
rect 2834 250 2844 420
rect 2792 240 2844 250
rect 3048 626 3100 640
rect 3048 460 3058 626
rect 3058 460 3092 626
rect 3092 460 3100 626
rect 3816 626 3868 640
rect 3816 460 3826 626
rect 3826 460 3860 626
rect 3860 460 3868 626
rect 3308 250 3316 420
rect 3316 250 3350 420
rect 3350 250 3360 420
rect 3308 240 3360 250
rect 3512 64 3692 276
rect 4076 250 4084 420
rect 4084 250 4118 420
rect 4118 250 4128 420
rect 4076 240 4128 250
rect 4332 626 4384 640
rect 4332 460 4342 626
rect 4342 460 4376 626
rect 4376 460 4384 626
rect 4592 250 4600 420
rect 4600 250 4634 420
rect 4634 250 4644 420
rect 4592 240 4644 250
rect 4848 626 4900 640
rect 4848 460 4858 626
rect 4858 460 4892 626
rect 4892 460 4900 626
rect 5616 626 5668 640
rect 5616 460 5626 626
rect 5626 460 5660 626
rect 5660 460 5668 626
rect 5108 250 5116 420
rect 5116 250 5150 420
rect 5150 250 5160 420
rect 5108 240 5160 250
rect 5288 64 5468 276
rect 5876 250 5884 420
rect 5884 250 5918 420
rect 5918 250 5928 420
rect 5876 240 5928 250
rect 6132 626 6184 640
rect 6132 460 6142 626
rect 6142 460 6176 626
rect 6176 460 6184 626
rect 6392 250 6400 420
rect 6400 250 6434 420
rect 6434 250 6444 420
rect 6392 240 6444 250
rect 6648 626 6700 640
rect 6648 460 6658 626
rect 6658 460 6692 626
rect 6692 460 6700 626
rect 14616 626 14668 640
rect 14616 460 14626 626
rect 14626 460 14660 626
rect 14660 460 14668 626
rect 6908 250 6916 420
rect 6916 250 6950 420
rect 6950 250 6960 420
rect 6908 240 6960 250
rect 14876 250 14884 420
rect 14884 250 14918 420
rect 14918 250 14928 420
rect 14876 240 14928 250
rect 15132 626 15184 640
rect 15132 460 15142 626
rect 15142 460 15176 626
rect 15176 460 15184 626
rect 15392 250 15400 420
rect 15400 250 15434 420
rect 15434 250 15444 420
rect 15392 240 15444 250
rect 15648 626 15700 640
rect 15648 460 15658 626
rect 15658 460 15692 626
rect 15692 460 15700 626
rect 16416 626 16468 640
rect 16416 460 16426 626
rect 16426 460 16460 626
rect 16460 460 16468 626
rect 15908 250 15916 420
rect 15916 250 15950 420
rect 15950 250 15960 420
rect 15908 240 15960 250
rect 16096 68 16276 268
rect 16676 250 16684 420
rect 16684 250 16718 420
rect 16718 250 16728 420
rect 16676 240 16728 250
rect 16932 626 16984 640
rect 16932 460 16942 626
rect 16942 460 16976 626
rect 16976 460 16984 626
rect 17192 250 17200 420
rect 17200 250 17234 420
rect 17234 250 17244 420
rect 17192 240 17244 250
rect 17448 626 17500 640
rect 17448 460 17458 626
rect 17458 460 17492 626
rect 17492 460 17500 626
rect 18216 626 18268 640
rect 18216 460 18226 626
rect 18226 460 18260 626
rect 18260 460 18268 626
rect 17708 250 17716 420
rect 17716 250 17750 420
rect 17750 250 17760 420
rect 17708 240 17760 250
rect 17912 64 18092 276
rect 18476 250 18484 420
rect 18484 250 18518 420
rect 18518 250 18528 420
rect 18476 240 18528 250
rect 18732 626 18784 640
rect 18732 460 18742 626
rect 18742 460 18776 626
rect 18776 460 18784 626
rect 18992 250 19000 420
rect 19000 250 19034 420
rect 19034 250 19044 420
rect 18992 240 19044 250
rect 19248 626 19300 640
rect 19248 460 19258 626
rect 19258 460 19292 626
rect 19292 460 19300 626
rect 20016 626 20068 640
rect 20016 460 20026 626
rect 20026 460 20060 626
rect 20060 460 20068 626
rect 19508 250 19516 420
rect 19516 250 19550 420
rect 19550 250 19560 420
rect 19508 240 19560 250
rect 19688 64 19868 276
rect 20276 250 20284 420
rect 20284 250 20318 420
rect 20318 250 20328 420
rect 20276 240 20328 250
rect 20532 626 20584 640
rect 20532 460 20542 626
rect 20542 460 20576 626
rect 20576 460 20584 626
rect 20792 250 20800 420
rect 20800 250 20834 420
rect 20834 250 20844 420
rect 20792 240 20844 250
rect 21048 626 21100 640
rect 21048 460 21058 626
rect 21058 460 21092 626
rect 21092 460 21100 626
rect 21308 250 21316 420
rect 21316 250 21350 420
rect 21350 250 21360 420
rect 21308 240 21360 250
rect -2768 -1188 -1960 -382
rect 11632 -1188 12440 -382
<< metal2 >>
rect 7440 27436 7540 27446
rect 7440 27326 7540 27336
rect 6632 27182 7960 27184
rect 8852 27182 10180 27184
rect 11032 27182 12360 27184
rect 13212 27182 14540 27184
rect 15412 27182 16740 27184
rect 6632 27172 8240 27182
rect 6632 27092 7384 27172
rect 6696 26916 6948 27092
rect 6632 26902 6696 26912
rect 7012 26916 7264 27092
rect 6948 26902 7012 26912
rect 7328 26928 7384 27092
rect 7328 26916 7580 26928
rect 7264 26902 7328 26912
rect 7644 26916 7896 26928
rect 7580 26902 7644 26912
rect 7960 26918 8240 26928
rect 8852 27172 10460 27182
rect 8852 27092 9604 27172
rect 7896 26902 7960 26912
rect 8916 26916 9168 27092
rect 8852 26902 8916 26912
rect 9232 26916 9484 27092
rect 9168 26902 9232 26912
rect 9548 26928 9604 27092
rect 9548 26916 9800 26928
rect 9484 26902 9548 26912
rect 9864 26916 10116 26928
rect 9800 26902 9864 26912
rect 10180 26918 10460 26928
rect 11032 27172 12640 27182
rect 11032 27092 11784 27172
rect 10116 26902 10180 26912
rect 11096 26916 11348 27092
rect 11032 26902 11096 26912
rect 11412 26916 11664 27092
rect 11348 26902 11412 26912
rect 11728 26928 11784 27092
rect 11728 26916 11980 26928
rect 11664 26902 11728 26912
rect 12044 26916 12296 26928
rect 11980 26902 12044 26912
rect 12360 26918 12640 26928
rect 13212 27172 14820 27182
rect 13212 27092 13964 27172
rect 12296 26902 12360 26912
rect 13276 26916 13528 27092
rect 13212 26902 13276 26912
rect 13592 26916 13844 27092
rect 13528 26902 13592 26912
rect 13908 26928 13964 27092
rect 13908 26916 14160 26928
rect 13844 26902 13908 26912
rect 14224 26916 14476 26928
rect 14160 26902 14224 26912
rect 14540 26918 14820 26928
rect 15412 27172 17020 27182
rect 15412 27092 16164 27172
rect 14476 26902 14540 26912
rect 15476 26916 15728 27092
rect 15412 26902 15476 26912
rect 15792 26916 16044 27092
rect 15728 26902 15792 26912
rect 16108 26928 16164 27092
rect 16108 26916 16360 26928
rect 16044 26902 16108 26912
rect 16424 26916 16676 26928
rect 16360 26902 16424 26912
rect 16740 26918 17020 26928
rect 16676 26902 16740 26912
rect 6476 26868 6540 26878
rect 6792 26868 6856 26878
rect 6540 26852 6792 26862
rect 7108 26868 7172 26878
rect 6856 26852 7108 26862
rect 7424 26868 7488 26878
rect 7172 26860 7268 26862
rect 7172 26852 7424 26860
rect 7268 26688 7424 26852
rect 7740 26868 7804 26878
rect 7488 26688 7740 26860
rect 8056 26868 8120 26878
rect 7804 26688 8056 26860
rect 6476 26608 6488 26688
rect 7268 26608 8120 26688
rect 6476 26592 8120 26608
rect 8696 26868 8760 26878
rect 9012 26868 9076 26878
rect 8760 26852 9012 26862
rect 9328 26868 9392 26878
rect 9076 26852 9328 26862
rect 9644 26868 9708 26878
rect 9392 26860 9488 26862
rect 9392 26852 9644 26860
rect 9488 26688 9644 26852
rect 9960 26868 10024 26878
rect 9708 26688 9960 26860
rect 10276 26868 10340 26878
rect 10024 26688 10276 26860
rect 8696 26608 8708 26688
rect 9488 26608 10340 26688
rect 8696 26592 10340 26608
rect 10876 26868 10940 26878
rect 11192 26868 11256 26878
rect 10940 26852 11192 26862
rect 11508 26868 11572 26878
rect 11256 26852 11508 26862
rect 11824 26868 11888 26878
rect 11572 26860 11668 26862
rect 11572 26852 11824 26860
rect 11668 26688 11824 26852
rect 12140 26868 12204 26878
rect 11888 26688 12140 26860
rect 12456 26868 12520 26878
rect 12204 26688 12456 26860
rect 10876 26608 10888 26688
rect 11668 26608 12520 26688
rect 10876 26592 12520 26608
rect 13056 26868 13120 26878
rect 13372 26868 13436 26878
rect 13120 26852 13372 26862
rect 13688 26868 13752 26878
rect 13436 26852 13688 26862
rect 14004 26868 14068 26878
rect 13752 26860 13848 26862
rect 13752 26852 14004 26860
rect 13848 26688 14004 26852
rect 14320 26868 14384 26878
rect 14068 26688 14320 26860
rect 14636 26868 14700 26878
rect 14384 26688 14636 26860
rect 13056 26608 13068 26688
rect 13848 26608 14700 26688
rect 13056 26592 14700 26608
rect 15256 26868 15320 26878
rect 15572 26868 15636 26878
rect 15320 26852 15572 26862
rect 15888 26868 15952 26878
rect 15636 26852 15888 26862
rect 16204 26868 16268 26878
rect 15952 26860 16048 26862
rect 15952 26852 16204 26860
rect 16048 26688 16204 26852
rect 16520 26868 16584 26878
rect 16268 26688 16520 26860
rect 16836 26868 16900 26878
rect 16584 26688 16836 26860
rect 15256 26608 15268 26688
rect 16048 26608 16900 26688
rect 15256 26592 16900 26608
rect 7384 26548 8240 26550
rect 9604 26548 10460 26550
rect 11784 26548 12640 26550
rect 13964 26548 14820 26550
rect 16164 26548 17020 26550
rect 6632 26540 8240 26548
rect 6632 26456 7384 26540
rect 6696 26280 6948 26456
rect 6632 26266 6696 26276
rect 7012 26280 7264 26456
rect 6948 26266 7012 26276
rect 7328 26296 7384 26456
rect 7328 26280 7580 26296
rect 7264 26266 7328 26276
rect 7644 26280 7896 26296
rect 7580 26266 7644 26276
rect 7960 26286 8240 26296
rect 8852 26540 10460 26548
rect 8852 26456 9604 26540
rect 7896 26266 7960 26276
rect 8916 26280 9168 26456
rect 8852 26266 8916 26276
rect 9232 26280 9484 26456
rect 9168 26266 9232 26276
rect 9548 26296 9604 26456
rect 9548 26280 9800 26296
rect 9484 26266 9548 26276
rect 9864 26280 10116 26296
rect 9800 26266 9864 26276
rect 10180 26286 10460 26296
rect 11032 26540 12640 26548
rect 11032 26456 11784 26540
rect 10116 26266 10180 26276
rect 11096 26280 11348 26456
rect 11032 26266 11096 26276
rect 11412 26280 11664 26456
rect 11348 26266 11412 26276
rect 11728 26296 11784 26456
rect 11728 26280 11980 26296
rect 11664 26266 11728 26276
rect 12044 26280 12296 26296
rect 11980 26266 12044 26276
rect 12360 26286 12640 26296
rect 13212 26540 14820 26548
rect 13212 26456 13964 26540
rect 12296 26266 12360 26276
rect 13276 26280 13528 26456
rect 13212 26266 13276 26276
rect 13592 26280 13844 26456
rect 13528 26266 13592 26276
rect 13908 26296 13964 26456
rect 13908 26280 14160 26296
rect 13844 26266 13908 26276
rect 14224 26280 14476 26296
rect 14160 26266 14224 26276
rect 14540 26286 14820 26296
rect 15412 26540 17020 26548
rect 15412 26456 16164 26540
rect 14476 26266 14540 26276
rect 15476 26280 15728 26456
rect 15412 26266 15476 26276
rect 15792 26280 16044 26456
rect 15728 26266 15792 26276
rect 16108 26296 16164 26456
rect 16108 26280 16360 26296
rect 16044 26266 16108 26276
rect 16424 26280 16676 26296
rect 16360 26266 16424 26276
rect 16740 26286 17020 26296
rect 16676 26266 16740 26276
rect 6476 26232 6540 26242
rect 6792 26232 6856 26242
rect 6540 26216 6792 26226
rect 7108 26232 7172 26242
rect 6856 26216 7108 26226
rect 7424 26232 7488 26242
rect 7172 26224 7268 26226
rect 7172 26216 7424 26224
rect 7268 26052 7424 26216
rect 7740 26232 7804 26242
rect 7488 26052 7740 26224
rect 8056 26232 8120 26242
rect 7804 26052 8056 26224
rect 6476 25972 6488 26052
rect 7268 25972 8120 26052
rect 6476 25956 8120 25972
rect 8696 26232 8760 26242
rect 9012 26232 9076 26242
rect 8760 26216 9012 26226
rect 9328 26232 9392 26242
rect 9076 26216 9328 26226
rect 9644 26232 9708 26242
rect 9392 26224 9488 26226
rect 9392 26216 9644 26224
rect 9488 26052 9644 26216
rect 9960 26232 10024 26242
rect 9708 26052 9960 26224
rect 10276 26232 10340 26242
rect 10024 26052 10276 26224
rect 8696 25972 8708 26052
rect 9488 25972 10340 26052
rect 8696 25956 10340 25972
rect 10876 26232 10940 26242
rect 11192 26232 11256 26242
rect 10940 26216 11192 26226
rect 11508 26232 11572 26242
rect 11256 26216 11508 26226
rect 11824 26232 11888 26242
rect 11572 26224 11668 26226
rect 11572 26216 11824 26224
rect 11668 26052 11824 26216
rect 12140 26232 12204 26242
rect 11888 26052 12140 26224
rect 12456 26232 12520 26242
rect 12204 26052 12456 26224
rect 10876 25972 10888 26052
rect 11668 25972 12520 26052
rect 10876 25956 12520 25972
rect 13056 26232 13120 26242
rect 13372 26232 13436 26242
rect 13120 26216 13372 26226
rect 13688 26232 13752 26242
rect 13436 26216 13688 26226
rect 14004 26232 14068 26242
rect 13752 26224 13848 26226
rect 13752 26216 14004 26224
rect 13848 26052 14004 26216
rect 14320 26232 14384 26242
rect 14068 26052 14320 26224
rect 14636 26232 14700 26242
rect 14384 26052 14636 26224
rect 13056 25972 13068 26052
rect 13848 25972 14700 26052
rect 13056 25956 14700 25972
rect 15256 26232 15320 26242
rect 15572 26232 15636 26242
rect 15320 26216 15572 26226
rect 15888 26232 15952 26242
rect 15636 26216 15888 26226
rect 16204 26232 16268 26242
rect 15952 26224 16048 26226
rect 15952 26216 16204 26224
rect 16048 26052 16204 26216
rect 16520 26232 16584 26242
rect 16268 26052 16520 26224
rect 16836 26232 16900 26242
rect 16584 26052 16836 26224
rect 15256 25972 15268 26052
rect 16048 25972 16900 26052
rect 15256 25956 16900 25972
rect 7384 25908 8240 25914
rect 9604 25908 10460 25914
rect 11784 25908 12640 25914
rect 13964 25908 14820 25914
rect 16164 25908 17020 25914
rect 6632 25904 8240 25908
rect 6632 25816 7384 25904
rect 6696 25640 6948 25816
rect 6632 25626 6696 25636
rect 7012 25640 7264 25816
rect 6948 25626 7012 25636
rect 7328 25660 7384 25816
rect 7328 25640 7580 25660
rect 7264 25626 7328 25636
rect 7644 25640 7896 25660
rect 7580 25626 7644 25636
rect 7960 25650 8240 25660
rect 8852 25904 10460 25908
rect 8852 25816 9604 25904
rect 7896 25626 7960 25636
rect 8916 25640 9168 25816
rect 8852 25626 8916 25636
rect 9232 25640 9484 25816
rect 9168 25626 9232 25636
rect 9548 25660 9604 25816
rect 9548 25640 9800 25660
rect 9484 25626 9548 25636
rect 9864 25640 10116 25660
rect 9800 25626 9864 25636
rect 10180 25650 10460 25660
rect 11032 25904 12640 25908
rect 11032 25816 11784 25904
rect 10116 25626 10180 25636
rect 11096 25640 11348 25816
rect 11032 25626 11096 25636
rect 11412 25640 11664 25816
rect 11348 25626 11412 25636
rect 11728 25660 11784 25816
rect 11728 25640 11980 25660
rect 11664 25626 11728 25636
rect 12044 25640 12296 25660
rect 11980 25626 12044 25636
rect 12360 25650 12640 25660
rect 13212 25904 14820 25908
rect 13212 25816 13964 25904
rect 12296 25626 12360 25636
rect 13276 25640 13528 25816
rect 13212 25626 13276 25636
rect 13592 25640 13844 25816
rect 13528 25626 13592 25636
rect 13908 25660 13964 25816
rect 13908 25640 14160 25660
rect 13844 25626 13908 25636
rect 14224 25640 14476 25660
rect 14160 25626 14224 25636
rect 14540 25650 14820 25660
rect 15412 25904 17020 25908
rect 15412 25816 16164 25904
rect 14476 25626 14540 25636
rect 15476 25640 15728 25816
rect 15412 25626 15476 25636
rect 15792 25640 16044 25816
rect 15728 25626 15792 25636
rect 16108 25660 16164 25816
rect 16108 25640 16360 25660
rect 16044 25626 16108 25636
rect 16424 25640 16676 25660
rect 16360 25626 16424 25636
rect 16740 25650 17020 25660
rect 16676 25626 16740 25636
rect 6476 25592 6540 25602
rect 6792 25592 6856 25602
rect 6540 25576 6792 25588
rect 7108 25592 7172 25602
rect 6856 25576 7108 25588
rect 7424 25592 7488 25602
rect 7172 25576 7424 25588
rect 7268 25412 7424 25576
rect 7740 25592 7804 25602
rect 7488 25412 7740 25588
rect 8056 25592 8120 25602
rect 7804 25412 8056 25588
rect 6476 25332 6488 25412
rect 7268 25332 8120 25412
rect 6476 25320 8120 25332
rect 8696 25592 8760 25602
rect 9012 25592 9076 25602
rect 8760 25576 9012 25588
rect 9328 25592 9392 25602
rect 9076 25576 9328 25588
rect 9644 25592 9708 25602
rect 9392 25576 9644 25588
rect 9488 25412 9644 25576
rect 9960 25592 10024 25602
rect 9708 25412 9960 25588
rect 10276 25592 10340 25602
rect 10024 25412 10276 25588
rect 8696 25332 8708 25412
rect 9488 25332 10340 25412
rect 8696 25320 10340 25332
rect 10876 25592 10940 25602
rect 11192 25592 11256 25602
rect 10940 25576 11192 25588
rect 11508 25592 11572 25602
rect 11256 25576 11508 25588
rect 11824 25592 11888 25602
rect 11572 25576 11824 25588
rect 11668 25412 11824 25576
rect 12140 25592 12204 25602
rect 11888 25412 12140 25588
rect 12456 25592 12520 25602
rect 12204 25412 12456 25588
rect 10876 25332 10888 25412
rect 11668 25332 12520 25412
rect 10876 25320 12520 25332
rect 13056 25592 13120 25602
rect 13372 25592 13436 25602
rect 13120 25576 13372 25588
rect 13688 25592 13752 25602
rect 13436 25576 13688 25588
rect 14004 25592 14068 25602
rect 13752 25576 14004 25588
rect 13848 25412 14004 25576
rect 14320 25592 14384 25602
rect 14068 25412 14320 25588
rect 14636 25592 14700 25602
rect 14384 25412 14636 25588
rect 13056 25332 13068 25412
rect 13848 25332 14700 25412
rect 13056 25320 14700 25332
rect 15256 25592 15320 25602
rect 15572 25592 15636 25602
rect 15320 25576 15572 25588
rect 15888 25592 15952 25602
rect 15636 25576 15888 25588
rect 16204 25592 16268 25602
rect 15952 25576 16204 25588
rect 16048 25412 16204 25576
rect 16520 25592 16584 25602
rect 16268 25412 16520 25588
rect 16836 25592 16900 25602
rect 16584 25412 16836 25588
rect 15256 25332 15268 25412
rect 16048 25332 16900 25412
rect 15256 25320 16900 25332
rect 18940 25260 19360 25280
rect 6492 25084 7276 25086
rect 8712 25084 9496 25086
rect 10100 25084 16760 25140
rect 6492 25076 7980 25084
rect 7276 24992 7980 25076
rect 7276 24828 7340 24992
rect 6492 24818 6572 24828
rect 6636 24816 6764 24828
rect 6572 24802 6636 24812
rect 6828 24816 6956 24828
rect 6764 24802 6828 24812
rect 7020 24816 7148 24828
rect 6956 24802 7020 24812
rect 7212 24816 7340 24828
rect 7148 24802 7212 24812
rect 7404 24816 7532 24992
rect 7340 24802 7404 24812
rect 7596 24816 7724 24992
rect 7532 24802 7596 24812
rect 7788 24816 7916 24992
rect 7724 24802 7788 24812
rect 8712 25076 16760 25084
rect 9496 24992 10892 25076
rect 11676 24992 13072 25076
rect 13856 24992 15272 25076
rect 16056 24992 16760 25076
rect 9496 24828 9560 24992
rect 8712 24818 8792 24828
rect 7916 24802 7980 24812
rect 8856 24816 8984 24828
rect 8792 24802 8856 24812
rect 9048 24816 9176 24828
rect 8984 24802 9048 24812
rect 9240 24816 9368 24828
rect 9176 24802 9240 24812
rect 9432 24816 9560 24828
rect 9368 24802 9432 24812
rect 9624 24816 9752 24992
rect 9560 24802 9624 24812
rect 9816 24816 9944 24992
rect 9752 24802 9816 24812
rect 10008 24816 10136 24992
rect 9944 24802 10008 24812
rect 10200 24828 10892 24992
rect 11676 24828 11740 24992
rect 10200 24816 10972 24828
rect 10136 24802 10200 24812
rect 11036 24816 11164 24828
rect 10972 24802 11036 24812
rect 11228 24816 11356 24828
rect 11164 24802 11228 24812
rect 11420 24816 11548 24828
rect 11356 24802 11420 24812
rect 11612 24816 11740 24828
rect 11548 24802 11612 24812
rect 11804 24816 11932 24992
rect 11740 24802 11804 24812
rect 11996 24816 12124 24992
rect 11932 24802 11996 24812
rect 12188 24816 12316 24992
rect 12124 24802 12188 24812
rect 12380 24828 13072 24992
rect 13856 24828 13920 24992
rect 12380 24816 13152 24828
rect 12316 24802 12380 24812
rect 13216 24816 13344 24828
rect 13152 24802 13216 24812
rect 13408 24816 13536 24828
rect 13344 24802 13408 24812
rect 13600 24816 13728 24828
rect 13536 24802 13600 24812
rect 13792 24816 13920 24828
rect 13728 24802 13792 24812
rect 13984 24816 14112 24992
rect 13920 24802 13984 24812
rect 14176 24816 14304 24992
rect 14112 24802 14176 24812
rect 14368 24816 14496 24992
rect 14304 24802 14368 24812
rect 14560 24828 15272 24992
rect 16056 24828 16120 24992
rect 14560 24816 15352 24828
rect 14496 24802 14560 24812
rect 15416 24816 15544 24828
rect 15352 24802 15416 24812
rect 15608 24816 15736 24828
rect 15544 24802 15608 24812
rect 15800 24816 15928 24828
rect 15736 24802 15800 24812
rect 15992 24816 16120 24828
rect 15928 24802 15992 24812
rect 16184 24816 16312 24992
rect 16120 24802 16184 24812
rect 16376 24816 16504 24992
rect 16312 24802 16376 24812
rect 16568 24816 16696 24992
rect 16504 24802 16568 24812
rect 16696 24802 16760 24812
rect 18280 25120 18640 25130
rect 6476 24768 6540 24778
rect 6664 24768 6728 24778
rect 6540 24588 6664 24764
rect 6856 24768 6920 24778
rect 6728 24588 6856 24764
rect 7052 24768 7116 24778
rect 6920 24588 7052 24764
rect 7244 24768 7308 24778
rect 7116 24588 7244 24764
rect 7436 24768 7500 24778
rect 7308 24748 7436 24764
rect 7628 24768 7692 24778
rect 7500 24748 7628 24764
rect 7820 24768 7884 24778
rect 7692 24748 7820 24764
rect 8696 24768 8760 24778
rect 7884 24748 8240 24758
rect 7308 24588 7388 24748
rect 6476 24508 7388 24588
rect 6476 24498 8240 24508
rect 8884 24768 8948 24778
rect 8760 24588 8884 24764
rect 9076 24768 9140 24778
rect 8948 24588 9076 24764
rect 9272 24768 9336 24778
rect 9140 24588 9272 24764
rect 9464 24768 9528 24778
rect 9336 24588 9464 24764
rect 9656 24768 9720 24778
rect 9528 24748 9656 24764
rect 9848 24768 9912 24778
rect 9720 24748 9848 24764
rect 10040 24768 10104 24778
rect 9912 24748 10040 24764
rect 10876 24768 10940 24778
rect 10104 24748 10460 24758
rect 9528 24588 9608 24748
rect 8696 24508 9608 24588
rect 8696 24498 10460 24508
rect 11064 24768 11128 24778
rect 10940 24588 11064 24764
rect 11256 24768 11320 24778
rect 11128 24588 11256 24764
rect 11452 24768 11516 24778
rect 11320 24588 11452 24764
rect 11644 24768 11708 24778
rect 11516 24588 11644 24764
rect 11836 24768 11900 24778
rect 11708 24748 11836 24764
rect 12028 24768 12092 24778
rect 11900 24748 12028 24764
rect 12220 24768 12284 24778
rect 12092 24748 12220 24764
rect 13056 24768 13120 24778
rect 12284 24748 12640 24758
rect 11708 24588 11788 24748
rect 10876 24508 11788 24588
rect 10876 24498 12640 24508
rect 13244 24768 13308 24778
rect 13120 24588 13244 24764
rect 13436 24768 13500 24778
rect 13308 24588 13436 24764
rect 13632 24768 13696 24778
rect 13500 24588 13632 24764
rect 13824 24768 13888 24778
rect 13696 24588 13824 24764
rect 14016 24768 14080 24778
rect 13888 24748 14016 24764
rect 14208 24768 14272 24778
rect 14080 24748 14208 24764
rect 14400 24768 14464 24778
rect 14272 24748 14400 24764
rect 15256 24768 15320 24778
rect 14464 24748 14820 24758
rect 13888 24588 13968 24748
rect 13056 24508 13968 24588
rect 13056 24498 14820 24508
rect 15444 24768 15508 24778
rect 15320 24588 15444 24764
rect 15636 24768 15700 24778
rect 15508 24588 15636 24764
rect 15832 24768 15896 24778
rect 15700 24588 15832 24764
rect 16024 24768 16088 24778
rect 15896 24588 16024 24764
rect 16216 24768 16280 24778
rect 16088 24748 16216 24764
rect 16408 24768 16472 24778
rect 16280 24748 16408 24764
rect 16600 24768 16664 24778
rect 16472 24748 16600 24764
rect 16664 24748 17020 24758
rect 16088 24588 16168 24748
rect 18280 24590 18640 24600
rect 18940 25040 19040 25260
rect 19240 25040 19360 25260
rect 15256 24508 16168 24588
rect 15256 24498 17020 24508
rect 6476 24496 7884 24498
rect 8696 24496 10104 24498
rect 10876 24496 12284 24498
rect 13056 24496 14464 24498
rect 15256 24496 16664 24498
rect 6572 24446 7980 24448
rect 8792 24446 10200 24448
rect 10972 24446 12380 24448
rect 13152 24446 14560 24448
rect 15352 24446 16760 24448
rect 6492 24436 7980 24446
rect 7276 24356 7980 24436
rect 7276 24188 7340 24356
rect 6492 24178 6572 24188
rect 6636 24178 6764 24188
rect 6572 24166 6636 24176
rect 6828 24178 6956 24188
rect 6764 24166 6828 24176
rect 7020 24178 7148 24188
rect 6956 24166 7020 24176
rect 7212 24180 7340 24188
rect 7212 24178 7276 24180
rect 7148 24166 7212 24176
rect 7404 24180 7532 24356
rect 7340 24166 7404 24176
rect 7596 24180 7724 24356
rect 7532 24166 7596 24176
rect 7788 24180 7916 24356
rect 7724 24166 7788 24176
rect 8156 24436 8328 24446
rect 8156 24202 8328 24212
rect 8712 24436 10200 24446
rect 9496 24356 10200 24436
rect 9496 24188 9560 24356
rect 8712 24178 8792 24188
rect 7916 24166 7980 24176
rect 8856 24178 8984 24188
rect 8792 24166 8856 24176
rect 9048 24178 9176 24188
rect 8984 24166 9048 24176
rect 9240 24178 9368 24188
rect 9176 24166 9240 24176
rect 9432 24180 9560 24188
rect 9432 24178 9496 24180
rect 9368 24166 9432 24176
rect 9624 24180 9752 24356
rect 9560 24166 9624 24176
rect 9816 24180 9944 24356
rect 9752 24166 9816 24176
rect 10008 24180 10136 24356
rect 9944 24166 10008 24176
rect 10892 24436 12380 24446
rect 11676 24356 12380 24436
rect 11676 24188 11740 24356
rect 10892 24178 10972 24188
rect 10136 24166 10200 24176
rect 11036 24178 11164 24188
rect 10972 24166 11036 24176
rect 11228 24178 11356 24188
rect 11164 24166 11228 24176
rect 11420 24178 11548 24188
rect 11356 24166 11420 24176
rect 11612 24180 11740 24188
rect 11612 24178 11676 24180
rect 11548 24166 11612 24176
rect 11804 24180 11932 24356
rect 11740 24166 11804 24176
rect 11996 24180 12124 24356
rect 11932 24166 11996 24176
rect 12188 24180 12316 24356
rect 12124 24166 12188 24176
rect 13072 24436 14560 24446
rect 13856 24356 14560 24436
rect 13856 24188 13920 24356
rect 13072 24178 13152 24188
rect 12316 24166 12380 24176
rect 13216 24178 13344 24188
rect 13152 24166 13216 24176
rect 13408 24178 13536 24188
rect 13344 24166 13408 24176
rect 13600 24178 13728 24188
rect 13536 24166 13600 24176
rect 13792 24180 13920 24188
rect 13792 24178 13856 24180
rect 13728 24166 13792 24176
rect 13984 24180 14112 24356
rect 13920 24166 13984 24176
rect 14176 24180 14304 24356
rect 14112 24166 14176 24176
rect 14368 24180 14496 24356
rect 14304 24166 14368 24176
rect 15272 24436 16760 24446
rect 16056 24356 16760 24436
rect 18940 24420 19360 25040
rect 16056 24188 16120 24356
rect 15272 24178 15352 24188
rect 14496 24166 14560 24176
rect 15416 24178 15544 24188
rect 15352 24166 15416 24176
rect 15608 24178 15736 24188
rect 15544 24166 15608 24176
rect 15800 24178 15928 24188
rect 15736 24166 15800 24176
rect 15992 24180 16120 24188
rect 15992 24178 16056 24180
rect 15928 24166 15992 24176
rect 16184 24180 16312 24356
rect 16120 24166 16184 24176
rect 16376 24180 16504 24356
rect 16312 24166 16376 24176
rect 16568 24180 16696 24356
rect 16504 24166 16568 24176
rect 16696 24166 16760 24176
rect 6476 24132 6540 24142
rect 6664 24132 6728 24142
rect 6540 23952 6664 24128
rect 6856 24132 6920 24142
rect 6728 23952 6856 24128
rect 7052 24132 7116 24142
rect 6920 23952 7052 24128
rect 7244 24132 7308 24142
rect 7116 23952 7244 24128
rect 7436 24132 7500 24142
rect 7308 24116 7436 24128
rect 7628 24132 7692 24142
rect 7500 24116 7628 24128
rect 7820 24132 7884 24142
rect 7692 24116 7820 24128
rect 8696 24132 8760 24142
rect 7884 24116 8240 24126
rect 7308 23952 7388 24116
rect 6476 23876 7388 23952
rect 6476 23866 8240 23876
rect 8884 24132 8948 24142
rect 8760 23952 8884 24128
rect 9076 24132 9140 24142
rect 8948 23952 9076 24128
rect 9272 24132 9336 24142
rect 9140 23952 9272 24128
rect 9464 24132 9528 24142
rect 9336 23952 9464 24128
rect 9656 24132 9720 24142
rect 9528 24116 9656 24128
rect 9848 24132 9912 24142
rect 9720 24116 9848 24128
rect 10040 24132 10104 24142
rect 9912 24116 10040 24128
rect 10876 24132 10940 24142
rect 10104 24116 10460 24126
rect 9528 23952 9608 24116
rect 8696 23876 9608 23952
rect 8696 23866 10460 23876
rect 11064 24132 11128 24142
rect 10940 23952 11064 24128
rect 11256 24132 11320 24142
rect 11128 23952 11256 24128
rect 11452 24132 11516 24142
rect 11320 23952 11452 24128
rect 11644 24132 11708 24142
rect 11516 23952 11644 24128
rect 11836 24132 11900 24142
rect 11708 24116 11836 24128
rect 12028 24132 12092 24142
rect 11900 24116 12028 24128
rect 12220 24132 12284 24142
rect 12092 24116 12220 24128
rect 13056 24132 13120 24142
rect 12284 24116 12640 24126
rect 11708 23952 11788 24116
rect 10876 23876 11788 23952
rect 10876 23866 12640 23876
rect 13244 24132 13308 24142
rect 13120 23952 13244 24128
rect 13436 24132 13500 24142
rect 13308 23952 13436 24128
rect 13632 24132 13696 24142
rect 13500 23952 13632 24128
rect 13824 24132 13888 24142
rect 13696 23952 13824 24128
rect 14016 24132 14080 24142
rect 13888 24116 14016 24128
rect 14208 24132 14272 24142
rect 14080 24116 14208 24128
rect 14400 24132 14464 24142
rect 14272 24116 14400 24128
rect 15256 24132 15320 24142
rect 14464 24116 14820 24126
rect 13888 23952 13968 24116
rect 13056 23876 13968 23952
rect 13056 23866 14820 23876
rect 15444 24132 15508 24142
rect 15320 23952 15444 24128
rect 15636 24132 15700 24142
rect 15508 23952 15636 24128
rect 15832 24132 15896 24142
rect 15700 23952 15832 24128
rect 16024 24132 16088 24142
rect 15896 23952 16024 24128
rect 16216 24132 16280 24142
rect 16088 24116 16216 24128
rect 16408 24132 16472 24142
rect 16280 24116 16408 24128
rect 16600 24132 16664 24142
rect 16472 24116 16600 24128
rect 16664 24116 17020 24126
rect 16088 23952 16168 24116
rect 15256 23876 16168 23952
rect 15256 23866 17020 23876
rect 17480 24040 19360 24420
rect 6476 23860 7884 23866
rect 8696 23860 10104 23866
rect 10876 23860 12284 23866
rect 13056 23860 14464 23866
rect 15256 23860 16664 23866
rect 6688 23680 9676 23704
rect 6688 23424 7408 23680
rect 8236 23424 9676 23680
rect 6688 23244 6696 23424
rect 6748 23244 6888 23424
rect 6940 23244 7080 23424
rect 7132 23244 7272 23424
rect 7324 23272 7408 23424
rect 8236 23272 8416 23424
rect 7324 23244 7464 23272
rect 7516 23244 8416 23272
rect 8468 23244 8608 23424
rect 8660 23244 8800 23424
rect 8852 23244 8992 23424
rect 9044 23244 9184 23424
rect 9236 23244 9676 23424
rect 17480 23300 17840 24040
rect 18328 23852 18688 23862
rect 18688 23420 18700 23852
rect 18328 23410 18700 23420
rect 6696 23234 6748 23244
rect 6888 23234 6940 23244
rect 7080 23234 7132 23244
rect 7272 23234 7324 23244
rect 7464 23234 7516 23244
rect 6600 23202 6652 23210
rect 6792 23202 6844 23210
rect 6984 23202 7036 23210
rect 7176 23202 7228 23210
rect 6596 23200 7228 23202
rect 7368 23200 7420 23210
rect 7560 23200 7612 23210
rect 6596 23192 6600 23200
rect 6652 23192 6792 23200
rect 6844 23192 6984 23200
rect 7036 23192 7176 23200
rect 7228 23020 7368 23200
rect 7420 23020 7560 23200
rect 7200 23012 7612 23020
rect 7200 23010 7228 23012
rect 7368 23010 7420 23012
rect 7560 23010 7612 23012
rect 6596 22998 7200 23008
rect 6696 22816 7516 22820
rect 7644 22816 7956 23244
rect 8416 23234 8468 23244
rect 8608 23234 8660 23244
rect 8800 23234 8852 23244
rect 8992 23234 9044 23244
rect 9184 23234 9236 23244
rect 8320 23202 8372 23210
rect 8512 23202 8564 23210
rect 8704 23202 8756 23210
rect 8896 23202 8948 23210
rect 8316 23200 8948 23202
rect 9088 23200 9140 23210
rect 9280 23200 9332 23210
rect 8316 23192 8320 23200
rect 8372 23192 8512 23200
rect 8564 23192 8704 23200
rect 8756 23192 8896 23200
rect 8948 23020 9088 23200
rect 9140 23020 9280 23200
rect 8920 23012 9332 23020
rect 8920 23010 8948 23012
rect 9088 23010 9140 23012
rect 9280 23010 9332 23012
rect 8316 22998 8920 23008
rect 6696 22808 7956 22816
rect 6748 22628 6888 22808
rect 6940 22628 7080 22808
rect 7132 22628 7272 22808
rect 7324 22628 7464 22808
rect 7516 22628 7956 22808
rect 6696 22618 6748 22628
rect 6888 22618 6940 22628
rect 7080 22618 7132 22628
rect 7272 22618 7324 22628
rect 7464 22618 7516 22628
rect 6600 22586 6652 22594
rect 6792 22586 6844 22594
rect 6984 22586 7036 22594
rect 7176 22586 7228 22594
rect 6596 22584 7228 22586
rect 7368 22584 7420 22594
rect 7560 22584 7612 22594
rect 6596 22576 6600 22584
rect 6652 22576 6792 22584
rect 6844 22576 6984 22584
rect 7036 22576 7176 22584
rect 7228 22404 7368 22584
rect 7420 22404 7560 22584
rect 7200 22396 7612 22404
rect 7200 22394 7228 22396
rect 7368 22394 7420 22396
rect 7560 22394 7612 22396
rect 6596 22382 7200 22392
rect 6696 22192 6748 22198
rect 6888 22192 6940 22198
rect 7080 22192 7132 22198
rect 7272 22192 7324 22198
rect 7464 22192 7516 22198
rect 7644 22192 7956 22628
rect 8416 22816 9236 22820
rect 9364 22816 9676 23244
rect 8416 22808 9676 22816
rect 8468 22628 8608 22808
rect 8660 22628 8800 22808
rect 8852 22628 8992 22808
rect 9044 22628 9184 22808
rect 9236 22628 9676 22808
rect 8416 22618 8468 22628
rect 8608 22618 8660 22628
rect 8800 22618 8852 22628
rect 8992 22618 9044 22628
rect 9184 22618 9236 22628
rect 8320 22586 8372 22594
rect 8512 22586 8564 22594
rect 8704 22586 8756 22594
rect 8896 22586 8948 22594
rect 8316 22584 8948 22586
rect 9088 22584 9140 22594
rect 9280 22584 9332 22594
rect 8316 22576 8320 22584
rect 8372 22576 8512 22584
rect 8564 22576 8704 22584
rect 8756 22576 8896 22584
rect 8948 22404 9088 22584
rect 9140 22404 9280 22584
rect 8920 22396 9332 22404
rect 8920 22394 8948 22396
rect 9088 22394 9140 22396
rect 9280 22394 9332 22396
rect 8316 22382 8920 22392
rect 6696 22188 7956 22192
rect 6748 22008 6888 22188
rect 6940 22008 7080 22188
rect 7132 22008 7272 22188
rect 7324 22008 7464 22188
rect 7516 22008 7956 22188
rect 6696 22004 7956 22008
rect 8416 22192 8468 22198
rect 8608 22192 8660 22198
rect 8800 22192 8852 22198
rect 8992 22192 9044 22198
rect 9184 22192 9236 22198
rect 9364 22192 9676 22628
rect 8416 22188 9676 22192
rect 8468 22008 8608 22188
rect 8660 22008 8800 22188
rect 8852 22008 8992 22188
rect 9044 22008 9184 22188
rect 9236 22008 9676 22188
rect 8416 22004 9676 22008
rect 15900 22940 17840 23300
rect 18336 23156 18700 23410
rect 19044 23448 19232 23458
rect 19044 23354 19232 23364
rect 18336 23024 19408 23156
rect 15900 22180 16300 22940
rect 18336 22848 18396 23024
rect 18448 22848 18588 23024
rect 18396 22834 18448 22844
rect 18640 22848 18780 23024
rect 18588 22834 18640 22844
rect 18832 22848 18972 23024
rect 18780 22834 18832 22844
rect 19024 22848 19164 23024
rect 18972 22834 19024 22844
rect 19216 22848 19408 23024
rect 19164 22834 19216 22844
rect 18300 22800 18352 22810
rect 18272 22784 18300 22794
rect 18492 22800 18544 22810
rect 18352 22784 18492 22796
rect 18684 22800 18736 22810
rect 18544 22784 18684 22796
rect 18876 22800 18928 22810
rect 18736 22784 18876 22796
rect 18860 22620 18876 22784
rect 19068 22800 19120 22810
rect 18928 22620 19068 22796
rect 19260 22800 19312 22810
rect 19120 22620 19260 22796
rect 18860 22488 19312 22620
rect 18272 22462 18860 22472
rect 18392 22238 19212 22336
rect 6696 21998 6748 22004
rect 6888 21998 6940 22004
rect 7080 21998 7132 22004
rect 7272 21998 7324 22004
rect 7464 21998 7516 22004
rect 8416 21998 8468 22004
rect 8608 21998 8660 22004
rect 8800 21998 8852 22004
rect 8992 21998 9044 22004
rect 9184 21998 9236 22004
rect 6600 21966 6652 21974
rect 6792 21966 6844 21974
rect 6984 21966 7036 21974
rect 7176 21966 7228 21974
rect 6592 21964 7228 21966
rect 7368 21964 7420 21974
rect 7560 21964 7612 21974
rect 8320 21966 8372 21974
rect 8512 21966 8564 21974
rect 8704 21966 8756 21974
rect 8896 21966 8948 21974
rect 6592 21956 6600 21964
rect 6652 21956 6792 21964
rect 6844 21956 6984 21964
rect 7036 21956 7176 21964
rect 7228 21784 7368 21964
rect 7420 21784 7560 21964
rect 7196 21776 7612 21784
rect 7196 21774 7228 21776
rect 7368 21774 7420 21776
rect 7560 21774 7612 21776
rect 8312 21964 8948 21966
rect 9088 21964 9140 21974
rect 9280 21964 9332 21974
rect 8312 21956 8320 21964
rect 8372 21956 8512 21964
rect 8564 21956 8704 21964
rect 8756 21956 8896 21964
rect 8948 21784 9088 21964
rect 9140 21784 9280 21964
rect 6592 21762 7196 21772
rect 8916 21776 9332 21784
rect 8916 21774 8948 21776
rect 9088 21774 9140 21776
rect 9280 21774 9332 21776
rect 8312 21762 8916 21772
rect 18284 22228 19212 22238
rect 18864 22168 19212 22228
rect 18864 21996 18968 22168
rect 18284 21988 18392 21996
rect 18444 21988 18584 21996
rect 18636 21988 18776 21996
rect 18828 21992 18968 21996
rect 18828 21988 18864 21992
rect 18284 21986 18864 21988
rect 19020 21992 19160 22168
rect 18392 21978 18444 21986
rect 18584 21978 18636 21986
rect 18776 21978 18828 21986
rect 18968 21978 19020 21988
rect 19160 21978 19212 21988
rect 15900 21730 16300 21740
rect 18300 21944 18352 21954
rect 18488 21944 18540 21954
rect 18352 21764 18488 21940
rect 18680 21944 18732 21954
rect 18540 21764 18680 21940
rect 18872 21944 18924 21954
rect 18732 21764 18872 21940
rect 19064 21944 19116 21954
rect 18924 21916 19064 21940
rect 19256 21944 19308 21954
rect 19116 21916 19256 21940
rect 19308 21926 19312 21940
rect 19308 21916 19628 21926
rect 18924 21764 18996 21916
rect 18300 21688 18996 21764
rect 18300 21678 19628 21688
rect 18300 21676 19312 21678
rect 18284 21616 19216 21640
rect 18864 21548 19216 21616
rect 18864 21384 18972 21548
rect 18284 21374 18396 21384
rect 18448 21372 18588 21384
rect 18396 21358 18448 21368
rect 18640 21372 18780 21384
rect 18588 21358 18640 21368
rect 18832 21372 18972 21384
rect 18780 21358 18832 21368
rect 19024 21372 19164 21548
rect 18972 21358 19024 21368
rect 19164 21358 19216 21368
rect 24560 21500 24880 21510
rect 18304 21328 18356 21334
rect 18492 21328 18544 21334
rect 18684 21328 18736 21334
rect 18876 21328 18928 21334
rect 19068 21330 19120 21334
rect 19260 21330 19312 21334
rect 19000 21328 19632 21330
rect 18304 21324 19636 21328
rect 6600 21288 7200 21298
rect 8320 21288 8920 21298
rect 7200 21276 8320 21288
rect 8920 21276 9404 21288
rect 7200 21104 7632 21276
rect 6652 21096 7116 21104
rect 7168 21096 7632 21104
rect 7684 21096 8320 21276
rect 8920 21104 9352 21276
rect 8372 21096 8836 21104
rect 8888 21096 9352 21104
rect 6600 21094 7200 21096
rect 6600 21086 6652 21094
rect 7116 21086 7168 21094
rect 7632 21086 7684 21096
rect 8320 21094 8920 21096
rect 8320 21086 8372 21094
rect 8836 21086 8888 21094
rect 9352 21086 9404 21096
rect 10380 21220 10840 21230
rect 6860 21056 6912 21066
rect 7376 21058 7428 21066
rect 7892 21058 7944 21066
rect 7344 21056 7944 21058
rect 6912 21048 7376 21056
rect 7428 21048 7892 21056
rect 6912 20876 7344 21048
rect 6860 20864 7344 20876
rect 8580 21056 8632 21066
rect 9096 21058 9148 21066
rect 9612 21058 9664 21066
rect 9064 21056 9664 21058
rect 8632 21048 9096 21056
rect 9148 21048 9612 21056
rect 8632 20876 9064 21048
rect 8580 20864 9064 20876
rect 7344 20854 7944 20864
rect 9064 20854 9664 20864
rect 18356 21144 18492 21324
rect 18544 21144 18684 21324
rect 18736 21144 18876 21324
rect 18928 21320 19068 21324
rect 19120 21320 19260 21324
rect 19312 21320 19636 21324
rect 18928 21144 19000 21320
rect 18304 21092 19000 21144
rect 19632 21092 19636 21320
rect 24880 21140 25620 21500
rect 24560 21130 24880 21140
rect 18304 21080 19636 21092
rect 10380 20850 10840 20860
rect 18996 20752 19628 20762
rect 18560 20684 18996 20752
rect 19628 20684 19644 20752
rect 6600 20672 7200 20682
rect 8320 20672 8920 20682
rect 7200 20660 7684 20672
rect 7200 20488 7632 20660
rect 6652 20480 7116 20488
rect 7168 20480 7632 20488
rect 6600 20478 7200 20480
rect 6600 20470 6652 20478
rect 7116 20470 7168 20478
rect 7632 20470 7684 20480
rect 8920 20660 9404 20672
rect 8920 20488 9352 20660
rect 8372 20480 8836 20488
rect 8888 20480 9352 20488
rect 18612 20524 18996 20684
rect 18612 20508 19076 20524
rect 18560 20494 18612 20504
rect 19128 20508 19592 20524
rect 19076 20494 19128 20504
rect 19592 20494 19644 20504
rect 8320 20478 8920 20480
rect 8320 20470 8372 20478
rect 8836 20470 8888 20478
rect 9352 20470 9404 20480
rect 18300 20460 18352 20470
rect 6860 20440 6912 20450
rect 7376 20442 7428 20450
rect 7892 20442 7944 20450
rect 7344 20440 7944 20442
rect 6912 20432 7376 20440
rect 7428 20432 7892 20440
rect 6912 20260 7344 20432
rect 6860 20248 7344 20260
rect 8580 20440 8632 20450
rect 9096 20442 9148 20450
rect 9612 20442 9664 20450
rect 9064 20440 9664 20442
rect 8632 20432 9096 20440
rect 9148 20432 9612 20440
rect 8632 20260 9064 20432
rect 8580 20248 9064 20260
rect 7344 20238 7944 20248
rect 9064 20238 9664 20248
rect 18816 20460 18868 20470
rect 18352 20448 18816 20458
rect 19332 20460 19384 20470
rect 18868 20456 18888 20458
rect 18868 20448 19332 20456
rect 18888 20280 19332 20448
rect 18300 20220 18308 20280
rect 18888 20220 19384 20280
rect 18300 20212 19384 20220
rect 18308 20210 18888 20212
rect 18996 20132 19628 20138
rect 18560 20128 19644 20132
rect 18560 20064 18996 20128
rect 19628 20064 19644 20128
rect 6600 20052 7200 20062
rect 8320 20052 8920 20062
rect 7200 20040 7684 20052
rect 7200 19868 7632 20040
rect 6652 19860 7116 19868
rect 7168 19860 7632 19868
rect 6600 19858 7200 19860
rect 6600 19850 6652 19858
rect 7116 19850 7168 19858
rect 7632 19850 7684 19860
rect 8920 20040 9404 20052
rect 8920 19868 9352 20040
rect 8372 19860 8836 19868
rect 8888 19860 9352 19868
rect 8320 19858 8920 19860
rect 8320 19850 8372 19858
rect 8836 19850 8888 19858
rect 9352 19850 9404 19860
rect 10252 19868 10900 19892
rect 18612 19900 18996 20064
rect 18612 19888 19076 19900
rect 18560 19874 18612 19884
rect 19128 19888 19592 19900
rect 19076 19874 19128 19884
rect 19592 19874 19644 19884
rect 10252 19846 10276 19868
rect 10188 19836 10276 19846
rect 6860 19820 6912 19830
rect 7376 19822 7428 19830
rect 7892 19822 7944 19830
rect 7344 19820 7944 19822
rect 6912 19812 7376 19820
rect 7428 19812 7892 19820
rect 6912 19640 7344 19812
rect 6860 19628 7344 19640
rect 8580 19820 8632 19830
rect 9096 19822 9148 19830
rect 9612 19822 9664 19830
rect 9064 19820 9664 19822
rect 8632 19812 9096 19820
rect 9148 19812 9612 19820
rect 8632 19640 9064 19812
rect 10260 19768 10276 19836
rect 10188 19758 10276 19768
rect 8580 19628 9064 19640
rect 7344 19618 7944 19628
rect 9064 19618 9664 19628
rect 10252 19728 10276 19758
rect 10876 19728 10900 19868
rect 10312 19556 10444 19580
rect 10252 19538 10312 19548
rect 10504 19556 10636 19580
rect 10444 19538 10504 19548
rect 10696 19556 10828 19580
rect 10636 19538 10696 19548
rect 10888 19556 10900 19728
rect 18300 19840 18352 19850
rect 18816 19840 18868 19850
rect 18352 19828 18816 19838
rect 19332 19840 19384 19850
rect 18868 19836 18888 19838
rect 18868 19828 19332 19836
rect 18888 19660 19332 19828
rect 18300 19600 18308 19660
rect 18888 19600 19384 19660
rect 18300 19592 19384 19600
rect 18308 19590 18888 19592
rect 10828 19538 10888 19548
rect 18996 19516 19628 19522
rect 10160 19504 10220 19514
rect 10040 19478 10160 19498
rect 10024 19468 10160 19478
rect 10348 19504 10408 19514
rect 10220 19468 10348 19498
rect 10540 19504 10600 19514
rect 10408 19468 10540 19498
rect 10732 19504 10792 19514
rect 10600 19496 10624 19498
rect 10600 19468 10732 19496
rect 6600 19436 7200 19446
rect 8320 19436 8920 19446
rect 7200 19424 7684 19436
rect 7200 19252 7632 19424
rect 6652 19244 7116 19252
rect 7168 19244 7632 19252
rect 6600 19242 7200 19244
rect 6600 19234 6652 19242
rect 7116 19234 7168 19242
rect 7632 19234 7684 19244
rect 8920 19424 9404 19436
rect 8920 19252 9352 19424
rect 8372 19244 8836 19252
rect 8888 19244 9352 19252
rect 8320 19242 8920 19244
rect 8320 19234 8372 19242
rect 8836 19234 8888 19242
rect 9352 19234 9404 19244
rect 10640 19324 10732 19468
rect 6860 19204 6912 19214
rect 7376 19206 7428 19214
rect 7892 19206 7944 19214
rect 7344 19204 7944 19206
rect 6912 19196 7376 19204
rect 7428 19196 7892 19204
rect 6912 19024 7344 19196
rect 6860 19012 7344 19024
rect 8580 19204 8632 19214
rect 9096 19206 9148 19214
rect 9612 19206 9664 19214
rect 9064 19204 9664 19206
rect 8632 19196 9096 19204
rect 9148 19196 9612 19204
rect 8632 19024 9064 19196
rect 10640 19284 10792 19324
rect 18560 19512 19644 19516
rect 18560 19448 18996 19512
rect 19628 19448 19644 19512
rect 18612 19284 18996 19448
rect 18612 19272 19076 19284
rect 18560 19258 18612 19268
rect 19128 19272 19592 19284
rect 19076 19258 19128 19268
rect 19592 19258 19644 19268
rect 10024 19162 10640 19172
rect 18300 19224 18352 19234
rect 18816 19224 18868 19234
rect 18352 19212 18816 19222
rect 19332 19224 19384 19234
rect 18868 19220 18888 19222
rect 18868 19212 19332 19220
rect 8580 19012 9064 19024
rect 7344 19002 7944 19012
rect 9064 19002 9664 19012
rect 18888 19044 19332 19212
rect 18300 18984 18308 19044
rect 18888 18984 19384 19044
rect 18300 18976 19384 18984
rect 18308 18974 18888 18976
rect 19000 18916 19632 18926
rect 10252 18886 11080 18888
rect 10040 18876 11080 18886
rect 6600 18816 7200 18826
rect 8320 18816 8920 18826
rect 7200 18804 7684 18816
rect 7200 18632 7632 18804
rect 6652 18624 7116 18632
rect 7168 18624 7632 18632
rect 6600 18622 7200 18624
rect 6600 18614 6652 18622
rect 7116 18614 7168 18622
rect 7632 18614 7684 18624
rect 8920 18804 9404 18816
rect 8920 18632 9352 18804
rect 8372 18624 8836 18632
rect 8888 18624 9352 18632
rect 10624 18804 11080 18876
rect 10624 18644 10636 18804
rect 10040 18634 10252 18644
rect 8320 18622 8920 18624
rect 8320 18614 8372 18622
rect 8836 18614 8888 18622
rect 9352 18614 9404 18624
rect 10312 18632 10444 18644
rect 10252 18614 10312 18624
rect 10504 18632 10636 18644
rect 10444 18614 10504 18624
rect 10696 18632 10828 18804
rect 10636 18614 10696 18624
rect 10888 18632 11020 18804
rect 10828 18614 10888 18624
rect 11020 18614 11080 18624
rect 15580 18860 15980 18870
rect 6860 18584 6912 18594
rect 7376 18586 7428 18594
rect 7892 18586 7944 18594
rect 7344 18584 7944 18586
rect 6912 18576 7376 18584
rect 7428 18576 7892 18584
rect 6912 18404 7344 18576
rect 6860 18392 7344 18404
rect 8580 18584 8632 18594
rect 9096 18586 9148 18594
rect 9612 18586 9664 18594
rect 9064 18584 9664 18586
rect 8632 18576 9096 18584
rect 9148 18576 9612 18584
rect 8632 18404 9064 18576
rect 8580 18392 9064 18404
rect 7344 18382 7944 18392
rect 9064 18382 9664 18392
rect 10160 18584 10220 18594
rect 10348 18584 10408 18594
rect 10220 18404 10348 18576
rect 10540 18584 10600 18594
rect 10408 18404 10540 18576
rect 10732 18584 10792 18594
rect 10600 18404 10732 18576
rect 10924 18584 10984 18594
rect 10792 18560 10924 18576
rect 11116 18584 11176 18594
rect 10984 18560 11116 18576
rect 11176 18560 11296 18570
rect 15580 18410 15980 18420
rect 10160 18336 10768 18404
rect 10160 18326 11296 18336
rect 10160 18320 11176 18326
rect 10252 18266 11080 18272
rect 10040 18256 11080 18266
rect 6600 18200 7200 18210
rect 8320 18200 8920 18210
rect 7200 18188 7684 18200
rect 7200 18016 7632 18188
rect 6652 18008 7116 18016
rect 7168 18008 7632 18016
rect 6600 18006 7200 18008
rect 6600 17998 6652 18006
rect 7116 17998 7168 18006
rect 7632 17998 7684 18008
rect 8920 18188 9404 18200
rect 8920 18016 9352 18188
rect 8372 18008 8836 18016
rect 8888 18008 9352 18016
rect 10624 18188 11080 18256
rect 10624 18032 10636 18188
rect 10040 18022 10252 18032
rect 8320 18006 8920 18008
rect 8320 17998 8372 18006
rect 8836 17998 8888 18006
rect 9352 17998 9404 18008
rect 10312 18016 10444 18032
rect 10252 17998 10312 18008
rect 10504 18016 10636 18032
rect 10444 17998 10504 18008
rect 10696 18016 10828 18188
rect 10636 17998 10696 18008
rect 10888 18016 11020 18188
rect 10828 17998 10888 18008
rect 11020 17998 11080 18008
rect 6860 17968 6912 17978
rect 7376 17970 7428 17978
rect 7892 17970 7944 17978
rect 7344 17968 7944 17970
rect 6912 17960 7376 17968
rect 7428 17960 7892 17968
rect 6912 17788 7344 17960
rect 6860 17776 7344 17788
rect 8580 17968 8632 17978
rect 9096 17970 9148 17978
rect 9612 17970 9664 17978
rect 9064 17968 9664 17970
rect 8632 17960 9096 17968
rect 9148 17960 9612 17968
rect 8632 17788 9064 17960
rect 7344 17766 7944 17776
rect 8040 17776 8220 17786
rect 8580 17776 9064 17788
rect 9064 17766 9664 17776
rect 10160 17964 10220 17974
rect 10348 17964 10408 17974
rect 10220 17784 10348 17956
rect 10540 17964 10600 17974
rect 10408 17784 10540 17956
rect 10732 17964 10792 17974
rect 10600 17784 10732 17956
rect 10924 17964 10984 17974
rect 10792 17940 10924 17956
rect 11116 17964 11176 17974
rect 10984 17940 11116 17956
rect 11176 17940 11292 17950
rect 10160 17716 10764 17784
rect 10160 17706 11292 17716
rect 10160 17700 11176 17706
rect 8040 17606 8220 17616
rect 15620 11760 15980 18410
rect 1980 11400 15980 11760
rect 16220 18860 16620 18870
rect 18560 18828 19000 18896
rect 19632 18828 19644 18896
rect 18612 18688 19000 18828
rect 18612 18652 19076 18688
rect 18560 18638 18612 18648
rect 19128 18652 19592 18688
rect 19076 18638 19128 18648
rect 19592 18638 19644 18648
rect 1300 10768 1568 10778
rect 1300 10522 1568 10532
rect 1980 9800 2300 11400
rect 2588 11148 4792 11158
rect 2588 10650 4792 10660
rect 6096 10808 6276 10818
rect 6096 10598 6276 10608
rect 15700 10768 15968 10778
rect 15700 10522 15968 10532
rect 5208 10364 7200 10380
rect 5208 10284 6212 10364
rect 5208 10108 5212 10284
rect 5268 10108 5404 10284
rect 5212 10094 5268 10104
rect 5460 10108 5596 10284
rect 5404 10094 5460 10104
rect 5652 10108 5788 10284
rect 5596 10094 5652 10104
rect 5844 10108 5980 10284
rect 5788 10094 5844 10104
rect 6036 10108 6172 10284
rect 7188 10120 7200 10364
rect 8760 10292 9632 10302
rect 5980 10094 6036 10104
rect 6228 10108 6364 10120
rect 6172 10094 6228 10104
rect 6420 10108 6556 10120
rect 6364 10094 6420 10104
rect 6612 10108 6748 10120
rect 6556 10094 6612 10104
rect 6804 10108 6940 10120
rect 6748 10094 6804 10104
rect 6996 10108 7200 10120
rect 7708 10264 8760 10276
rect 6940 10094 6996 10104
rect 7708 10084 7712 10264
rect 7768 10084 7904 10264
rect 7712 10070 7768 10080
rect 7960 10084 8096 10264
rect 7904 10070 7960 10080
rect 8152 10084 8288 10264
rect 8096 10070 8152 10080
rect 8344 10084 8480 10264
rect 8288 10070 8344 10080
rect 8536 10084 8672 10264
rect 8480 10070 8536 10080
rect 8728 10092 8760 10264
rect 8728 10084 8864 10092
rect 8760 10082 8864 10084
rect 8672 10070 8728 10080
rect 8920 10082 9056 10092
rect 8864 10070 8920 10080
rect 9112 10082 9248 10092
rect 9056 10070 9112 10080
rect 9304 10082 9440 10092
rect 9248 10070 9304 10080
rect 9496 10082 9632 10092
rect 9440 10070 9496 10080
rect 5116 10062 5172 10070
rect 5308 10062 5364 10070
rect 5500 10062 5556 10070
rect 5692 10062 5748 10070
rect 5884 10062 5940 10070
rect 6076 10062 6132 10070
rect 5112 10060 6132 10062
rect 5112 10052 5116 10060
rect 5172 10052 5308 10060
rect 5364 10052 5500 10060
rect 5556 10052 5692 10060
rect 5748 10052 5884 10060
rect 5940 10052 6076 10060
rect 6268 10060 6324 10070
rect 2588 9908 4780 9918
rect -3300 9796 2320 9800
rect -3300 9440 2588 9796
rect 6132 9880 6268 10056
rect 6460 10060 6516 10070
rect 6324 9880 6460 10056
rect 6652 10060 6708 10070
rect 6516 9880 6652 10056
rect 6844 10060 6900 10070
rect 6708 9880 6844 10056
rect 7036 10060 7092 10070
rect 6900 9880 7036 10056
rect 7092 9880 7104 10056
rect 7616 10044 7672 10054
rect 6088 9796 7104 9880
rect 7608 10032 7616 10042
rect 7808 10044 7864 10054
rect 7672 10032 7808 10042
rect 8000 10044 8056 10054
rect 7864 10032 8000 10042
rect 8192 10044 8248 10054
rect 8056 10032 8192 10042
rect 8384 10044 8440 10054
rect 8248 10032 8384 10042
rect 8576 10044 8632 10054
rect 8440 10032 8576 10042
rect 8768 10044 8824 10054
rect 8632 9860 8768 10040
rect 8960 10044 9016 10054
rect 8824 9860 8960 10040
rect 9152 10044 9208 10054
rect 9016 9860 9152 10040
rect 9344 10044 9400 10054
rect 9208 9860 9344 10040
rect 9536 10044 9592 10054
rect 9400 9860 9536 10040
rect 8592 9848 9592 9860
rect 7608 9834 8592 9844
rect 16220 9796 16620 18420
rect 18300 18604 18352 18614
rect 18816 18604 18868 18614
rect 18352 18592 18816 18602
rect 19332 18604 19384 18614
rect 18868 18600 18888 18602
rect 18868 18592 19332 18600
rect 18888 18424 19332 18592
rect 18300 18364 18308 18424
rect 18888 18364 19384 18424
rect 18300 18356 19384 18364
rect 18308 18354 18888 18356
rect 18480 18156 18680 18166
rect 18480 18046 18680 18056
rect 16988 11148 19192 11158
rect 16988 10650 19192 10660
rect 20496 10808 20676 10818
rect 20496 10598 20676 10608
rect 19608 10364 21600 10380
rect 19608 10284 20612 10364
rect 19608 10108 19612 10284
rect 19668 10108 19804 10284
rect 19612 10094 19668 10104
rect 19860 10108 19996 10284
rect 19804 10094 19860 10104
rect 20052 10108 20188 10284
rect 19996 10094 20052 10104
rect 20244 10108 20380 10284
rect 20188 10094 20244 10104
rect 20436 10108 20572 10284
rect 21588 10120 21600 10364
rect 23160 10292 24032 10302
rect 20380 10094 20436 10104
rect 20628 10108 20764 10120
rect 20572 10094 20628 10104
rect 20820 10108 20956 10120
rect 20764 10094 20820 10104
rect 21012 10108 21148 10120
rect 20956 10094 21012 10104
rect 21204 10108 21340 10120
rect 21148 10094 21204 10104
rect 21396 10108 21600 10120
rect 22108 10264 23160 10276
rect 21340 10094 21396 10104
rect 22108 10084 22112 10264
rect 22168 10084 22304 10264
rect 22112 10070 22168 10080
rect 22360 10084 22496 10264
rect 22304 10070 22360 10080
rect 22552 10084 22688 10264
rect 22496 10070 22552 10080
rect 22744 10084 22880 10264
rect 22688 10070 22744 10080
rect 22936 10084 23072 10264
rect 22880 10070 22936 10080
rect 23128 10092 23160 10264
rect 23128 10084 23264 10092
rect 23160 10082 23264 10084
rect 23072 10070 23128 10080
rect 23320 10082 23456 10092
rect 23264 10070 23320 10080
rect 23512 10082 23648 10092
rect 23456 10070 23512 10080
rect 23704 10082 23840 10092
rect 23648 10070 23704 10080
rect 23896 10082 24032 10092
rect 23840 10070 23896 10080
rect 19516 10062 19572 10070
rect 19708 10062 19764 10070
rect 19900 10062 19956 10070
rect 20092 10062 20148 10070
rect 20284 10062 20340 10070
rect 20476 10062 20532 10070
rect 19512 10060 20532 10062
rect 19512 10052 19516 10060
rect 19572 10052 19708 10060
rect 19764 10052 19900 10060
rect 19956 10052 20092 10060
rect 20148 10052 20284 10060
rect 20340 10052 20476 10060
rect 20668 10060 20724 10070
rect 16988 9908 19180 9918
rect 4780 9440 4784 9796
rect 5112 9784 7104 9796
rect 5200 9732 7192 9748
rect 5200 9652 6212 9732
rect 5200 9476 5212 9652
rect 5268 9476 5404 9652
rect 5212 9462 5268 9472
rect 5460 9476 5596 9652
rect 5404 9462 5460 9472
rect 5652 9476 5788 9652
rect 5596 9462 5652 9472
rect 5844 9476 5980 9652
rect 5788 9462 5844 9472
rect 6036 9476 6172 9652
rect 7188 9488 7192 9732
rect 8764 9676 9636 9686
rect 5980 9462 6036 9472
rect 6228 9476 6364 9488
rect 6172 9462 6228 9472
rect 6420 9476 6556 9488
rect 6364 9462 6420 9472
rect 6612 9476 6748 9488
rect 6556 9462 6612 9472
rect 6804 9476 6940 9488
rect 6748 9462 6804 9472
rect 6996 9476 7192 9488
rect 7708 9648 8764 9660
rect 6940 9462 6996 9472
rect 7708 9468 7712 9648
rect 7768 9468 7904 9648
rect 7712 9454 7768 9464
rect 7960 9468 8096 9648
rect 7904 9454 7960 9464
rect 8152 9468 8288 9648
rect 8096 9454 8152 9464
rect 8344 9468 8480 9648
rect 8288 9454 8344 9464
rect 8536 9468 8672 9648
rect 8480 9454 8536 9464
rect 8728 9476 8764 9648
rect 8728 9468 8864 9476
rect 8764 9466 8864 9468
rect 8672 9454 8728 9464
rect 8920 9466 9056 9476
rect 8864 9454 8920 9464
rect 9112 9466 9248 9476
rect 9056 9454 9112 9464
rect 9304 9466 9440 9476
rect 9248 9454 9304 9464
rect 9496 9466 9636 9476
rect 9440 9454 9496 9464
rect -10000 8800 -8800 9400
rect -3300 9124 4784 9440
rect 15388 9440 16988 9796
rect 20532 9880 20668 10056
rect 20860 10060 20916 10070
rect 20724 9880 20860 10056
rect 21052 10060 21108 10070
rect 20916 9880 21052 10056
rect 21244 10060 21300 10070
rect 21108 9880 21244 10056
rect 21436 10060 21492 10070
rect 21300 9880 21436 10056
rect 21492 9880 21504 10056
rect 22016 10044 22072 10054
rect 20488 9796 21504 9880
rect 22008 10032 22016 10042
rect 22208 10044 22264 10054
rect 22072 10032 22208 10042
rect 22400 10044 22456 10054
rect 22264 10032 22400 10042
rect 22592 10044 22648 10054
rect 22456 10032 22592 10042
rect 22784 10044 22840 10054
rect 22648 10032 22784 10042
rect 22976 10044 23032 10054
rect 22840 10032 22976 10042
rect 23168 10044 23224 10054
rect 23032 9860 23168 10040
rect 23360 10044 23416 10054
rect 23224 9860 23360 10040
rect 23552 10044 23608 10054
rect 23416 9860 23552 10040
rect 23744 10044 23800 10054
rect 23608 9860 23744 10040
rect 23936 10044 23992 10054
rect 23800 9860 23936 10040
rect 22992 9848 23992 9860
rect 22008 9834 22992 9844
rect 19180 9440 19184 9796
rect 19512 9784 21504 9796
rect 21460 9780 21490 9784
rect 19600 9732 21592 9748
rect 19600 9652 20612 9732
rect 19600 9476 19612 9652
rect 19668 9476 19804 9652
rect 19612 9462 19668 9472
rect 19860 9476 19996 9652
rect 19804 9462 19860 9472
rect 20052 9476 20188 9652
rect 19996 9462 20052 9472
rect 20244 9476 20380 9652
rect 20188 9462 20244 9472
rect 20436 9476 20572 9652
rect 21588 9488 21592 9732
rect 23164 9676 24036 9686
rect 20380 9462 20436 9472
rect 20628 9476 20764 9488
rect 20572 9462 20628 9472
rect 20820 9476 20956 9488
rect 20764 9462 20820 9472
rect 21012 9476 21148 9488
rect 20956 9462 21012 9472
rect 21204 9476 21340 9488
rect 21148 9462 21204 9472
rect 21396 9476 21592 9488
rect 22108 9648 23164 9660
rect 21340 9462 21396 9472
rect 22108 9468 22112 9648
rect 22168 9468 22304 9648
rect 22112 9454 22168 9464
rect 22360 9468 22496 9648
rect 22304 9454 22360 9464
rect 22552 9468 22688 9648
rect 22496 9454 22552 9464
rect 22744 9468 22880 9648
rect 22688 9454 22744 9464
rect 22936 9468 23072 9648
rect 22880 9454 22936 9464
rect 23128 9476 23164 9648
rect 23128 9468 23264 9476
rect 23164 9466 23264 9468
rect 23072 9454 23128 9464
rect 23320 9466 23456 9476
rect 23264 9454 23320 9464
rect 23512 9466 23648 9476
rect 23456 9454 23512 9464
rect 23704 9466 23840 9476
rect 23648 9454 23704 9464
rect 23896 9466 24036 9476
rect 23840 9454 23896 9464
rect 5116 9430 5172 9438
rect 5308 9430 5364 9438
rect 5500 9430 5556 9438
rect 5692 9430 5748 9438
rect 5884 9430 5940 9438
rect 6076 9430 6132 9438
rect 5112 9428 6132 9430
rect 5112 9420 5116 9428
rect 5172 9420 5308 9428
rect 5364 9420 5500 9428
rect 5556 9420 5692 9428
rect 5748 9420 5884 9428
rect 5940 9420 6076 9428
rect 6268 9428 6324 9438
rect 6132 9248 6268 9424
rect 6460 9428 6516 9438
rect 6324 9248 6460 9424
rect 6652 9428 6708 9438
rect 6516 9248 6652 9424
rect 6844 9428 6900 9438
rect 6708 9248 6844 9424
rect 7036 9428 7092 9438
rect 6900 9248 7036 9424
rect 7616 9428 7672 9438
rect 7092 9248 7104 9424
rect 6088 9160 7104 9248
rect 7612 9412 7616 9424
rect 7808 9428 7864 9438
rect 7672 9412 7808 9424
rect 8000 9428 8056 9438
rect 7864 9412 8000 9424
rect 8192 9428 8248 9438
rect 8056 9412 8192 9424
rect 8384 9428 8440 9438
rect 8248 9412 8384 9424
rect 8576 9428 8632 9438
rect 8440 9412 8576 9424
rect 8768 9428 8824 9438
rect 8632 9244 8768 9424
rect 8960 9428 9016 9438
rect 8824 9244 8960 9424
rect 9152 9428 9208 9438
rect 9016 9244 9152 9424
rect 9344 9428 9400 9438
rect 9208 9244 9344 9424
rect 9536 9428 9592 9438
rect 9400 9244 9536 9424
rect 8596 9232 9592 9244
rect 7612 9214 8596 9224
rect 5112 9152 7104 9160
rect 5112 9150 6088 9152
rect 15388 9124 19184 9440
rect 19516 9430 19572 9438
rect 19708 9430 19764 9438
rect 19900 9430 19956 9438
rect 20092 9430 20148 9438
rect 20284 9430 20340 9438
rect 20476 9430 20532 9438
rect 19512 9428 20532 9430
rect 19512 9420 19516 9428
rect 19572 9420 19708 9428
rect 19764 9420 19900 9428
rect 19956 9420 20092 9428
rect 20148 9420 20284 9428
rect 20340 9420 20476 9428
rect 20668 9428 20724 9438
rect 20532 9248 20668 9424
rect 20860 9428 20916 9438
rect 20724 9248 20860 9424
rect 21052 9428 21108 9438
rect 20916 9248 21052 9424
rect 21244 9428 21300 9438
rect 21108 9248 21244 9424
rect 21436 9428 21492 9438
rect 21300 9248 21436 9424
rect 22016 9428 22072 9438
rect 21492 9248 21504 9424
rect 20488 9160 21504 9248
rect 22012 9412 22016 9424
rect 22208 9428 22264 9438
rect 22072 9412 22208 9424
rect 22400 9428 22456 9438
rect 22264 9412 22400 9424
rect 22592 9428 22648 9438
rect 22456 9412 22592 9424
rect 22784 9428 22840 9438
rect 22648 9412 22784 9424
rect 22976 9428 23032 9438
rect 22840 9412 22976 9424
rect 23168 9428 23224 9438
rect 23032 9244 23168 9424
rect 23360 9428 23416 9438
rect 23224 9244 23360 9424
rect 23552 9428 23608 9438
rect 23416 9244 23552 9424
rect 23744 9428 23800 9438
rect 23608 9244 23744 9424
rect 23936 9428 23992 9438
rect 23800 9244 23936 9424
rect 22996 9232 23992 9244
rect 22012 9214 22996 9224
rect 19512 9152 21504 9160
rect 19512 9150 20488 9152
rect -3300 9120 2320 9124
rect -9960 8360 -9690 8608
rect -9200 8360 -8860 8800
rect 988 8518 1688 9120
rect 8764 9060 9636 9070
rect 7708 9028 8764 9040
rect 4588 8984 5008 8994
rect 1764 8964 2056 8974
rect 1764 8894 2056 8904
rect 1776 8820 2056 8894
rect 2540 8964 2832 8974
rect 3476 8968 3768 8974
rect 3476 8964 3772 8968
rect 2832 8904 2836 8960
rect 2540 8820 2836 8904
rect 3768 8904 3772 8964
rect 3476 8820 3772 8904
rect 1776 8732 4500 8820
rect 1828 8560 1968 8732
rect 1776 8542 1828 8552
rect 2020 8560 2160 8732
rect 1968 8542 2020 8552
rect 2212 8560 2352 8732
rect 2160 8542 2212 8552
rect 2404 8560 2544 8732
rect 2352 8542 2404 8552
rect 2596 8560 2736 8732
rect 2544 8542 2596 8552
rect 2788 8560 2928 8732
rect 2736 8542 2788 8552
rect 2980 8560 3120 8732
rect 2928 8542 2980 8552
rect 3172 8560 3312 8732
rect 3120 8542 3172 8552
rect 3364 8560 3504 8732
rect 3312 8542 3364 8552
rect 3556 8672 4500 8732
rect 3556 8560 3740 8672
rect 3504 8542 3556 8552
rect 988 8508 1732 8518
rect -9964 8356 -8716 8360
rect -9964 8280 -9044 8356
rect -8904 8280 -8716 8356
rect 988 8328 1680 8508
rect 1872 8508 1924 8518
rect 1732 8328 1872 8500
rect 2064 8508 2116 8518
rect 1924 8328 2064 8500
rect 2256 8508 2308 8518
rect 2116 8328 2256 8500
rect 2448 8508 2500 8518
rect 2308 8328 2448 8500
rect 2640 8508 2692 8518
rect 2500 8328 2640 8500
rect 2832 8508 2884 8518
rect 2692 8328 2832 8500
rect 3024 8508 3076 8518
rect 2884 8328 3024 8500
rect 3216 8508 3268 8518
rect 3076 8328 3216 8500
rect 3408 8508 3460 8518
rect 3268 8328 3408 8500
rect 3600 8508 3652 8518
rect 3460 8328 3600 8500
rect 3800 8560 4500 8672
rect 3740 8406 3800 8416
rect -9964 8236 -8716 8280
rect -9912 8060 -9772 8236
rect -9964 8046 -9912 8056
rect -9720 8060 -9580 8236
rect -9772 8046 -9720 8056
rect -9528 8060 -9388 8236
rect -9580 8046 -9528 8056
rect -9336 8060 -9196 8236
rect -9388 8046 -9336 8056
rect -9144 8060 -8716 8236
rect -8660 8296 -8480 8306
rect -8660 8186 -8480 8196
rect 988 8240 3652 8328
rect 4124 8356 4500 8560
rect 7708 8848 7712 9028
rect 7768 8848 7904 9028
rect 7712 8834 7768 8844
rect 7960 8848 8096 9028
rect 7904 8834 7960 8844
rect 8152 8848 8288 9028
rect 8096 8834 8152 8844
rect 8344 8848 8480 9028
rect 8288 8834 8344 8844
rect 8536 8848 8672 9028
rect 8480 8834 8536 8844
rect 8728 8860 8764 9028
rect 8728 8848 8864 8860
rect 8672 8834 8728 8844
rect 8920 8848 9056 8860
rect 8864 8834 8920 8844
rect 9112 8848 9248 8860
rect 9056 8834 9112 8844
rect 9304 8848 9440 8860
rect 9248 8834 9304 8844
rect 9496 8850 9636 8860
rect 9496 8848 9500 8850
rect 9440 8834 9496 8844
rect 7616 8808 7672 8818
rect 7608 8796 7616 8806
rect 7808 8808 7864 8818
rect 7672 8796 7808 8806
rect 8000 8808 8056 8818
rect 7864 8796 8000 8806
rect 8192 8808 8248 8818
rect 8056 8796 8192 8806
rect 8384 8808 8440 8818
rect 8248 8796 8384 8806
rect 8576 8808 8632 8818
rect 8440 8796 8576 8806
rect 8768 8808 8824 8818
rect 5208 8784 7200 8796
rect 5208 8700 6224 8784
rect 5208 8524 5212 8700
rect 5268 8524 5404 8700
rect 5212 8510 5268 8520
rect 5460 8524 5596 8700
rect 5404 8510 5460 8520
rect 5652 8524 5788 8700
rect 5596 8510 5652 8520
rect 5844 8524 5980 8700
rect 5788 8510 5844 8520
rect 6036 8524 6172 8700
rect 8632 8624 8768 8804
rect 8960 8808 9016 8818
rect 8824 8624 8960 8804
rect 9152 8808 9208 8818
rect 9016 8624 9152 8804
rect 9344 8808 9400 8818
rect 9208 8624 9344 8804
rect 9536 8808 9592 8818
rect 9400 8624 9536 8804
rect 8592 8612 9592 8624
rect 7608 8598 8592 8608
rect 5980 8510 6036 8520
rect 6228 8524 6364 8536
rect 6172 8510 6228 8520
rect 6420 8524 6556 8536
rect 6364 8510 6420 8520
rect 6612 8524 6748 8536
rect 6556 8510 6612 8520
rect 6804 8524 6940 8536
rect 6748 8510 6804 8520
rect 6996 8524 7200 8536
rect 6940 8510 6996 8520
rect 15388 8518 16088 9124
rect 16220 9120 16620 9124
rect 23164 9060 24036 9070
rect 22108 9028 23164 9040
rect 18988 8984 19408 8994
rect 16164 8964 16456 8974
rect 16164 8894 16456 8904
rect 16176 8820 16456 8894
rect 16940 8964 17232 8974
rect 17876 8968 18168 8974
rect 17876 8964 18172 8968
rect 17232 8904 17236 8960
rect 16940 8820 17236 8904
rect 18168 8904 18172 8964
rect 17876 8820 18172 8904
rect 16176 8732 18900 8820
rect 16228 8560 16368 8732
rect 16176 8542 16228 8552
rect 16420 8560 16560 8732
rect 16368 8542 16420 8552
rect 16612 8560 16752 8732
rect 16560 8542 16612 8552
rect 16804 8560 16944 8732
rect 16752 8542 16804 8552
rect 16996 8560 17136 8732
rect 16944 8542 16996 8552
rect 17188 8560 17328 8732
rect 17136 8542 17188 8552
rect 17380 8560 17520 8732
rect 17328 8542 17380 8552
rect 17572 8560 17712 8732
rect 17520 8542 17572 8552
rect 17764 8560 17904 8732
rect 17712 8542 17764 8552
rect 17956 8672 18900 8732
rect 17956 8560 18140 8672
rect 17904 8542 17956 8552
rect 15388 8508 16132 8518
rect 5116 8482 5172 8486
rect 5308 8482 5364 8486
rect 5500 8482 5556 8486
rect 5692 8482 5748 8486
rect 5884 8482 5940 8486
rect 6076 8482 6132 8486
rect 5104 8476 6132 8482
rect 5104 8472 5116 8476
rect 5172 8472 5308 8476
rect 5364 8472 5500 8476
rect 5556 8472 5692 8476
rect 5748 8472 5884 8476
rect 5940 8472 6076 8476
rect 6268 8476 6324 8486
rect 4588 8422 5008 8432
rect -9196 8046 -9144 8056
rect -10060 8012 -10008 8022
rect -9868 8012 -9816 8022
rect -10008 7852 -9868 8008
rect -9676 8012 -9624 8022
rect -9816 7852 -9676 8008
rect -9484 8012 -9432 8022
rect -9624 7852 -9484 8008
rect -9292 8012 -9240 8022
rect -9432 7852 -9292 8008
rect -10008 7832 -9968 7852
rect -9316 7832 -9292 7852
rect -9100 8012 -9048 8022
rect -9240 7832 -9100 8008
rect -10060 7584 -9968 7832
rect -9316 7620 -9048 7832
rect -9316 7584 -9196 7620
rect -10060 7448 -9964 7584
rect -9912 7448 -9772 7584
rect -9964 7430 -9912 7440
rect -9720 7448 -9580 7584
rect -9772 7430 -9720 7440
rect -9528 7448 -9388 7584
rect -9580 7430 -9528 7440
rect -9336 7448 -9196 7584
rect -9388 7430 -9336 7440
rect -9144 7448 -9048 7620
rect -9196 7430 -9144 7440
rect -10060 7396 -10008 7406
rect -10064 7216 -10060 7392
rect -9868 7396 -9816 7406
rect -10008 7216 -9868 7392
rect -9676 7396 -9624 7406
rect -9816 7216 -9676 7392
rect -9484 7396 -9432 7406
rect -9624 7216 -9484 7392
rect -9292 7396 -9240 7406
rect -9432 7216 -9292 7392
rect -9100 7396 -9048 7406
rect -9240 7216 -9100 7392
rect -8996 7392 -8716 8060
rect -9048 7216 -8716 7392
rect -10064 7050 -8716 7216
rect 988 7652 1620 8240
rect 1776 8162 2072 8164
rect 1764 8152 2072 8162
rect 2056 8088 2072 8152
rect 1764 8060 2072 8088
rect 1776 7936 2072 8060
rect 2540 8152 2860 8162
rect 2540 8078 2860 8088
rect 3476 8152 3768 8162
rect 3768 8092 3776 8144
rect 3476 8082 3776 8092
rect 2540 8000 2836 8078
rect 3480 8000 3776 8082
rect 4124 8000 4928 8356
rect 2540 7936 4928 8000
rect 1776 7912 4928 7936
rect 1828 7740 1968 7912
rect 1776 7722 1828 7732
rect 2020 7740 2160 7912
rect 1968 7722 2020 7732
rect 2212 7740 2352 7912
rect 2160 7722 2212 7732
rect 2404 7740 2544 7912
rect 2352 7722 2404 7732
rect 2596 7740 2736 7912
rect 2544 7722 2596 7732
rect 2788 7740 2928 7912
rect 2736 7722 2788 7732
rect 2980 7740 3120 7912
rect 2928 7722 2980 7732
rect 3172 7740 3312 7912
rect 3120 7722 3172 7732
rect 3364 7740 3504 7912
rect 3312 7722 3364 7732
rect 3556 7824 4928 7912
rect 3556 7740 3740 7824
rect 3504 7722 3556 7732
rect 1680 7688 1732 7698
rect 988 7508 1680 7652
rect 1872 7688 1924 7698
rect 1732 7508 1872 7652
rect 2064 7688 2116 7698
rect 1924 7508 2064 7680
rect 2256 7688 2308 7698
rect 2116 7508 2256 7680
rect 2448 7688 2500 7698
rect 2308 7508 2448 7680
rect 2640 7688 2692 7698
rect 2500 7508 2640 7680
rect 2832 7688 2884 7698
rect 2692 7508 2832 7680
rect 3024 7688 3076 7698
rect 2884 7508 3024 7680
rect 3216 7688 3268 7698
rect 3076 7508 3216 7680
rect 3408 7688 3460 7698
rect 3268 7508 3408 7680
rect 3600 7688 3652 7698
rect 3460 7508 3600 7680
rect 3800 7740 4928 7824
rect 3740 7558 3800 7568
rect 988 7420 3652 7508
rect -10064 7040 -8680 7050
rect -8456 7044 -8380 7054
rect -10064 7000 -8756 7040
rect -10064 6828 -9964 7000
rect -9912 6828 -9772 7000
rect -9964 6810 -9912 6820
rect -9720 6828 -9580 7000
rect -9772 6810 -9720 6820
rect -9528 6828 -9388 7000
rect -9580 6810 -9528 6820
rect -9336 6828 -9196 7000
rect -9388 6810 -9336 6820
rect -9144 6828 -8756 7000
rect -8680 6832 -8456 7040
rect -8680 6828 -8380 6832
rect -9196 6810 -9144 6820
rect -8756 6818 -8680 6828
rect -8456 6822 -8380 6828
rect -10060 6776 -10008 6786
rect -9868 6776 -9816 6786
rect -10008 6740 -9868 6772
rect -9676 6776 -9624 6786
rect -9816 6740 -9676 6772
rect -9484 6776 -9432 6786
rect -9624 6740 -9484 6772
rect -9292 6776 -9240 6786
rect -9432 6740 -9292 6772
rect -10008 6596 -9968 6740
rect -9316 6596 -9292 6740
rect -9100 6776 -9048 6786
rect -9240 6596 -9100 6772
rect -9048 6596 -9020 6772
rect -10060 6508 -9968 6596
rect -9316 6472 -9020 6596
rect -8660 6576 -8480 6582
rect -9968 6462 -9020 6472
rect -9324 6256 -9020 6462
rect -8720 6572 -8460 6576
rect -8720 6492 -8660 6572
rect -8480 6492 -8460 6572
rect -8720 6256 -8460 6492
rect -3090 6468 -2352 6910
rect 988 6878 1688 7420
rect 1764 7328 2056 7338
rect 2536 7328 2828 7338
rect 2056 7268 2060 7316
rect 1764 7180 2060 7268
rect 3476 7328 3768 7338
rect 2828 7268 2832 7320
rect 2536 7180 2832 7268
rect 3768 7268 3772 7292
rect 3476 7180 3772 7268
rect 4124 7180 4928 7740
rect 5076 8224 5104 8472
rect 6132 8296 6268 8472
rect 6460 8476 6516 8486
rect 6324 8296 6460 8472
rect 6652 8476 6708 8486
rect 6516 8296 6652 8472
rect 6844 8476 6900 8486
rect 6708 8296 6844 8472
rect 7036 8476 7092 8486
rect 6900 8296 7036 8472
rect 8764 8440 9636 8450
rect 6080 8224 7092 8296
rect 7708 8412 8764 8424
rect 7708 8232 7712 8412
rect 5076 8212 7092 8224
rect 7768 8232 7904 8412
rect 7712 8218 7768 8228
rect 7960 8232 8096 8412
rect 7904 8218 7960 8228
rect 8152 8232 8288 8412
rect 8096 8218 8152 8228
rect 8344 8232 8480 8412
rect 8288 8218 8344 8228
rect 8536 8232 8672 8412
rect 8480 8218 8536 8228
rect 8728 8240 8764 8412
rect 8728 8232 8864 8240
rect 8764 8230 8864 8232
rect 8672 8218 8728 8228
rect 8920 8230 9056 8240
rect 8864 8218 8920 8228
rect 9112 8230 9248 8240
rect 9056 8218 9112 8228
rect 9304 8230 9440 8240
rect 9248 8218 9304 8228
rect 9496 8230 9636 8240
rect 15388 8328 16080 8508
rect 16272 8508 16324 8518
rect 16132 8328 16272 8500
rect 16464 8508 16516 8518
rect 16324 8328 16464 8500
rect 16656 8508 16708 8518
rect 16516 8328 16656 8500
rect 16848 8508 16900 8518
rect 16708 8328 16848 8500
rect 17040 8508 17092 8518
rect 16900 8328 17040 8500
rect 17232 8508 17284 8518
rect 17092 8328 17232 8500
rect 17424 8508 17476 8518
rect 17284 8328 17424 8500
rect 17616 8508 17668 8518
rect 17476 8328 17616 8500
rect 17808 8508 17860 8518
rect 17668 8328 17808 8500
rect 18000 8508 18052 8518
rect 17860 8328 18000 8500
rect 18200 8560 18900 8672
rect 18140 8406 18200 8416
rect 15388 8240 18052 8328
rect 18524 8356 18900 8560
rect 22108 8848 22112 9028
rect 22168 8848 22304 9028
rect 22112 8834 22168 8844
rect 22360 8848 22496 9028
rect 22304 8834 22360 8844
rect 22552 8848 22688 9028
rect 22496 8834 22552 8844
rect 22744 8848 22880 9028
rect 22688 8834 22744 8844
rect 22936 8848 23072 9028
rect 22880 8834 22936 8844
rect 23128 8860 23164 9028
rect 23128 8848 23264 8860
rect 23072 8834 23128 8844
rect 23320 8848 23456 8860
rect 23264 8834 23320 8844
rect 23512 8848 23648 8860
rect 23456 8834 23512 8844
rect 23704 8848 23840 8860
rect 23648 8834 23704 8844
rect 23896 8850 24036 8860
rect 23896 8848 23900 8850
rect 23840 8834 23896 8844
rect 22016 8808 22072 8818
rect 22008 8796 22016 8806
rect 22208 8808 22264 8818
rect 22072 8796 22208 8806
rect 22400 8808 22456 8818
rect 22264 8796 22400 8806
rect 22592 8808 22648 8818
rect 22456 8796 22592 8806
rect 22784 8808 22840 8818
rect 22648 8796 22784 8806
rect 22976 8808 23032 8818
rect 22840 8796 22976 8806
rect 23168 8808 23224 8818
rect 19608 8784 21600 8796
rect 19608 8700 20624 8784
rect 19608 8524 19612 8700
rect 19668 8524 19804 8700
rect 19612 8510 19668 8520
rect 19860 8524 19996 8700
rect 19804 8510 19860 8520
rect 20052 8524 20188 8700
rect 19996 8510 20052 8520
rect 20244 8524 20380 8700
rect 20188 8510 20244 8520
rect 20436 8524 20572 8700
rect 23032 8624 23168 8804
rect 23360 8808 23416 8818
rect 23224 8624 23360 8804
rect 23552 8808 23608 8818
rect 23416 8624 23552 8804
rect 23744 8808 23800 8818
rect 23608 8624 23744 8804
rect 23936 8808 23992 8818
rect 23800 8624 23936 8804
rect 22992 8612 23992 8624
rect 22008 8598 22992 8608
rect 20380 8510 20436 8520
rect 20628 8524 20764 8536
rect 20572 8510 20628 8520
rect 20820 8524 20956 8536
rect 20764 8510 20820 8520
rect 21012 8524 21148 8536
rect 20956 8510 21012 8520
rect 21204 8524 21340 8536
rect 21148 8510 21204 8520
rect 21396 8524 21600 8536
rect 21340 8510 21396 8520
rect 19516 8482 19572 8486
rect 19708 8482 19764 8486
rect 19900 8482 19956 8486
rect 20092 8482 20148 8486
rect 20284 8482 20340 8486
rect 20476 8482 20532 8486
rect 19504 8476 20532 8482
rect 19504 8472 19516 8476
rect 19572 8472 19708 8476
rect 19764 8472 19900 8476
rect 19956 8472 20092 8476
rect 20148 8472 20284 8476
rect 20340 8472 20476 8476
rect 20668 8476 20724 8486
rect 18988 8422 19408 8432
rect 9440 8218 9496 8228
rect 5076 7858 5176 8212
rect 7616 8192 7672 8202
rect 7604 8180 7616 8190
rect 7808 8192 7864 8202
rect 7672 8180 7808 8190
rect 8000 8192 8056 8202
rect 7864 8180 8000 8190
rect 8192 8192 8248 8202
rect 8056 8180 8192 8190
rect 8384 8192 8440 8202
rect 8248 8180 8384 8190
rect 8576 8192 8632 8202
rect 8440 8180 8576 8190
rect 8768 8192 8824 8202
rect 5208 8164 7200 8176
rect 5208 8080 6224 8164
rect 5208 7904 5212 8080
rect 5268 7904 5404 8080
rect 5212 7890 5268 7900
rect 5460 7904 5596 8080
rect 5404 7890 5460 7900
rect 5652 7904 5788 8080
rect 5596 7890 5652 7900
rect 5844 7904 5980 8080
rect 5788 7890 5844 7900
rect 6036 7904 6172 8080
rect 8632 8008 8768 8188
rect 8960 8192 9016 8202
rect 8824 8008 8960 8188
rect 9152 8192 9208 8202
rect 9016 8008 9152 8188
rect 9344 8192 9400 8202
rect 9208 8008 9344 8188
rect 9536 8192 9592 8202
rect 9400 8008 9536 8188
rect 8588 7996 9592 8008
rect 7604 7982 8588 7992
rect 5980 7890 6036 7900
rect 6228 7904 6364 7916
rect 6172 7890 6228 7900
rect 6420 7904 6556 7916
rect 6364 7890 6420 7900
rect 6612 7904 6748 7916
rect 6556 7890 6612 7900
rect 6804 7904 6940 7916
rect 6748 7890 6804 7900
rect 6996 7904 7200 7916
rect 10800 7928 11300 7938
rect 6940 7890 6996 7900
rect 5308 7858 5364 7866
rect 5500 7858 5556 7866
rect 5692 7858 5748 7866
rect 5884 7858 5940 7866
rect 6076 7858 6132 7866
rect 5076 7856 6132 7858
rect 6268 7856 6324 7866
rect 6460 7856 6516 7866
rect 6652 7856 6708 7866
rect 6844 7856 6900 7866
rect 7036 7856 7092 7866
rect 5076 7848 5116 7856
rect 5172 7848 5308 7856
rect 5364 7848 5500 7856
rect 5556 7848 5692 7856
rect 5748 7848 5884 7856
rect 5940 7848 6076 7856
rect 5076 7600 5104 7848
rect 6132 7676 6268 7856
rect 6324 7676 6460 7856
rect 6516 7676 6652 7856
rect 6708 7676 6844 7856
rect 6900 7676 7036 7856
rect 7092 7676 7096 7856
rect 8764 7820 9636 7830
rect 6080 7600 7096 7676
rect 7708 7792 8764 7804
rect 7708 7612 7712 7792
rect 5076 7584 7096 7600
rect 7768 7612 7904 7792
rect 7712 7598 7768 7608
rect 7960 7612 8096 7792
rect 7904 7598 7960 7608
rect 8152 7612 8288 7792
rect 8096 7598 8152 7608
rect 8344 7612 8480 7792
rect 8288 7598 8344 7608
rect 8536 7612 8672 7792
rect 8480 7598 8536 7608
rect 8728 7620 8764 7792
rect 8728 7612 8864 7620
rect 8764 7610 8864 7612
rect 8672 7598 8728 7608
rect 8920 7610 9056 7620
rect 8864 7598 8920 7608
rect 9112 7610 9248 7620
rect 9056 7598 9112 7608
rect 9304 7610 9440 7620
rect 9248 7598 9304 7608
rect 9496 7610 9636 7620
rect 9440 7598 9496 7608
rect 5136 7572 5364 7584
rect 7616 7572 7672 7582
rect 7612 7566 7616 7568
rect 7608 7556 7616 7566
rect 7808 7572 7864 7582
rect 7672 7556 7808 7568
rect 8000 7572 8056 7582
rect 7864 7556 8000 7568
rect 8192 7572 8248 7582
rect 8056 7556 8192 7568
rect 8384 7572 8440 7582
rect 8248 7556 8384 7568
rect 8576 7572 8632 7582
rect 8440 7556 8576 7568
rect 8768 7572 8824 7582
rect 1764 7124 4928 7180
rect 1776 7092 4928 7124
rect 1828 6920 1968 7092
rect 1776 6902 1828 6912
rect 2020 6920 2160 7092
rect 1968 6902 2020 6912
rect 2212 6920 2352 7092
rect 2160 6902 2212 6912
rect 2404 6920 2544 7092
rect 2352 6902 2404 6912
rect 2596 6920 2736 7092
rect 2544 6902 2596 6912
rect 2788 6920 2928 7092
rect 2736 6902 2788 6912
rect 2980 6920 3120 7092
rect 2928 6902 2980 6912
rect 3172 6920 3312 7092
rect 3120 6902 3172 6912
rect 3364 6920 3504 7092
rect 3312 6902 3364 6912
rect 3556 7012 4928 7092
rect 3556 6920 3740 7012
rect 3504 6902 3556 6912
rect 988 6868 1732 6878
rect 988 6688 1680 6868
rect 1872 6868 1924 6878
rect 1732 6688 1872 6860
rect 2064 6868 2116 6878
rect 1924 6688 2064 6860
rect 2256 6868 2308 6878
rect 2116 6688 2256 6860
rect 2448 6868 2500 6878
rect 2308 6688 2448 6860
rect 2640 6868 2692 6878
rect 2500 6688 2640 6860
rect 2832 6868 2884 6878
rect 2692 6688 2832 6860
rect 3024 6868 3076 6878
rect 2884 6688 3024 6860
rect 3216 6868 3268 6878
rect 3076 6688 3216 6860
rect 3408 6868 3460 6878
rect 3268 6688 3408 6860
rect 3600 6868 3652 6878
rect 3460 6688 3600 6860
rect 3800 6928 4928 7012
rect 6384 7512 7076 7522
rect 8632 7388 8768 7568
rect 8960 7572 9016 7582
rect 8824 7388 8960 7568
rect 9152 7572 9208 7582
rect 9016 7388 9152 7568
rect 9344 7572 9400 7582
rect 9208 7388 9344 7568
rect 9536 7572 9592 7582
rect 9400 7388 9536 7568
rect 8592 7376 9592 7388
rect 10580 7472 10800 7600
rect 15388 7652 16020 8240
rect 16176 8162 16472 8164
rect 16164 8152 16472 8162
rect 16456 8088 16472 8152
rect 16164 8060 16472 8088
rect 16176 7936 16472 8060
rect 16940 8152 17260 8162
rect 16940 8078 17260 8088
rect 17876 8152 18168 8162
rect 18168 8092 18176 8144
rect 17876 8082 18176 8092
rect 16940 8000 17236 8078
rect 17880 8000 18176 8082
rect 18524 8000 19328 8356
rect 16940 7936 19328 8000
rect 16176 7912 19328 7936
rect 16228 7740 16368 7912
rect 16176 7722 16228 7732
rect 16420 7740 16560 7912
rect 16368 7722 16420 7732
rect 16612 7740 16752 7912
rect 16560 7722 16612 7732
rect 16804 7740 16944 7912
rect 16752 7722 16804 7732
rect 16996 7740 17136 7912
rect 16944 7722 16996 7732
rect 17188 7740 17328 7912
rect 17136 7722 17188 7732
rect 17380 7740 17520 7912
rect 17328 7722 17380 7732
rect 17572 7740 17712 7912
rect 17520 7722 17572 7732
rect 17764 7740 17904 7912
rect 17712 7722 17764 7732
rect 17956 7824 19328 7912
rect 17956 7740 18140 7824
rect 17904 7722 17956 7732
rect 16080 7688 16132 7698
rect 11300 7472 12028 7580
rect 7608 7358 8592 7368
rect 8764 7204 9636 7214
rect 6384 6990 7076 7000
rect 7708 7176 8764 7188
rect 7708 6996 7712 7176
rect 7768 6996 7904 7176
rect 7712 6982 7768 6992
rect 7960 6996 8096 7176
rect 7904 6982 7960 6992
rect 8152 6996 8288 7176
rect 8096 6982 8152 6992
rect 8344 6996 8480 7176
rect 8288 6982 8344 6992
rect 8536 6996 8672 7176
rect 8480 6982 8536 6992
rect 8728 7004 8764 7176
rect 8728 6996 8864 7004
rect 8764 6994 8864 6996
rect 8672 6982 8728 6992
rect 8920 6994 9056 7004
rect 8864 6982 8920 6992
rect 9112 6994 9248 7004
rect 9056 6982 9112 6992
rect 9304 6994 9440 7004
rect 9248 6982 9304 6992
rect 9496 6994 9636 7004
rect 9440 6982 9496 6992
rect 7616 6956 7672 6966
rect 7608 6944 7616 6954
rect 7808 6956 7864 6966
rect 7672 6944 7808 6954
rect 8000 6956 8056 6966
rect 7864 6944 8000 6954
rect 8192 6956 8248 6966
rect 8056 6944 8192 6954
rect 8384 6956 8440 6966
rect 8248 6944 8384 6954
rect 8576 6956 8632 6966
rect 8440 6944 8576 6954
rect 8768 6956 8824 6966
rect 7000 6928 7528 6938
rect 3800 6920 7000 6928
rect 3740 6746 3800 6756
rect 988 6600 3652 6688
rect 4124 6600 7000 6920
rect 8632 6772 8768 6952
rect 8960 6956 9016 6966
rect 8824 6772 8960 6952
rect 9152 6956 9208 6966
rect 9016 6772 9152 6952
rect 9344 6956 9400 6966
rect 9208 6772 9344 6952
rect 9536 6956 9592 6966
rect 9400 6772 9536 6952
rect 8592 6760 9592 6772
rect 7608 6746 8592 6756
rect 4124 6590 7528 6600
rect 1672 6516 1964 6526
rect -9972 6164 -8460 6256
rect -9972 6156 -8992 6164
rect -9972 5988 -9964 6156
rect -9912 5976 -9772 6156
rect -9720 5976 -9580 6156
rect -9528 5976 -9388 6156
rect -9336 5976 -9196 6156
rect -9144 5988 -8992 6156
rect -8824 5988 -8460 6164
rect -3092 6456 1672 6468
rect 2540 6516 2832 6526
rect 1964 6456 2540 6468
rect 3476 6512 3768 6522
rect 2832 6456 3476 6468
rect -3092 6452 3476 6456
rect 4124 6482 7204 6590
rect 8764 6588 9636 6598
rect 7708 6556 8764 6568
rect 4124 6472 7456 6482
rect 4124 6468 6960 6472
rect 3768 6452 6960 6468
rect -3092 6156 6960 6452
rect 7708 6376 7712 6556
rect 7768 6376 7904 6556
rect 7712 6362 7768 6372
rect 7960 6376 8096 6556
rect 7904 6362 7960 6372
rect 8152 6376 8288 6556
rect 8096 6362 8152 6372
rect 8344 6376 8480 6556
rect 8288 6362 8344 6372
rect 8536 6376 8672 6556
rect 8480 6362 8536 6372
rect 8728 6388 8764 6556
rect 8728 6376 8864 6388
rect 8672 6362 8728 6372
rect 8920 6376 9056 6388
rect 8864 6362 8920 6372
rect 9112 6376 9248 6388
rect 9056 6362 9112 6372
rect 9304 6376 9440 6388
rect 9248 6362 9304 6372
rect 9496 6378 9636 6388
rect 10580 6468 12028 7472
rect 15388 7508 16080 7652
rect 16272 7688 16324 7698
rect 16132 7508 16272 7652
rect 16464 7688 16516 7698
rect 16324 7508 16464 7680
rect 16656 7688 16708 7698
rect 16516 7508 16656 7680
rect 16848 7688 16900 7698
rect 16708 7508 16848 7680
rect 17040 7688 17092 7698
rect 16900 7508 17040 7680
rect 17232 7688 17284 7698
rect 17092 7508 17232 7680
rect 17424 7688 17476 7698
rect 17284 7508 17424 7680
rect 17616 7688 17668 7698
rect 17476 7508 17616 7680
rect 17808 7688 17860 7698
rect 17668 7508 17808 7680
rect 18000 7688 18052 7698
rect 17860 7508 18000 7680
rect 18200 7740 19328 7824
rect 18140 7558 18200 7568
rect 15388 7420 18052 7508
rect 15388 6878 16088 7420
rect 16164 7328 16456 7338
rect 16936 7328 17228 7338
rect 16456 7268 16460 7316
rect 16164 7180 16460 7268
rect 17876 7328 18168 7338
rect 17228 7268 17232 7320
rect 16936 7180 17232 7268
rect 18168 7268 18172 7292
rect 17876 7180 18172 7268
rect 18524 7180 19328 7740
rect 19476 8224 19504 8472
rect 20532 8296 20668 8472
rect 20860 8476 20916 8486
rect 20724 8296 20860 8472
rect 21052 8476 21108 8486
rect 20916 8296 21052 8472
rect 21244 8476 21300 8486
rect 21108 8296 21244 8472
rect 21436 8476 21492 8486
rect 21300 8296 21436 8472
rect 23164 8440 24036 8450
rect 20480 8224 21492 8296
rect 22108 8412 23164 8424
rect 22108 8232 22112 8412
rect 19476 8212 21492 8224
rect 22168 8232 22304 8412
rect 22112 8218 22168 8228
rect 22360 8232 22496 8412
rect 22304 8218 22360 8228
rect 22552 8232 22688 8412
rect 22496 8218 22552 8228
rect 22744 8232 22880 8412
rect 22688 8218 22744 8228
rect 22936 8232 23072 8412
rect 22880 8218 22936 8228
rect 23128 8240 23164 8412
rect 23128 8232 23264 8240
rect 23164 8230 23264 8232
rect 23072 8218 23128 8228
rect 23320 8230 23456 8240
rect 23264 8218 23320 8228
rect 23512 8230 23648 8240
rect 23456 8218 23512 8228
rect 23704 8230 23840 8240
rect 23648 8218 23704 8228
rect 23896 8230 24036 8240
rect 23840 8218 23896 8228
rect 19476 7858 19576 8212
rect 22016 8192 22072 8202
rect 22004 8180 22016 8190
rect 22208 8192 22264 8202
rect 22072 8180 22208 8190
rect 22400 8192 22456 8202
rect 22264 8180 22400 8190
rect 22592 8192 22648 8202
rect 22456 8180 22592 8190
rect 22784 8192 22840 8202
rect 22648 8180 22784 8190
rect 22976 8192 23032 8202
rect 22840 8180 22976 8190
rect 23168 8192 23224 8202
rect 19608 8164 21600 8176
rect 19608 8080 20624 8164
rect 19608 7904 19612 8080
rect 19668 7904 19804 8080
rect 19612 7890 19668 7900
rect 19860 7904 19996 8080
rect 19804 7890 19860 7900
rect 20052 7904 20188 8080
rect 19996 7890 20052 7900
rect 20244 7904 20380 8080
rect 20188 7890 20244 7900
rect 20436 7904 20572 8080
rect 23032 8008 23168 8188
rect 23360 8192 23416 8202
rect 23224 8008 23360 8188
rect 23552 8192 23608 8202
rect 23416 8008 23552 8188
rect 23744 8192 23800 8202
rect 23608 8008 23744 8188
rect 23936 8192 23992 8202
rect 23800 8008 23936 8188
rect 22988 7996 23992 8008
rect 22004 7982 22988 7992
rect 20380 7890 20436 7900
rect 20628 7904 20764 7916
rect 20572 7890 20628 7900
rect 20820 7904 20956 7916
rect 20764 7890 20820 7900
rect 21012 7904 21148 7916
rect 20956 7890 21012 7900
rect 21204 7904 21340 7916
rect 21148 7890 21204 7900
rect 21396 7904 21600 7916
rect 21340 7890 21396 7900
rect 19708 7858 19764 7866
rect 19900 7858 19956 7866
rect 20092 7858 20148 7866
rect 20284 7858 20340 7866
rect 20476 7858 20532 7866
rect 19476 7856 20532 7858
rect 20668 7856 20724 7866
rect 20860 7856 20916 7866
rect 21052 7856 21108 7866
rect 21244 7856 21300 7866
rect 21436 7856 21492 7866
rect 19476 7848 19516 7856
rect 19572 7848 19708 7856
rect 19764 7848 19900 7856
rect 19956 7848 20092 7856
rect 20148 7848 20284 7856
rect 20340 7848 20476 7856
rect 19476 7600 19504 7848
rect 20532 7676 20668 7856
rect 20724 7676 20860 7856
rect 20916 7676 21052 7856
rect 21108 7676 21244 7856
rect 21300 7676 21436 7856
rect 21492 7676 21496 7856
rect 23164 7820 24036 7830
rect 20480 7600 21496 7676
rect 22108 7792 23164 7804
rect 22108 7612 22112 7792
rect 19476 7584 21496 7600
rect 22168 7612 22304 7792
rect 22112 7598 22168 7608
rect 22360 7612 22496 7792
rect 22304 7598 22360 7608
rect 22552 7612 22688 7792
rect 22496 7598 22552 7608
rect 22744 7612 22880 7792
rect 22688 7598 22744 7608
rect 22936 7612 23072 7792
rect 22880 7598 22936 7608
rect 23128 7620 23164 7792
rect 23128 7612 23264 7620
rect 23164 7610 23264 7612
rect 23072 7598 23128 7608
rect 23320 7610 23456 7620
rect 23264 7598 23320 7608
rect 23512 7610 23648 7620
rect 23456 7598 23512 7608
rect 23704 7610 23840 7620
rect 23648 7598 23704 7608
rect 23896 7610 24036 7620
rect 23840 7598 23896 7608
rect 19536 7572 19764 7584
rect 22016 7572 22072 7582
rect 22012 7566 22016 7568
rect 22008 7556 22016 7566
rect 22208 7572 22264 7582
rect 22072 7556 22208 7568
rect 22400 7572 22456 7582
rect 22264 7556 22400 7568
rect 22592 7572 22648 7582
rect 22456 7556 22592 7568
rect 22784 7572 22840 7582
rect 22648 7556 22784 7568
rect 22976 7572 23032 7582
rect 22840 7556 22976 7568
rect 23168 7572 23224 7582
rect 16164 7124 19328 7180
rect 16176 7092 19328 7124
rect 16228 6920 16368 7092
rect 16176 6902 16228 6912
rect 16420 6920 16560 7092
rect 16368 6902 16420 6912
rect 16612 6920 16752 7092
rect 16560 6902 16612 6912
rect 16804 6920 16944 7092
rect 16752 6902 16804 6912
rect 16996 6920 17136 7092
rect 16944 6902 16996 6912
rect 17188 6920 17328 7092
rect 17136 6902 17188 6912
rect 17380 6920 17520 7092
rect 17328 6902 17380 6912
rect 17572 6920 17712 7092
rect 17520 6902 17572 6912
rect 17764 6920 17904 7092
rect 17712 6902 17764 6912
rect 17956 7012 19328 7092
rect 17956 6920 18140 7012
rect 17904 6902 17956 6912
rect 15388 6868 16132 6878
rect 15388 6688 16080 6868
rect 16272 6868 16324 6878
rect 16132 6688 16272 6860
rect 16464 6868 16516 6878
rect 16324 6688 16464 6860
rect 16656 6868 16708 6878
rect 16516 6688 16656 6860
rect 16848 6868 16900 6878
rect 16708 6688 16848 6860
rect 17040 6868 17092 6878
rect 16900 6688 17040 6860
rect 17232 6868 17284 6878
rect 17092 6688 17232 6860
rect 17424 6868 17476 6878
rect 17284 6688 17424 6860
rect 17616 6868 17668 6878
rect 17476 6688 17616 6860
rect 17808 6868 17860 6878
rect 17668 6688 17808 6860
rect 18000 6868 18052 6878
rect 17860 6688 18000 6860
rect 18200 6928 19328 7012
rect 20784 7512 21476 7522
rect 23032 7388 23168 7568
rect 23360 7572 23416 7582
rect 23224 7388 23360 7568
rect 23552 7572 23608 7582
rect 23416 7388 23552 7568
rect 23744 7572 23800 7582
rect 23608 7388 23744 7568
rect 23936 7572 23992 7582
rect 23800 7388 23936 7568
rect 22992 7376 23992 7388
rect 22008 7358 22992 7368
rect 23164 7204 24036 7214
rect 20784 6990 21476 7000
rect 22108 7176 23164 7188
rect 22108 6996 22112 7176
rect 22168 6996 22304 7176
rect 22112 6982 22168 6992
rect 22360 6996 22496 7176
rect 22304 6982 22360 6992
rect 22552 6996 22688 7176
rect 22496 6982 22552 6992
rect 22744 6996 22880 7176
rect 22688 6982 22744 6992
rect 22936 6996 23072 7176
rect 22880 6982 22936 6992
rect 23128 7004 23164 7176
rect 23128 6996 23264 7004
rect 23164 6994 23264 6996
rect 23072 6982 23128 6992
rect 23320 6994 23456 7004
rect 23264 6982 23320 6992
rect 23512 6994 23648 7004
rect 23456 6982 23512 6992
rect 23704 6994 23840 7004
rect 23648 6982 23704 6992
rect 23896 6994 24036 7004
rect 23840 6982 23896 6992
rect 22016 6956 22072 6966
rect 22008 6944 22016 6954
rect 22208 6956 22264 6966
rect 22072 6944 22208 6954
rect 22400 6956 22456 6966
rect 22264 6944 22400 6954
rect 22592 6956 22648 6966
rect 22456 6944 22592 6954
rect 22784 6956 22840 6966
rect 22648 6944 22784 6954
rect 22976 6956 23032 6966
rect 22840 6944 22976 6954
rect 23168 6956 23224 6966
rect 21400 6928 21928 6938
rect 18200 6920 21400 6928
rect 18140 6746 18200 6756
rect 15388 6600 18052 6688
rect 18524 6600 21400 6920
rect 23032 6772 23168 6952
rect 23360 6956 23416 6966
rect 23224 6772 23360 6952
rect 23552 6956 23608 6966
rect 23416 6772 23552 6952
rect 23744 6956 23800 6966
rect 23608 6772 23744 6952
rect 23936 6956 23992 6966
rect 23800 6772 23936 6952
rect 22992 6760 23992 6772
rect 22008 6746 22992 6756
rect 18524 6590 21928 6600
rect 16072 6516 16364 6526
rect 10580 6456 16072 6468
rect 16940 6516 17232 6526
rect 16364 6456 16940 6468
rect 17876 6512 18168 6522
rect 17232 6456 17876 6468
rect 10580 6452 17876 6456
rect 18524 6482 21604 6590
rect 23164 6588 24036 6598
rect 22108 6556 23164 6568
rect 18524 6472 21856 6482
rect 18524 6468 21360 6472
rect 18168 6452 21360 6468
rect 9496 6376 9500 6378
rect 9440 6362 9496 6372
rect 7616 6336 7672 6346
rect 7612 6330 7616 6332
rect -3092 6146 7456 6156
rect 7604 6320 7616 6330
rect 7808 6336 7864 6346
rect 7672 6320 7808 6332
rect 8000 6336 8056 6346
rect 7864 6320 8000 6332
rect 8192 6336 8248 6346
rect 8056 6320 8192 6332
rect 8384 6336 8440 6346
rect 8248 6320 8384 6332
rect 8576 6336 8632 6346
rect 8440 6320 8576 6332
rect 8768 6336 8824 6346
rect 8632 6152 8768 6332
rect 8960 6336 9016 6346
rect 8824 6152 8960 6332
rect 9152 6336 9208 6346
rect 9016 6152 9152 6332
rect 9344 6336 9400 6346
rect 9208 6152 9344 6332
rect 9536 6336 9592 6346
rect 9400 6152 9536 6332
rect -3092 6084 6972 6146
rect 8588 6140 9592 6152
rect 10580 6156 21360 6452
rect 22108 6376 22112 6556
rect 22168 6376 22304 6556
rect 22112 6362 22168 6372
rect 22360 6376 22496 6556
rect 22304 6362 22360 6372
rect 22552 6376 22688 6556
rect 22496 6362 22552 6372
rect 22744 6376 22880 6556
rect 22688 6362 22744 6372
rect 22936 6376 23072 6556
rect 22880 6362 22936 6372
rect 23128 6388 23164 6556
rect 23128 6376 23264 6388
rect 23072 6362 23128 6372
rect 23320 6376 23456 6388
rect 23264 6362 23320 6372
rect 23512 6376 23648 6388
rect 23456 6362 23512 6372
rect 23704 6376 23840 6388
rect 23648 6362 23704 6372
rect 23896 6378 24036 6388
rect 23896 6376 23900 6378
rect 23840 6362 23896 6372
rect 22016 6336 22072 6346
rect 22012 6330 22016 6332
rect 10580 6146 21856 6156
rect 22004 6320 22016 6330
rect 22208 6336 22264 6346
rect 22072 6320 22208 6332
rect 22400 6336 22456 6346
rect 22264 6320 22400 6332
rect 22592 6336 22648 6346
rect 22456 6320 22592 6332
rect 22784 6336 22840 6346
rect 22648 6320 22784 6332
rect 22976 6336 23032 6346
rect 22840 6320 22976 6332
rect 23168 6336 23224 6346
rect 23032 6152 23168 6332
rect 23360 6336 23416 6346
rect 23224 6152 23360 6332
rect 23552 6336 23608 6346
rect 23416 6152 23552 6332
rect 23744 6336 23800 6346
rect 23608 6152 23744 6332
rect 23936 6336 23992 6346
rect 23800 6152 23936 6332
rect 10580 6140 21372 6146
rect 7604 6122 8588 6132
rect 11130 6130 21372 6140
rect 7088 6084 7372 6090
rect -3092 6080 7372 6084
rect -3092 6052 7088 6080
rect -3092 5996 5172 6052
rect -9144 5976 -8704 5988
rect -9964 5966 -9912 5976
rect -9772 5966 -9720 5976
rect -9580 5966 -9528 5976
rect -9388 5966 -9336 5976
rect -9196 5966 -9144 5976
rect -10060 5934 -10008 5942
rect -9868 5934 -9816 5942
rect -9676 5934 -9624 5942
rect -9484 5934 -9432 5942
rect -10064 5932 -9432 5934
rect -9292 5932 -9240 5942
rect -9100 5932 -9048 5942
rect -10064 5924 -10060 5932
rect -10008 5924 -9868 5932
rect -9816 5924 -9676 5932
rect -9624 5924 -9484 5932
rect -9432 5752 -9292 5932
rect -9240 5752 -9100 5932
rect -9460 5744 -9048 5752
rect -9460 5742 -9432 5744
rect -9292 5742 -9240 5744
rect -9100 5742 -9048 5744
rect -10064 5730 -9460 5740
rect -9964 5548 -9144 5552
rect -9016 5548 -8704 5976
rect 312 5884 1132 5888
rect 1260 5884 1572 5996
rect 312 5876 1572 5884
rect 364 5696 504 5876
rect 556 5696 696 5876
rect 748 5696 888 5876
rect 940 5696 1080 5876
rect 1132 5696 1572 5876
rect 312 5686 364 5696
rect 504 5686 556 5696
rect 696 5686 748 5696
rect 888 5686 940 5696
rect 1080 5686 1132 5696
rect 216 5654 268 5662
rect 408 5654 460 5662
rect 600 5654 652 5662
rect 792 5654 844 5662
rect -9964 5540 -8704 5548
rect -9912 5360 -9772 5540
rect -9720 5360 -9580 5540
rect -9528 5360 -9388 5540
rect -9336 5360 -9196 5540
rect -9144 5360 -8704 5540
rect 212 5652 844 5654
rect 984 5652 1036 5662
rect 1176 5652 1228 5662
rect 212 5644 216 5652
rect 268 5644 408 5652
rect 460 5644 600 5652
rect 652 5644 792 5652
rect 844 5472 984 5652
rect 1036 5472 1176 5652
rect 816 5464 1228 5472
rect 816 5462 844 5464
rect 984 5462 1036 5464
rect 1176 5462 1228 5464
rect 212 5450 816 5460
rect -9964 5350 -9912 5360
rect -9772 5350 -9720 5360
rect -9580 5350 -9528 5360
rect -9388 5350 -9336 5360
rect -9196 5350 -9144 5360
rect -10060 5318 -10008 5326
rect -9868 5318 -9816 5326
rect -9676 5318 -9624 5326
rect -9484 5318 -9432 5326
rect -10064 5316 -9432 5318
rect -9292 5316 -9240 5326
rect -9100 5316 -9048 5326
rect -10064 5308 -10060 5316
rect -10008 5308 -9868 5316
rect -9816 5308 -9676 5316
rect -9624 5308 -9484 5316
rect -9432 5136 -9292 5316
rect -9240 5136 -9100 5316
rect -9460 5128 -9048 5136
rect -9460 5126 -9432 5128
rect -9292 5126 -9240 5128
rect -9100 5126 -9048 5128
rect -10064 5114 -9460 5124
rect -9964 4924 -9912 4930
rect -9772 4924 -9720 4930
rect -9580 4924 -9528 4930
rect -9388 4924 -9336 4930
rect -9196 4924 -9144 4930
rect -9016 4924 -8704 5360
rect 312 5268 1132 5272
rect 1260 5268 1572 5696
rect 2112 5884 2932 5888
rect 3060 5884 3372 5996
rect 2112 5876 3372 5884
rect 2164 5696 2304 5876
rect 2356 5696 2496 5876
rect 2548 5696 2688 5876
rect 2740 5696 2880 5876
rect 2932 5696 3372 5876
rect 2112 5686 2164 5696
rect 2304 5686 2356 5696
rect 2496 5686 2548 5696
rect 2688 5686 2740 5696
rect 2880 5686 2932 5696
rect 2016 5654 2068 5662
rect 2208 5654 2260 5662
rect 2400 5654 2452 5662
rect 2592 5654 2644 5662
rect 2012 5652 2644 5654
rect 2784 5652 2836 5662
rect 2976 5652 3028 5662
rect 2012 5644 2016 5652
rect 2068 5644 2208 5652
rect 2260 5644 2400 5652
rect 2452 5644 2592 5652
rect 2644 5472 2784 5652
rect 2836 5472 2976 5652
rect 2616 5464 3028 5472
rect 2616 5462 2644 5464
rect 2784 5462 2836 5464
rect 2976 5462 3028 5464
rect 2012 5450 2616 5460
rect 312 5260 1572 5268
rect -9964 4920 -8704 4924
rect -9912 4740 -9772 4920
rect -9720 4740 -9580 4920
rect -9528 4740 -9388 4920
rect -9336 4740 -9196 4920
rect -9144 4740 -8704 4920
rect -404 5092 28 5102
rect -9964 4736 -8704 4740
rect -808 4816 -404 4826
rect 364 5080 504 5260
rect 556 5080 696 5260
rect 748 5080 888 5260
rect 940 5080 1080 5260
rect 1132 5080 1572 5260
rect 312 5070 364 5080
rect 504 5070 556 5080
rect 696 5070 748 5080
rect 888 5070 940 5080
rect 1080 5070 1132 5080
rect 216 5038 268 5046
rect 408 5038 460 5046
rect 600 5038 652 5046
rect 792 5038 844 5046
rect 212 5036 844 5038
rect 984 5036 1036 5046
rect 1176 5036 1228 5046
rect 212 5028 216 5036
rect 268 5028 408 5036
rect 460 5028 600 5036
rect 652 5028 792 5036
rect 844 4856 984 5036
rect 1036 4856 1176 5036
rect 816 4848 1228 4856
rect 816 4846 844 4848
rect 984 4846 1036 4848
rect 1176 4846 1228 4848
rect 212 4834 816 4844
rect -9964 4730 -9912 4736
rect -9772 4730 -9720 4736
rect -9580 4730 -9528 4736
rect -9388 4730 -9336 4736
rect -9196 4730 -9144 4736
rect -10060 4698 -10008 4706
rect -9868 4698 -9816 4706
rect -9676 4698 -9624 4706
rect -9484 4698 -9432 4706
rect -10068 4696 -9432 4698
rect -9292 4696 -9240 4706
rect -9100 4696 -9048 4706
rect -10068 4688 -10060 4696
rect -10008 4688 -9868 4696
rect -9816 4688 -9676 4696
rect -9624 4688 -9484 4696
rect -9432 4516 -9292 4696
rect -9240 4516 -9100 4696
rect -9464 4508 -9048 4516
rect -9464 4506 -9432 4508
rect -9292 4506 -9240 4508
rect -9100 4506 -9048 4508
rect -3172 4532 -3028 4542
rect -10068 4494 -9464 4504
rect -3172 4410 -3028 4420
rect 312 4644 364 4650
rect 504 4644 556 4650
rect 696 4644 748 4650
rect 888 4644 940 4650
rect 1080 4644 1132 4650
rect 1260 4644 1572 5080
rect 2112 5268 2932 5272
rect 3060 5268 3372 5696
rect 3912 5884 4732 5888
rect 4860 5884 5172 5996
rect 3912 5876 5172 5884
rect 3964 5696 4104 5876
rect 4156 5696 4296 5876
rect 4348 5696 4488 5876
rect 4540 5696 4680 5876
rect 4732 5696 5172 5876
rect 3912 5686 3964 5696
rect 4104 5686 4156 5696
rect 4296 5686 4348 5696
rect 4488 5686 4540 5696
rect 4680 5686 4732 5696
rect 3816 5654 3868 5662
rect 4008 5654 4060 5662
rect 4200 5654 4252 5662
rect 4392 5654 4444 5662
rect 3812 5652 4444 5654
rect 4584 5652 4636 5662
rect 4776 5652 4828 5662
rect 3812 5644 3816 5652
rect 3868 5644 4008 5652
rect 4060 5644 4200 5652
rect 4252 5644 4392 5652
rect 4444 5472 4584 5652
rect 4636 5472 4776 5652
rect 4416 5464 4828 5472
rect 4416 5462 4444 5464
rect 4584 5462 4636 5464
rect 4776 5462 4828 5464
rect 3812 5450 4416 5460
rect 2112 5260 3372 5268
rect 2164 5080 2304 5260
rect 2356 5080 2496 5260
rect 2548 5080 2688 5260
rect 2740 5080 2880 5260
rect 2932 5080 3372 5260
rect 2112 5070 2164 5080
rect 2304 5070 2356 5080
rect 2496 5070 2548 5080
rect 2688 5070 2740 5080
rect 2880 5070 2932 5080
rect 2016 5038 2068 5046
rect 2208 5038 2260 5046
rect 2400 5038 2452 5046
rect 2592 5038 2644 5046
rect 2012 5036 2644 5038
rect 2784 5036 2836 5046
rect 2976 5036 3028 5046
rect 2012 5028 2016 5036
rect 2068 5028 2208 5036
rect 2260 5028 2400 5036
rect 2452 5028 2592 5036
rect 2644 4856 2784 5036
rect 2836 4856 2976 5036
rect 2616 4848 3028 4856
rect 2616 4846 2644 4848
rect 2784 4846 2836 4848
rect 2976 4846 3028 4848
rect 2012 4834 2616 4844
rect 312 4640 1572 4644
rect 364 4460 504 4640
rect 556 4460 696 4640
rect 748 4460 888 4640
rect 940 4460 1080 4640
rect 1132 4460 1572 4640
rect 312 4456 1572 4460
rect 2112 4644 2164 4650
rect 2304 4644 2356 4650
rect 2496 4644 2548 4650
rect 2688 4644 2740 4650
rect 2880 4644 2932 4650
rect 3060 4644 3372 5080
rect 3912 5268 4732 5272
rect 4860 5268 5172 5696
rect 5712 5884 6532 5888
rect 6660 5884 7088 6052
rect 5712 5876 7088 5884
rect 5764 5696 5904 5876
rect 5956 5696 6096 5876
rect 6148 5696 6288 5876
rect 6340 5696 6480 5876
rect 6532 5696 7088 5876
rect 5712 5686 5764 5696
rect 5904 5686 5956 5696
rect 6096 5686 6148 5696
rect 6288 5686 6340 5696
rect 6480 5686 6532 5696
rect 5616 5654 5668 5662
rect 5808 5654 5860 5662
rect 6000 5654 6052 5662
rect 6192 5654 6244 5662
rect 5612 5652 6244 5654
rect 6384 5652 6436 5662
rect 6576 5652 6628 5662
rect 5612 5644 5616 5652
rect 5668 5644 5808 5652
rect 5860 5644 6000 5652
rect 6052 5644 6192 5652
rect 6244 5472 6384 5652
rect 6436 5472 6576 5652
rect 6216 5464 6628 5472
rect 6216 5462 6244 5464
rect 6384 5462 6436 5464
rect 6576 5462 6628 5464
rect 6660 5584 7088 5696
rect 5612 5450 6216 5460
rect 3912 5260 5172 5268
rect 3964 5080 4104 5260
rect 4156 5080 4296 5260
rect 4348 5080 4488 5260
rect 4540 5080 4680 5260
rect 4732 5080 5172 5260
rect 3912 5070 3964 5080
rect 4104 5070 4156 5080
rect 4296 5070 4348 5080
rect 4488 5070 4540 5080
rect 4680 5070 4732 5080
rect 3816 5038 3868 5046
rect 4008 5038 4060 5046
rect 4200 5038 4252 5046
rect 4392 5038 4444 5046
rect 3812 5036 4444 5038
rect 4584 5036 4636 5046
rect 4776 5036 4828 5046
rect 3812 5028 3816 5036
rect 3868 5028 4008 5036
rect 4060 5028 4200 5036
rect 4252 5028 4392 5036
rect 4444 4856 4584 5036
rect 4636 4856 4776 5036
rect 4416 4848 4828 4856
rect 4416 4846 4444 4848
rect 4584 4846 4636 4848
rect 4776 4846 4828 4848
rect 3812 4834 4416 4844
rect 2112 4640 3372 4644
rect 2164 4460 2304 4640
rect 2356 4460 2496 4640
rect 2548 4460 2688 4640
rect 2740 4460 2880 4640
rect 2932 4460 3372 4640
rect 2112 4456 3372 4460
rect 3912 4644 3964 4650
rect 4104 4644 4156 4650
rect 4296 4644 4348 4650
rect 4488 4644 4540 4650
rect 4680 4644 4732 4650
rect 4860 4644 5172 5080
rect 5712 5268 6532 5272
rect 6660 5268 6972 5584
rect 11308 6084 21372 6130
rect 22988 6140 23992 6152
rect 22004 6122 22988 6132
rect 21488 6084 21772 6090
rect 11308 6080 21772 6084
rect 11308 6052 21488 6080
rect 11308 5996 19572 6052
rect 8760 5968 9632 5978
rect 7708 5940 8760 5952
rect 7708 5760 7712 5940
rect 7768 5760 7904 5940
rect 7712 5746 7768 5756
rect 7960 5760 8096 5940
rect 7904 5746 7960 5756
rect 8152 5760 8288 5940
rect 8096 5746 8152 5756
rect 8344 5760 8480 5940
rect 8288 5746 8344 5756
rect 8536 5760 8672 5940
rect 8480 5746 8536 5756
rect 8728 5768 8760 5940
rect 8728 5760 8864 5768
rect 8760 5758 8864 5760
rect 8672 5746 8728 5756
rect 8920 5758 9056 5768
rect 8864 5746 8920 5756
rect 9112 5758 9248 5768
rect 9056 5746 9112 5756
rect 9304 5758 9440 5768
rect 9248 5746 9304 5756
rect 9496 5758 9632 5768
rect 14712 5884 15532 5888
rect 15660 5884 15972 5996
rect 14712 5876 15972 5884
rect 9440 5746 9496 5756
rect 7616 5720 7672 5730
rect 7088 5570 7372 5580
rect 7604 5708 7616 5718
rect 7808 5720 7864 5730
rect 7672 5708 7808 5718
rect 8000 5720 8056 5730
rect 7864 5708 8000 5718
rect 8192 5720 8248 5730
rect 8056 5708 8192 5718
rect 8384 5720 8440 5730
rect 8248 5708 8384 5718
rect 8576 5720 8632 5730
rect 8440 5708 8576 5718
rect 8768 5720 8824 5730
rect 8632 5536 8768 5716
rect 8960 5720 9016 5730
rect 8824 5536 8960 5716
rect 9152 5720 9208 5730
rect 9016 5536 9152 5716
rect 9344 5720 9400 5730
rect 9208 5536 9344 5716
rect 9536 5720 9592 5730
rect 9400 5536 9536 5716
rect 14764 5696 14904 5876
rect 14956 5696 15096 5876
rect 15148 5696 15288 5876
rect 15340 5696 15480 5876
rect 15532 5696 15972 5876
rect 14712 5686 14764 5696
rect 14904 5686 14956 5696
rect 15096 5686 15148 5696
rect 15288 5686 15340 5696
rect 15480 5686 15532 5696
rect 14616 5654 14668 5662
rect 14808 5654 14860 5662
rect 15000 5654 15052 5662
rect 15192 5654 15244 5662
rect 8588 5524 9592 5536
rect 14612 5652 15244 5654
rect 15384 5652 15436 5662
rect 15576 5652 15628 5662
rect 14612 5644 14616 5652
rect 14668 5644 14808 5652
rect 14860 5644 15000 5652
rect 15052 5644 15192 5652
rect 7604 5510 8588 5520
rect 15244 5472 15384 5652
rect 15436 5472 15576 5652
rect 15216 5464 15628 5472
rect 15216 5462 15244 5464
rect 15384 5462 15436 5464
rect 15576 5462 15628 5464
rect 14612 5450 15216 5460
rect 8760 5348 9632 5358
rect 5712 5260 6972 5268
rect 5764 5080 5904 5260
rect 5956 5080 6096 5260
rect 6148 5080 6288 5260
rect 6340 5080 6480 5260
rect 6532 5080 6972 5260
rect 7708 5320 8760 5332
rect 7708 5140 7712 5320
rect 7768 5140 7904 5320
rect 7712 5126 7768 5136
rect 7960 5140 8096 5320
rect 7904 5126 7960 5136
rect 8152 5140 8288 5320
rect 8096 5126 8152 5136
rect 8344 5140 8480 5320
rect 8288 5126 8344 5136
rect 8536 5140 8672 5320
rect 8480 5126 8536 5136
rect 8728 5148 8760 5320
rect 8728 5140 8864 5148
rect 8760 5138 8864 5140
rect 8672 5126 8728 5136
rect 8920 5138 9056 5148
rect 8864 5126 8920 5136
rect 9112 5138 9248 5148
rect 9056 5126 9112 5136
rect 9304 5138 9440 5148
rect 9248 5126 9304 5136
rect 9496 5138 9632 5148
rect 14712 5268 15532 5272
rect 15660 5268 15972 5696
rect 16512 5884 17332 5888
rect 17460 5884 17772 5996
rect 16512 5876 17772 5884
rect 16564 5696 16704 5876
rect 16756 5696 16896 5876
rect 16948 5696 17088 5876
rect 17140 5696 17280 5876
rect 17332 5696 17772 5876
rect 16512 5686 16564 5696
rect 16704 5686 16756 5696
rect 16896 5686 16948 5696
rect 17088 5686 17140 5696
rect 17280 5686 17332 5696
rect 16416 5654 16468 5662
rect 16608 5654 16660 5662
rect 16800 5654 16852 5662
rect 16992 5654 17044 5662
rect 16412 5652 17044 5654
rect 17184 5652 17236 5662
rect 17376 5652 17428 5662
rect 16412 5644 16416 5652
rect 16468 5644 16608 5652
rect 16660 5644 16800 5652
rect 16852 5644 16992 5652
rect 17044 5472 17184 5652
rect 17236 5472 17376 5652
rect 17016 5464 17428 5472
rect 17016 5462 17044 5464
rect 17184 5462 17236 5464
rect 17376 5462 17428 5464
rect 16412 5450 17016 5460
rect 14712 5260 15972 5268
rect 9440 5126 9496 5136
rect 7616 5100 7672 5110
rect 7612 5094 7616 5096
rect 5712 5070 5764 5080
rect 5904 5070 5956 5080
rect 6096 5070 6148 5080
rect 6288 5070 6340 5080
rect 6480 5070 6532 5080
rect 5616 5038 5668 5046
rect 5808 5038 5860 5046
rect 6000 5038 6052 5046
rect 6192 5038 6244 5046
rect 5612 5036 6244 5038
rect 6384 5036 6436 5046
rect 6576 5036 6628 5046
rect 5612 5028 5616 5036
rect 5668 5028 5808 5036
rect 5860 5028 6000 5036
rect 6052 5028 6192 5036
rect 6244 4856 6384 5036
rect 6436 4856 6576 5036
rect 6216 4848 6628 4856
rect 6216 4846 6244 4848
rect 6384 4846 6436 4848
rect 6576 4846 6628 4848
rect 5612 4834 6216 4844
rect 3912 4640 5172 4644
rect 3964 4460 4104 4640
rect 4156 4460 4296 4640
rect 4348 4460 4488 4640
rect 4540 4460 4680 4640
rect 4732 4460 5172 4640
rect 3912 4456 5172 4460
rect 5712 4644 5764 4650
rect 5904 4644 5956 4650
rect 6096 4644 6148 4650
rect 6288 4644 6340 4650
rect 6480 4644 6532 4650
rect 6660 4644 6972 5080
rect 7604 5084 7616 5094
rect 7808 5100 7864 5110
rect 7672 5084 7808 5096
rect 8000 5100 8056 5110
rect 7864 5084 8000 5096
rect 8192 5100 8248 5110
rect 8056 5084 8192 5096
rect 8384 5100 8440 5110
rect 8248 5084 8384 5096
rect 8576 5100 8632 5110
rect 8440 5084 8576 5096
rect 8768 5100 8824 5110
rect 8632 4916 8768 5096
rect 8960 5100 9016 5110
rect 8824 4916 8960 5096
rect 9152 5100 9208 5110
rect 9016 4916 9152 5096
rect 9344 5100 9400 5110
rect 9208 4916 9344 5096
rect 9536 5100 9592 5110
rect 9400 4916 9536 5096
rect 8588 4904 9592 4916
rect 13996 5092 14428 5102
rect 7604 4886 8588 4896
rect 5712 4640 6972 4644
rect 5764 4460 5904 4640
rect 5956 4460 6096 4640
rect 6148 4460 6288 4640
rect 6340 4460 6480 4640
rect 6532 4460 6972 4640
rect 11480 4860 11820 4870
rect 11480 4570 11820 4580
rect 13592 4816 13996 4826
rect 14764 5080 14904 5260
rect 14956 5080 15096 5260
rect 15148 5080 15288 5260
rect 15340 5080 15480 5260
rect 15532 5080 15972 5260
rect 14712 5070 14764 5080
rect 14904 5070 14956 5080
rect 15096 5070 15148 5080
rect 15288 5070 15340 5080
rect 15480 5070 15532 5080
rect 14616 5038 14668 5046
rect 14808 5038 14860 5046
rect 15000 5038 15052 5046
rect 15192 5038 15244 5046
rect 14612 5036 15244 5038
rect 15384 5036 15436 5046
rect 15576 5036 15628 5046
rect 14612 5028 14616 5036
rect 14668 5028 14808 5036
rect 14860 5028 15000 5036
rect 15052 5028 15192 5036
rect 15244 4856 15384 5036
rect 15436 4856 15576 5036
rect 15216 4848 15628 4856
rect 15216 4846 15244 4848
rect 15384 4846 15436 4848
rect 15576 4846 15628 4848
rect 14612 4834 15216 4844
rect 5712 4456 6972 4460
rect 312 4450 364 4456
rect 504 4450 556 4456
rect 696 4450 748 4456
rect 888 4450 940 4456
rect 1080 4450 1132 4456
rect 2112 4450 2164 4456
rect 2304 4450 2356 4456
rect 2496 4450 2548 4456
rect 2688 4450 2740 4456
rect 2880 4450 2932 4456
rect 3912 4450 3964 4456
rect 4104 4450 4156 4456
rect 4296 4450 4348 4456
rect 4488 4450 4540 4456
rect 4680 4450 4732 4456
rect 5712 4450 5764 4456
rect 5904 4450 5956 4456
rect 6096 4450 6148 4456
rect 6288 4450 6340 4456
rect 6480 4450 6532 4456
rect 216 4418 268 4426
rect 408 4418 460 4426
rect 600 4418 652 4426
rect 792 4418 844 4426
rect -808 4400 -404 4404
rect -808 4394 28 4400
rect -404 4390 28 4394
rect 208 4416 844 4418
rect 984 4416 1036 4426
rect 1176 4416 1228 4426
rect 2016 4418 2068 4426
rect 2208 4418 2260 4426
rect 2400 4418 2452 4426
rect 2592 4418 2644 4426
rect 208 4408 216 4416
rect 268 4408 408 4416
rect 460 4408 600 4416
rect 652 4408 792 4416
rect 844 4236 984 4416
rect 1036 4236 1176 4416
rect 812 4228 1228 4236
rect 812 4226 844 4228
rect 984 4226 1036 4228
rect 1176 4226 1228 4228
rect 2008 4416 2644 4418
rect 2784 4416 2836 4426
rect 2976 4416 3028 4426
rect 3816 4418 3868 4426
rect 4008 4418 4060 4426
rect 4200 4418 4252 4426
rect 4392 4418 4444 4426
rect 2008 4408 2016 4416
rect 2068 4408 2208 4416
rect 2260 4408 2400 4416
rect 2452 4408 2592 4416
rect 2644 4236 2784 4416
rect 2836 4236 2976 4416
rect 208 4214 812 4224
rect 2612 4228 3028 4236
rect 2612 4226 2644 4228
rect 2784 4226 2836 4228
rect 2976 4226 3028 4228
rect 3808 4416 4444 4418
rect 4584 4416 4636 4426
rect 4776 4416 4828 4426
rect 5616 4418 5668 4426
rect 5808 4418 5860 4426
rect 6000 4418 6052 4426
rect 6192 4418 6244 4426
rect 3808 4408 3816 4416
rect 3868 4408 4008 4416
rect 4060 4408 4200 4416
rect 4252 4408 4392 4416
rect 4444 4236 4584 4416
rect 4636 4236 4776 4416
rect 2008 4214 2612 4224
rect 4412 4228 4828 4236
rect 4412 4226 4444 4228
rect 4584 4226 4636 4228
rect 4776 4226 4828 4228
rect 5608 4416 6244 4418
rect 6384 4416 6436 4426
rect 6576 4416 6628 4426
rect 5608 4408 5616 4416
rect 5668 4408 5808 4416
rect 5860 4408 6000 4416
rect 6052 4408 6192 4416
rect 6244 4236 6384 4416
rect 6436 4236 6576 4416
rect 14712 4644 14764 4650
rect 14904 4644 14956 4650
rect 15096 4644 15148 4650
rect 15288 4644 15340 4650
rect 15480 4644 15532 4650
rect 15660 4644 15972 5080
rect 16512 5268 17332 5272
rect 17460 5268 17772 5696
rect 18312 5884 19132 5888
rect 19260 5884 19572 5996
rect 18312 5876 19572 5884
rect 18364 5696 18504 5876
rect 18556 5696 18696 5876
rect 18748 5696 18888 5876
rect 18940 5696 19080 5876
rect 19132 5696 19572 5876
rect 18312 5686 18364 5696
rect 18504 5686 18556 5696
rect 18696 5686 18748 5696
rect 18888 5686 18940 5696
rect 19080 5686 19132 5696
rect 18216 5654 18268 5662
rect 18408 5654 18460 5662
rect 18600 5654 18652 5662
rect 18792 5654 18844 5662
rect 18212 5652 18844 5654
rect 18984 5652 19036 5662
rect 19176 5652 19228 5662
rect 18212 5644 18216 5652
rect 18268 5644 18408 5652
rect 18460 5644 18600 5652
rect 18652 5644 18792 5652
rect 18844 5472 18984 5652
rect 19036 5472 19176 5652
rect 18816 5464 19228 5472
rect 18816 5462 18844 5464
rect 18984 5462 19036 5464
rect 19176 5462 19228 5464
rect 18212 5450 18816 5460
rect 16512 5260 17772 5268
rect 16564 5080 16704 5260
rect 16756 5080 16896 5260
rect 16948 5080 17088 5260
rect 17140 5080 17280 5260
rect 17332 5080 17772 5260
rect 16512 5070 16564 5080
rect 16704 5070 16756 5080
rect 16896 5070 16948 5080
rect 17088 5070 17140 5080
rect 17280 5070 17332 5080
rect 16416 5038 16468 5046
rect 16608 5038 16660 5046
rect 16800 5038 16852 5046
rect 16992 5038 17044 5046
rect 16412 5036 17044 5038
rect 17184 5036 17236 5046
rect 17376 5036 17428 5046
rect 16412 5028 16416 5036
rect 16468 5028 16608 5036
rect 16660 5028 16800 5036
rect 16852 5028 16992 5036
rect 17044 4856 17184 5036
rect 17236 4856 17376 5036
rect 17016 4848 17428 4856
rect 17016 4846 17044 4848
rect 17184 4846 17236 4848
rect 17376 4846 17428 4848
rect 16412 4834 17016 4844
rect 14712 4640 15972 4644
rect 14764 4460 14904 4640
rect 14956 4460 15096 4640
rect 15148 4460 15288 4640
rect 15340 4460 15480 4640
rect 15532 4460 15972 4640
rect 14712 4456 15972 4460
rect 16512 4644 16564 4650
rect 16704 4644 16756 4650
rect 16896 4644 16948 4650
rect 17088 4644 17140 4650
rect 17280 4644 17332 4650
rect 17460 4644 17772 5080
rect 18312 5268 19132 5272
rect 19260 5268 19572 5696
rect 20112 5884 20932 5888
rect 21060 5884 21488 6052
rect 20112 5876 21488 5884
rect 20164 5696 20304 5876
rect 20356 5696 20496 5876
rect 20548 5696 20688 5876
rect 20740 5696 20880 5876
rect 20932 5696 21488 5876
rect 20112 5686 20164 5696
rect 20304 5686 20356 5696
rect 20496 5686 20548 5696
rect 20688 5686 20740 5696
rect 20880 5686 20932 5696
rect 20016 5654 20068 5662
rect 20208 5654 20260 5662
rect 20400 5654 20452 5662
rect 20592 5654 20644 5662
rect 20012 5652 20644 5654
rect 20784 5652 20836 5662
rect 20976 5652 21028 5662
rect 20012 5644 20016 5652
rect 20068 5644 20208 5652
rect 20260 5644 20400 5652
rect 20452 5644 20592 5652
rect 20644 5472 20784 5652
rect 20836 5472 20976 5652
rect 20616 5464 21028 5472
rect 20616 5462 20644 5464
rect 20784 5462 20836 5464
rect 20976 5462 21028 5464
rect 21060 5584 21488 5696
rect 20012 5450 20616 5460
rect 18312 5260 19572 5268
rect 18364 5080 18504 5260
rect 18556 5080 18696 5260
rect 18748 5080 18888 5260
rect 18940 5080 19080 5260
rect 19132 5080 19572 5260
rect 18312 5070 18364 5080
rect 18504 5070 18556 5080
rect 18696 5070 18748 5080
rect 18888 5070 18940 5080
rect 19080 5070 19132 5080
rect 18216 5038 18268 5046
rect 18408 5038 18460 5046
rect 18600 5038 18652 5046
rect 18792 5038 18844 5046
rect 18212 5036 18844 5038
rect 18984 5036 19036 5046
rect 19176 5036 19228 5046
rect 18212 5028 18216 5036
rect 18268 5028 18408 5036
rect 18460 5028 18600 5036
rect 18652 5028 18792 5036
rect 18844 4856 18984 5036
rect 19036 4856 19176 5036
rect 18816 4848 19228 4856
rect 18816 4846 18844 4848
rect 18984 4846 19036 4848
rect 19176 4846 19228 4848
rect 18212 4834 18816 4844
rect 16512 4640 17772 4644
rect 16564 4460 16704 4640
rect 16756 4460 16896 4640
rect 16948 4460 17088 4640
rect 17140 4460 17280 4640
rect 17332 4460 17772 4640
rect 16512 4456 17772 4460
rect 18312 4644 18364 4650
rect 18504 4644 18556 4650
rect 18696 4644 18748 4650
rect 18888 4644 18940 4650
rect 19080 4644 19132 4650
rect 19260 4644 19572 5080
rect 20112 5268 20932 5272
rect 21060 5268 21372 5584
rect 23160 5968 24032 5978
rect 22108 5940 23160 5952
rect 22108 5760 22112 5940
rect 22168 5760 22304 5940
rect 22112 5746 22168 5756
rect 22360 5760 22496 5940
rect 22304 5746 22360 5756
rect 22552 5760 22688 5940
rect 22496 5746 22552 5756
rect 22744 5760 22880 5940
rect 22688 5746 22744 5756
rect 22936 5760 23072 5940
rect 22880 5746 22936 5756
rect 23128 5768 23160 5940
rect 23128 5760 23264 5768
rect 23160 5758 23264 5760
rect 23072 5746 23128 5756
rect 23320 5758 23456 5768
rect 23264 5746 23320 5756
rect 23512 5758 23648 5768
rect 23456 5746 23512 5756
rect 23704 5758 23840 5768
rect 23648 5746 23704 5756
rect 23896 5758 24032 5768
rect 23840 5746 23896 5756
rect 22016 5720 22072 5730
rect 21488 5570 21772 5580
rect 22004 5708 22016 5718
rect 22208 5720 22264 5730
rect 22072 5708 22208 5718
rect 22400 5720 22456 5730
rect 22264 5708 22400 5718
rect 22592 5720 22648 5730
rect 22456 5708 22592 5718
rect 22784 5720 22840 5730
rect 22648 5708 22784 5718
rect 22976 5720 23032 5730
rect 22840 5708 22976 5718
rect 23168 5720 23224 5730
rect 23032 5536 23168 5716
rect 23360 5720 23416 5730
rect 23224 5536 23360 5716
rect 23552 5720 23608 5730
rect 23416 5536 23552 5716
rect 23744 5720 23800 5730
rect 23608 5536 23744 5716
rect 23936 5720 23992 5730
rect 23800 5536 23936 5716
rect 22988 5524 23992 5536
rect 22004 5510 22988 5520
rect 23160 5348 24032 5358
rect 20112 5260 21372 5268
rect 20164 5080 20304 5260
rect 20356 5080 20496 5260
rect 20548 5080 20688 5260
rect 20740 5080 20880 5260
rect 20932 5080 21372 5260
rect 22108 5320 23160 5332
rect 22108 5140 22112 5320
rect 22168 5140 22304 5320
rect 22112 5126 22168 5136
rect 22360 5140 22496 5320
rect 22304 5126 22360 5136
rect 22552 5140 22688 5320
rect 22496 5126 22552 5136
rect 22744 5140 22880 5320
rect 22688 5126 22744 5136
rect 22936 5140 23072 5320
rect 22880 5126 22936 5136
rect 23128 5148 23160 5320
rect 23128 5140 23264 5148
rect 23160 5138 23264 5140
rect 23072 5126 23128 5136
rect 23320 5138 23456 5148
rect 23264 5126 23320 5136
rect 23512 5138 23648 5148
rect 23456 5126 23512 5136
rect 23704 5138 23840 5148
rect 23648 5126 23704 5136
rect 23896 5138 24032 5148
rect 23840 5126 23896 5136
rect 22016 5100 22072 5110
rect 22012 5094 22016 5096
rect 20112 5070 20164 5080
rect 20304 5070 20356 5080
rect 20496 5070 20548 5080
rect 20688 5070 20740 5080
rect 20880 5070 20932 5080
rect 20016 5038 20068 5046
rect 20208 5038 20260 5046
rect 20400 5038 20452 5046
rect 20592 5038 20644 5046
rect 20012 5036 20644 5038
rect 20784 5036 20836 5046
rect 20976 5036 21028 5046
rect 20012 5028 20016 5036
rect 20068 5028 20208 5036
rect 20260 5028 20400 5036
rect 20452 5028 20592 5036
rect 20644 4856 20784 5036
rect 20836 4856 20976 5036
rect 20616 4848 21028 4856
rect 20616 4846 20644 4848
rect 20784 4846 20836 4848
rect 20976 4846 21028 4848
rect 20012 4834 20616 4844
rect 18312 4640 19572 4644
rect 18364 4460 18504 4640
rect 18556 4460 18696 4640
rect 18748 4460 18888 4640
rect 18940 4460 19080 4640
rect 19132 4460 19572 4640
rect 18312 4456 19572 4460
rect 20112 4644 20164 4650
rect 20304 4644 20356 4650
rect 20496 4644 20548 4650
rect 20688 4644 20740 4650
rect 20880 4644 20932 4650
rect 21060 4644 21372 5080
rect 22004 5084 22016 5094
rect 22208 5100 22264 5110
rect 22072 5084 22208 5096
rect 22400 5100 22456 5110
rect 22264 5084 22400 5096
rect 22592 5100 22648 5110
rect 22456 5084 22592 5096
rect 22784 5100 22840 5110
rect 22648 5084 22784 5096
rect 22976 5100 23032 5110
rect 22840 5084 22976 5096
rect 23168 5100 23224 5110
rect 23032 4916 23168 5096
rect 23360 5100 23416 5110
rect 23224 4916 23360 5096
rect 23552 5100 23608 5110
rect 23416 4916 23552 5096
rect 23744 5100 23800 5110
rect 23608 4916 23744 5096
rect 23936 5100 23992 5110
rect 23800 4916 23936 5096
rect 22988 4904 23992 4916
rect 22004 4886 22988 4896
rect 20112 4640 21372 4644
rect 20164 4460 20304 4640
rect 20356 4460 20496 4640
rect 20548 4460 20688 4640
rect 20740 4460 20880 4640
rect 20932 4460 21372 4640
rect 20112 4456 21372 4460
rect 24520 4700 24900 4710
rect 14712 4450 14764 4456
rect 14904 4450 14956 4456
rect 15096 4450 15148 4456
rect 15288 4450 15340 4456
rect 15480 4450 15532 4456
rect 16512 4450 16564 4456
rect 16704 4450 16756 4456
rect 16896 4450 16948 4456
rect 17088 4450 17140 4456
rect 17280 4450 17332 4456
rect 18312 4450 18364 4456
rect 18504 4450 18556 4456
rect 18696 4450 18748 4456
rect 18888 4450 18940 4456
rect 19080 4450 19132 4456
rect 20112 4450 20164 4456
rect 20304 4450 20356 4456
rect 20496 4450 20548 4456
rect 20688 4450 20740 4456
rect 20880 4450 20932 4456
rect 14616 4418 14668 4426
rect 14808 4418 14860 4426
rect 15000 4418 15052 4426
rect 15192 4418 15244 4426
rect 13592 4400 13996 4404
rect 13592 4394 14428 4400
rect 13996 4390 14428 4394
rect 14608 4416 15244 4418
rect 15384 4416 15436 4426
rect 15576 4416 15628 4426
rect 16416 4418 16468 4426
rect 16608 4418 16660 4426
rect 16800 4418 16852 4426
rect 16992 4418 17044 4426
rect 14608 4408 14616 4416
rect 14668 4408 14808 4416
rect 14860 4408 15000 4416
rect 15052 4408 15192 4416
rect 3808 4214 4412 4224
rect 6212 4228 6628 4236
rect 6212 4226 6244 4228
rect 6384 4226 6436 4228
rect 6576 4226 6628 4228
rect 15244 4236 15384 4416
rect 15436 4236 15576 4416
rect 5608 4214 6212 4224
rect 15212 4228 15628 4236
rect 15212 4226 15244 4228
rect 15384 4226 15436 4228
rect 15576 4226 15628 4228
rect 16408 4416 17044 4418
rect 17184 4416 17236 4426
rect 17376 4416 17428 4426
rect 18216 4418 18268 4426
rect 18408 4418 18460 4426
rect 18600 4418 18652 4426
rect 18792 4418 18844 4426
rect 16408 4408 16416 4416
rect 16468 4408 16608 4416
rect 16660 4408 16800 4416
rect 16852 4408 16992 4416
rect 17044 4236 17184 4416
rect 17236 4236 17376 4416
rect 14608 4214 15212 4224
rect 17012 4228 17428 4236
rect 17012 4226 17044 4228
rect 17184 4226 17236 4228
rect 17376 4226 17428 4228
rect 18208 4416 18844 4418
rect 18984 4416 19036 4426
rect 19176 4416 19228 4426
rect 20016 4418 20068 4426
rect 20208 4418 20260 4426
rect 20400 4418 20452 4426
rect 20592 4418 20644 4426
rect 18208 4408 18216 4416
rect 18268 4408 18408 4416
rect 18460 4408 18600 4416
rect 18652 4408 18792 4416
rect 18844 4236 18984 4416
rect 19036 4236 19176 4416
rect 16408 4214 17012 4224
rect 18812 4228 19228 4236
rect 18812 4226 18844 4228
rect 18984 4226 19036 4228
rect 19176 4226 19228 4228
rect 20008 4416 20644 4418
rect 20784 4416 20836 4426
rect 20976 4416 21028 4426
rect 20008 4408 20016 4416
rect 20068 4408 20208 4416
rect 20260 4408 20400 4416
rect 20452 4408 20592 4416
rect 20644 4236 20784 4416
rect 20836 4236 20976 4416
rect 24520 4350 24900 4360
rect 18208 4214 18812 4224
rect 20612 4228 21028 4236
rect 20612 4226 20644 4228
rect 20784 4226 20836 4228
rect 20976 4226 21028 4228
rect 20008 4214 20612 4224
rect -10060 4020 -9460 4030
rect -9460 4008 -8976 4020
rect -9460 3836 -9028 4008
rect -10008 3828 -9544 3836
rect -9492 3828 -9028 3836
rect -10060 3826 -9460 3828
rect -10060 3818 -10008 3826
rect -9544 3818 -9492 3826
rect -9028 3818 -8976 3828
rect -9800 3788 -9748 3798
rect -9284 3790 -9232 3798
rect -8768 3790 -8716 3798
rect -9316 3788 -8716 3790
rect -9748 3780 -9284 3788
rect -9232 3780 -8768 3788
rect -9748 3608 -9316 3780
rect -9800 3596 -9316 3608
rect -9316 3586 -8716 3596
rect 216 3740 816 3750
rect 1236 3740 6712 3764
rect 816 3728 2016 3740
rect 2616 3728 3816 3740
rect 4416 3728 5616 3740
rect 6216 3728 6712 3740
rect 816 3556 1248 3728
rect 268 3548 732 3556
rect 784 3548 1248 3556
rect 1300 3548 2016 3728
rect 2616 3556 3048 3728
rect 2068 3548 2532 3556
rect 2584 3548 3048 3556
rect 3100 3548 3816 3728
rect 4416 3556 4848 3728
rect 3868 3548 4332 3556
rect 4384 3548 4848 3556
rect 4900 3548 5616 3728
rect 6216 3556 6648 3728
rect 5668 3548 6132 3556
rect 6184 3548 6648 3556
rect 6700 3548 6712 3728
rect 14616 3740 15216 3750
rect 15636 3740 21112 3764
rect 15216 3728 16416 3740
rect 17016 3728 18216 3740
rect 18816 3728 20016 3740
rect 20616 3728 21112 3740
rect 15216 3556 15648 3728
rect 14668 3548 15132 3556
rect 15184 3548 15648 3556
rect 15700 3548 16416 3728
rect 17016 3556 17448 3728
rect 16468 3548 16932 3556
rect 16984 3548 17448 3556
rect 17500 3548 18216 3728
rect 18816 3556 19248 3728
rect 18268 3548 18732 3556
rect 18784 3548 19248 3556
rect 19300 3548 20016 3728
rect 20616 3556 21048 3728
rect 20068 3548 20532 3556
rect 20584 3548 21048 3556
rect 21100 3548 21112 3728
rect 216 3546 816 3548
rect 216 3538 268 3546
rect 732 3538 784 3546
rect 1248 3538 1300 3548
rect 2016 3546 2616 3548
rect 2016 3538 2068 3546
rect 2532 3538 2584 3546
rect 3048 3538 3100 3548
rect 3816 3546 4416 3548
rect 3816 3538 3868 3546
rect 4332 3538 4384 3546
rect 4848 3538 4900 3548
rect 5616 3546 6216 3548
rect 5616 3538 5668 3546
rect 6132 3538 6184 3546
rect 6648 3538 6700 3548
rect 14616 3546 15216 3548
rect 14616 3538 14668 3546
rect 15132 3538 15184 3546
rect 15648 3538 15700 3548
rect 16416 3546 17016 3548
rect 16416 3538 16468 3546
rect 16932 3538 16984 3546
rect 17448 3538 17500 3548
rect 18216 3546 18816 3548
rect 18216 3538 18268 3546
rect 18732 3538 18784 3546
rect 19248 3538 19300 3548
rect 20016 3546 20616 3548
rect 20016 3538 20068 3546
rect 20532 3538 20584 3546
rect 21048 3538 21100 3548
rect 476 3508 528 3518
rect 992 3510 1044 3518
rect 1508 3510 1560 3518
rect 960 3508 1560 3510
rect -10060 3404 -9460 3414
rect -9460 3392 -8976 3404
rect -9460 3220 -9028 3392
rect -10008 3212 -9544 3220
rect -9492 3212 -9028 3220
rect 528 3500 992 3508
rect 1044 3500 1508 3508
rect 528 3328 960 3500
rect 476 3316 960 3328
rect 2276 3508 2328 3518
rect 2792 3510 2844 3518
rect 3308 3510 3360 3518
rect 2760 3508 3360 3510
rect 2328 3500 2792 3508
rect 2844 3500 3308 3508
rect 2328 3328 2760 3500
rect 2276 3316 2760 3328
rect 4076 3508 4128 3518
rect 4592 3510 4644 3518
rect 5108 3510 5160 3518
rect 4560 3508 5160 3510
rect 4128 3500 4592 3508
rect 4644 3500 5108 3508
rect 4128 3328 4560 3500
rect 4076 3316 4560 3328
rect 5876 3508 5928 3518
rect 6392 3510 6444 3518
rect 6908 3510 6960 3518
rect 6360 3508 6960 3510
rect 5928 3500 6392 3508
rect 6444 3500 6908 3508
rect 5928 3328 6360 3500
rect 5876 3316 6360 3328
rect 14876 3508 14928 3518
rect 15392 3510 15444 3518
rect 15908 3510 15960 3518
rect 15360 3508 15960 3510
rect 14928 3500 15392 3508
rect 15444 3500 15908 3508
rect 14928 3328 15360 3500
rect 14876 3316 15360 3328
rect 16676 3508 16728 3518
rect 17192 3510 17244 3518
rect 17708 3510 17760 3518
rect 17160 3508 17760 3510
rect 16728 3500 17192 3508
rect 17244 3500 17708 3508
rect 16728 3328 17160 3500
rect 16676 3316 17160 3328
rect 18476 3508 18528 3518
rect 18992 3510 19044 3518
rect 19508 3510 19560 3518
rect 18960 3508 19560 3510
rect 18528 3500 18992 3508
rect 19044 3500 19508 3508
rect 18528 3328 18960 3500
rect 18476 3316 18960 3328
rect 20276 3508 20328 3518
rect 20792 3510 20844 3518
rect 21308 3510 21360 3518
rect 20760 3508 21360 3510
rect 20328 3500 20792 3508
rect 20844 3500 21308 3508
rect 20328 3328 20760 3500
rect 20276 3316 20760 3328
rect 960 3306 1560 3316
rect 2760 3306 3360 3316
rect 4560 3306 5160 3316
rect 6360 3306 6960 3316
rect 15360 3306 15960 3316
rect 17160 3306 17760 3316
rect 18960 3306 19560 3316
rect 20760 3306 21360 3316
rect -10060 3210 -9460 3212
rect -10060 3202 -10008 3210
rect -9544 3202 -9492 3210
rect -9028 3202 -8976 3212
rect -9800 3172 -9748 3182
rect -9284 3174 -9232 3182
rect -8768 3174 -8716 3182
rect -9316 3172 -8716 3174
rect -9748 3164 -9284 3172
rect -9232 3164 -8768 3172
rect -9748 2992 -9316 3164
rect -9800 2980 -9316 2992
rect -9316 2970 -8716 2980
rect 216 3124 816 3134
rect 2016 3124 2616 3134
rect 3816 3124 4416 3134
rect 5616 3124 6216 3134
rect 14616 3124 15216 3134
rect 16416 3124 17016 3134
rect 18216 3124 18816 3134
rect 20016 3124 20616 3134
rect 816 3112 1300 3124
rect 816 2940 1248 3112
rect 268 2932 732 2940
rect 784 2932 1248 2940
rect 216 2930 816 2932
rect 216 2922 268 2930
rect 732 2922 784 2930
rect 1248 2922 1300 2932
rect 2616 3112 3100 3124
rect 2616 2940 3048 3112
rect 2068 2932 2532 2940
rect 2584 2932 3048 2940
rect 2016 2930 2616 2932
rect 2016 2922 2068 2930
rect 2532 2922 2584 2930
rect 3048 2922 3100 2932
rect 4416 3112 4900 3124
rect 4416 2940 4848 3112
rect 3868 2932 4332 2940
rect 4384 2932 4848 2940
rect 3816 2930 4416 2932
rect 3816 2922 3868 2930
rect 4332 2922 4384 2930
rect 4848 2922 4900 2932
rect 6216 3112 6700 3124
rect 6216 2940 6648 3112
rect 5668 2932 6132 2940
rect 6184 2932 6648 2940
rect 5616 2930 6216 2932
rect 5616 2922 5668 2930
rect 6132 2922 6184 2930
rect 6648 2922 6700 2932
rect 15216 3112 15700 3124
rect 15216 2940 15648 3112
rect 14668 2932 15132 2940
rect 15184 2932 15648 2940
rect 14616 2930 15216 2932
rect 14616 2922 14668 2930
rect 15132 2922 15184 2930
rect 15648 2922 15700 2932
rect 17016 3112 17500 3124
rect 17016 2940 17448 3112
rect 16468 2932 16932 2940
rect 16984 2932 17448 2940
rect 16416 2930 17016 2932
rect 16416 2922 16468 2930
rect 16932 2922 16984 2930
rect 17448 2922 17500 2932
rect 18816 3112 19300 3124
rect 18816 2940 19248 3112
rect 18268 2932 18732 2940
rect 18784 2932 19248 2940
rect 18216 2930 18816 2932
rect 18216 2922 18268 2930
rect 18732 2922 18784 2930
rect 19248 2922 19300 2932
rect 20616 3112 21100 3124
rect 20616 2940 21048 3112
rect 20068 2932 20532 2940
rect 20584 2932 21048 2940
rect 20016 2930 20616 2932
rect 20016 2922 20068 2930
rect 20532 2922 20584 2930
rect 21048 2922 21100 2932
rect 476 2892 528 2902
rect 992 2894 1044 2902
rect 1508 2894 1560 2902
rect 960 2892 1560 2894
rect -10060 2784 -9460 2794
rect -9460 2772 -8976 2784
rect -9460 2600 -9028 2772
rect -10008 2592 -9544 2600
rect -9492 2592 -9028 2600
rect 528 2884 992 2892
rect 1044 2884 1508 2892
rect 528 2712 960 2884
rect 476 2700 960 2712
rect 2276 2892 2328 2902
rect 2792 2894 2844 2902
rect 3308 2894 3360 2902
rect 2760 2892 3360 2894
rect 2328 2884 2792 2892
rect 2844 2884 3308 2892
rect 2328 2712 2760 2884
rect 2276 2700 2760 2712
rect 4076 2892 4128 2902
rect 4592 2894 4644 2902
rect 5108 2894 5160 2902
rect 4560 2892 5160 2894
rect 4128 2884 4592 2892
rect 4644 2884 5108 2892
rect 4128 2712 4560 2884
rect 4076 2700 4560 2712
rect 5876 2892 5928 2902
rect 6392 2894 6444 2902
rect 6908 2894 6960 2902
rect 6360 2892 6960 2894
rect 5928 2884 6392 2892
rect 6444 2884 6908 2892
rect 5928 2712 6360 2884
rect 5876 2700 6360 2712
rect 14876 2892 14928 2902
rect 15392 2894 15444 2902
rect 15908 2894 15960 2902
rect 15360 2892 15960 2894
rect 14928 2884 15392 2892
rect 15444 2884 15908 2892
rect 14928 2712 15360 2884
rect 14876 2700 15360 2712
rect 16676 2892 16728 2902
rect 17192 2894 17244 2902
rect 17708 2894 17760 2902
rect 17160 2892 17760 2894
rect 16728 2884 17192 2892
rect 17244 2884 17708 2892
rect 16728 2712 17160 2884
rect 16676 2700 17160 2712
rect 18476 2892 18528 2902
rect 18992 2894 19044 2902
rect 19508 2894 19560 2902
rect 18960 2892 19560 2894
rect 18528 2884 18992 2892
rect 19044 2884 19508 2892
rect 18528 2712 18960 2884
rect 18476 2700 18960 2712
rect 20276 2892 20328 2902
rect 20792 2894 20844 2902
rect 21308 2894 21360 2902
rect 20760 2892 21360 2894
rect 20328 2884 20792 2892
rect 20844 2884 21308 2892
rect 20328 2712 20760 2884
rect 20276 2700 20760 2712
rect 960 2690 1560 2700
rect 2760 2690 3360 2700
rect 4560 2690 5160 2700
rect 6360 2690 6960 2700
rect 15360 2690 15960 2700
rect 17160 2690 17760 2700
rect 18960 2690 19560 2700
rect 20760 2690 21360 2700
rect -10060 2590 -9460 2592
rect -10060 2582 -10008 2590
rect -9544 2582 -9492 2590
rect -9028 2582 -8976 2592
rect -9800 2552 -9748 2562
rect -9284 2554 -9232 2562
rect -8768 2554 -8716 2562
rect -9316 2552 -8716 2554
rect -9748 2544 -9284 2552
rect -9232 2544 -8768 2552
rect -9748 2372 -9316 2544
rect -9800 2360 -9316 2372
rect -9316 2350 -8716 2360
rect 216 2504 816 2514
rect 2016 2504 2616 2514
rect 3816 2504 4416 2514
rect 5616 2504 6216 2514
rect 14616 2504 15216 2514
rect 16416 2504 17016 2514
rect 18216 2504 18816 2514
rect 20016 2504 20616 2514
rect 816 2492 1300 2504
rect 816 2320 1248 2492
rect 268 2312 732 2320
rect 784 2312 1248 2320
rect 216 2310 816 2312
rect 216 2302 268 2310
rect 732 2302 784 2310
rect 1248 2302 1300 2312
rect 2616 2492 3100 2504
rect 2616 2320 3048 2492
rect 2068 2312 2532 2320
rect 2584 2312 3048 2320
rect 2016 2310 2616 2312
rect 2016 2302 2068 2310
rect 2532 2302 2584 2310
rect 3048 2302 3100 2312
rect 4416 2492 4900 2504
rect 4416 2320 4848 2492
rect 3868 2312 4332 2320
rect 4384 2312 4848 2320
rect 3816 2310 4416 2312
rect 3816 2302 3868 2310
rect 4332 2302 4384 2310
rect 4848 2302 4900 2312
rect 6216 2492 6700 2504
rect 6216 2320 6648 2492
rect 5668 2312 6132 2320
rect 6184 2312 6648 2320
rect 5616 2310 6216 2312
rect 5616 2302 5668 2310
rect 6132 2302 6184 2310
rect 6648 2302 6700 2312
rect 15216 2492 15700 2504
rect 15216 2320 15648 2492
rect 14668 2312 15132 2320
rect 15184 2312 15648 2320
rect 14616 2310 15216 2312
rect 14616 2302 14668 2310
rect 15132 2302 15184 2310
rect 15648 2302 15700 2312
rect 17016 2492 17500 2504
rect 17016 2320 17448 2492
rect 16468 2312 16932 2320
rect 16984 2312 17448 2320
rect 16416 2310 17016 2312
rect 16416 2302 16468 2310
rect 16932 2302 16984 2310
rect 17448 2302 17500 2312
rect 18816 2492 19300 2504
rect 18816 2320 19248 2492
rect 18268 2312 18732 2320
rect 18784 2312 19248 2320
rect 18216 2310 18816 2312
rect 18216 2302 18268 2310
rect 18732 2302 18784 2310
rect 19248 2302 19300 2312
rect 20616 2492 21100 2504
rect 20616 2320 21048 2492
rect 20068 2312 20532 2320
rect 20584 2312 21048 2320
rect 20016 2310 20616 2312
rect 20016 2302 20068 2310
rect 20532 2302 20584 2310
rect 21048 2302 21100 2312
rect 476 2272 528 2282
rect 992 2274 1044 2282
rect 1508 2274 1560 2282
rect 960 2272 1560 2274
rect -10060 2168 -9460 2178
rect -9460 2156 -8976 2168
rect -9460 1984 -9028 2156
rect -10008 1976 -9544 1984
rect -9492 1976 -9028 1984
rect 528 2264 992 2272
rect 1044 2264 1508 2272
rect 528 2092 960 2264
rect 476 2080 960 2092
rect 2276 2272 2328 2282
rect 2792 2274 2844 2282
rect 3308 2274 3360 2282
rect 2760 2272 3360 2274
rect 2328 2264 2792 2272
rect 2844 2264 3308 2272
rect 2328 2092 2760 2264
rect 2276 2080 2760 2092
rect 4076 2272 4128 2282
rect 4592 2274 4644 2282
rect 5108 2274 5160 2282
rect 4560 2272 5160 2274
rect 4128 2264 4592 2272
rect 4644 2264 5108 2272
rect 4128 2092 4560 2264
rect 4076 2080 4560 2092
rect 5876 2272 5928 2282
rect 6392 2274 6444 2282
rect 6908 2274 6960 2282
rect 6360 2272 6960 2274
rect 5928 2264 6392 2272
rect 6444 2264 6908 2272
rect 5928 2092 6360 2264
rect 5876 2080 6360 2092
rect 14876 2272 14928 2282
rect 15392 2274 15444 2282
rect 15908 2274 15960 2282
rect 15360 2272 15960 2274
rect 14928 2264 15392 2272
rect 15444 2264 15908 2272
rect 14928 2092 15360 2264
rect 14876 2080 15360 2092
rect 16676 2272 16728 2282
rect 17192 2274 17244 2282
rect 17708 2274 17760 2282
rect 17160 2272 17760 2274
rect 16728 2264 17192 2272
rect 17244 2264 17708 2272
rect 16728 2092 17160 2264
rect 16676 2080 17160 2092
rect 18476 2272 18528 2282
rect 18992 2274 19044 2282
rect 19508 2274 19560 2282
rect 18960 2272 19560 2274
rect 18528 2264 18992 2272
rect 19044 2264 19508 2272
rect 18528 2092 18960 2264
rect 18476 2080 18960 2092
rect 20276 2272 20328 2282
rect 20792 2274 20844 2282
rect 21308 2274 21360 2282
rect 20760 2272 21360 2274
rect 20328 2264 20792 2272
rect 20844 2264 21308 2272
rect 20328 2092 20760 2264
rect 20276 2080 20760 2092
rect 960 2070 1560 2080
rect 2760 2070 3360 2080
rect 4560 2070 5160 2080
rect 6360 2070 6960 2080
rect 15360 2070 15960 2080
rect 17160 2070 17760 2080
rect 18960 2070 19560 2080
rect 20760 2070 21360 2080
rect -10060 1974 -9460 1976
rect -10060 1966 -10008 1974
rect -9544 1966 -9492 1974
rect -9028 1966 -8976 1976
rect -9800 1936 -9748 1946
rect -9284 1938 -9232 1946
rect -8768 1938 -8716 1946
rect -9316 1936 -8716 1938
rect -9748 1928 -9284 1936
rect -9232 1928 -8768 1936
rect -9748 1756 -9316 1928
rect -9800 1744 -9316 1756
rect -9316 1734 -8716 1744
rect 216 1888 816 1898
rect 2016 1888 2616 1898
rect 3816 1888 4416 1898
rect 5616 1888 6216 1898
rect 14616 1888 15216 1898
rect 16416 1888 17016 1898
rect 18216 1888 18816 1898
rect 20016 1888 20616 1898
rect 816 1876 1300 1888
rect 816 1704 1248 1876
rect 268 1696 732 1704
rect 784 1696 1248 1704
rect 216 1694 816 1696
rect 216 1686 268 1694
rect 732 1686 784 1694
rect 1248 1686 1300 1696
rect 2616 1876 3100 1888
rect 2616 1704 3048 1876
rect 2068 1696 2532 1704
rect 2584 1696 3048 1704
rect 2016 1694 2616 1696
rect 2016 1686 2068 1694
rect 2532 1686 2584 1694
rect 3048 1686 3100 1696
rect 4416 1876 4900 1888
rect 4416 1704 4848 1876
rect 3868 1696 4332 1704
rect 4384 1696 4848 1704
rect 3816 1694 4416 1696
rect 3816 1686 3868 1694
rect 4332 1686 4384 1694
rect 4848 1686 4900 1696
rect 6216 1876 6700 1888
rect 6216 1704 6648 1876
rect 5668 1696 6132 1704
rect 6184 1696 6648 1704
rect 5616 1694 6216 1696
rect 5616 1686 5668 1694
rect 6132 1686 6184 1694
rect 6648 1686 6700 1696
rect 15216 1876 15700 1888
rect 15216 1704 15648 1876
rect 14668 1696 15132 1704
rect 15184 1696 15648 1704
rect 14616 1694 15216 1696
rect 14616 1686 14668 1694
rect 15132 1686 15184 1694
rect 15648 1686 15700 1696
rect 17016 1876 17500 1888
rect 17016 1704 17448 1876
rect 16468 1696 16932 1704
rect 16984 1696 17448 1704
rect 16416 1694 17016 1696
rect 16416 1686 16468 1694
rect 16932 1686 16984 1694
rect 17448 1686 17500 1696
rect 18816 1876 19300 1888
rect 18816 1704 19248 1876
rect 18268 1696 18732 1704
rect 18784 1696 19248 1704
rect 18216 1694 18816 1696
rect 18216 1686 18268 1694
rect 18732 1686 18784 1694
rect 19248 1686 19300 1696
rect 20616 1876 21100 1888
rect 20616 1704 21048 1876
rect 20068 1696 20532 1704
rect 20584 1696 21048 1704
rect 20016 1694 20616 1696
rect 20016 1686 20068 1694
rect 20532 1686 20584 1694
rect 21048 1686 21100 1696
rect 476 1656 528 1666
rect 992 1658 1044 1666
rect 1508 1658 1560 1666
rect 960 1656 1560 1658
rect -10060 1548 -9460 1558
rect -9460 1536 -8976 1548
rect -9460 1364 -9028 1536
rect -10008 1356 -9544 1364
rect -9492 1356 -9028 1364
rect 528 1648 992 1656
rect 1044 1648 1508 1656
rect 528 1476 960 1648
rect 476 1464 960 1476
rect 2276 1656 2328 1666
rect 2792 1658 2844 1666
rect 3308 1658 3360 1666
rect 2760 1656 3360 1658
rect 2328 1648 2792 1656
rect 2844 1648 3308 1656
rect 2328 1476 2760 1648
rect 2276 1464 2760 1476
rect 4076 1656 4128 1666
rect 4592 1658 4644 1666
rect 5108 1658 5160 1666
rect 4560 1656 5160 1658
rect 4128 1648 4592 1656
rect 4644 1648 5108 1656
rect 4128 1476 4560 1648
rect 4076 1464 4560 1476
rect 5876 1656 5928 1666
rect 6392 1658 6444 1666
rect 6908 1658 6960 1666
rect 6360 1656 6960 1658
rect 5928 1648 6392 1656
rect 6444 1648 6908 1656
rect 5928 1476 6360 1648
rect 5876 1464 6360 1476
rect 14876 1656 14928 1666
rect 15392 1658 15444 1666
rect 15908 1658 15960 1666
rect 15360 1656 15960 1658
rect 14928 1648 15392 1656
rect 15444 1648 15908 1656
rect 14928 1476 15360 1648
rect 14876 1464 15360 1476
rect 16676 1656 16728 1666
rect 17192 1658 17244 1666
rect 17708 1658 17760 1666
rect 17160 1656 17760 1658
rect 16728 1648 17192 1656
rect 17244 1648 17708 1656
rect 16728 1476 17160 1648
rect 16676 1464 17160 1476
rect 18476 1656 18528 1666
rect 18992 1658 19044 1666
rect 19508 1658 19560 1666
rect 18960 1656 19560 1658
rect 18528 1648 18992 1656
rect 19044 1648 19508 1656
rect 18528 1476 18960 1648
rect 18476 1464 18960 1476
rect 20276 1656 20328 1666
rect 20792 1658 20844 1666
rect 21308 1658 21360 1666
rect 20760 1656 21360 1658
rect 20328 1648 20792 1656
rect 20844 1648 21308 1656
rect 20328 1476 20760 1648
rect 20276 1464 20760 1476
rect 960 1454 1560 1464
rect 2760 1454 3360 1464
rect 4560 1454 5160 1464
rect 6360 1454 6960 1464
rect 15360 1454 15960 1464
rect 17160 1454 17760 1464
rect 18960 1454 19560 1464
rect 20760 1454 21360 1464
rect -10060 1354 -9460 1356
rect -10060 1346 -10008 1354
rect -9544 1346 -9492 1354
rect -9028 1346 -8976 1356
rect -9800 1316 -9748 1326
rect -9284 1318 -9232 1326
rect -8768 1318 -8716 1326
rect -9316 1316 -8716 1318
rect -9748 1308 -9284 1316
rect -9232 1308 -8768 1316
rect -9748 1136 -9316 1308
rect -9800 1124 -9316 1136
rect -9316 1114 -8716 1124
rect 216 1268 816 1278
rect 2016 1268 2616 1278
rect 3816 1268 4416 1278
rect 5616 1268 6216 1278
rect 14616 1268 15216 1278
rect 16416 1268 17016 1278
rect 18216 1268 18816 1278
rect 20016 1268 20616 1278
rect 816 1256 1300 1268
rect 816 1084 1248 1256
rect 268 1076 732 1084
rect 784 1076 1248 1084
rect 216 1074 816 1076
rect 216 1066 268 1074
rect 732 1066 784 1074
rect 1248 1066 1300 1076
rect 2616 1256 3100 1268
rect 2616 1084 3048 1256
rect 2068 1076 2532 1084
rect 2584 1076 3048 1084
rect 2016 1074 2616 1076
rect 2016 1066 2068 1074
rect 2532 1066 2584 1074
rect 3048 1066 3100 1076
rect 4416 1256 4900 1268
rect 4416 1084 4848 1256
rect 3868 1076 4332 1084
rect 4384 1076 4848 1084
rect 3816 1074 4416 1076
rect 3816 1066 3868 1074
rect 4332 1066 4384 1074
rect 4848 1066 4900 1076
rect 6216 1256 6700 1268
rect 6216 1084 6648 1256
rect 5668 1076 6132 1084
rect 6184 1076 6648 1084
rect 5616 1074 6216 1076
rect 5616 1066 5668 1074
rect 6132 1066 6184 1074
rect 6648 1066 6700 1076
rect 15216 1256 15700 1268
rect 15216 1084 15648 1256
rect 14668 1076 15132 1084
rect 15184 1076 15648 1084
rect 14616 1074 15216 1076
rect 14616 1066 14668 1074
rect 15132 1066 15184 1074
rect 15648 1066 15700 1076
rect 17016 1256 17500 1268
rect 17016 1084 17448 1256
rect 16468 1076 16932 1084
rect 16984 1076 17448 1084
rect 16416 1074 17016 1076
rect 16416 1066 16468 1074
rect 16932 1066 16984 1074
rect 17448 1066 17500 1076
rect 18816 1256 19300 1268
rect 18816 1084 19248 1256
rect 18268 1076 18732 1084
rect 18784 1076 19248 1084
rect 18216 1074 18816 1076
rect 18216 1066 18268 1074
rect 18732 1066 18784 1074
rect 19248 1066 19300 1076
rect 20616 1256 21100 1268
rect 20616 1084 21048 1256
rect 20068 1076 20532 1084
rect 20584 1076 21048 1084
rect 20016 1074 20616 1076
rect 20016 1066 20068 1074
rect 20532 1066 20584 1074
rect 21048 1066 21100 1076
rect 476 1036 528 1046
rect 992 1038 1044 1046
rect 1508 1038 1560 1046
rect 960 1036 1560 1038
rect -10060 932 -9460 942
rect -9460 920 -8976 932
rect -9460 748 -9028 920
rect -10008 740 -9544 748
rect -9492 740 -9028 748
rect 528 1028 992 1036
rect 1044 1028 1508 1036
rect 528 856 960 1028
rect 476 844 960 856
rect 2276 1036 2328 1046
rect 2792 1038 2844 1046
rect 3308 1038 3360 1046
rect 2760 1036 3360 1038
rect 2328 1028 2792 1036
rect 2844 1028 3308 1036
rect 2328 856 2760 1028
rect 2276 844 2760 856
rect 4076 1036 4128 1046
rect 4592 1038 4644 1046
rect 5108 1038 5160 1046
rect 4560 1036 5160 1038
rect 4128 1028 4592 1036
rect 4644 1028 5108 1036
rect 4128 856 4560 1028
rect 4076 844 4560 856
rect 5876 1036 5928 1046
rect 6392 1038 6444 1046
rect 6908 1038 6960 1046
rect 6360 1036 6960 1038
rect 5928 1028 6392 1036
rect 6444 1028 6908 1036
rect 5928 856 6360 1028
rect 5876 844 6360 856
rect 14876 1036 14928 1046
rect 15392 1038 15444 1046
rect 15908 1038 15960 1046
rect 15360 1036 15960 1038
rect 14928 1028 15392 1036
rect 15444 1028 15908 1036
rect 14928 856 15360 1028
rect 14876 844 15360 856
rect 16676 1036 16728 1046
rect 17192 1038 17244 1046
rect 17708 1038 17760 1046
rect 17160 1036 17760 1038
rect 16728 1028 17192 1036
rect 17244 1028 17708 1036
rect 16728 856 17160 1028
rect 16676 844 17160 856
rect 18476 1036 18528 1046
rect 18992 1038 19044 1046
rect 19508 1038 19560 1046
rect 18960 1036 19560 1038
rect 18528 1028 18992 1036
rect 19044 1028 19508 1036
rect 18528 856 18960 1028
rect 18476 844 18960 856
rect 20276 1036 20328 1046
rect 20792 1038 20844 1046
rect 21308 1038 21360 1046
rect 20760 1036 21360 1038
rect 20328 1028 20792 1036
rect 20844 1028 21308 1036
rect 20328 856 20760 1028
rect 20276 844 20760 856
rect 960 834 1560 844
rect 2760 834 3360 844
rect 4560 834 5160 844
rect 6360 834 6960 844
rect 15360 834 15960 844
rect 17160 834 17760 844
rect 18960 834 19560 844
rect 20760 834 21360 844
rect -10060 738 -9460 740
rect -10060 730 -10008 738
rect -9544 730 -9492 738
rect -9028 730 -8976 740
rect -9800 700 -9748 710
rect -9284 702 -9232 710
rect -8768 702 -8716 710
rect -9316 700 -8716 702
rect -9748 692 -9284 700
rect -9232 692 -8768 700
rect -9748 520 -9316 692
rect -9800 508 -9316 520
rect 216 652 816 662
rect 2016 652 2616 662
rect 3816 652 4416 662
rect 5616 652 6216 662
rect 14616 652 15216 662
rect 16416 652 17016 662
rect 18216 652 18816 662
rect 20016 652 20616 662
rect 816 640 1300 652
rect -9316 498 -8716 508
rect -8500 508 -8360 518
rect 816 468 1248 640
rect 268 460 732 468
rect 784 460 1248 468
rect 216 458 816 460
rect 216 450 268 458
rect 732 450 784 458
rect 1248 450 1300 460
rect 2616 640 3100 652
rect 2616 468 3048 640
rect 2068 460 2532 468
rect 2584 460 3048 468
rect 2016 458 2616 460
rect 2016 450 2068 458
rect 2532 450 2584 458
rect 3048 450 3100 460
rect 4416 640 4900 652
rect 4416 468 4848 640
rect 3868 460 4332 468
rect 4384 460 4848 468
rect 3816 458 4416 460
rect 3816 450 3868 458
rect 4332 450 4384 458
rect 4848 450 4900 460
rect 6216 640 6700 652
rect 6216 468 6648 640
rect 5668 460 6132 468
rect 6184 460 6648 468
rect 5616 458 6216 460
rect 5616 450 5668 458
rect 6132 450 6184 458
rect 6648 450 6700 460
rect 15216 640 15700 652
rect 15216 468 15648 640
rect 14668 460 15132 468
rect 15184 460 15648 468
rect 14616 458 15216 460
rect 14616 450 14668 458
rect 15132 450 15184 458
rect 15648 450 15700 460
rect 17016 640 17500 652
rect 17016 468 17448 640
rect 16468 460 16932 468
rect 16984 460 17448 468
rect 16416 458 17016 460
rect 16416 450 16468 458
rect 16932 450 16984 458
rect 17448 450 17500 460
rect 18816 640 19300 652
rect 18816 468 19248 640
rect 18268 460 18732 468
rect 18784 460 19248 468
rect 18216 458 18816 460
rect 18216 450 18268 458
rect 18732 450 18784 458
rect 19248 450 19300 460
rect 20616 640 21100 652
rect 20616 468 21048 640
rect 20068 460 20532 468
rect 20584 460 21048 468
rect 20016 458 20616 460
rect 20016 450 20068 458
rect 20532 450 20584 458
rect 21048 450 21100 460
rect -8500 338 -8360 348
rect 476 420 528 430
rect 992 422 1044 430
rect 1508 422 1560 430
rect 960 420 1560 422
rect 528 412 992 420
rect 1044 412 1508 420
rect 528 240 960 412
rect 2276 420 2328 430
rect 2792 422 2844 430
rect 3308 422 3360 430
rect 2760 420 3360 422
rect 476 228 960 240
rect 960 218 1560 228
rect 1696 268 1876 278
rect 2328 412 2792 420
rect 2844 412 3308 420
rect 2328 240 2760 412
rect 4076 420 4128 430
rect 4592 422 4644 430
rect 5108 422 5160 430
rect 4560 420 5160 422
rect 2276 228 2760 240
rect 2760 218 3360 228
rect 3512 276 3692 286
rect 1696 58 1876 68
rect 4128 412 4592 420
rect 4644 412 5108 420
rect 4128 240 4560 412
rect 5876 420 5928 430
rect 6392 422 6444 430
rect 6908 422 6960 430
rect 6360 420 6960 422
rect 4076 228 4560 240
rect 4560 218 5160 228
rect 5288 276 5468 286
rect 3512 54 3692 64
rect 5928 412 6392 420
rect 6444 412 6908 420
rect 5928 240 6360 412
rect 5876 228 6360 240
rect 14876 420 14928 430
rect 15392 422 15444 430
rect 15908 422 15960 430
rect 15360 420 15960 422
rect 14928 412 15392 420
rect 15444 412 15908 420
rect 14928 240 15360 412
rect 16676 420 16728 430
rect 17192 422 17244 430
rect 17708 422 17760 430
rect 17160 420 17760 422
rect 14876 228 15360 240
rect 6360 218 6960 228
rect 15360 218 15960 228
rect 16096 268 16276 278
rect 5288 54 5468 64
rect 16728 412 17192 420
rect 17244 412 17708 420
rect 16728 240 17160 412
rect 18476 420 18528 430
rect 18992 422 19044 430
rect 19508 422 19560 430
rect 18960 420 19560 422
rect 16676 228 17160 240
rect 17160 218 17760 228
rect 17912 276 18092 286
rect 16096 58 16276 68
rect 18528 412 18992 420
rect 19044 412 19508 420
rect 18528 240 18960 412
rect 20276 420 20328 430
rect 20792 422 20844 430
rect 21308 422 21360 430
rect 20760 420 21360 422
rect 18476 228 18960 240
rect 18960 218 19560 228
rect 19688 276 19868 286
rect 17912 54 18092 64
rect 20328 412 20792 420
rect 20844 412 21308 420
rect 20328 240 20760 412
rect 20276 228 20760 240
rect 20760 218 21360 228
rect 19688 54 19868 64
rect -2768 -382 -1960 -372
rect -2768 -1198 -1960 -1188
rect 11632 -382 12440 -372
rect 11632 -1198 12440 -1188
<< via2 >>
rect 7440 27336 7540 27436
rect 7384 27092 8240 27172
rect 7384 26928 7580 27092
rect 7580 26928 7644 27092
rect 7644 26928 7896 27092
rect 7896 26928 7960 27092
rect 7960 26928 8240 27092
rect 9604 27092 10460 27172
rect 9604 26928 9800 27092
rect 9800 26928 9864 27092
rect 9864 26928 10116 27092
rect 10116 26928 10180 27092
rect 10180 26928 10460 27092
rect 11784 27092 12640 27172
rect 11784 26928 11980 27092
rect 11980 26928 12044 27092
rect 12044 26928 12296 27092
rect 12296 26928 12360 27092
rect 12360 26928 12640 27092
rect 13964 27092 14820 27172
rect 13964 26928 14160 27092
rect 14160 26928 14224 27092
rect 14224 26928 14476 27092
rect 14476 26928 14540 27092
rect 14540 26928 14820 27092
rect 16164 27092 17020 27172
rect 16164 26928 16360 27092
rect 16360 26928 16424 27092
rect 16424 26928 16676 27092
rect 16676 26928 16740 27092
rect 16740 26928 17020 27092
rect 6488 26688 6540 26852
rect 6540 26688 6792 26852
rect 6792 26688 6856 26852
rect 6856 26688 7108 26852
rect 7108 26688 7172 26852
rect 7172 26688 7268 26852
rect 6488 26608 7268 26688
rect 8708 26688 8760 26852
rect 8760 26688 9012 26852
rect 9012 26688 9076 26852
rect 9076 26688 9328 26852
rect 9328 26688 9392 26852
rect 9392 26688 9488 26852
rect 8708 26608 9488 26688
rect 10888 26688 10940 26852
rect 10940 26688 11192 26852
rect 11192 26688 11256 26852
rect 11256 26688 11508 26852
rect 11508 26688 11572 26852
rect 11572 26688 11668 26852
rect 10888 26608 11668 26688
rect 13068 26688 13120 26852
rect 13120 26688 13372 26852
rect 13372 26688 13436 26852
rect 13436 26688 13688 26852
rect 13688 26688 13752 26852
rect 13752 26688 13848 26852
rect 13068 26608 13848 26688
rect 15268 26688 15320 26852
rect 15320 26688 15572 26852
rect 15572 26688 15636 26852
rect 15636 26688 15888 26852
rect 15888 26688 15952 26852
rect 15952 26688 16048 26852
rect 15268 26608 16048 26688
rect 7384 26456 8240 26540
rect 7384 26296 7580 26456
rect 7580 26296 7644 26456
rect 7644 26296 7896 26456
rect 7896 26296 7960 26456
rect 7960 26296 8240 26456
rect 9604 26456 10460 26540
rect 9604 26296 9800 26456
rect 9800 26296 9864 26456
rect 9864 26296 10116 26456
rect 10116 26296 10180 26456
rect 10180 26296 10460 26456
rect 11784 26456 12640 26540
rect 11784 26296 11980 26456
rect 11980 26296 12044 26456
rect 12044 26296 12296 26456
rect 12296 26296 12360 26456
rect 12360 26296 12640 26456
rect 13964 26456 14820 26540
rect 13964 26296 14160 26456
rect 14160 26296 14224 26456
rect 14224 26296 14476 26456
rect 14476 26296 14540 26456
rect 14540 26296 14820 26456
rect 16164 26456 17020 26540
rect 16164 26296 16360 26456
rect 16360 26296 16424 26456
rect 16424 26296 16676 26456
rect 16676 26296 16740 26456
rect 16740 26296 17020 26456
rect 6488 26052 6540 26216
rect 6540 26052 6792 26216
rect 6792 26052 6856 26216
rect 6856 26052 7108 26216
rect 7108 26052 7172 26216
rect 7172 26052 7268 26216
rect 6488 25972 7268 26052
rect 8708 26052 8760 26216
rect 8760 26052 9012 26216
rect 9012 26052 9076 26216
rect 9076 26052 9328 26216
rect 9328 26052 9392 26216
rect 9392 26052 9488 26216
rect 8708 25972 9488 26052
rect 10888 26052 10940 26216
rect 10940 26052 11192 26216
rect 11192 26052 11256 26216
rect 11256 26052 11508 26216
rect 11508 26052 11572 26216
rect 11572 26052 11668 26216
rect 10888 25972 11668 26052
rect 13068 26052 13120 26216
rect 13120 26052 13372 26216
rect 13372 26052 13436 26216
rect 13436 26052 13688 26216
rect 13688 26052 13752 26216
rect 13752 26052 13848 26216
rect 13068 25972 13848 26052
rect 15268 26052 15320 26216
rect 15320 26052 15572 26216
rect 15572 26052 15636 26216
rect 15636 26052 15888 26216
rect 15888 26052 15952 26216
rect 15952 26052 16048 26216
rect 15268 25972 16048 26052
rect 7384 25816 8240 25904
rect 7384 25660 7580 25816
rect 7580 25660 7644 25816
rect 7644 25660 7896 25816
rect 7896 25660 7960 25816
rect 7960 25660 8240 25816
rect 9604 25816 10460 25904
rect 9604 25660 9800 25816
rect 9800 25660 9864 25816
rect 9864 25660 10116 25816
rect 10116 25660 10180 25816
rect 10180 25660 10460 25816
rect 11784 25816 12640 25904
rect 11784 25660 11980 25816
rect 11980 25660 12044 25816
rect 12044 25660 12296 25816
rect 12296 25660 12360 25816
rect 12360 25660 12640 25816
rect 13964 25816 14820 25904
rect 13964 25660 14160 25816
rect 14160 25660 14224 25816
rect 14224 25660 14476 25816
rect 14476 25660 14540 25816
rect 14540 25660 14820 25816
rect 16164 25816 17020 25904
rect 16164 25660 16360 25816
rect 16360 25660 16424 25816
rect 16424 25660 16676 25816
rect 16676 25660 16740 25816
rect 16740 25660 17020 25816
rect 6488 25412 6540 25576
rect 6540 25412 6792 25576
rect 6792 25412 6856 25576
rect 6856 25412 7108 25576
rect 7108 25412 7172 25576
rect 7172 25412 7268 25576
rect 6488 25332 7268 25412
rect 8708 25412 8760 25576
rect 8760 25412 9012 25576
rect 9012 25412 9076 25576
rect 9076 25412 9328 25576
rect 9328 25412 9392 25576
rect 9392 25412 9488 25576
rect 8708 25332 9488 25412
rect 10888 25412 10940 25576
rect 10940 25412 11192 25576
rect 11192 25412 11256 25576
rect 11256 25412 11508 25576
rect 11508 25412 11572 25576
rect 11572 25412 11668 25576
rect 10888 25332 11668 25412
rect 13068 25412 13120 25576
rect 13120 25412 13372 25576
rect 13372 25412 13436 25576
rect 13436 25412 13688 25576
rect 13688 25412 13752 25576
rect 13752 25412 13848 25576
rect 13068 25332 13848 25412
rect 15268 25412 15320 25576
rect 15320 25412 15572 25576
rect 15572 25412 15636 25576
rect 15636 25412 15888 25576
rect 15888 25412 15952 25576
rect 15952 25412 16048 25576
rect 15268 25332 16048 25412
rect 6492 24992 7276 25076
rect 6492 24828 6572 24992
rect 6572 24828 6636 24992
rect 6636 24828 6764 24992
rect 6764 24828 6828 24992
rect 6828 24828 6956 24992
rect 6956 24828 7020 24992
rect 7020 24828 7148 24992
rect 7148 24828 7212 24992
rect 7212 24828 7276 24992
rect 8712 24992 9496 25076
rect 10892 24992 11676 25076
rect 13072 24992 13856 25076
rect 15272 24992 16056 25076
rect 8712 24828 8792 24992
rect 8792 24828 8856 24992
rect 8856 24828 8984 24992
rect 8984 24828 9048 24992
rect 9048 24828 9176 24992
rect 9176 24828 9240 24992
rect 9240 24828 9368 24992
rect 9368 24828 9432 24992
rect 9432 24828 9496 24992
rect 10892 24828 10972 24992
rect 10972 24828 11036 24992
rect 11036 24828 11164 24992
rect 11164 24828 11228 24992
rect 11228 24828 11356 24992
rect 11356 24828 11420 24992
rect 11420 24828 11548 24992
rect 11548 24828 11612 24992
rect 11612 24828 11676 24992
rect 13072 24828 13152 24992
rect 13152 24828 13216 24992
rect 13216 24828 13344 24992
rect 13344 24828 13408 24992
rect 13408 24828 13536 24992
rect 13536 24828 13600 24992
rect 13600 24828 13728 24992
rect 13728 24828 13792 24992
rect 13792 24828 13856 24992
rect 15272 24828 15352 24992
rect 15352 24828 15416 24992
rect 15416 24828 15544 24992
rect 15544 24828 15608 24992
rect 15608 24828 15736 24992
rect 15736 24828 15800 24992
rect 15800 24828 15928 24992
rect 15928 24828 15992 24992
rect 15992 24828 16056 24992
rect 7388 24588 7436 24748
rect 7436 24588 7500 24748
rect 7500 24588 7628 24748
rect 7628 24588 7692 24748
rect 7692 24588 7820 24748
rect 7820 24588 7884 24748
rect 7884 24588 8240 24748
rect 7388 24508 8240 24588
rect 9608 24588 9656 24748
rect 9656 24588 9720 24748
rect 9720 24588 9848 24748
rect 9848 24588 9912 24748
rect 9912 24588 10040 24748
rect 10040 24588 10104 24748
rect 10104 24588 10460 24748
rect 9608 24508 10460 24588
rect 11788 24588 11836 24748
rect 11836 24588 11900 24748
rect 11900 24588 12028 24748
rect 12028 24588 12092 24748
rect 12092 24588 12220 24748
rect 12220 24588 12284 24748
rect 12284 24588 12640 24748
rect 11788 24508 12640 24588
rect 13968 24588 14016 24748
rect 14016 24588 14080 24748
rect 14080 24588 14208 24748
rect 14208 24588 14272 24748
rect 14272 24588 14400 24748
rect 14400 24588 14464 24748
rect 14464 24588 14820 24748
rect 13968 24508 14820 24588
rect 16168 24588 16216 24748
rect 16216 24588 16280 24748
rect 16280 24588 16408 24748
rect 16408 24588 16472 24748
rect 16472 24588 16600 24748
rect 16600 24588 16664 24748
rect 16664 24588 17020 24748
rect 18280 24600 18640 25120
rect 16168 24508 17020 24588
rect 6492 24356 7276 24436
rect 6492 24188 6572 24356
rect 6572 24188 6636 24356
rect 6636 24188 6764 24356
rect 6764 24188 6828 24356
rect 6828 24188 6956 24356
rect 6956 24188 7020 24356
rect 7020 24188 7148 24356
rect 7148 24188 7212 24356
rect 7212 24188 7276 24356
rect 8156 24212 8328 24436
rect 8712 24356 9496 24436
rect 8712 24188 8792 24356
rect 8792 24188 8856 24356
rect 8856 24188 8984 24356
rect 8984 24188 9048 24356
rect 9048 24188 9176 24356
rect 9176 24188 9240 24356
rect 9240 24188 9368 24356
rect 9368 24188 9432 24356
rect 9432 24188 9496 24356
rect 10892 24356 11676 24436
rect 10892 24188 10972 24356
rect 10972 24188 11036 24356
rect 11036 24188 11164 24356
rect 11164 24188 11228 24356
rect 11228 24188 11356 24356
rect 11356 24188 11420 24356
rect 11420 24188 11548 24356
rect 11548 24188 11612 24356
rect 11612 24188 11676 24356
rect 13072 24356 13856 24436
rect 13072 24188 13152 24356
rect 13152 24188 13216 24356
rect 13216 24188 13344 24356
rect 13344 24188 13408 24356
rect 13408 24188 13536 24356
rect 13536 24188 13600 24356
rect 13600 24188 13728 24356
rect 13728 24188 13792 24356
rect 13792 24188 13856 24356
rect 15272 24356 16056 24436
rect 15272 24188 15352 24356
rect 15352 24188 15416 24356
rect 15416 24188 15544 24356
rect 15544 24188 15608 24356
rect 15608 24188 15736 24356
rect 15736 24188 15800 24356
rect 15800 24188 15928 24356
rect 15928 24188 15992 24356
rect 15992 24188 16056 24356
rect 7388 23952 7436 24116
rect 7436 23952 7500 24116
rect 7500 23952 7628 24116
rect 7628 23952 7692 24116
rect 7692 23952 7820 24116
rect 7820 23952 7884 24116
rect 7884 23952 8240 24116
rect 7388 23876 8240 23952
rect 9608 23952 9656 24116
rect 9656 23952 9720 24116
rect 9720 23952 9848 24116
rect 9848 23952 9912 24116
rect 9912 23952 10040 24116
rect 10040 23952 10104 24116
rect 10104 23952 10460 24116
rect 9608 23876 10460 23952
rect 11788 23952 11836 24116
rect 11836 23952 11900 24116
rect 11900 23952 12028 24116
rect 12028 23952 12092 24116
rect 12092 23952 12220 24116
rect 12220 23952 12284 24116
rect 12284 23952 12640 24116
rect 11788 23876 12640 23952
rect 13968 23952 14016 24116
rect 14016 23952 14080 24116
rect 14080 23952 14208 24116
rect 14208 23952 14272 24116
rect 14272 23952 14400 24116
rect 14400 23952 14464 24116
rect 14464 23952 14820 24116
rect 13968 23876 14820 23952
rect 16168 23952 16216 24116
rect 16216 23952 16280 24116
rect 16280 23952 16408 24116
rect 16408 23952 16472 24116
rect 16472 23952 16600 24116
rect 16600 23952 16664 24116
rect 16664 23952 17020 24116
rect 16168 23876 17020 23952
rect 7408 23424 8236 23680
rect 7408 23272 7464 23424
rect 7464 23272 7516 23424
rect 7516 23272 8236 23424
rect 6596 23020 6600 23192
rect 6600 23020 6652 23192
rect 6652 23020 6792 23192
rect 6792 23020 6844 23192
rect 6844 23020 6984 23192
rect 6984 23020 7036 23192
rect 7036 23020 7176 23192
rect 7176 23020 7200 23192
rect 6596 23008 7200 23020
rect 8316 23020 8320 23192
rect 8320 23020 8372 23192
rect 8372 23020 8512 23192
rect 8512 23020 8564 23192
rect 8564 23020 8704 23192
rect 8704 23020 8756 23192
rect 8756 23020 8896 23192
rect 8896 23020 8920 23192
rect 8316 23008 8920 23020
rect 6596 22404 6600 22576
rect 6600 22404 6652 22576
rect 6652 22404 6792 22576
rect 6792 22404 6844 22576
rect 6844 22404 6984 22576
rect 6984 22404 7036 22576
rect 7036 22404 7176 22576
rect 7176 22404 7200 22576
rect 6596 22392 7200 22404
rect 8316 22404 8320 22576
rect 8320 22404 8372 22576
rect 8372 22404 8512 22576
rect 8512 22404 8564 22576
rect 8564 22404 8704 22576
rect 8704 22404 8756 22576
rect 8756 22404 8896 22576
rect 8896 22404 8920 22576
rect 8316 22392 8920 22404
rect 19044 23364 19232 23448
rect 18272 22620 18300 22784
rect 18300 22620 18352 22784
rect 18352 22620 18492 22784
rect 18492 22620 18544 22784
rect 18544 22620 18684 22784
rect 18684 22620 18736 22784
rect 18736 22620 18860 22784
rect 18272 22572 18860 22620
rect 18272 22484 18860 22572
rect 6592 21784 6600 21956
rect 6600 21784 6652 21956
rect 6652 21784 6792 21956
rect 6792 21784 6844 21956
rect 6844 21784 6984 21956
rect 6984 21784 7036 21956
rect 7036 21784 7176 21956
rect 7176 21784 7196 21956
rect 6592 21772 7196 21784
rect 8312 21784 8320 21956
rect 8320 21784 8372 21956
rect 8372 21784 8512 21956
rect 8512 21784 8564 21956
rect 8564 21784 8704 21956
rect 8704 21784 8756 21956
rect 8756 21784 8896 21956
rect 8896 21784 8916 21956
rect 8312 21772 8916 21784
rect 15900 21740 16300 22180
rect 18284 22168 18864 22228
rect 18284 21996 18392 22168
rect 18392 21996 18444 22168
rect 18444 21996 18584 22168
rect 18584 21996 18636 22168
rect 18636 21996 18776 22168
rect 18776 21996 18828 22168
rect 18828 21996 18864 22168
rect 18996 21764 19064 21916
rect 19064 21764 19116 21916
rect 19116 21764 19256 21916
rect 19256 21764 19308 21916
rect 19308 21764 19628 21916
rect 18996 21688 19628 21764
rect 18284 21548 18864 21616
rect 18284 21384 18396 21548
rect 18396 21384 18448 21548
rect 18448 21384 18588 21548
rect 18588 21384 18640 21548
rect 18640 21384 18780 21548
rect 18780 21384 18832 21548
rect 18832 21384 18864 21548
rect 6600 21276 7200 21288
rect 8320 21276 8920 21288
rect 6600 21104 6652 21276
rect 6652 21104 7116 21276
rect 7116 21104 7168 21276
rect 7168 21104 7200 21276
rect 8320 21104 8372 21276
rect 8372 21104 8836 21276
rect 8836 21104 8888 21276
rect 8888 21104 8920 21276
rect 7344 20876 7376 21048
rect 7376 20876 7428 21048
rect 7428 20876 7892 21048
rect 7892 20876 7944 21048
rect 7344 20864 7944 20876
rect 9064 20876 9096 21048
rect 9096 20876 9148 21048
rect 9148 20876 9612 21048
rect 9612 20876 9664 21048
rect 9064 20864 9664 20876
rect 10380 20860 10840 21220
rect 19000 21144 19068 21320
rect 19068 21144 19120 21320
rect 19120 21144 19260 21320
rect 19260 21144 19312 21320
rect 19312 21144 19632 21320
rect 19000 21092 19632 21144
rect 24560 21140 24880 21500
rect 18996 20684 19628 20752
rect 6600 20660 7200 20672
rect 6600 20488 6652 20660
rect 6652 20488 7116 20660
rect 7116 20488 7168 20660
rect 7168 20488 7200 20660
rect 8320 20660 8920 20672
rect 8320 20488 8372 20660
rect 8372 20488 8836 20660
rect 8836 20488 8888 20660
rect 8888 20488 8920 20660
rect 18996 20524 19076 20684
rect 19076 20524 19128 20684
rect 19128 20524 19592 20684
rect 19592 20524 19628 20684
rect 7344 20260 7376 20432
rect 7376 20260 7428 20432
rect 7428 20260 7892 20432
rect 7892 20260 7944 20432
rect 7344 20248 7944 20260
rect 9064 20260 9096 20432
rect 9096 20260 9148 20432
rect 9148 20260 9612 20432
rect 9612 20260 9664 20432
rect 9064 20248 9664 20260
rect 18308 20280 18352 20448
rect 18352 20280 18816 20448
rect 18816 20280 18868 20448
rect 18868 20280 18888 20448
rect 18308 20220 18888 20280
rect 18996 20064 19628 20128
rect 6600 20040 7200 20052
rect 6600 19868 6652 20040
rect 6652 19868 7116 20040
rect 7116 19868 7168 20040
rect 7168 19868 7200 20040
rect 8320 20040 8920 20052
rect 8320 19868 8372 20040
rect 8372 19868 8836 20040
rect 8836 19868 8888 20040
rect 8888 19868 8920 20040
rect 18996 19900 19076 20064
rect 19076 19900 19128 20064
rect 19128 19900 19592 20064
rect 19592 19900 19628 20064
rect 7344 19640 7376 19812
rect 7376 19640 7428 19812
rect 7428 19640 7892 19812
rect 7892 19640 7944 19812
rect 7344 19628 7944 19640
rect 9064 19640 9096 19812
rect 9096 19640 9148 19812
rect 9148 19640 9612 19812
rect 9612 19640 9664 19812
rect 9064 19628 9664 19640
rect 10276 19728 10876 19868
rect 10276 19580 10312 19728
rect 10312 19580 10444 19728
rect 10444 19580 10504 19728
rect 10504 19580 10636 19728
rect 10636 19580 10696 19728
rect 10696 19580 10828 19728
rect 10828 19580 10876 19728
rect 18308 19660 18352 19828
rect 18352 19660 18816 19828
rect 18816 19660 18868 19828
rect 18868 19660 18888 19828
rect 18308 19600 18888 19660
rect 6600 19424 7200 19436
rect 6600 19252 6652 19424
rect 6652 19252 7116 19424
rect 7116 19252 7168 19424
rect 7168 19252 7200 19424
rect 8320 19424 8920 19436
rect 8320 19252 8372 19424
rect 8372 19252 8836 19424
rect 8836 19252 8888 19424
rect 8888 19252 8920 19424
rect 10024 19324 10160 19468
rect 10160 19324 10220 19468
rect 10220 19324 10348 19468
rect 10348 19324 10408 19468
rect 10408 19324 10540 19468
rect 10540 19324 10600 19468
rect 10600 19324 10640 19468
rect 7344 19024 7376 19196
rect 7376 19024 7428 19196
rect 7428 19024 7892 19196
rect 7892 19024 7944 19196
rect 7344 19012 7944 19024
rect 9064 19024 9096 19196
rect 9096 19024 9148 19196
rect 9148 19024 9612 19196
rect 9612 19024 9664 19196
rect 10024 19172 10640 19324
rect 18996 19448 19628 19512
rect 18996 19284 19076 19448
rect 19076 19284 19128 19448
rect 19128 19284 19592 19448
rect 19592 19284 19628 19448
rect 9064 19012 9664 19024
rect 18308 19044 18352 19212
rect 18352 19044 18816 19212
rect 18816 19044 18868 19212
rect 18868 19044 18888 19212
rect 18308 18984 18888 19044
rect 6600 18804 7200 18816
rect 6600 18632 6652 18804
rect 6652 18632 7116 18804
rect 7116 18632 7168 18804
rect 7168 18632 7200 18804
rect 8320 18804 8920 18816
rect 8320 18632 8372 18804
rect 8372 18632 8836 18804
rect 8836 18632 8888 18804
rect 8888 18632 8920 18804
rect 10040 18804 10624 18876
rect 10040 18644 10252 18804
rect 10252 18644 10312 18804
rect 10312 18644 10444 18804
rect 10444 18644 10504 18804
rect 10504 18644 10624 18804
rect 7344 18404 7376 18576
rect 7376 18404 7428 18576
rect 7428 18404 7892 18576
rect 7892 18404 7944 18576
rect 7344 18392 7944 18404
rect 9064 18404 9096 18576
rect 9096 18404 9148 18576
rect 9148 18404 9612 18576
rect 9612 18404 9664 18576
rect 9064 18392 9664 18404
rect 10768 18404 10792 18560
rect 10792 18404 10924 18560
rect 10924 18404 10984 18560
rect 10984 18404 11116 18560
rect 11116 18404 11176 18560
rect 11176 18404 11296 18560
rect 15580 18420 15980 18860
rect 10768 18336 11296 18404
rect 6600 18188 7200 18200
rect 6600 18016 6652 18188
rect 6652 18016 7116 18188
rect 7116 18016 7168 18188
rect 7168 18016 7200 18188
rect 8320 18188 8920 18200
rect 8320 18016 8372 18188
rect 8372 18016 8836 18188
rect 8836 18016 8888 18188
rect 8888 18016 8920 18188
rect 10040 18188 10624 18256
rect 10040 18032 10252 18188
rect 10252 18032 10312 18188
rect 10312 18032 10444 18188
rect 10444 18032 10504 18188
rect 10504 18032 10624 18188
rect 7344 17788 7376 17960
rect 7376 17788 7428 17960
rect 7428 17788 7892 17960
rect 7892 17788 7944 17960
rect 7344 17776 7944 17788
rect 9064 17788 9096 17960
rect 9096 17788 9148 17960
rect 9148 17788 9612 17960
rect 9612 17788 9664 17960
rect 9064 17776 9664 17788
rect 8040 17616 8220 17776
rect 10764 17784 10792 17940
rect 10792 17784 10924 17940
rect 10924 17784 10984 17940
rect 10984 17784 11116 17940
rect 11116 17784 11176 17940
rect 11176 17784 11292 17940
rect 10764 17716 11292 17784
rect 16220 18420 16620 18860
rect 19000 18828 19632 18916
rect 19000 18688 19076 18828
rect 19076 18688 19128 18828
rect 19128 18688 19592 18828
rect 19592 18688 19632 18828
rect 1300 10532 1568 10768
rect 2588 10660 4792 11148
rect 6096 10608 6276 10808
rect 15700 10532 15968 10768
rect 6212 10284 7188 10364
rect 6212 10120 6228 10284
rect 6228 10120 6364 10284
rect 6364 10120 6420 10284
rect 6420 10120 6556 10284
rect 6556 10120 6612 10284
rect 6612 10120 6748 10284
rect 6748 10120 6804 10284
rect 6804 10120 6940 10284
rect 6940 10120 6996 10284
rect 6996 10120 7188 10284
rect 8760 10264 9632 10292
rect 8760 10092 8864 10264
rect 8864 10092 8920 10264
rect 8920 10092 9056 10264
rect 9056 10092 9112 10264
rect 9112 10092 9248 10264
rect 9248 10092 9304 10264
rect 9304 10092 9440 10264
rect 9440 10092 9496 10264
rect 9496 10092 9632 10264
rect 5112 9880 5116 10052
rect 5116 9880 5172 10052
rect 5172 9880 5308 10052
rect 5308 9880 5364 10052
rect 5364 9880 5500 10052
rect 5500 9880 5556 10052
rect 5556 9880 5692 10052
rect 5692 9880 5748 10052
rect 5748 9880 5884 10052
rect 5884 9880 5940 10052
rect 5940 9880 6076 10052
rect 6076 9880 6088 10052
rect 5112 9796 6088 9880
rect 7608 9860 7616 10032
rect 7616 9860 7672 10032
rect 7672 9860 7808 10032
rect 7808 9860 7864 10032
rect 7864 9860 8000 10032
rect 8000 9860 8056 10032
rect 8056 9860 8192 10032
rect 8192 9860 8248 10032
rect 8248 9860 8384 10032
rect 8384 9860 8440 10032
rect 8440 9860 8576 10032
rect 8576 9860 8592 10032
rect 7608 9844 8592 9860
rect 18308 18424 18352 18592
rect 18352 18424 18816 18592
rect 18816 18424 18868 18592
rect 18868 18424 18888 18592
rect 18308 18364 18888 18424
rect 18480 18056 18680 18156
rect 16988 10660 19192 11148
rect 20496 10608 20676 10808
rect 20612 10284 21588 10364
rect 20612 10120 20628 10284
rect 20628 10120 20764 10284
rect 20764 10120 20820 10284
rect 20820 10120 20956 10284
rect 20956 10120 21012 10284
rect 21012 10120 21148 10284
rect 21148 10120 21204 10284
rect 21204 10120 21340 10284
rect 21340 10120 21396 10284
rect 21396 10120 21588 10284
rect 23160 10264 24032 10292
rect 23160 10092 23264 10264
rect 23264 10092 23320 10264
rect 23320 10092 23456 10264
rect 23456 10092 23512 10264
rect 23512 10092 23648 10264
rect 23648 10092 23704 10264
rect 23704 10092 23840 10264
rect 23840 10092 23896 10264
rect 23896 10092 24032 10264
rect 6212 9652 7188 9732
rect 6212 9488 6228 9652
rect 6228 9488 6364 9652
rect 6364 9488 6420 9652
rect 6420 9488 6556 9652
rect 6556 9488 6612 9652
rect 6612 9488 6748 9652
rect 6748 9488 6804 9652
rect 6804 9488 6940 9652
rect 6940 9488 6996 9652
rect 6996 9488 7188 9652
rect 8764 9648 9636 9676
rect 8764 9476 8864 9648
rect 8864 9476 8920 9648
rect 8920 9476 9056 9648
rect 9056 9476 9112 9648
rect 9112 9476 9248 9648
rect 9248 9476 9304 9648
rect 9304 9476 9440 9648
rect 9440 9476 9496 9648
rect 9496 9476 9636 9648
rect 19512 9880 19516 10052
rect 19516 9880 19572 10052
rect 19572 9880 19708 10052
rect 19708 9880 19764 10052
rect 19764 9880 19900 10052
rect 19900 9880 19956 10052
rect 19956 9880 20092 10052
rect 20092 9880 20148 10052
rect 20148 9880 20284 10052
rect 20284 9880 20340 10052
rect 20340 9880 20476 10052
rect 20476 9880 20488 10052
rect 19512 9796 20488 9880
rect 22008 9860 22016 10032
rect 22016 9860 22072 10032
rect 22072 9860 22208 10032
rect 22208 9860 22264 10032
rect 22264 9860 22400 10032
rect 22400 9860 22456 10032
rect 22456 9860 22592 10032
rect 22592 9860 22648 10032
rect 22648 9860 22784 10032
rect 22784 9860 22840 10032
rect 22840 9860 22976 10032
rect 22976 9860 22992 10032
rect 22008 9844 22992 9860
rect 20612 9652 21588 9732
rect 20612 9488 20628 9652
rect 20628 9488 20764 9652
rect 20764 9488 20820 9652
rect 20820 9488 20956 9652
rect 20956 9488 21012 9652
rect 21012 9488 21148 9652
rect 21148 9488 21204 9652
rect 21204 9488 21340 9652
rect 21340 9488 21396 9652
rect 21396 9488 21588 9652
rect 23164 9648 24036 9676
rect 23164 9476 23264 9648
rect 23264 9476 23320 9648
rect 23320 9476 23456 9648
rect 23456 9476 23512 9648
rect 23512 9476 23648 9648
rect 23648 9476 23704 9648
rect 23704 9476 23840 9648
rect 23840 9476 23896 9648
rect 23896 9476 24036 9648
rect 5112 9248 5116 9420
rect 5116 9248 5172 9420
rect 5172 9248 5308 9420
rect 5308 9248 5364 9420
rect 5364 9248 5500 9420
rect 5500 9248 5556 9420
rect 5556 9248 5692 9420
rect 5692 9248 5748 9420
rect 5748 9248 5884 9420
rect 5884 9248 5940 9420
rect 5940 9248 6076 9420
rect 6076 9248 6088 9420
rect 5112 9160 6088 9248
rect 7612 9244 7616 9412
rect 7616 9244 7672 9412
rect 7672 9244 7808 9412
rect 7808 9244 7864 9412
rect 7864 9244 8000 9412
rect 8000 9244 8056 9412
rect 8056 9244 8192 9412
rect 8192 9244 8248 9412
rect 8248 9244 8384 9412
rect 8384 9244 8440 9412
rect 8440 9244 8576 9412
rect 8576 9244 8596 9412
rect 7612 9224 8596 9244
rect 19512 9248 19516 9420
rect 19516 9248 19572 9420
rect 19572 9248 19708 9420
rect 19708 9248 19764 9420
rect 19764 9248 19900 9420
rect 19900 9248 19956 9420
rect 19956 9248 20092 9420
rect 20092 9248 20148 9420
rect 20148 9248 20284 9420
rect 20284 9248 20340 9420
rect 20340 9248 20476 9420
rect 20476 9248 20488 9420
rect 19512 9160 20488 9248
rect 22012 9244 22016 9412
rect 22016 9244 22072 9412
rect 22072 9244 22208 9412
rect 22208 9244 22264 9412
rect 22264 9244 22400 9412
rect 22400 9244 22456 9412
rect 22456 9244 22592 9412
rect 22592 9244 22648 9412
rect 22648 9244 22784 9412
rect 22784 9244 22840 9412
rect 22840 9244 22976 9412
rect 22976 9244 22996 9412
rect 22012 9224 22996 9244
rect 8764 9028 9636 9060
rect -8660 8196 -8480 8296
rect 4588 8432 5008 8984
rect 8764 8860 8864 9028
rect 8864 8860 8920 9028
rect 8920 8860 9056 9028
rect 9056 8860 9112 9028
rect 9112 8860 9248 9028
rect 9248 8860 9304 9028
rect 9304 8860 9440 9028
rect 9440 8860 9496 9028
rect 9496 8860 9636 9028
rect 6224 8700 7200 8784
rect 6224 8536 6228 8700
rect 6228 8536 6364 8700
rect 6364 8536 6420 8700
rect 6420 8536 6556 8700
rect 6556 8536 6612 8700
rect 6612 8536 6748 8700
rect 6748 8536 6804 8700
rect 6804 8536 6940 8700
rect 6940 8536 6996 8700
rect 6996 8536 7200 8700
rect 7608 8624 7616 8796
rect 7616 8624 7672 8796
rect 7672 8624 7808 8796
rect 7808 8624 7864 8796
rect 7864 8624 8000 8796
rect 8000 8624 8056 8796
rect 8056 8624 8192 8796
rect 8192 8624 8248 8796
rect 8248 8624 8384 8796
rect 8384 8624 8440 8796
rect 8440 8624 8576 8796
rect 8576 8624 8592 8796
rect 7608 8608 8592 8624
rect 23164 9028 24036 9060
rect -9968 7832 -9868 7852
rect -9868 7832 -9816 7852
rect -9816 7832 -9676 7852
rect -9676 7832 -9624 7852
rect -9624 7832 -9484 7852
rect -9484 7832 -9432 7852
rect -9432 7832 -9316 7852
rect -9968 7620 -9316 7832
rect -9968 7584 -9964 7620
rect -9964 7584 -9912 7620
rect -9912 7584 -9772 7620
rect -9772 7584 -9720 7620
rect -9720 7584 -9580 7620
rect -9580 7584 -9528 7620
rect -9528 7584 -9388 7620
rect -9388 7584 -9336 7620
rect -9336 7584 -9316 7620
rect -9968 6596 -9868 6740
rect -9868 6596 -9816 6740
rect -9816 6596 -9676 6740
rect -9676 6596 -9624 6740
rect -9624 6596 -9484 6740
rect -9484 6596 -9432 6740
rect -9432 6596 -9316 6740
rect -9968 6472 -9316 6596
rect 5104 8296 5116 8472
rect 5116 8296 5172 8472
rect 5172 8296 5308 8472
rect 5308 8296 5364 8472
rect 5364 8296 5500 8472
rect 5500 8296 5556 8472
rect 5556 8296 5692 8472
rect 5692 8296 5748 8472
rect 5748 8296 5884 8472
rect 5884 8296 5940 8472
rect 5940 8296 6076 8472
rect 6076 8296 6080 8472
rect 5104 8224 6080 8296
rect 8764 8412 9636 8440
rect 8764 8240 8864 8412
rect 8864 8240 8920 8412
rect 8920 8240 9056 8412
rect 9056 8240 9112 8412
rect 9112 8240 9248 8412
rect 9248 8240 9304 8412
rect 9304 8240 9440 8412
rect 9440 8240 9496 8412
rect 9496 8240 9636 8412
rect 18988 8432 19408 8984
rect 23164 8860 23264 9028
rect 23264 8860 23320 9028
rect 23320 8860 23456 9028
rect 23456 8860 23512 9028
rect 23512 8860 23648 9028
rect 23648 8860 23704 9028
rect 23704 8860 23840 9028
rect 23840 8860 23896 9028
rect 23896 8860 24036 9028
rect 20624 8700 21600 8784
rect 20624 8536 20628 8700
rect 20628 8536 20764 8700
rect 20764 8536 20820 8700
rect 20820 8536 20956 8700
rect 20956 8536 21012 8700
rect 21012 8536 21148 8700
rect 21148 8536 21204 8700
rect 21204 8536 21340 8700
rect 21340 8536 21396 8700
rect 21396 8536 21600 8700
rect 22008 8624 22016 8796
rect 22016 8624 22072 8796
rect 22072 8624 22208 8796
rect 22208 8624 22264 8796
rect 22264 8624 22400 8796
rect 22400 8624 22456 8796
rect 22456 8624 22592 8796
rect 22592 8624 22648 8796
rect 22648 8624 22784 8796
rect 22784 8624 22840 8796
rect 22840 8624 22976 8796
rect 22976 8624 22992 8796
rect 22008 8608 22992 8624
rect 6224 8080 7200 8164
rect 6224 7916 6228 8080
rect 6228 7916 6364 8080
rect 6364 7916 6420 8080
rect 6420 7916 6556 8080
rect 6556 7916 6612 8080
rect 6612 7916 6748 8080
rect 6748 7916 6804 8080
rect 6804 7916 6940 8080
rect 6940 7916 6996 8080
rect 6996 7916 7200 8080
rect 7604 8008 7616 8180
rect 7616 8008 7672 8180
rect 7672 8008 7808 8180
rect 7808 8008 7864 8180
rect 7864 8008 8000 8180
rect 8000 8008 8056 8180
rect 8056 8008 8192 8180
rect 8192 8008 8248 8180
rect 8248 8008 8384 8180
rect 8384 8008 8440 8180
rect 8440 8008 8576 8180
rect 8576 8008 8588 8180
rect 7604 7992 8588 8008
rect 5104 7676 5116 7848
rect 5116 7676 5172 7848
rect 5172 7676 5308 7848
rect 5308 7676 5364 7848
rect 5364 7676 5500 7848
rect 5500 7676 5556 7848
rect 5556 7676 5692 7848
rect 5692 7676 5748 7848
rect 5748 7676 5884 7848
rect 5884 7676 5940 7848
rect 5940 7676 6076 7848
rect 6076 7676 6080 7848
rect 5104 7600 6080 7676
rect 8764 7792 9636 7820
rect 8764 7620 8864 7792
rect 8864 7620 8920 7792
rect 8920 7620 9056 7792
rect 9056 7620 9112 7792
rect 9112 7620 9248 7792
rect 9248 7620 9304 7792
rect 9304 7620 9440 7792
rect 9440 7620 9496 7792
rect 9496 7620 9636 7792
rect 6384 7000 7076 7512
rect 7608 7388 7616 7556
rect 7616 7388 7672 7556
rect 7672 7388 7808 7556
rect 7808 7388 7864 7556
rect 7864 7388 8000 7556
rect 8000 7388 8056 7556
rect 8056 7388 8192 7556
rect 8192 7388 8248 7556
rect 8248 7388 8384 7556
rect 8384 7388 8440 7556
rect 8440 7388 8576 7556
rect 8576 7388 8592 7556
rect 7608 7368 8592 7388
rect 8764 7176 9636 7204
rect 8764 7004 8864 7176
rect 8864 7004 8920 7176
rect 8920 7004 9056 7176
rect 9056 7004 9112 7176
rect 9112 7004 9248 7176
rect 9248 7004 9304 7176
rect 9304 7004 9440 7176
rect 9440 7004 9496 7176
rect 9496 7004 9636 7176
rect 7608 6772 7616 6944
rect 7616 6772 7672 6944
rect 7672 6772 7808 6944
rect 7808 6772 7864 6944
rect 7864 6772 8000 6944
rect 8000 6772 8056 6944
rect 8056 6772 8192 6944
rect 8192 6772 8248 6944
rect 8248 6772 8384 6944
rect 8384 6772 8440 6944
rect 8440 6772 8576 6944
rect 8576 6772 8592 6944
rect 7608 6756 8592 6772
rect 8764 6556 9636 6588
rect 8764 6388 8864 6556
rect 8864 6388 8920 6556
rect 8920 6388 9056 6556
rect 9056 6388 9112 6556
rect 9112 6388 9248 6556
rect 9248 6388 9304 6556
rect 9304 6388 9440 6556
rect 9440 6388 9496 6556
rect 9496 6388 9636 6556
rect 19504 8296 19516 8472
rect 19516 8296 19572 8472
rect 19572 8296 19708 8472
rect 19708 8296 19764 8472
rect 19764 8296 19900 8472
rect 19900 8296 19956 8472
rect 19956 8296 20092 8472
rect 20092 8296 20148 8472
rect 20148 8296 20284 8472
rect 20284 8296 20340 8472
rect 20340 8296 20476 8472
rect 20476 8296 20480 8472
rect 19504 8224 20480 8296
rect 23164 8412 24036 8440
rect 23164 8240 23264 8412
rect 23264 8240 23320 8412
rect 23320 8240 23456 8412
rect 23456 8240 23512 8412
rect 23512 8240 23648 8412
rect 23648 8240 23704 8412
rect 23704 8240 23840 8412
rect 23840 8240 23896 8412
rect 23896 8240 24036 8412
rect 20624 8080 21600 8164
rect 20624 7916 20628 8080
rect 20628 7916 20764 8080
rect 20764 7916 20820 8080
rect 20820 7916 20956 8080
rect 20956 7916 21012 8080
rect 21012 7916 21148 8080
rect 21148 7916 21204 8080
rect 21204 7916 21340 8080
rect 21340 7916 21396 8080
rect 21396 7916 21600 8080
rect 22004 8008 22016 8180
rect 22016 8008 22072 8180
rect 22072 8008 22208 8180
rect 22208 8008 22264 8180
rect 22264 8008 22400 8180
rect 22400 8008 22456 8180
rect 22456 8008 22592 8180
rect 22592 8008 22648 8180
rect 22648 8008 22784 8180
rect 22784 8008 22840 8180
rect 22840 8008 22976 8180
rect 22976 8008 22988 8180
rect 22004 7992 22988 8008
rect 19504 7676 19516 7848
rect 19516 7676 19572 7848
rect 19572 7676 19708 7848
rect 19708 7676 19764 7848
rect 19764 7676 19900 7848
rect 19900 7676 19956 7848
rect 19956 7676 20092 7848
rect 20092 7676 20148 7848
rect 20148 7676 20284 7848
rect 20284 7676 20340 7848
rect 20340 7676 20476 7848
rect 20476 7676 20480 7848
rect 19504 7600 20480 7676
rect 23164 7792 24036 7820
rect 23164 7620 23264 7792
rect 23264 7620 23320 7792
rect 23320 7620 23456 7792
rect 23456 7620 23512 7792
rect 23512 7620 23648 7792
rect 23648 7620 23704 7792
rect 23704 7620 23840 7792
rect 23840 7620 23896 7792
rect 23896 7620 24036 7792
rect 20784 7000 21476 7512
rect 22008 7388 22016 7556
rect 22016 7388 22072 7556
rect 22072 7388 22208 7556
rect 22208 7388 22264 7556
rect 22264 7388 22400 7556
rect 22400 7388 22456 7556
rect 22456 7388 22592 7556
rect 22592 7388 22648 7556
rect 22648 7388 22784 7556
rect 22784 7388 22840 7556
rect 22840 7388 22976 7556
rect 22976 7388 22992 7556
rect 22008 7368 22992 7388
rect 23164 7176 24036 7204
rect 23164 7004 23264 7176
rect 23264 7004 23320 7176
rect 23320 7004 23456 7176
rect 23456 7004 23512 7176
rect 23512 7004 23648 7176
rect 23648 7004 23704 7176
rect 23704 7004 23840 7176
rect 23840 7004 23896 7176
rect 23896 7004 24036 7176
rect 22008 6772 22016 6944
rect 22016 6772 22072 6944
rect 22072 6772 22208 6944
rect 22208 6772 22264 6944
rect 22264 6772 22400 6944
rect 22400 6772 22456 6944
rect 22456 6772 22592 6944
rect 22592 6772 22648 6944
rect 22648 6772 22784 6944
rect 22784 6772 22840 6944
rect 22840 6772 22976 6944
rect 22976 6772 22992 6944
rect 22008 6756 22992 6772
rect 23164 6556 24036 6588
rect 7604 6152 7616 6320
rect 7616 6152 7672 6320
rect 7672 6152 7808 6320
rect 7808 6152 7864 6320
rect 7864 6152 8000 6320
rect 8000 6152 8056 6320
rect 8056 6152 8192 6320
rect 8192 6152 8248 6320
rect 8248 6152 8384 6320
rect 8384 6152 8440 6320
rect 8440 6152 8576 6320
rect 8576 6152 8588 6320
rect 7604 6132 8588 6152
rect 23164 6388 23264 6556
rect 23264 6388 23320 6556
rect 23320 6388 23456 6556
rect 23456 6388 23512 6556
rect 23512 6388 23648 6556
rect 23648 6388 23704 6556
rect 23704 6388 23840 6556
rect 23840 6388 23896 6556
rect 23896 6388 24036 6556
rect 22004 6152 22016 6320
rect 22016 6152 22072 6320
rect 22072 6152 22208 6320
rect 22208 6152 22264 6320
rect 22264 6152 22400 6320
rect 22400 6152 22456 6320
rect 22456 6152 22592 6320
rect 22592 6152 22648 6320
rect 22648 6152 22784 6320
rect 22784 6152 22840 6320
rect 22840 6152 22976 6320
rect 22976 6152 22988 6320
rect -10064 5752 -10060 5924
rect -10060 5752 -10008 5924
rect -10008 5752 -9868 5924
rect -9868 5752 -9816 5924
rect -9816 5752 -9676 5924
rect -9676 5752 -9624 5924
rect -9624 5752 -9484 5924
rect -9484 5752 -9460 5924
rect -10064 5740 -9460 5752
rect 212 5472 216 5644
rect 216 5472 268 5644
rect 268 5472 408 5644
rect 408 5472 460 5644
rect 460 5472 600 5644
rect 600 5472 652 5644
rect 652 5472 792 5644
rect 792 5472 816 5644
rect 212 5460 816 5472
rect -10064 5136 -10060 5308
rect -10060 5136 -10008 5308
rect -10008 5136 -9868 5308
rect -9868 5136 -9816 5308
rect -9816 5136 -9676 5308
rect -9676 5136 -9624 5308
rect -9624 5136 -9484 5308
rect -9484 5136 -9460 5308
rect -10064 5124 -9460 5136
rect 2012 5472 2016 5644
rect 2016 5472 2068 5644
rect 2068 5472 2208 5644
rect 2208 5472 2260 5644
rect 2260 5472 2400 5644
rect 2400 5472 2452 5644
rect 2452 5472 2592 5644
rect 2592 5472 2616 5644
rect 2012 5460 2616 5472
rect 212 4856 216 5028
rect 216 4856 268 5028
rect 268 4856 408 5028
rect 408 4856 460 5028
rect 460 4856 600 5028
rect 600 4856 652 5028
rect 652 4856 792 5028
rect 792 4856 816 5028
rect 212 4844 816 4856
rect -10068 4516 -10060 4688
rect -10060 4516 -10008 4688
rect -10008 4516 -9868 4688
rect -9868 4516 -9816 4688
rect -9816 4516 -9676 4688
rect -9676 4516 -9624 4688
rect -9624 4516 -9484 4688
rect -9484 4516 -9464 4688
rect -10068 4504 -9464 4516
rect -3172 4420 -3028 4532
rect -808 4404 -404 4816
rect -404 4404 -32 4816
rect 3812 5472 3816 5644
rect 3816 5472 3868 5644
rect 3868 5472 4008 5644
rect 4008 5472 4060 5644
rect 4060 5472 4200 5644
rect 4200 5472 4252 5644
rect 4252 5472 4392 5644
rect 4392 5472 4416 5644
rect 3812 5460 4416 5472
rect 2012 4856 2016 5028
rect 2016 4856 2068 5028
rect 2068 4856 2208 5028
rect 2208 4856 2260 5028
rect 2260 4856 2400 5028
rect 2400 4856 2452 5028
rect 2452 4856 2592 5028
rect 2592 4856 2616 5028
rect 2012 4844 2616 4856
rect 5612 5472 5616 5644
rect 5616 5472 5668 5644
rect 5668 5472 5808 5644
rect 5808 5472 5860 5644
rect 5860 5472 6000 5644
rect 6000 5472 6052 5644
rect 6052 5472 6192 5644
rect 6192 5472 6216 5644
rect 5612 5460 6216 5472
rect 3812 4856 3816 5028
rect 3816 4856 3868 5028
rect 3868 4856 4008 5028
rect 4008 4856 4060 5028
rect 4060 4856 4200 5028
rect 4200 4856 4252 5028
rect 4252 4856 4392 5028
rect 4392 4856 4416 5028
rect 3812 4844 4416 4856
rect 22004 6132 22988 6152
rect 8760 5940 9632 5968
rect 8760 5768 8864 5940
rect 8864 5768 8920 5940
rect 8920 5768 9056 5940
rect 9056 5768 9112 5940
rect 9112 5768 9248 5940
rect 9248 5768 9304 5940
rect 9304 5768 9440 5940
rect 9440 5768 9496 5940
rect 9496 5768 9632 5940
rect 7604 5536 7616 5708
rect 7616 5536 7672 5708
rect 7672 5536 7808 5708
rect 7808 5536 7864 5708
rect 7864 5536 8000 5708
rect 8000 5536 8056 5708
rect 8056 5536 8192 5708
rect 8192 5536 8248 5708
rect 8248 5536 8384 5708
rect 8384 5536 8440 5708
rect 8440 5536 8576 5708
rect 8576 5536 8588 5708
rect 7604 5520 8588 5536
rect 14612 5472 14616 5644
rect 14616 5472 14668 5644
rect 14668 5472 14808 5644
rect 14808 5472 14860 5644
rect 14860 5472 15000 5644
rect 15000 5472 15052 5644
rect 15052 5472 15192 5644
rect 15192 5472 15216 5644
rect 14612 5460 15216 5472
rect 8760 5320 9632 5348
rect 8760 5148 8864 5320
rect 8864 5148 8920 5320
rect 8920 5148 9056 5320
rect 9056 5148 9112 5320
rect 9112 5148 9248 5320
rect 9248 5148 9304 5320
rect 9304 5148 9440 5320
rect 9440 5148 9496 5320
rect 9496 5148 9632 5320
rect 16412 5472 16416 5644
rect 16416 5472 16468 5644
rect 16468 5472 16608 5644
rect 16608 5472 16660 5644
rect 16660 5472 16800 5644
rect 16800 5472 16852 5644
rect 16852 5472 16992 5644
rect 16992 5472 17016 5644
rect 16412 5460 17016 5472
rect 5612 4856 5616 5028
rect 5616 4856 5668 5028
rect 5668 4856 5808 5028
rect 5808 4856 5860 5028
rect 5860 4856 6000 5028
rect 6000 4856 6052 5028
rect 6052 4856 6192 5028
rect 6192 4856 6216 5028
rect 5612 4844 6216 4856
rect 7604 4916 7616 5084
rect 7616 4916 7672 5084
rect 7672 4916 7808 5084
rect 7808 4916 7864 5084
rect 7864 4916 8000 5084
rect 8000 4916 8056 5084
rect 8056 4916 8192 5084
rect 8192 4916 8248 5084
rect 8248 4916 8384 5084
rect 8384 4916 8440 5084
rect 8440 4916 8576 5084
rect 8576 4916 8588 5084
rect 7604 4896 8588 4916
rect 11480 4580 11820 4860
rect 14612 4856 14616 5028
rect 14616 4856 14668 5028
rect 14668 4856 14808 5028
rect 14808 4856 14860 5028
rect 14860 4856 15000 5028
rect 15000 4856 15052 5028
rect 15052 4856 15192 5028
rect 15192 4856 15216 5028
rect 14612 4844 15216 4856
rect 208 4236 216 4408
rect 216 4236 268 4408
rect 268 4236 408 4408
rect 408 4236 460 4408
rect 460 4236 600 4408
rect 600 4236 652 4408
rect 652 4236 792 4408
rect 792 4236 812 4408
rect 208 4224 812 4236
rect 2008 4236 2016 4408
rect 2016 4236 2068 4408
rect 2068 4236 2208 4408
rect 2208 4236 2260 4408
rect 2260 4236 2400 4408
rect 2400 4236 2452 4408
rect 2452 4236 2592 4408
rect 2592 4236 2612 4408
rect 2008 4224 2612 4236
rect 3808 4236 3816 4408
rect 3816 4236 3868 4408
rect 3868 4236 4008 4408
rect 4008 4236 4060 4408
rect 4060 4236 4200 4408
rect 4200 4236 4252 4408
rect 4252 4236 4392 4408
rect 4392 4236 4412 4408
rect 3808 4224 4412 4236
rect 5608 4236 5616 4408
rect 5616 4236 5668 4408
rect 5668 4236 5808 4408
rect 5808 4236 5860 4408
rect 5860 4236 6000 4408
rect 6000 4236 6052 4408
rect 6052 4236 6192 4408
rect 6192 4236 6212 4408
rect 13592 4404 13996 4816
rect 13996 4404 14368 4816
rect 18212 5472 18216 5644
rect 18216 5472 18268 5644
rect 18268 5472 18408 5644
rect 18408 5472 18460 5644
rect 18460 5472 18600 5644
rect 18600 5472 18652 5644
rect 18652 5472 18792 5644
rect 18792 5472 18816 5644
rect 18212 5460 18816 5472
rect 16412 4856 16416 5028
rect 16416 4856 16468 5028
rect 16468 4856 16608 5028
rect 16608 4856 16660 5028
rect 16660 4856 16800 5028
rect 16800 4856 16852 5028
rect 16852 4856 16992 5028
rect 16992 4856 17016 5028
rect 16412 4844 17016 4856
rect 20012 5472 20016 5644
rect 20016 5472 20068 5644
rect 20068 5472 20208 5644
rect 20208 5472 20260 5644
rect 20260 5472 20400 5644
rect 20400 5472 20452 5644
rect 20452 5472 20592 5644
rect 20592 5472 20616 5644
rect 20012 5460 20616 5472
rect 18212 4856 18216 5028
rect 18216 4856 18268 5028
rect 18268 4856 18408 5028
rect 18408 4856 18460 5028
rect 18460 4856 18600 5028
rect 18600 4856 18652 5028
rect 18652 4856 18792 5028
rect 18792 4856 18816 5028
rect 18212 4844 18816 4856
rect 23160 5940 24032 5968
rect 23160 5768 23264 5940
rect 23264 5768 23320 5940
rect 23320 5768 23456 5940
rect 23456 5768 23512 5940
rect 23512 5768 23648 5940
rect 23648 5768 23704 5940
rect 23704 5768 23840 5940
rect 23840 5768 23896 5940
rect 23896 5768 24032 5940
rect 22004 5536 22016 5708
rect 22016 5536 22072 5708
rect 22072 5536 22208 5708
rect 22208 5536 22264 5708
rect 22264 5536 22400 5708
rect 22400 5536 22456 5708
rect 22456 5536 22592 5708
rect 22592 5536 22648 5708
rect 22648 5536 22784 5708
rect 22784 5536 22840 5708
rect 22840 5536 22976 5708
rect 22976 5536 22988 5708
rect 22004 5520 22988 5536
rect 23160 5320 24032 5348
rect 23160 5148 23264 5320
rect 23264 5148 23320 5320
rect 23320 5148 23456 5320
rect 23456 5148 23512 5320
rect 23512 5148 23648 5320
rect 23648 5148 23704 5320
rect 23704 5148 23840 5320
rect 23840 5148 23896 5320
rect 23896 5148 24032 5320
rect 20012 4856 20016 5028
rect 20016 4856 20068 5028
rect 20068 4856 20208 5028
rect 20208 4856 20260 5028
rect 20260 4856 20400 5028
rect 20400 4856 20452 5028
rect 20452 4856 20592 5028
rect 20592 4856 20616 5028
rect 20012 4844 20616 4856
rect 22004 4916 22016 5084
rect 22016 4916 22072 5084
rect 22072 4916 22208 5084
rect 22208 4916 22264 5084
rect 22264 4916 22400 5084
rect 22400 4916 22456 5084
rect 22456 4916 22592 5084
rect 22592 4916 22648 5084
rect 22648 4916 22784 5084
rect 22784 4916 22840 5084
rect 22840 4916 22976 5084
rect 22976 4916 22988 5084
rect 22004 4896 22988 4916
rect 5608 4224 6212 4236
rect 14608 4236 14616 4408
rect 14616 4236 14668 4408
rect 14668 4236 14808 4408
rect 14808 4236 14860 4408
rect 14860 4236 15000 4408
rect 15000 4236 15052 4408
rect 15052 4236 15192 4408
rect 15192 4236 15212 4408
rect 14608 4224 15212 4236
rect 16408 4236 16416 4408
rect 16416 4236 16468 4408
rect 16468 4236 16608 4408
rect 16608 4236 16660 4408
rect 16660 4236 16800 4408
rect 16800 4236 16852 4408
rect 16852 4236 16992 4408
rect 16992 4236 17012 4408
rect 16408 4224 17012 4236
rect 18208 4236 18216 4408
rect 18216 4236 18268 4408
rect 18268 4236 18408 4408
rect 18408 4236 18460 4408
rect 18460 4236 18600 4408
rect 18600 4236 18652 4408
rect 18652 4236 18792 4408
rect 18792 4236 18812 4408
rect 18208 4224 18812 4236
rect 20008 4236 20016 4408
rect 20016 4236 20068 4408
rect 20068 4236 20208 4408
rect 20208 4236 20260 4408
rect 20260 4236 20400 4408
rect 20400 4236 20452 4408
rect 20452 4236 20592 4408
rect 20592 4236 20612 4408
rect 24520 4360 24900 4700
rect 20008 4224 20612 4236
rect -10060 4008 -9460 4020
rect -10060 3836 -10008 4008
rect -10008 3836 -9544 4008
rect -9544 3836 -9492 4008
rect -9492 3836 -9460 4008
rect -9316 3608 -9284 3780
rect -9284 3608 -9232 3780
rect -9232 3608 -8768 3780
rect -8768 3608 -8716 3780
rect -9316 3596 -8716 3608
rect 216 3728 816 3740
rect 2016 3728 2616 3740
rect 3816 3728 4416 3740
rect 5616 3728 6216 3740
rect 216 3556 268 3728
rect 268 3556 732 3728
rect 732 3556 784 3728
rect 784 3556 816 3728
rect 2016 3556 2068 3728
rect 2068 3556 2532 3728
rect 2532 3556 2584 3728
rect 2584 3556 2616 3728
rect 3816 3556 3868 3728
rect 3868 3556 4332 3728
rect 4332 3556 4384 3728
rect 4384 3556 4416 3728
rect 5616 3556 5668 3728
rect 5668 3556 6132 3728
rect 6132 3556 6184 3728
rect 6184 3556 6216 3728
rect 14616 3728 15216 3740
rect 16416 3728 17016 3740
rect 18216 3728 18816 3740
rect 20016 3728 20616 3740
rect 14616 3556 14668 3728
rect 14668 3556 15132 3728
rect 15132 3556 15184 3728
rect 15184 3556 15216 3728
rect 16416 3556 16468 3728
rect 16468 3556 16932 3728
rect 16932 3556 16984 3728
rect 16984 3556 17016 3728
rect 18216 3556 18268 3728
rect 18268 3556 18732 3728
rect 18732 3556 18784 3728
rect 18784 3556 18816 3728
rect 20016 3556 20068 3728
rect 20068 3556 20532 3728
rect 20532 3556 20584 3728
rect 20584 3556 20616 3728
rect -10060 3392 -9460 3404
rect -10060 3220 -10008 3392
rect -10008 3220 -9544 3392
rect -9544 3220 -9492 3392
rect -9492 3220 -9460 3392
rect 960 3328 992 3500
rect 992 3328 1044 3500
rect 1044 3328 1508 3500
rect 1508 3328 1560 3500
rect 960 3316 1560 3328
rect 2760 3328 2792 3500
rect 2792 3328 2844 3500
rect 2844 3328 3308 3500
rect 3308 3328 3360 3500
rect 2760 3316 3360 3328
rect 4560 3328 4592 3500
rect 4592 3328 4644 3500
rect 4644 3328 5108 3500
rect 5108 3328 5160 3500
rect 4560 3316 5160 3328
rect 6360 3328 6392 3500
rect 6392 3328 6444 3500
rect 6444 3328 6908 3500
rect 6908 3328 6960 3500
rect 6360 3316 6960 3328
rect 15360 3328 15392 3500
rect 15392 3328 15444 3500
rect 15444 3328 15908 3500
rect 15908 3328 15960 3500
rect 15360 3316 15960 3328
rect 17160 3328 17192 3500
rect 17192 3328 17244 3500
rect 17244 3328 17708 3500
rect 17708 3328 17760 3500
rect 17160 3316 17760 3328
rect 18960 3328 18992 3500
rect 18992 3328 19044 3500
rect 19044 3328 19508 3500
rect 19508 3328 19560 3500
rect 18960 3316 19560 3328
rect 20760 3328 20792 3500
rect 20792 3328 20844 3500
rect 20844 3328 21308 3500
rect 21308 3328 21360 3500
rect 20760 3316 21360 3328
rect -9316 2992 -9284 3164
rect -9284 2992 -9232 3164
rect -9232 2992 -8768 3164
rect -8768 2992 -8716 3164
rect -9316 2980 -8716 2992
rect 216 3112 816 3124
rect 216 2940 268 3112
rect 268 2940 732 3112
rect 732 2940 784 3112
rect 784 2940 816 3112
rect 2016 3112 2616 3124
rect 2016 2940 2068 3112
rect 2068 2940 2532 3112
rect 2532 2940 2584 3112
rect 2584 2940 2616 3112
rect 3816 3112 4416 3124
rect 3816 2940 3868 3112
rect 3868 2940 4332 3112
rect 4332 2940 4384 3112
rect 4384 2940 4416 3112
rect 5616 3112 6216 3124
rect 5616 2940 5668 3112
rect 5668 2940 6132 3112
rect 6132 2940 6184 3112
rect 6184 2940 6216 3112
rect 14616 3112 15216 3124
rect 14616 2940 14668 3112
rect 14668 2940 15132 3112
rect 15132 2940 15184 3112
rect 15184 2940 15216 3112
rect 16416 3112 17016 3124
rect 16416 2940 16468 3112
rect 16468 2940 16932 3112
rect 16932 2940 16984 3112
rect 16984 2940 17016 3112
rect 18216 3112 18816 3124
rect 18216 2940 18268 3112
rect 18268 2940 18732 3112
rect 18732 2940 18784 3112
rect 18784 2940 18816 3112
rect 20016 3112 20616 3124
rect 20016 2940 20068 3112
rect 20068 2940 20532 3112
rect 20532 2940 20584 3112
rect 20584 2940 20616 3112
rect -10060 2772 -9460 2784
rect -10060 2600 -10008 2772
rect -10008 2600 -9544 2772
rect -9544 2600 -9492 2772
rect -9492 2600 -9460 2772
rect 960 2712 992 2884
rect 992 2712 1044 2884
rect 1044 2712 1508 2884
rect 1508 2712 1560 2884
rect 960 2700 1560 2712
rect 2760 2712 2792 2884
rect 2792 2712 2844 2884
rect 2844 2712 3308 2884
rect 3308 2712 3360 2884
rect 2760 2700 3360 2712
rect 4560 2712 4592 2884
rect 4592 2712 4644 2884
rect 4644 2712 5108 2884
rect 5108 2712 5160 2884
rect 4560 2700 5160 2712
rect 6360 2712 6392 2884
rect 6392 2712 6444 2884
rect 6444 2712 6908 2884
rect 6908 2712 6960 2884
rect 6360 2700 6960 2712
rect 15360 2712 15392 2884
rect 15392 2712 15444 2884
rect 15444 2712 15908 2884
rect 15908 2712 15960 2884
rect 15360 2700 15960 2712
rect 17160 2712 17192 2884
rect 17192 2712 17244 2884
rect 17244 2712 17708 2884
rect 17708 2712 17760 2884
rect 17160 2700 17760 2712
rect 18960 2712 18992 2884
rect 18992 2712 19044 2884
rect 19044 2712 19508 2884
rect 19508 2712 19560 2884
rect 18960 2700 19560 2712
rect 20760 2712 20792 2884
rect 20792 2712 20844 2884
rect 20844 2712 21308 2884
rect 21308 2712 21360 2884
rect 20760 2700 21360 2712
rect -9316 2372 -9284 2544
rect -9284 2372 -9232 2544
rect -9232 2372 -8768 2544
rect -8768 2372 -8716 2544
rect -9316 2360 -8716 2372
rect 216 2492 816 2504
rect 216 2320 268 2492
rect 268 2320 732 2492
rect 732 2320 784 2492
rect 784 2320 816 2492
rect 2016 2492 2616 2504
rect 2016 2320 2068 2492
rect 2068 2320 2532 2492
rect 2532 2320 2584 2492
rect 2584 2320 2616 2492
rect 3816 2492 4416 2504
rect 3816 2320 3868 2492
rect 3868 2320 4332 2492
rect 4332 2320 4384 2492
rect 4384 2320 4416 2492
rect 5616 2492 6216 2504
rect 5616 2320 5668 2492
rect 5668 2320 6132 2492
rect 6132 2320 6184 2492
rect 6184 2320 6216 2492
rect 14616 2492 15216 2504
rect 14616 2320 14668 2492
rect 14668 2320 15132 2492
rect 15132 2320 15184 2492
rect 15184 2320 15216 2492
rect 16416 2492 17016 2504
rect 16416 2320 16468 2492
rect 16468 2320 16932 2492
rect 16932 2320 16984 2492
rect 16984 2320 17016 2492
rect 18216 2492 18816 2504
rect 18216 2320 18268 2492
rect 18268 2320 18732 2492
rect 18732 2320 18784 2492
rect 18784 2320 18816 2492
rect 20016 2492 20616 2504
rect 20016 2320 20068 2492
rect 20068 2320 20532 2492
rect 20532 2320 20584 2492
rect 20584 2320 20616 2492
rect -10060 2156 -9460 2168
rect -10060 1984 -10008 2156
rect -10008 1984 -9544 2156
rect -9544 1984 -9492 2156
rect -9492 1984 -9460 2156
rect 960 2092 992 2264
rect 992 2092 1044 2264
rect 1044 2092 1508 2264
rect 1508 2092 1560 2264
rect 960 2080 1560 2092
rect 2760 2092 2792 2264
rect 2792 2092 2844 2264
rect 2844 2092 3308 2264
rect 3308 2092 3360 2264
rect 2760 2080 3360 2092
rect 4560 2092 4592 2264
rect 4592 2092 4644 2264
rect 4644 2092 5108 2264
rect 5108 2092 5160 2264
rect 4560 2080 5160 2092
rect 6360 2092 6392 2264
rect 6392 2092 6444 2264
rect 6444 2092 6908 2264
rect 6908 2092 6960 2264
rect 6360 2080 6960 2092
rect 15360 2092 15392 2264
rect 15392 2092 15444 2264
rect 15444 2092 15908 2264
rect 15908 2092 15960 2264
rect 15360 2080 15960 2092
rect 17160 2092 17192 2264
rect 17192 2092 17244 2264
rect 17244 2092 17708 2264
rect 17708 2092 17760 2264
rect 17160 2080 17760 2092
rect 18960 2092 18992 2264
rect 18992 2092 19044 2264
rect 19044 2092 19508 2264
rect 19508 2092 19560 2264
rect 18960 2080 19560 2092
rect 20760 2092 20792 2264
rect 20792 2092 20844 2264
rect 20844 2092 21308 2264
rect 21308 2092 21360 2264
rect 20760 2080 21360 2092
rect -9316 1756 -9284 1928
rect -9284 1756 -9232 1928
rect -9232 1756 -8768 1928
rect -8768 1756 -8716 1928
rect -9316 1744 -8716 1756
rect 216 1876 816 1888
rect 216 1704 268 1876
rect 268 1704 732 1876
rect 732 1704 784 1876
rect 784 1704 816 1876
rect 2016 1876 2616 1888
rect 2016 1704 2068 1876
rect 2068 1704 2532 1876
rect 2532 1704 2584 1876
rect 2584 1704 2616 1876
rect 3816 1876 4416 1888
rect 3816 1704 3868 1876
rect 3868 1704 4332 1876
rect 4332 1704 4384 1876
rect 4384 1704 4416 1876
rect 5616 1876 6216 1888
rect 5616 1704 5668 1876
rect 5668 1704 6132 1876
rect 6132 1704 6184 1876
rect 6184 1704 6216 1876
rect 14616 1876 15216 1888
rect 14616 1704 14668 1876
rect 14668 1704 15132 1876
rect 15132 1704 15184 1876
rect 15184 1704 15216 1876
rect 16416 1876 17016 1888
rect 16416 1704 16468 1876
rect 16468 1704 16932 1876
rect 16932 1704 16984 1876
rect 16984 1704 17016 1876
rect 18216 1876 18816 1888
rect 18216 1704 18268 1876
rect 18268 1704 18732 1876
rect 18732 1704 18784 1876
rect 18784 1704 18816 1876
rect 20016 1876 20616 1888
rect 20016 1704 20068 1876
rect 20068 1704 20532 1876
rect 20532 1704 20584 1876
rect 20584 1704 20616 1876
rect -10060 1536 -9460 1548
rect -10060 1364 -10008 1536
rect -10008 1364 -9544 1536
rect -9544 1364 -9492 1536
rect -9492 1364 -9460 1536
rect 960 1476 992 1648
rect 992 1476 1044 1648
rect 1044 1476 1508 1648
rect 1508 1476 1560 1648
rect 960 1464 1560 1476
rect 2760 1476 2792 1648
rect 2792 1476 2844 1648
rect 2844 1476 3308 1648
rect 3308 1476 3360 1648
rect 2760 1464 3360 1476
rect 4560 1476 4592 1648
rect 4592 1476 4644 1648
rect 4644 1476 5108 1648
rect 5108 1476 5160 1648
rect 4560 1464 5160 1476
rect 6360 1476 6392 1648
rect 6392 1476 6444 1648
rect 6444 1476 6908 1648
rect 6908 1476 6960 1648
rect 6360 1464 6960 1476
rect 15360 1476 15392 1648
rect 15392 1476 15444 1648
rect 15444 1476 15908 1648
rect 15908 1476 15960 1648
rect 15360 1464 15960 1476
rect 17160 1476 17192 1648
rect 17192 1476 17244 1648
rect 17244 1476 17708 1648
rect 17708 1476 17760 1648
rect 17160 1464 17760 1476
rect 18960 1476 18992 1648
rect 18992 1476 19044 1648
rect 19044 1476 19508 1648
rect 19508 1476 19560 1648
rect 18960 1464 19560 1476
rect 20760 1476 20792 1648
rect 20792 1476 20844 1648
rect 20844 1476 21308 1648
rect 21308 1476 21360 1648
rect 20760 1464 21360 1476
rect -9316 1136 -9284 1308
rect -9284 1136 -9232 1308
rect -9232 1136 -8768 1308
rect -8768 1136 -8716 1308
rect -9316 1124 -8716 1136
rect 216 1256 816 1268
rect 216 1084 268 1256
rect 268 1084 732 1256
rect 732 1084 784 1256
rect 784 1084 816 1256
rect 2016 1256 2616 1268
rect 2016 1084 2068 1256
rect 2068 1084 2532 1256
rect 2532 1084 2584 1256
rect 2584 1084 2616 1256
rect 3816 1256 4416 1268
rect 3816 1084 3868 1256
rect 3868 1084 4332 1256
rect 4332 1084 4384 1256
rect 4384 1084 4416 1256
rect 5616 1256 6216 1268
rect 5616 1084 5668 1256
rect 5668 1084 6132 1256
rect 6132 1084 6184 1256
rect 6184 1084 6216 1256
rect 14616 1256 15216 1268
rect 14616 1084 14668 1256
rect 14668 1084 15132 1256
rect 15132 1084 15184 1256
rect 15184 1084 15216 1256
rect 16416 1256 17016 1268
rect 16416 1084 16468 1256
rect 16468 1084 16932 1256
rect 16932 1084 16984 1256
rect 16984 1084 17016 1256
rect 18216 1256 18816 1268
rect 18216 1084 18268 1256
rect 18268 1084 18732 1256
rect 18732 1084 18784 1256
rect 18784 1084 18816 1256
rect 20016 1256 20616 1268
rect 20016 1084 20068 1256
rect 20068 1084 20532 1256
rect 20532 1084 20584 1256
rect 20584 1084 20616 1256
rect -10060 920 -9460 932
rect -10060 748 -10008 920
rect -10008 748 -9544 920
rect -9544 748 -9492 920
rect -9492 748 -9460 920
rect 960 856 992 1028
rect 992 856 1044 1028
rect 1044 856 1508 1028
rect 1508 856 1560 1028
rect 960 844 1560 856
rect 2760 856 2792 1028
rect 2792 856 2844 1028
rect 2844 856 3308 1028
rect 3308 856 3360 1028
rect 2760 844 3360 856
rect 4560 856 4592 1028
rect 4592 856 4644 1028
rect 4644 856 5108 1028
rect 5108 856 5160 1028
rect 4560 844 5160 856
rect 6360 856 6392 1028
rect 6392 856 6444 1028
rect 6444 856 6908 1028
rect 6908 856 6960 1028
rect 6360 844 6960 856
rect 15360 856 15392 1028
rect 15392 856 15444 1028
rect 15444 856 15908 1028
rect 15908 856 15960 1028
rect 15360 844 15960 856
rect 17160 856 17192 1028
rect 17192 856 17244 1028
rect 17244 856 17708 1028
rect 17708 856 17760 1028
rect 17160 844 17760 856
rect 18960 856 18992 1028
rect 18992 856 19044 1028
rect 19044 856 19508 1028
rect 19508 856 19560 1028
rect 18960 844 19560 856
rect 20760 856 20792 1028
rect 20792 856 20844 1028
rect 20844 856 21308 1028
rect 21308 856 21360 1028
rect 20760 844 21360 856
rect -9316 520 -9284 692
rect -9284 520 -9232 692
rect -9232 520 -8768 692
rect -8768 520 -8716 692
rect -9316 508 -8716 520
rect 216 640 816 652
rect -8500 348 -8360 508
rect 216 468 268 640
rect 268 468 732 640
rect 732 468 784 640
rect 784 468 816 640
rect 2016 640 2616 652
rect 2016 468 2068 640
rect 2068 468 2532 640
rect 2532 468 2584 640
rect 2584 468 2616 640
rect 3816 640 4416 652
rect 3816 468 3868 640
rect 3868 468 4332 640
rect 4332 468 4384 640
rect 4384 468 4416 640
rect 5616 640 6216 652
rect 5616 468 5668 640
rect 5668 468 6132 640
rect 6132 468 6184 640
rect 6184 468 6216 640
rect 14616 640 15216 652
rect 14616 468 14668 640
rect 14668 468 15132 640
rect 15132 468 15184 640
rect 15184 468 15216 640
rect 16416 640 17016 652
rect 16416 468 16468 640
rect 16468 468 16932 640
rect 16932 468 16984 640
rect 16984 468 17016 640
rect 18216 640 18816 652
rect 18216 468 18268 640
rect 18268 468 18732 640
rect 18732 468 18784 640
rect 18784 468 18816 640
rect 20016 640 20616 652
rect 20016 468 20068 640
rect 20068 468 20532 640
rect 20532 468 20584 640
rect 20584 468 20616 640
rect 960 240 992 412
rect 992 240 1044 412
rect 1044 240 1508 412
rect 1508 240 1560 412
rect 960 228 1560 240
rect 1696 68 1876 268
rect 2760 240 2792 412
rect 2792 240 2844 412
rect 2844 240 3308 412
rect 3308 240 3360 412
rect 2760 228 3360 240
rect 4560 240 4592 412
rect 4592 240 4644 412
rect 4644 240 5108 412
rect 5108 240 5160 412
rect 4560 228 5160 240
rect 5288 64 5468 276
rect 6360 240 6392 412
rect 6392 240 6444 412
rect 6444 240 6908 412
rect 6908 240 6960 412
rect 6360 228 6960 240
rect 15360 240 15392 412
rect 15392 240 15444 412
rect 15444 240 15908 412
rect 15908 240 15960 412
rect 15360 228 15960 240
rect 16096 68 16276 268
rect 17160 240 17192 412
rect 17192 240 17244 412
rect 17244 240 17708 412
rect 17708 240 17760 412
rect 17160 228 17760 240
rect 18960 240 18992 412
rect 18992 240 19044 412
rect 19044 240 19508 412
rect 19508 240 19560 412
rect 18960 228 19560 240
rect 19688 64 19868 276
rect 20760 240 20792 412
rect 20792 240 20844 412
rect 20844 240 21308 412
rect 21308 240 21360 412
rect 20760 228 21360 240
rect -2768 -1188 -1960 -382
rect 11632 -1188 12440 -382
<< metal3 >>
rect 6460 27860 28460 29380
rect 6452 27440 28460 27860
rect 6452 27436 17036 27440
rect 6452 27360 7440 27436
rect 7372 27336 7440 27360
rect 7540 27360 17036 27436
rect 7540 27336 8256 27360
rect 7372 27172 8256 27336
rect 7372 26928 7384 27172
rect 8240 26928 8256 27172
rect 6476 26852 7288 26868
rect 6476 26608 6488 26852
rect 7268 26608 7288 26852
rect 6476 26216 7288 26608
rect 6476 25972 6488 26216
rect 7268 25972 7288 26216
rect 6476 25576 7288 25972
rect 7372 26540 8256 26928
rect 9592 27172 10476 27360
rect 9592 26928 9604 27172
rect 10460 26928 10476 27172
rect 7372 26296 7384 26540
rect 8240 26296 8256 26540
rect 7372 25904 8256 26296
rect 7372 25660 7384 25904
rect 8240 25660 8256 25904
rect 7372 25644 8256 25660
rect 8696 26852 9508 26868
rect 8696 26608 8708 26852
rect 9488 26608 9508 26852
rect 8696 26216 9508 26608
rect 8696 25972 8708 26216
rect 9488 25972 9508 26216
rect 6476 25332 6488 25576
rect 7268 25332 7288 25576
rect 6476 25076 7288 25332
rect 6476 24828 6492 25076
rect 7276 24828 7288 25076
rect 6476 24436 7288 24828
rect 8696 25576 9508 25972
rect 9592 26540 10476 26928
rect 11772 27172 12656 27360
rect 11772 26928 11784 27172
rect 12640 26928 12656 27172
rect 9592 26296 9604 26540
rect 10460 26296 10476 26540
rect 9592 25904 10476 26296
rect 9592 25660 9604 25904
rect 10460 25660 10476 25904
rect 9592 25644 10476 25660
rect 10876 26852 11688 26868
rect 10876 26608 10888 26852
rect 11668 26608 11688 26852
rect 10876 26216 11688 26608
rect 10876 25972 10888 26216
rect 11668 25972 11688 26216
rect 8696 25332 8708 25576
rect 9488 25332 9508 25576
rect 8696 25076 9508 25332
rect 8696 24828 8712 25076
rect 9496 24828 9508 25076
rect 6476 24188 6492 24436
rect 7276 24188 7288 24436
rect 6476 24160 7288 24188
rect 7372 24748 8256 24764
rect 7372 24508 7388 24748
rect 8240 24508 8256 24748
rect 7372 24441 8256 24508
rect 7372 24436 8338 24441
rect 7372 24212 8156 24436
rect 8328 24212 8338 24436
rect 7372 24207 8338 24212
rect 8696 24436 9508 24828
rect 10876 25576 11688 25972
rect 11772 26540 12656 26928
rect 13952 27172 14836 27360
rect 13952 26928 13964 27172
rect 14820 26928 14836 27172
rect 11772 26296 11784 26540
rect 12640 26296 12656 26540
rect 11772 25904 12656 26296
rect 11772 25660 11784 25904
rect 12640 25660 12656 25904
rect 11772 25644 12656 25660
rect 13056 26852 13868 26868
rect 13056 26608 13068 26852
rect 13848 26608 13868 26852
rect 13056 26216 13868 26608
rect 13056 25972 13068 26216
rect 13848 25972 13868 26216
rect 10876 25332 10888 25576
rect 11668 25332 11688 25576
rect 10876 25076 11688 25332
rect 10876 24828 10892 25076
rect 11676 24828 11688 25076
rect 7372 24116 8256 24207
rect 8696 24188 8712 24436
rect 9496 24188 9508 24436
rect 8696 24160 9508 24188
rect 9592 24748 10476 24764
rect 9592 24508 9608 24748
rect 10460 24508 10476 24748
rect 7372 23876 7388 24116
rect 8240 23876 8256 24116
rect 7372 23744 8256 23876
rect 9592 24116 10476 24508
rect 10876 24436 11688 24828
rect 13056 25576 13868 25972
rect 13952 26540 14836 26928
rect 16152 27172 17036 27360
rect 16152 26928 16164 27172
rect 17020 26928 17036 27172
rect 13952 26296 13964 26540
rect 14820 26296 14836 26540
rect 13952 25904 14836 26296
rect 13952 25660 13964 25904
rect 14820 25660 14836 25904
rect 13952 25644 14836 25660
rect 15256 26852 16068 26868
rect 15256 26608 15268 26852
rect 16048 26608 16068 26852
rect 15256 26216 16068 26608
rect 15256 25972 15268 26216
rect 16048 25972 16068 26216
rect 13056 25332 13068 25576
rect 13848 25332 13868 25576
rect 13056 25076 13868 25332
rect 13056 24828 13072 25076
rect 13856 24828 13868 25076
rect 10876 24188 10892 24436
rect 11676 24188 11688 24436
rect 10876 24160 11688 24188
rect 11772 24748 12656 24764
rect 11772 24508 11788 24748
rect 12640 24508 12656 24748
rect 9592 23876 9608 24116
rect 10460 24060 10476 24116
rect 11772 24116 12656 24508
rect 13056 24436 13868 24828
rect 15256 25576 16068 25972
rect 16152 26540 17036 26928
rect 16152 26296 16164 26540
rect 17020 26296 17036 26540
rect 16152 25904 17036 26296
rect 16152 25660 16164 25904
rect 17020 25660 17036 25904
rect 16152 25644 17036 25660
rect 15256 25332 15268 25576
rect 16048 25332 16068 25576
rect 15256 25076 16068 25332
rect 15256 24828 15272 25076
rect 16056 24828 16068 25076
rect 13056 24188 13072 24436
rect 13856 24188 13868 24436
rect 13056 24160 13868 24188
rect 13952 24748 14836 24764
rect 13952 24508 13968 24748
rect 14820 24508 14836 24748
rect 11772 24060 11788 24116
rect 10460 23876 11788 24060
rect 12640 24060 12656 24116
rect 13952 24116 14836 24508
rect 15256 24436 16068 24828
rect 18220 25120 18680 27440
rect 15256 24188 15272 24436
rect 16056 24188 16068 24436
rect 15256 24160 16068 24188
rect 16152 24748 17036 24764
rect 16152 24508 16168 24748
rect 17020 24508 17036 24748
rect 18220 24600 18280 25120
rect 18640 24600 18680 25120
rect 18220 24560 18680 24600
rect 19860 27108 24232 27136
rect 13952 24060 13968 24116
rect 12640 23876 13968 24060
rect 14820 24060 14836 24116
rect 16152 24116 17036 24508
rect 16152 24060 16168 24116
rect 14820 23876 16168 24060
rect 17020 23876 17036 24116
rect 9592 23744 17036 23876
rect 7392 23680 8256 23744
rect 7392 23376 7408 23680
rect 7398 23272 7408 23376
rect 8236 23376 8256 23680
rect 9604 23588 17024 23744
rect 8236 23272 8246 23376
rect 7398 23267 8246 23272
rect 6596 23197 7200 23200
rect 8316 23197 8920 23200
rect 6586 23192 7210 23197
rect 6586 23008 6596 23192
rect 7200 23008 7210 23192
rect 6586 23003 7210 23008
rect 8306 23192 8930 23197
rect 8306 23008 8316 23192
rect 8920 23008 8930 23192
rect 8306 23003 8930 23008
rect 6596 22581 7200 23003
rect 8316 22581 8920 23003
rect 6586 22576 7210 22581
rect 6586 22392 6596 22576
rect 7200 22392 7210 22576
rect 6586 22387 7210 22392
rect 8306 22576 8930 22581
rect 8306 22392 8316 22576
rect 8920 22392 8930 22576
rect 8306 22387 8930 22392
rect 6596 21961 7200 22387
rect 8316 21961 8920 22387
rect 6582 21956 7206 21961
rect 6582 21772 6592 21956
rect 7196 21772 7206 21956
rect 6582 21767 7206 21772
rect 8302 21956 8926 21961
rect 8302 21772 8312 21956
rect 8916 21772 8926 21956
rect 8302 21767 8926 21772
rect 6596 21293 7200 21767
rect 8316 21293 8920 21767
rect 6590 21288 7210 21293
rect 6590 21104 6600 21288
rect 7200 21104 7210 21288
rect 6590 21099 7210 21104
rect 8310 21288 8930 21293
rect 8310 21104 8320 21288
rect 8920 21104 8930 21288
rect 8310 21099 8930 21104
rect 10268 21220 10908 23588
rect 19860 23536 24148 27108
rect 19020 23448 24148 23536
rect 19020 23364 19044 23448
rect 19232 23364 24148 23448
rect 19020 23316 24148 23364
rect 19860 23084 24148 23316
rect 24212 23084 24232 27108
rect 19860 23056 24232 23084
rect 18262 22784 18870 22789
rect 18262 22484 18272 22784
rect 18860 22484 18870 22784
rect 18262 22479 18870 22484
rect 18272 22233 18860 22479
rect 19860 22296 20120 23056
rect 19860 22268 24232 22296
rect 18272 22228 18874 22233
rect 15890 22180 16310 22185
rect 15890 21740 15900 22180
rect 16300 21740 16310 22180
rect 15890 21735 16310 21740
rect 18272 21996 18284 22228
rect 18864 21996 18874 22228
rect 18272 21991 18874 21996
rect 18272 21621 18860 21991
rect 18984 21916 19640 21932
rect 18984 21688 18996 21916
rect 19628 21688 19640 21916
rect 18272 21616 18874 21621
rect 18272 21384 18284 21616
rect 18864 21384 18874 21616
rect 18272 21379 18874 21384
rect 18272 21376 18860 21379
rect 6596 20677 7200 21099
rect 7334 21048 7954 21053
rect 7334 20864 7344 21048
rect 7944 20864 7954 21048
rect 7334 20859 7954 20864
rect 6590 20672 7210 20677
rect 6590 20488 6600 20672
rect 7200 20488 7210 20672
rect 6590 20483 7210 20488
rect 6596 20057 7200 20483
rect 7344 20437 7944 20859
rect 8316 20677 8920 21099
rect 9054 21048 9674 21053
rect 9054 20864 9064 21048
rect 9664 20864 9674 21048
rect 9054 20859 9674 20864
rect 10268 20860 10380 21220
rect 10840 20860 10908 21220
rect 8310 20672 8930 20677
rect 8310 20488 8320 20672
rect 8920 20488 8930 20672
rect 8310 20483 8930 20488
rect 7334 20432 7954 20437
rect 7334 20248 7344 20432
rect 7944 20248 7954 20432
rect 7334 20243 7954 20248
rect 6590 20052 7210 20057
rect 6590 19868 6600 20052
rect 7200 19868 7210 20052
rect 6590 19863 7210 19868
rect 6596 19441 7200 19863
rect 7344 19817 7944 20243
rect 8316 20057 8920 20483
rect 9064 20437 9664 20859
rect 9054 20432 9674 20437
rect 9054 20248 9064 20432
rect 9664 20248 9674 20432
rect 9054 20243 9674 20248
rect 8310 20052 8930 20057
rect 8310 19868 8320 20052
rect 8920 19868 8930 20052
rect 8310 19863 8930 19868
rect 7334 19812 7954 19817
rect 7334 19628 7344 19812
rect 7944 19628 7954 19812
rect 7334 19623 7954 19628
rect 6590 19436 7210 19441
rect 6590 19252 6600 19436
rect 7200 19252 7210 19436
rect 6590 19247 7210 19252
rect 6596 18821 7200 19247
rect 7344 19201 7944 19623
rect 8316 19441 8920 19863
rect 9064 19817 9664 20243
rect 10268 19873 10908 20860
rect 18984 21325 19640 21688
rect 18984 21320 19642 21325
rect 18984 21092 19000 21320
rect 19632 21092 19642 21320
rect 18984 21087 19642 21092
rect 18984 20752 19640 21087
rect 18984 20524 18996 20752
rect 19628 20524 19640 20752
rect 18300 20453 18896 20456
rect 18298 20448 18898 20453
rect 18298 20220 18308 20448
rect 18888 20220 18898 20448
rect 18298 20215 18898 20220
rect 10266 19868 10908 19873
rect 9054 19812 9674 19817
rect 9054 19628 9064 19812
rect 9664 19628 9674 19812
rect 9054 19623 9674 19628
rect 8310 19436 8930 19441
rect 8310 19252 8320 19436
rect 8920 19252 8930 19436
rect 8310 19247 8930 19252
rect 7334 19196 7954 19201
rect 7334 19012 7344 19196
rect 7944 19012 7954 19196
rect 7334 19007 7954 19012
rect 6590 18816 7210 18821
rect 6590 18632 6600 18816
rect 7200 18632 7210 18816
rect 6590 18627 7210 18632
rect 6596 18205 7200 18627
rect 7344 18581 7944 19007
rect 8316 18821 8920 19247
rect 9064 19201 9664 19623
rect 10266 19580 10276 19868
rect 10876 19580 10908 19868
rect 18300 19833 18896 20215
rect 18984 20128 19640 20524
rect 18984 19900 18996 20128
rect 19628 19900 19640 20128
rect 18298 19828 18898 19833
rect 18298 19600 18308 19828
rect 18888 19600 18898 19828
rect 18298 19595 18898 19600
rect 10266 19576 10908 19580
rect 10266 19575 10886 19576
rect 10024 19473 10640 19484
rect 10014 19468 10650 19473
rect 9054 19196 9674 19201
rect 9054 19012 9064 19196
rect 9664 19012 9674 19196
rect 10014 19172 10024 19468
rect 10640 19172 10650 19468
rect 18300 19217 18896 19595
rect 18984 19512 19640 19900
rect 18984 19284 18996 19512
rect 19628 19284 19640 19512
rect 10014 19167 10650 19172
rect 18298 19212 18898 19217
rect 9054 19007 9674 19012
rect 8310 18816 8930 18821
rect 8310 18632 8320 18816
rect 8920 18632 8930 18816
rect 8310 18627 8930 18632
rect 7334 18576 7954 18581
rect 7334 18392 7344 18576
rect 7944 18392 7954 18576
rect 7334 18387 7954 18392
rect 7344 18220 7944 18387
rect 6590 18200 7210 18205
rect 6590 18016 6600 18200
rect 7200 18016 7210 18200
rect 6590 18011 7210 18016
rect 6596 17992 7200 18011
rect 7344 17965 7356 18220
rect 7334 17960 7356 17965
rect 7888 17965 7944 18220
rect 8316 18205 8920 18627
rect 9064 18581 9664 19007
rect 10024 18876 10640 19167
rect 18298 18984 18308 19212
rect 18888 18984 18898 19212
rect 18298 18979 18898 18984
rect 10024 18644 10040 18876
rect 10624 18644 10640 18876
rect 9054 18576 9674 18581
rect 9054 18392 9064 18576
rect 9664 18392 9674 18576
rect 9054 18387 9674 18392
rect 8310 18200 8930 18205
rect 8310 18016 8320 18200
rect 8920 18016 8930 18200
rect 8310 18011 8930 18016
rect 9064 18200 9664 18387
rect 8316 17992 8920 18011
rect 9064 17965 9076 18200
rect 7888 17960 7954 17965
rect 7334 17776 7344 17960
rect 7944 17776 7954 17960
rect 9054 17960 9076 17965
rect 9608 17965 9664 18200
rect 10024 18256 10640 18644
rect 15570 18860 15990 18865
rect 10024 18032 10040 18256
rect 10624 18032 10640 18256
rect 10024 18016 10640 18032
rect 10748 18560 11316 18576
rect 10748 18336 10768 18560
rect 11296 18336 11316 18560
rect 15570 18420 15580 18860
rect 15980 18420 15990 18860
rect 15570 18415 15990 18420
rect 16210 18860 16630 18865
rect 16210 18420 16220 18860
rect 16620 18420 16630 18860
rect 18300 18597 18896 18979
rect 18984 18921 19640 19284
rect 18984 18916 19642 18921
rect 18984 18688 19000 18916
rect 19632 18688 19642 18916
rect 18984 18683 19642 18688
rect 18984 18676 19640 18683
rect 16210 18415 16630 18420
rect 18298 18592 18898 18597
rect 18298 18364 18308 18592
rect 18888 18364 18898 18592
rect 18298 18359 18898 18364
rect 10748 18132 11316 18336
rect 18300 18180 18896 18359
rect 19860 18244 24148 22268
rect 24212 21500 24232 22268
rect 24550 21500 24890 21505
rect 24212 21140 24560 21500
rect 24880 21140 24890 21500
rect 24212 18244 24232 21140
rect 24550 21135 24890 21140
rect 19860 18216 24232 18244
rect 9608 17960 9674 17965
rect 7334 17771 7954 17776
rect 8030 17776 8230 17781
rect 8030 17616 8040 17776
rect 8220 17616 8230 17776
rect 9054 17776 9064 17960
rect 9664 17776 9674 17960
rect 9054 17771 9076 17776
rect 9066 17764 9076 17771
rect 9608 17771 9674 17776
rect 9608 17764 9618 17771
rect 8030 17611 8230 17616
rect 10748 17592 10764 18132
rect 11300 17592 11316 18132
rect 18290 17720 18300 18180
rect 18900 17720 18910 18180
rect 10748 17576 11316 17592
rect 26380 14740 28460 27440
rect -10460 11148 28460 14740
rect -10460 10768 2588 11148
rect -10460 10740 1300 10768
rect -1860 10532 1300 10740
rect 1568 10660 2588 10768
rect 4792 10808 16988 11148
rect 4792 10660 6096 10808
rect 1568 10608 6096 10660
rect 6276 10768 16988 10808
rect 6276 10740 15700 10768
rect 6276 10608 7320 10740
rect 1568 10532 7320 10608
rect -1860 10508 7320 10532
rect -1860 10180 -540 10508
rect 4904 10364 7320 10508
rect -2584 10160 1496 10180
rect -2584 10096 -2556 10160
rect 1468 10096 1496 10160
rect 4904 10160 6212 10364
rect 4904 10156 5304 10160
rect 6202 10120 6212 10160
rect 7188 10160 7320 10364
rect 12540 10532 15700 10740
rect 15968 10660 16988 10768
rect 19192 10808 28460 11148
rect 19192 10660 20496 10808
rect 15968 10608 20496 10660
rect 20676 10740 28460 10808
rect 20676 10608 21720 10740
rect 24540 10720 28460 10740
rect 15968 10532 21720 10608
rect 12540 10508 21720 10532
rect 8750 10292 9642 10297
rect 7188 10120 7228 10160
rect 6202 10115 7228 10120
rect -8160 8660 -3788 8688
rect -8160 8376 -3872 8660
rect -8660 8301 -3872 8376
rect -8670 8296 -3872 8301
rect -8670 8196 -8660 8296
rect -8480 8196 -3872 8296
rect -8670 8191 -8470 8196
rect -9984 7852 -9292 7876
rect -9984 7584 -9968 7852
rect -9316 7584 -9292 7852
rect -9984 6740 -9292 7584
rect -9984 6472 -9968 6740
rect -9316 6472 -9292 6740
rect -9984 6444 -9292 6472
rect -10064 5929 -9460 5932
rect -10074 5924 -9450 5929
rect -10074 5740 -10064 5924
rect -9460 5740 -9450 5924
rect -10074 5735 -9450 5740
rect -10064 5313 -9460 5735
rect -10074 5308 -9450 5313
rect -10074 5124 -10064 5308
rect -9460 5124 -9450 5308
rect -10074 5119 -9450 5124
rect -10064 4693 -9460 5119
rect -10078 4688 -9454 4693
rect -10078 4504 -10068 4688
rect -9464 4504 -9454 4688
rect -10078 4499 -9454 4504
rect -8160 4636 -3872 8196
rect -3808 4636 -3788 8660
rect -2584 5808 1496 10096
rect 5102 10056 6098 10057
rect 5092 10052 6098 10056
rect 5092 9796 5112 10052
rect 6088 9796 6098 10052
rect 5092 9791 6098 9796
rect 5092 9425 6088 9791
rect 6212 9737 7228 10115
rect 8750 10092 8760 10292
rect 9632 10092 9642 10292
rect 12540 10180 13920 10508
rect 19304 10364 21720 10508
rect 8750 10087 9642 10092
rect 11816 10160 15896 10180
rect 11816 10096 11844 10160
rect 15868 10096 15896 10160
rect 19304 10160 20612 10364
rect 19304 10156 19704 10160
rect 20602 10120 20612 10160
rect 21588 10160 21720 10364
rect 23150 10292 24042 10297
rect 21588 10120 21628 10160
rect 20602 10115 21628 10120
rect 7600 10037 8600 10040
rect 7598 10032 8602 10037
rect 7598 9844 7608 10032
rect 8592 9844 8602 10032
rect 7598 9839 8602 9844
rect 6202 9732 7228 9737
rect 6202 9488 6212 9732
rect 7188 9488 7228 9732
rect 6202 9483 7228 9488
rect 6212 9476 7228 9483
rect 5092 9420 6098 9425
rect 5092 9160 5112 9420
rect 6088 9160 6098 9420
rect 5092 9020 5120 9160
rect 4548 8984 5120 9020
rect 4548 8432 4588 8984
rect 5008 8740 5120 8984
rect 6060 9155 6098 9160
rect 7600 9417 8600 9839
rect 8760 9681 9636 10087
rect 8754 9676 9646 9681
rect 8754 9476 8764 9676
rect 9636 9476 9646 9676
rect 8754 9471 9646 9476
rect 7600 9412 8606 9417
rect 7600 9224 7612 9412
rect 8596 9224 8606 9412
rect 7600 9219 8606 9224
rect 6060 8740 6088 9155
rect 7600 8801 8600 9219
rect 8760 9065 9636 9471
rect 8754 9060 9646 9065
rect 8754 8860 8764 9060
rect 9636 8860 9646 9060
rect 8754 8855 9646 8860
rect 7598 8796 8602 8801
rect 5008 8477 6088 8740
rect 6214 8784 7210 8789
rect 6214 8536 6224 8784
rect 7200 8720 7210 8784
rect 7598 8720 7608 8796
rect 7200 8608 7608 8720
rect 8592 8608 8602 8796
rect 7200 8603 8602 8608
rect 7200 8536 8600 8603
rect 6214 8531 8600 8536
rect 5008 8472 6090 8477
rect 5008 8432 5104 8472
rect 4548 8376 5104 8432
rect 4940 8224 5104 8376
rect 6080 8224 6090 8472
rect 4940 8220 6090 8224
rect 5092 8219 6090 8220
rect 5092 7853 6088 8219
rect 6224 8180 8600 8531
rect 8760 8445 9636 8855
rect 8754 8440 9646 8445
rect 8754 8240 8764 8440
rect 9636 8240 9646 8440
rect 8754 8235 9646 8240
rect 6224 8169 7604 8180
rect 6214 8164 7604 8169
rect 6214 7916 6224 8164
rect 7200 7992 7604 8164
rect 8588 7992 8600 8180
rect 7200 7916 8600 7992
rect 6214 7911 8600 7916
rect 6224 7904 8600 7911
rect 5092 7848 6090 7853
rect 5092 7656 5104 7848
rect 5094 7600 5104 7656
rect 6080 7600 6090 7848
rect 5094 7595 6090 7600
rect 7600 7561 8600 7904
rect 8760 7825 9636 8235
rect 8754 7820 9646 7825
rect 8754 7620 8764 7820
rect 9636 7620 9646 7820
rect 8754 7615 9646 7620
rect 7598 7556 8602 7561
rect 6384 7517 7392 7552
rect 6374 7512 7392 7517
rect 6374 7000 6384 7512
rect 7076 7000 7392 7512
rect 7598 7368 7608 7556
rect 8592 7368 8602 7556
rect 7598 7363 8602 7368
rect 6374 6995 7392 7000
rect 212 5649 816 5652
rect 2012 5649 2616 5652
rect 3812 5649 4416 5652
rect 5612 5649 6216 5652
rect 202 5644 826 5649
rect 202 5460 212 5644
rect 816 5460 826 5644
rect 202 5455 826 5460
rect 2002 5644 2626 5649
rect 2002 5460 2012 5644
rect 2616 5460 2626 5644
rect 2002 5455 2626 5460
rect 3802 5644 4426 5649
rect 3802 5460 3812 5644
rect 4416 5460 4426 5644
rect 3802 5455 4426 5460
rect 5602 5644 6226 5649
rect 5602 5460 5612 5644
rect 6216 5460 6226 5644
rect 5602 5455 6226 5460
rect 212 5033 816 5455
rect 2012 5033 2616 5455
rect 3812 5033 4416 5455
rect 5612 5033 6216 5455
rect 202 5028 826 5033
rect 202 4844 212 5028
rect 816 4844 826 5028
rect 202 4839 826 4844
rect 2002 5028 2626 5033
rect 2002 4844 2012 5028
rect 2616 4844 2626 5028
rect 2002 4839 2626 4844
rect 3802 5028 4426 5033
rect 3802 4844 3812 5028
rect 4416 4844 4426 5028
rect 3802 4839 4426 4844
rect 5602 5028 6226 5033
rect 5602 4844 5612 5028
rect 6216 4844 6226 5028
rect 5602 4839 6226 4844
rect -8160 4608 -3788 4636
rect -818 4816 -22 4821
rect -10064 4025 -9460 4499
rect -8160 4368 -7992 4608
rect -3182 4532 -3018 4537
rect -3182 4420 -3172 4532
rect -3028 4420 -3018 4532
rect -3182 4415 -3018 4420
rect -818 4404 -808 4816
rect -32 4404 -22 4816
rect 212 4413 816 4839
rect 2012 4413 2616 4839
rect 3812 4413 4416 4839
rect 5612 4413 6216 4839
rect 6384 4456 7392 6995
rect 7600 6949 8600 7363
rect 8760 7209 9636 7615
rect 8754 7204 9646 7209
rect 8754 7004 8764 7204
rect 9636 7004 9646 7204
rect 8754 6999 9646 7004
rect 7598 6944 8602 6949
rect 7598 6756 7608 6944
rect 8592 6756 8602 6944
rect 7598 6751 8602 6756
rect 7600 6325 8600 6751
rect 8760 6593 9636 6999
rect 8754 6588 9646 6593
rect 8754 6388 8764 6588
rect 9636 6388 9646 6588
rect 8754 6383 9646 6388
rect 7594 6320 8600 6325
rect 7594 6132 7604 6320
rect 8588 6132 8600 6320
rect 7594 6127 8600 6132
rect 7600 5713 8600 6127
rect 8760 6020 9636 6383
rect 8760 5973 8772 6020
rect 8750 5968 8772 5973
rect 9616 5973 9636 6020
rect 9616 5968 9642 5973
rect 8750 5768 8760 5968
rect 9632 5768 9642 5968
rect 11816 5808 15896 10096
rect 19502 10056 20498 10057
rect 19492 10052 20498 10056
rect 19492 9796 19512 10052
rect 20488 9796 20498 10052
rect 19492 9791 20498 9796
rect 19492 9425 20488 9791
rect 20612 9737 21628 10115
rect 23150 10092 23160 10292
rect 24032 10092 24042 10292
rect 23150 10087 24042 10092
rect 22000 10037 23000 10040
rect 21998 10032 23002 10037
rect 21998 9844 22008 10032
rect 22992 9844 23002 10032
rect 21998 9839 23002 9844
rect 20602 9732 21628 9737
rect 20602 9488 20612 9732
rect 21588 9488 21628 9732
rect 20602 9483 21628 9488
rect 20612 9476 21628 9483
rect 19492 9420 20498 9425
rect 19492 9160 19512 9420
rect 20488 9160 20498 9420
rect 19492 9155 20498 9160
rect 22000 9417 23000 9839
rect 23160 9681 24036 10087
rect 23154 9676 24046 9681
rect 23154 9476 23164 9676
rect 24036 9476 24046 9676
rect 23154 9471 24046 9476
rect 22000 9412 23006 9417
rect 22000 9224 22012 9412
rect 22996 9224 23006 9412
rect 22000 9219 23006 9224
rect 19492 9020 20488 9155
rect 18948 8984 20488 9020
rect 18948 8432 18988 8984
rect 19408 8477 20488 8984
rect 22000 8801 23000 9219
rect 23160 9065 24036 9471
rect 23154 9060 24046 9065
rect 23154 8860 23164 9060
rect 24036 8860 24046 9060
rect 23154 8855 24046 8860
rect 21998 8796 23002 8801
rect 20614 8784 21610 8789
rect 20614 8536 20624 8784
rect 21600 8720 21610 8784
rect 21998 8720 22008 8796
rect 21600 8608 22008 8720
rect 22992 8608 23002 8796
rect 21600 8603 23002 8608
rect 21600 8536 23000 8603
rect 20614 8531 23000 8536
rect 19408 8472 20490 8477
rect 19408 8432 19504 8472
rect 18948 8376 19504 8432
rect 19340 8224 19504 8376
rect 20480 8224 20490 8472
rect 19340 8220 20490 8224
rect 19492 8219 20490 8220
rect 19492 7853 20488 8219
rect 20624 8180 23000 8531
rect 23160 8445 24036 8855
rect 23154 8440 24046 8445
rect 23154 8240 23164 8440
rect 24036 8240 24046 8440
rect 23154 8235 24046 8240
rect 20624 8169 22004 8180
rect 20614 8164 22004 8169
rect 20614 7916 20624 8164
rect 21600 7992 22004 8164
rect 22988 7992 23000 8180
rect 21600 7916 23000 7992
rect 20614 7911 23000 7916
rect 20624 7904 23000 7911
rect 19492 7848 20490 7853
rect 19492 7656 19504 7848
rect 19494 7600 19504 7656
rect 20480 7600 20490 7848
rect 19494 7595 20490 7600
rect 22000 7561 23000 7904
rect 23160 7825 24036 8235
rect 23154 7820 24046 7825
rect 23154 7620 23164 7820
rect 24036 7620 24046 7820
rect 23154 7615 24046 7620
rect 21998 7556 23002 7561
rect 20784 7517 21792 7552
rect 20774 7512 21792 7517
rect 20774 7000 20784 7512
rect 21476 7000 21792 7512
rect 21998 7368 22008 7556
rect 22992 7368 23002 7556
rect 21998 7363 23002 7368
rect 20774 6995 21792 7000
rect 8750 5763 8772 5768
rect 7594 5708 8600 5713
rect 7594 5520 7604 5708
rect 8588 5520 8600 5708
rect 7594 5515 8600 5520
rect 7600 5089 8600 5515
rect 8760 5353 8772 5763
rect 8750 5348 8772 5353
rect 9616 5763 9642 5768
rect 9616 5353 9636 5763
rect 14612 5649 15216 5652
rect 16412 5649 17016 5652
rect 18212 5649 18816 5652
rect 20012 5649 20616 5652
rect 14602 5644 15226 5649
rect 14602 5460 14612 5644
rect 15216 5460 15226 5644
rect 14602 5455 15226 5460
rect 16402 5644 17026 5649
rect 16402 5460 16412 5644
rect 17016 5460 17026 5644
rect 16402 5455 17026 5460
rect 18202 5644 18826 5649
rect 18202 5460 18212 5644
rect 18816 5460 18826 5644
rect 18202 5455 18826 5460
rect 20002 5644 20626 5649
rect 20002 5460 20012 5644
rect 20616 5460 20626 5644
rect 20002 5455 20626 5460
rect 9616 5348 9642 5353
rect 8750 5148 8760 5348
rect 9632 5148 9642 5348
rect 8750 5143 9642 5148
rect 8760 5140 9636 5143
rect 7594 5084 8600 5089
rect 7594 4896 7604 5084
rect 8588 4904 8600 5084
rect 14612 5033 15216 5455
rect 16412 5033 17016 5455
rect 18212 5033 18816 5455
rect 20012 5033 20616 5455
rect 14602 5028 15226 5033
rect 8588 4896 8598 4904
rect 7594 4891 8598 4896
rect 10200 4860 11860 4900
rect 10200 4580 11480 4860
rect 11820 4580 11860 4860
rect 14602 4844 14612 5028
rect 15216 4844 15226 5028
rect 14602 4839 15226 4844
rect 16402 5028 17026 5033
rect 16402 4844 16412 5028
rect 17016 4844 17026 5028
rect 16402 4839 17026 4844
rect 18202 5028 18826 5033
rect 18202 4844 18212 5028
rect 18816 4844 18826 5028
rect 18202 4839 18826 4844
rect 20002 5028 20626 5033
rect 20002 4844 20012 5028
rect 20616 4844 20626 5028
rect 20002 4839 20626 4844
rect 10200 4520 11860 4580
rect 13582 4816 14378 4821
rect -818 4399 -22 4404
rect 198 4408 822 4413
rect -8160 4340 -3788 4368
rect -10070 4020 -9450 4025
rect -10070 3836 -10060 4020
rect -9460 3836 -9450 4020
rect -10070 3831 -9450 3836
rect -10064 3409 -9460 3831
rect -9326 3780 -8706 3785
rect -9326 3596 -9316 3780
rect -8716 3596 -8706 3780
rect -9326 3591 -8706 3596
rect -10070 3404 -9450 3409
rect -10070 3220 -10060 3404
rect -9460 3220 -9450 3404
rect -10070 3215 -9450 3220
rect -10064 2789 -9460 3215
rect -9316 3169 -8716 3591
rect -9326 3164 -8706 3169
rect -9326 2980 -9316 3164
rect -8716 2980 -8706 3164
rect -9326 2975 -8706 2980
rect -10070 2784 -9450 2789
rect -10070 2600 -10060 2784
rect -9460 2600 -9450 2784
rect -10070 2595 -9450 2600
rect -10064 2173 -9460 2595
rect -9316 2549 -8716 2975
rect -9326 2544 -8706 2549
rect -9326 2360 -9316 2544
rect -8716 2360 -8706 2544
rect -9326 2355 -8706 2360
rect -10070 2168 -9450 2173
rect -10070 1984 -10060 2168
rect -9460 1984 -9450 2168
rect -10070 1979 -9450 1984
rect -10064 1553 -9460 1979
rect -9316 1933 -8716 2355
rect -9326 1928 -8706 1933
rect -9326 1744 -9316 1928
rect -8716 1744 -8706 1928
rect -9326 1739 -8706 1744
rect -10070 1548 -9450 1553
rect -10070 1364 -10060 1548
rect -9460 1364 -9450 1548
rect -10070 1359 -9450 1364
rect -10064 937 -9460 1359
rect -9316 1313 -8716 1739
rect -9326 1308 -8706 1313
rect -9326 1124 -9316 1308
rect -8716 1124 -8706 1308
rect -9326 1119 -8706 1124
rect -10070 932 -9450 937
rect -10070 748 -10060 932
rect -9460 748 -9450 932
rect -10070 743 -9450 748
rect -10064 724 -9460 743
rect -9316 697 -8716 1119
rect -9326 692 -8706 697
rect -9326 508 -9316 692
rect -8716 508 -8706 692
rect -9326 503 -8706 508
rect -8510 508 -8350 513
rect -9316 284 -8716 503
rect -8510 348 -8500 508
rect -8360 348 -8350 508
rect -8510 343 -8350 348
rect -8160 316 -3872 4340
rect -3808 316 -3788 4340
rect -804 4128 -28 4399
rect 198 4224 208 4408
rect 812 4224 822 4408
rect 198 4219 822 4224
rect 1998 4408 2622 4413
rect 1998 4224 2008 4408
rect 2612 4224 2622 4408
rect 1998 4219 2622 4224
rect 3798 4408 4422 4413
rect 3798 4224 3808 4408
rect 4412 4224 4422 4408
rect 3798 4219 4422 4224
rect 5598 4408 6222 4413
rect 5598 4224 5608 4408
rect 6212 4224 6222 4408
rect 5598 4219 6222 4224
rect -8160 288 -3788 316
rect -3400 4100 -28 4128
rect -9326 4 -9316 284
rect -8716 4 -8706 284
rect -3400 76 -112 4100
rect -48 76 -28 4100
rect 212 3745 816 4219
rect 2012 3745 2616 4219
rect 3812 3745 4416 4219
rect 5612 3745 6216 4219
rect 6384 4108 7396 4456
rect 10200 4108 10520 4520
rect 13582 4404 13592 4816
rect 14368 4404 14378 4816
rect 14612 4413 15216 4839
rect 16412 4413 17016 4839
rect 18212 4413 18816 4839
rect 20012 4413 20616 4839
rect 20784 4456 21792 6995
rect 22000 6949 23000 7363
rect 23160 7209 24036 7615
rect 23154 7204 24046 7209
rect 23154 7004 23164 7204
rect 24036 7004 24046 7204
rect 23154 6999 24046 7004
rect 21998 6944 23002 6949
rect 21998 6756 22008 6944
rect 22992 6756 23002 6944
rect 21998 6751 23002 6756
rect 22000 6325 23000 6751
rect 23160 6593 24036 6999
rect 23154 6588 24046 6593
rect 23154 6388 23164 6588
rect 24036 6388 24046 6588
rect 23154 6383 24046 6388
rect 21994 6320 23000 6325
rect 21994 6132 22004 6320
rect 22988 6132 23000 6320
rect 21994 6127 23000 6132
rect 22000 5713 23000 6127
rect 23160 6020 24036 6383
rect 23160 5973 23172 6020
rect 23150 5968 23172 5973
rect 24016 5973 24036 6020
rect 24016 5968 24042 5973
rect 23150 5768 23160 5968
rect 24032 5768 24042 5968
rect 23150 5763 23172 5768
rect 21994 5708 23000 5713
rect 21994 5520 22004 5708
rect 22988 5520 23000 5708
rect 21994 5515 23000 5520
rect 22000 5089 23000 5515
rect 23160 5353 23172 5763
rect 23150 5348 23172 5353
rect 24016 5763 24042 5768
rect 24016 5353 24036 5763
rect 24016 5348 24042 5353
rect 23150 5148 23160 5348
rect 24032 5148 24042 5348
rect 23150 5143 24042 5148
rect 23160 5140 24036 5143
rect 21994 5084 23000 5089
rect 21994 4896 22004 5084
rect 22988 4904 23000 5084
rect 22988 4896 22998 4904
rect 21994 4891 22998 4896
rect 24510 4700 24910 4705
rect 13582 4399 14378 4404
rect 14598 4408 15222 4413
rect 13596 4128 14372 4399
rect 14598 4224 14608 4408
rect 15212 4224 15222 4408
rect 14598 4219 15222 4224
rect 16398 4408 17022 4413
rect 16398 4224 16408 4408
rect 17012 4224 17022 4408
rect 16398 4219 17022 4224
rect 18198 4408 18822 4413
rect 18198 4224 18208 4408
rect 18812 4224 18822 4408
rect 18198 4219 18822 4224
rect 19998 4408 20622 4413
rect 19998 4224 20008 4408
rect 20612 4224 20622 4408
rect 19998 4219 20622 4224
rect 6384 4080 10552 4108
rect 6384 4052 10468 4080
rect 206 3740 826 3745
rect 206 3556 216 3740
rect 816 3556 826 3740
rect 206 3551 826 3556
rect 2006 3740 2626 3745
rect 2006 3556 2016 3740
rect 2616 3556 2626 3740
rect 2006 3551 2626 3556
rect 3806 3740 4426 3745
rect 3806 3556 3816 3740
rect 4416 3556 4426 3740
rect 3806 3551 4426 3556
rect 5606 3740 6226 3745
rect 6388 3740 10468 4052
rect 5606 3556 5616 3740
rect 6216 3556 6226 3740
rect 5606 3551 6226 3556
rect 212 3129 816 3551
rect 950 3500 1570 3505
rect 950 3316 960 3500
rect 1560 3316 1570 3500
rect 950 3311 1570 3316
rect 206 3124 826 3129
rect 206 2940 216 3124
rect 816 2940 826 3124
rect 206 2935 826 2940
rect 212 2509 816 2935
rect 960 2889 1560 3311
rect 2012 3129 2616 3551
rect 2750 3500 3370 3505
rect 2750 3316 2760 3500
rect 3360 3316 3370 3500
rect 2750 3311 3370 3316
rect 2006 3124 2626 3129
rect 2006 2940 2016 3124
rect 2616 2940 2626 3124
rect 2006 2935 2626 2940
rect 950 2884 1570 2889
rect 950 2700 960 2884
rect 1560 2700 1570 2884
rect 950 2695 1570 2700
rect 206 2504 826 2509
rect 206 2320 216 2504
rect 816 2320 826 2504
rect 206 2315 826 2320
rect 212 1893 816 2315
rect 960 2269 1560 2695
rect 2012 2509 2616 2935
rect 2760 2889 3360 3311
rect 3812 3129 4416 3551
rect 4550 3500 5170 3505
rect 4550 3316 4560 3500
rect 5160 3316 5170 3500
rect 4550 3311 5170 3316
rect 3806 3124 4426 3129
rect 3806 2940 3816 3124
rect 4416 2940 4426 3124
rect 3806 2935 4426 2940
rect 2750 2884 3370 2889
rect 2750 2700 2760 2884
rect 3360 2700 3370 2884
rect 2750 2695 3370 2700
rect 2006 2504 2626 2509
rect 2006 2320 2016 2504
rect 2616 2320 2626 2504
rect 2006 2315 2626 2320
rect 950 2264 1570 2269
rect 950 2080 960 2264
rect 1560 2080 1570 2264
rect 950 2075 1570 2080
rect 206 1888 826 1893
rect 206 1704 216 1888
rect 816 1704 826 1888
rect 206 1699 826 1704
rect 212 1273 816 1699
rect 960 1653 1560 2075
rect 2012 1893 2616 2315
rect 2760 2269 3360 2695
rect 3812 2509 4416 2935
rect 4560 2889 5160 3311
rect 5612 3129 6216 3551
rect 6350 3500 6970 3505
rect 6350 3316 6360 3500
rect 6960 3316 6970 3500
rect 6350 3311 6970 3316
rect 5606 3124 6226 3129
rect 5606 2940 5616 3124
rect 6216 2940 6226 3124
rect 5606 2935 6226 2940
rect 4550 2884 5170 2889
rect 4550 2700 4560 2884
rect 5160 2700 5170 2884
rect 4550 2695 5170 2700
rect 3806 2504 4426 2509
rect 3806 2320 3816 2504
rect 4416 2320 4426 2504
rect 3806 2315 4426 2320
rect 2750 2264 3370 2269
rect 2750 2080 2760 2264
rect 3360 2080 3370 2264
rect 2750 2075 3370 2080
rect 2006 1888 2626 1893
rect 2006 1704 2016 1888
rect 2616 1704 2626 1888
rect 2006 1699 2626 1704
rect 950 1648 1570 1653
rect 950 1464 960 1648
rect 1560 1464 1570 1648
rect 950 1459 1570 1464
rect 206 1268 826 1273
rect 206 1084 216 1268
rect 816 1084 826 1268
rect 206 1079 826 1084
rect 212 657 816 1079
rect 960 1033 1560 1459
rect 2012 1273 2616 1699
rect 2760 1653 3360 2075
rect 3812 1893 4416 2315
rect 4560 2269 5160 2695
rect 5612 2509 6216 2935
rect 6360 2889 6960 3311
rect 6350 2884 6970 2889
rect 6350 2700 6360 2884
rect 6960 2700 6970 2884
rect 6350 2695 6970 2700
rect 5606 2504 6226 2509
rect 5606 2320 5616 2504
rect 6216 2320 6226 2504
rect 5606 2315 6226 2320
rect 4550 2264 5170 2269
rect 4550 2080 4560 2264
rect 5160 2080 5170 2264
rect 4550 2075 5170 2080
rect 3806 1888 4426 1893
rect 3806 1704 3816 1888
rect 4416 1704 4426 1888
rect 3806 1699 4426 1704
rect 2750 1648 3370 1653
rect 2750 1464 2760 1648
rect 3360 1464 3370 1648
rect 2750 1459 3370 1464
rect 2006 1268 2626 1273
rect 2006 1084 2016 1268
rect 2616 1084 2626 1268
rect 2006 1079 2626 1084
rect 950 1028 1570 1033
rect 950 844 960 1028
rect 1560 844 1570 1028
rect 950 839 1570 844
rect 960 680 1560 839
rect 206 652 826 657
rect 206 468 216 652
rect 816 468 826 652
rect 206 463 826 468
rect 212 444 816 463
rect 960 417 976 680
rect 950 412 976 417
rect 1548 417 1560 680
rect 2012 657 2616 1079
rect 2760 1033 3360 1459
rect 3812 1273 4416 1699
rect 4560 1653 5160 2075
rect 5612 1893 6216 2315
rect 6360 2269 6960 2695
rect 6350 2264 6970 2269
rect 6350 2080 6360 2264
rect 6960 2080 6970 2264
rect 6350 2075 6970 2080
rect 5606 1888 6226 1893
rect 5606 1704 5616 1888
rect 6216 1704 6226 1888
rect 5606 1699 6226 1704
rect 4550 1648 5170 1653
rect 4550 1464 4560 1648
rect 5160 1464 5170 1648
rect 4550 1459 5170 1464
rect 3806 1268 4426 1273
rect 3806 1084 3816 1268
rect 4416 1084 4426 1268
rect 3806 1079 4426 1084
rect 2750 1028 3370 1033
rect 2750 844 2760 1028
rect 3360 844 3370 1028
rect 2750 839 3370 844
rect 2760 680 3360 839
rect 2006 652 2626 657
rect 2006 468 2016 652
rect 2616 468 2626 652
rect 2006 463 2626 468
rect 2012 444 2616 463
rect 2760 417 2776 680
rect 1548 412 1570 417
rect 950 228 960 412
rect 1560 228 1570 412
rect 2750 412 2776 417
rect 3348 417 3360 680
rect 3812 657 4416 1079
rect 4560 1033 5160 1459
rect 5612 1273 6216 1699
rect 6360 1653 6960 2075
rect 6350 1648 6970 1653
rect 6350 1464 6360 1648
rect 6960 1464 6970 1648
rect 6350 1459 6970 1464
rect 5606 1268 6226 1273
rect 5606 1084 5616 1268
rect 6216 1084 6226 1268
rect 5606 1079 6226 1084
rect 4550 1028 5170 1033
rect 4550 844 4560 1028
rect 5160 844 5170 1028
rect 4550 839 5170 844
rect 4560 676 5160 839
rect 3806 652 4426 657
rect 3806 468 3816 652
rect 4416 468 4426 652
rect 3806 463 4426 468
rect 3812 444 4416 463
rect 4560 417 4572 676
rect 3348 412 3370 417
rect 950 223 1570 228
rect 1686 268 1886 273
rect -3400 48 -28 76
rect 1686 68 1696 268
rect 1876 68 1886 268
rect 2750 228 2760 412
rect 3360 228 3370 412
rect 4550 412 4572 417
rect 5144 417 5160 676
rect 5612 657 6216 1079
rect 6360 1033 6960 1459
rect 6350 1028 6970 1033
rect 6350 844 6360 1028
rect 6960 844 6970 1028
rect 6350 839 6970 844
rect 6360 676 6960 839
rect 5606 652 6226 657
rect 5606 468 5616 652
rect 6216 468 6226 652
rect 5606 463 6226 468
rect 5612 444 6216 463
rect 6360 417 6372 676
rect 5144 412 5170 417
rect 2750 223 3370 228
rect 1686 63 1886 68
rect 3502 64 3512 276
rect 3692 64 3702 276
rect 4550 228 4560 412
rect 5160 228 5170 412
rect 6350 412 6372 417
rect 6944 417 6960 676
rect 6944 412 6970 417
rect 4550 223 5170 228
rect 5278 276 5478 281
rect 5278 64 5288 276
rect 5468 64 5478 276
rect 6350 228 6360 412
rect 6960 228 6970 412
rect 6350 223 6970 228
rect 5278 59 5478 64
rect 7180 56 10468 3740
rect 10532 56 10552 4080
rect 7180 28 10552 56
rect 11000 4100 14372 4128
rect 11000 76 14288 4100
rect 14352 76 14372 4100
rect 14612 3745 15216 4219
rect 16412 3745 17016 4219
rect 18212 3745 18816 4219
rect 20012 3745 20616 4219
rect 20784 4108 21796 4456
rect 24510 4360 24520 4700
rect 24900 4360 24910 4700
rect 24510 4355 24910 4360
rect 24520 4108 24900 4355
rect 20784 4080 24952 4108
rect 20784 4052 24868 4080
rect 14606 3740 15226 3745
rect 14606 3556 14616 3740
rect 15216 3556 15226 3740
rect 14606 3551 15226 3556
rect 16406 3740 17026 3745
rect 16406 3556 16416 3740
rect 17016 3556 17026 3740
rect 16406 3551 17026 3556
rect 18206 3740 18826 3745
rect 18206 3556 18216 3740
rect 18816 3556 18826 3740
rect 18206 3551 18826 3556
rect 20006 3740 20626 3745
rect 20788 3740 24868 4052
rect 20006 3556 20016 3740
rect 20616 3556 20626 3740
rect 20006 3551 20626 3556
rect 14612 3129 15216 3551
rect 15350 3500 15970 3505
rect 15350 3316 15360 3500
rect 15960 3316 15970 3500
rect 15350 3311 15970 3316
rect 14606 3124 15226 3129
rect 14606 2940 14616 3124
rect 15216 2940 15226 3124
rect 14606 2935 15226 2940
rect 14612 2509 15216 2935
rect 15360 2889 15960 3311
rect 16412 3129 17016 3551
rect 17150 3500 17770 3505
rect 17150 3316 17160 3500
rect 17760 3316 17770 3500
rect 17150 3311 17770 3316
rect 16406 3124 17026 3129
rect 16406 2940 16416 3124
rect 17016 2940 17026 3124
rect 16406 2935 17026 2940
rect 15350 2884 15970 2889
rect 15350 2700 15360 2884
rect 15960 2700 15970 2884
rect 15350 2695 15970 2700
rect 14606 2504 15226 2509
rect 14606 2320 14616 2504
rect 15216 2320 15226 2504
rect 14606 2315 15226 2320
rect 14612 1893 15216 2315
rect 15360 2269 15960 2695
rect 16412 2509 17016 2935
rect 17160 2889 17760 3311
rect 18212 3129 18816 3551
rect 18950 3500 19570 3505
rect 18950 3316 18960 3500
rect 19560 3316 19570 3500
rect 18950 3311 19570 3316
rect 18206 3124 18826 3129
rect 18206 2940 18216 3124
rect 18816 2940 18826 3124
rect 18206 2935 18826 2940
rect 17150 2884 17770 2889
rect 17150 2700 17160 2884
rect 17760 2700 17770 2884
rect 17150 2695 17770 2700
rect 16406 2504 17026 2509
rect 16406 2320 16416 2504
rect 17016 2320 17026 2504
rect 16406 2315 17026 2320
rect 15350 2264 15970 2269
rect 15350 2080 15360 2264
rect 15960 2080 15970 2264
rect 15350 2075 15970 2080
rect 14606 1888 15226 1893
rect 14606 1704 14616 1888
rect 15216 1704 15226 1888
rect 14606 1699 15226 1704
rect 14612 1273 15216 1699
rect 15360 1653 15960 2075
rect 16412 1893 17016 2315
rect 17160 2269 17760 2695
rect 18212 2509 18816 2935
rect 18960 2889 19560 3311
rect 20012 3129 20616 3551
rect 20750 3500 21370 3505
rect 20750 3316 20760 3500
rect 21360 3316 21370 3500
rect 20750 3311 21370 3316
rect 20006 3124 20626 3129
rect 20006 2940 20016 3124
rect 20616 2940 20626 3124
rect 20006 2935 20626 2940
rect 18950 2884 19570 2889
rect 18950 2700 18960 2884
rect 19560 2700 19570 2884
rect 18950 2695 19570 2700
rect 18206 2504 18826 2509
rect 18206 2320 18216 2504
rect 18816 2320 18826 2504
rect 18206 2315 18826 2320
rect 17150 2264 17770 2269
rect 17150 2080 17160 2264
rect 17760 2080 17770 2264
rect 17150 2075 17770 2080
rect 16406 1888 17026 1893
rect 16406 1704 16416 1888
rect 17016 1704 17026 1888
rect 16406 1699 17026 1704
rect 15350 1648 15970 1653
rect 15350 1464 15360 1648
rect 15960 1464 15970 1648
rect 15350 1459 15970 1464
rect 14606 1268 15226 1273
rect 14606 1084 14616 1268
rect 15216 1084 15226 1268
rect 14606 1079 15226 1084
rect 14612 657 15216 1079
rect 15360 1033 15960 1459
rect 16412 1273 17016 1699
rect 17160 1653 17760 2075
rect 18212 1893 18816 2315
rect 18960 2269 19560 2695
rect 20012 2509 20616 2935
rect 20760 2889 21360 3311
rect 20750 2884 21370 2889
rect 20750 2700 20760 2884
rect 21360 2700 21370 2884
rect 20750 2695 21370 2700
rect 20006 2504 20626 2509
rect 20006 2320 20016 2504
rect 20616 2320 20626 2504
rect 20006 2315 20626 2320
rect 18950 2264 19570 2269
rect 18950 2080 18960 2264
rect 19560 2080 19570 2264
rect 18950 2075 19570 2080
rect 18206 1888 18826 1893
rect 18206 1704 18216 1888
rect 18816 1704 18826 1888
rect 18206 1699 18826 1704
rect 17150 1648 17770 1653
rect 17150 1464 17160 1648
rect 17760 1464 17770 1648
rect 17150 1459 17770 1464
rect 16406 1268 17026 1273
rect 16406 1084 16416 1268
rect 17016 1084 17026 1268
rect 16406 1079 17026 1084
rect 15350 1028 15970 1033
rect 15350 844 15360 1028
rect 15960 844 15970 1028
rect 15350 839 15970 844
rect 15360 680 15960 839
rect 14606 652 15226 657
rect 14606 468 14616 652
rect 15216 468 15226 652
rect 14606 463 15226 468
rect 14612 444 15216 463
rect 15360 417 15376 680
rect 15350 412 15376 417
rect 15948 417 15960 680
rect 16412 657 17016 1079
rect 17160 1033 17760 1459
rect 18212 1273 18816 1699
rect 18960 1653 19560 2075
rect 20012 1893 20616 2315
rect 20760 2269 21360 2695
rect 20750 2264 21370 2269
rect 20750 2080 20760 2264
rect 21360 2080 21370 2264
rect 20750 2075 21370 2080
rect 20006 1888 20626 1893
rect 20006 1704 20016 1888
rect 20616 1704 20626 1888
rect 20006 1699 20626 1704
rect 18950 1648 19570 1653
rect 18950 1464 18960 1648
rect 19560 1464 19570 1648
rect 18950 1459 19570 1464
rect 18206 1268 18826 1273
rect 18206 1084 18216 1268
rect 18816 1084 18826 1268
rect 18206 1079 18826 1084
rect 17150 1028 17770 1033
rect 17150 844 17160 1028
rect 17760 844 17770 1028
rect 17150 839 17770 844
rect 17160 680 17760 839
rect 16406 652 17026 657
rect 16406 468 16416 652
rect 17016 468 17026 652
rect 16406 463 17026 468
rect 16412 444 17016 463
rect 17160 417 17176 680
rect 15948 412 15970 417
rect 15350 228 15360 412
rect 15960 228 15970 412
rect 17150 412 17176 417
rect 17748 417 17760 680
rect 18212 657 18816 1079
rect 18960 1033 19560 1459
rect 20012 1273 20616 1699
rect 20760 1653 21360 2075
rect 20750 1648 21370 1653
rect 20750 1464 20760 1648
rect 21360 1464 21370 1648
rect 20750 1459 21370 1464
rect 20006 1268 20626 1273
rect 20006 1084 20016 1268
rect 20616 1084 20626 1268
rect 20006 1079 20626 1084
rect 18950 1028 19570 1033
rect 18950 844 18960 1028
rect 19560 844 19570 1028
rect 18950 839 19570 844
rect 18960 676 19560 839
rect 18206 652 18826 657
rect 18206 468 18216 652
rect 18816 468 18826 652
rect 18206 463 18826 468
rect 18212 444 18816 463
rect 18960 417 18972 676
rect 17748 412 17770 417
rect 15350 223 15970 228
rect 16086 268 16286 273
rect 11000 48 14372 76
rect 16086 68 16096 268
rect 16276 68 16286 268
rect 17150 228 17160 412
rect 17760 228 17770 412
rect 18950 412 18972 417
rect 19544 417 19560 676
rect 20012 657 20616 1079
rect 20760 1033 21360 1459
rect 20750 1028 21370 1033
rect 20750 844 20760 1028
rect 21360 844 21370 1028
rect 20750 839 21370 844
rect 20760 676 21360 839
rect 20006 652 20626 657
rect 20006 468 20016 652
rect 20616 468 20626 652
rect 20006 463 20626 468
rect 20012 444 20616 463
rect 20760 417 20772 676
rect 19544 412 19570 417
rect 17150 223 17770 228
rect 16086 63 16286 68
rect 17902 64 17912 276
rect 18092 64 18102 276
rect 18950 228 18960 412
rect 19560 228 19570 412
rect 20750 412 20772 417
rect 21344 417 21360 676
rect 21344 412 21370 417
rect 18950 223 19570 228
rect 19678 276 19878 281
rect 19678 64 19688 276
rect 19868 64 19878 276
rect 20750 228 20760 412
rect 21360 228 21370 412
rect 20750 223 21370 228
rect 19678 59 19878 64
rect 21580 56 24868 3740
rect 24932 56 24952 4080
rect 21580 28 24952 56
rect -2778 -382 -1950 -377
rect -2778 -1188 -2768 -382
rect -1960 -1188 -1950 -382
rect -2778 -1193 -1950 -1188
rect 11622 -382 12450 -377
rect 11622 -1188 11632 -382
rect 12440 -1188 12450 -382
rect 11622 -1193 12450 -1188
<< via3 >>
rect 24148 23084 24212 27108
rect 15900 21740 16300 22180
rect 7356 17960 7888 18220
rect 7356 17784 7888 17960
rect 9076 17960 9608 18200
rect 15580 18420 15980 18860
rect 16220 18420 16620 18860
rect 24148 18244 24212 22268
rect 8040 17616 8220 17776
rect 9076 17776 9608 17960
rect 9076 17764 9608 17776
rect 10764 17940 11300 18132
rect 10764 17716 11292 17940
rect 11292 17716 11300 17940
rect 10764 17592 11300 17716
rect 18300 18156 18900 18180
rect 18300 18056 18480 18156
rect 18480 18056 18680 18156
rect 18680 18056 18900 18156
rect 18300 17720 18900 18056
rect -2556 10096 1468 10160
rect -3872 4636 -3808 8660
rect 11844 10096 15868 10160
rect 5120 9160 6060 9180
rect 5120 8740 6060 9160
rect -3172 4420 -3028 4532
rect 8772 5968 9616 6020
rect 8772 5768 9616 5968
rect 8772 5348 9616 5768
rect 8772 5160 9616 5348
rect -8500 348 -8360 508
rect -3872 316 -3808 4340
rect -9316 4 -8716 284
rect -112 76 -48 4100
rect 23172 5968 24016 6020
rect 23172 5768 24016 5968
rect 23172 5348 24016 5768
rect 23172 5160 24016 5348
rect 976 412 1548 680
rect 976 240 1548 412
rect 2776 412 3348 680
rect 1696 68 1876 268
rect 2776 240 3348 412
rect 4572 412 5144 676
rect 3512 64 3692 276
rect 4572 236 5144 412
rect 6372 412 6944 676
rect 5288 64 5468 276
rect 6372 236 6944 412
rect 10468 56 10532 4080
rect 14288 76 14352 4100
rect 15376 412 15948 680
rect 15376 240 15948 412
rect 17176 412 17748 680
rect 16096 68 16276 268
rect 17176 240 17748 412
rect 18972 412 19544 676
rect 17912 64 18092 276
rect 18972 236 19544 412
rect 20772 412 21344 676
rect 19688 64 19868 276
rect 20772 236 21344 412
rect 24868 56 24932 4080
rect -2768 -1188 -1960 -382
rect 11632 -1188 12440 -382
<< mimcap >>
rect 19900 27056 23900 27096
rect 19900 23136 19940 27056
rect 23860 23136 23900 27056
rect 19900 23096 23900 23136
rect 19900 22216 23900 22256
rect 19900 18296 19940 22216
rect 23860 18296 23900 22216
rect 19900 18256 23900 18296
rect -2544 9808 1456 9848
rect -8120 8608 -4120 8648
rect -8120 4688 -8080 8608
rect -4160 4688 -4120 8608
rect -2544 5888 -2504 9808
rect 1416 5888 1456 9808
rect -2544 5848 1456 5888
rect 11856 9808 15856 9848
rect 11856 5888 11896 9808
rect 15816 5888 15856 9808
rect 11856 5848 15856 5888
rect -8120 4648 -4120 4688
rect -8120 4288 -4120 4328
rect -8120 368 -8080 4288
rect -4160 368 -4120 4288
rect -8120 328 -4120 368
rect -3360 4048 -360 4088
rect -3360 128 -3320 4048
rect -400 128 -360 4048
rect -3360 88 -360 128
rect 7220 4028 10220 4068
rect 7220 108 7260 4028
rect 10180 108 10220 4028
rect 7220 68 10220 108
rect 11040 4048 14040 4088
rect 11040 128 11080 4048
rect 14000 128 14040 4048
rect 11040 88 14040 128
rect 21620 4028 24620 4068
rect 21620 108 21660 4028
rect 24580 108 24620 4028
rect 21620 68 24620 108
<< mimcapcontact >>
rect 19940 23136 23860 27056
rect 19940 18296 23860 22216
rect -8080 4688 -4160 8608
rect -2504 5888 1416 9808
rect 11896 5888 15816 9808
rect -8080 368 -4160 4288
rect -3320 128 -400 4048
rect 7260 108 10180 4028
rect 11080 128 14000 4048
rect 21660 108 24580 4028
<< metal4 >>
rect 24132 27108 24228 27124
rect 19939 27056 23861 27057
rect 19939 23136 19940 27056
rect 23860 23136 23861 27056
rect 19939 23135 23861 23136
rect 19940 22217 20160 23135
rect 24132 23084 24148 27108
rect 24212 23084 24228 27108
rect 24132 23068 24228 23084
rect 24132 22268 24228 22284
rect 19939 22216 23861 22217
rect 15899 22180 16301 22181
rect 15899 21740 15900 22180
rect 16300 21740 16301 22180
rect 15899 21739 16301 21740
rect 15900 20520 16300 21739
rect 15580 18861 15980 20000
rect 16220 18861 16620 20000
rect 15579 18860 15981 18861
rect 15579 18420 15580 18860
rect 15980 18420 15981 18860
rect 15579 18419 15981 18420
rect 16219 18860 16621 18861
rect 16219 18420 16220 18860
rect 16620 18420 16621 18860
rect 16219 18419 16621 18420
rect 19939 18296 19940 22216
rect 23860 18296 23861 22216
rect 19939 18295 23861 18296
rect 7344 18220 7896 18236
rect 7344 17784 7356 18220
rect 7888 17836 7896 18220
rect 9064 18200 9616 18212
rect 7888 17784 8260 17836
rect 7344 17776 8260 17784
rect 7344 17616 8040 17776
rect 8220 17616 8260 17776
rect 7344 17536 8260 17616
rect 9064 17764 9076 18200
rect 9608 17764 9616 18200
rect 18299 18180 18901 18181
rect 9064 17536 9616 17764
rect 10756 18132 11308 18144
rect 10756 17592 10764 18132
rect 11300 17592 11308 18132
rect 18299 17720 18300 18180
rect 18900 17720 18901 18180
rect 18299 17719 18901 17720
rect 10756 17536 11308 17592
rect 6652 17480 11508 17536
rect 18300 17480 18900 17719
rect 19992 17480 21096 18295
rect 24132 18244 24148 22268
rect 24212 18244 24228 22268
rect 24132 18228 24228 18244
rect 6652 16920 28600 17480
rect 6660 15540 28600 16920
rect -2572 10160 1484 10176
rect -2572 10096 -2556 10160
rect 1468 10096 1484 10160
rect -2572 10080 1484 10096
rect 11828 10160 15884 10176
rect 11828 10096 11844 10160
rect 15868 10096 15884 10160
rect 11828 10080 15884 10096
rect -2505 9808 1417 9809
rect -3888 8660 -3792 8676
rect -8081 8608 -4159 8609
rect -8081 4688 -8080 8608
rect -4160 4688 -4159 8608
rect -8081 4687 -4159 4688
rect -8080 4289 -7620 4687
rect -3888 4636 -3872 8660
rect -3808 4636 -3792 8660
rect -2505 5888 -2504 9808
rect 1416 5888 1417 9808
rect 11895 9808 15817 9809
rect 5120 9181 10640 9460
rect 5119 9180 10640 9181
rect 5119 8740 5120 9180
rect 6060 8740 10640 9180
rect 5119 8739 6061 8740
rect -2505 5887 1417 5888
rect 8760 6020 9636 6036
rect -3888 4620 -3792 4636
rect -3192 4532 -3008 4568
rect -3192 4420 -3172 4532
rect -3028 4420 -3008 4532
rect -3192 4368 -3008 4420
rect -3884 4356 -3008 4368
rect -3888 4340 -3008 4356
rect -8081 4288 -4159 4289
rect -8520 508 -8340 540
rect -8520 348 -8500 508
rect -8360 348 -8340 508
rect -8081 368 -8080 4288
rect -4160 368 -4159 4288
rect -8081 367 -4159 368
rect -9317 284 -8715 285
rect -8520 284 -8340 348
rect -8080 284 -7620 367
rect -3888 316 -3872 4340
rect -3808 4272 -3008 4340
rect -3808 316 -3792 4272
rect -2104 4049 -432 5887
rect 8760 5160 8772 6020
rect 9616 5160 9636 6020
rect 11895 5888 11896 9808
rect 15816 5888 15817 9808
rect 11895 5887 15817 5888
rect 23160 6020 24036 6036
rect -128 4100 -32 4116
rect -3888 300 -3792 316
rect -3321 4048 -399 4049
rect -9317 280 -9316 284
rect -9320 4 -9316 280
rect -8716 4 -7620 284
rect -3321 128 -3320 4048
rect -400 128 -399 4048
rect -3321 127 -399 128
rect -9320 -80 -7620 4
rect -2104 -80 -432 127
rect -128 76 -112 4100
rect -48 76 -32 4100
rect 8760 4029 9636 5160
rect 10452 4080 10548 4096
rect 7259 4028 10181 4029
rect -128 60 -32 76
rect 960 680 1560 688
rect 960 240 976 680
rect 1548 328 1560 680
rect 2760 680 3360 688
rect 1548 268 1936 328
rect 1548 240 1696 268
rect 960 68 1696 240
rect 1876 68 1936 268
rect 960 -80 1936 68
rect 2760 240 2776 680
rect 3348 324 3360 680
rect 4560 676 5160 688
rect 3348 276 3712 324
rect 3348 240 3512 276
rect 2760 64 3512 240
rect 3692 64 3712 276
rect 2760 -80 3712 64
rect 4560 236 4572 676
rect 5144 352 5160 676
rect 6360 676 6960 684
rect 5144 276 5496 352
rect 5144 236 5288 276
rect 4560 64 5288 236
rect 5468 64 5496 276
rect 4560 -80 5496 64
rect 6360 236 6372 676
rect 6944 236 6960 676
rect 6360 -80 6960 236
rect 7259 108 7260 4028
rect 10180 108 10181 4028
rect 7259 107 10181 108
rect 7716 -80 9092 107
rect 10452 56 10468 4080
rect 10532 56 10548 4080
rect 12296 4049 13968 5887
rect 23160 5160 23172 6020
rect 24016 5160 24036 6020
rect 14272 4100 14368 4116
rect 11079 4048 14001 4049
rect 11079 128 11080 4048
rect 14000 128 14001 4048
rect 11079 127 14001 128
rect 10452 40 10548 56
rect 12296 -80 13968 127
rect 14272 76 14288 4100
rect 14352 76 14368 4100
rect 23160 4029 24036 5160
rect 24852 4080 24948 4096
rect 21659 4028 24581 4029
rect 14272 60 14368 76
rect 15360 680 15960 688
rect 15360 240 15376 680
rect 15948 328 15960 680
rect 17160 680 17760 688
rect 15948 268 16336 328
rect 15948 240 16096 268
rect 15360 68 16096 240
rect 16276 68 16336 268
rect 15360 -80 16336 68
rect 17160 240 17176 680
rect 17748 324 17760 680
rect 18960 676 19560 688
rect 17748 276 18112 324
rect 17748 240 17912 276
rect 17160 64 17912 240
rect 18092 64 18112 276
rect 17160 -80 18112 64
rect 18960 236 18972 676
rect 19544 352 19560 676
rect 20760 676 21360 684
rect 19544 276 19896 352
rect 19544 236 19688 276
rect 18960 64 19688 236
rect 19868 64 19896 276
rect 18960 -80 19896 64
rect 20760 236 20772 676
rect 21344 236 21360 676
rect 20760 -80 21360 236
rect 21659 108 21660 4028
rect 24580 108 24581 4028
rect 21659 107 24581 108
rect 22116 -80 23492 107
rect 24852 56 24868 4080
rect 24932 56 24948 4080
rect 24852 40 24948 56
rect 26000 -80 28600 15540
rect -10640 -382 28600 -80
rect -10640 -1188 -2768 -382
rect -1960 -1188 11632 -382
rect 12440 -1188 28600 -382
rect -10640 -4080 28600 -1188
<< res1p41 >>
rect 18324 23852 18610 24656
rect 2600 9884 2886 10688
rect 2978 9884 3264 10688
rect 3356 9884 3642 10688
rect 3734 9884 4020 10688
rect 4112 9884 4398 10688
rect 4490 9884 4776 10688
rect 17000 9884 17286 10688
rect 17378 9884 17664 10688
rect 17756 9884 18042 10688
rect 18134 9884 18420 10688
rect 18512 9884 18798 10688
rect 18890 9884 19176 10688
<< labels >>
rlabel metal3 -10000 12200 -8800 13600 1 VP
port 1 n
rlabel metal2 -10000 8800 -9600 9400 1 I_Bias1
port 6 n
rlabel metal4 -10400 -2800 -9600 -1400 1 VN
port 7 n
rlabel metal2 10600 6400 11200 7400 1 Input_ref
port 4 n
rlabel metal2 -3020 6340 -2520 6830 1 Input
port 5 n
rlabel metal1 9884 5220 10104 5448 1 VM9G
rlabel metal2 -3220 9220 -2700 9740 1 Out_2
port 8 n
rlabel metal4 15940 20560 16260 21000 1 Filter_in
port 10 n
rlabel metal2 24960 21180 25560 21460 1 Filter_out
port 12 n
rlabel metal4 16260 19520 16580 19960 1 Out_ref
port 13 n
rlabel metal3 -1454 10898 -1084 11238 1 tia_core_1.VP
rlabel metal2 5606 6328 6076 6738 1 tia_core_1.Input
rlabel metal4 -1714 -1092 -1374 -522 1 tia_core_1.VN
rlabel metal1 -338 5428 -46 5900 1 tia_core_1.V_Bias1
rlabel metal3 7108 4336 7332 4620 1 tia_core_1.V_Bias2
rlabel metal3 12946 10898 13316 11238 1 tia_core_0.VP
rlabel metal2 20006 6328 20476 6738 1 tia_core_0.Input
rlabel metal4 12686 -1092 13026 -522 1 tia_core_0.VN
rlabel metal1 14062 5428 14354 5900 1 tia_core_0.V_Bias1
rlabel metal3 21508 4336 21732 4620 1 tia_core_0.V_Bias2
rlabel metal2 -9950 8458 -9710 8598 1 curr_filter_0.I_Bias1
rlabel metal3 -8150 4458 -8100 4558 1 curr_filter_0.Out
rlabel metal4 -8580 58 -8380 178 1 curr_filter_0.Vn
<< end >>
