magic
tech sky130A
magscale 1 2
timestamp 1683736937
<< pwell >>
rect -1063 -1482 1063 1482
<< psubdiff >>
rect -1027 1412 -931 1446
rect 931 1412 1027 1446
rect -1027 1350 -993 1412
rect 993 1350 1027 1412
rect -1027 -1412 -993 -1350
rect 993 -1412 1027 -1350
rect -1027 -1446 -931 -1412
rect 931 -1446 1027 -1412
<< psubdiffcont >>
rect -931 1412 931 1446
rect -1027 -1350 -993 1350
rect 993 -1350 1027 1350
rect -931 -1446 931 -1412
<< xpolycontact >>
rect -897 884 -615 1316
rect -897 52 -615 484
rect -519 884 -237 1316
rect -519 52 -237 484
rect -141 884 141 1316
rect -141 52 141 484
rect 237 884 519 1316
rect 237 52 519 484
rect 615 884 897 1316
rect 615 52 897 484
rect -897 -484 -615 -52
rect -897 -1316 -615 -884
rect -519 -484 -237 -52
rect -519 -1316 -237 -884
rect -141 -484 141 -52
rect -141 -1316 141 -884
rect 237 -484 519 -52
rect 237 -1316 519 -884
rect 615 -484 897 -52
rect 615 -1316 897 -884
<< xpolyres >>
rect -897 484 -615 884
rect -519 484 -237 884
rect -141 484 141 884
rect 237 484 519 884
rect 615 484 897 884
rect -897 -884 -615 -484
rect -519 -884 -237 -484
rect -141 -884 141 -484
rect 237 -884 519 -484
rect 615 -884 897 -484
<< locali >>
rect -1027 1412 -931 1446
rect 931 1412 1027 1446
rect -1027 1350 -993 1412
rect 993 1350 1027 1412
rect -1027 -1412 -993 -1350
rect 993 -1412 1027 -1350
rect -1027 -1446 -931 -1412
rect 931 -1446 1027 -1412
<< viali >>
rect -881 901 -631 1298
rect -503 901 -253 1298
rect -125 901 125 1298
rect 253 901 503 1298
rect 631 901 881 1298
rect -881 70 -631 467
rect -503 70 -253 467
rect -125 70 125 467
rect 253 70 503 467
rect 631 70 881 467
rect -881 -467 -631 -70
rect -503 -467 -253 -70
rect -125 -467 125 -70
rect 253 -467 503 -70
rect 631 -467 881 -70
rect -881 -1298 -631 -901
rect -503 -1298 -253 -901
rect -125 -1298 125 -901
rect 253 -1298 503 -901
rect 631 -1298 881 -901
<< metal1 >>
rect -887 1298 -625 1310
rect -887 901 -881 1298
rect -631 901 -625 1298
rect -887 889 -625 901
rect -509 1298 -247 1310
rect -509 901 -503 1298
rect -253 901 -247 1298
rect -509 889 -247 901
rect -131 1298 131 1310
rect -131 901 -125 1298
rect 125 901 131 1298
rect -131 889 131 901
rect 247 1298 509 1310
rect 247 901 253 1298
rect 503 901 509 1298
rect 247 889 509 901
rect 625 1298 887 1310
rect 625 901 631 1298
rect 881 901 887 1298
rect 625 889 887 901
rect -887 467 -625 479
rect -887 70 -881 467
rect -631 70 -625 467
rect -887 58 -625 70
rect -509 467 -247 479
rect -509 70 -503 467
rect -253 70 -247 467
rect -509 58 -247 70
rect -131 467 131 479
rect -131 70 -125 467
rect 125 70 131 467
rect -131 58 131 70
rect 247 467 509 479
rect 247 70 253 467
rect 503 70 509 467
rect 247 58 509 70
rect 625 467 887 479
rect 625 70 631 467
rect 881 70 887 467
rect 625 58 887 70
rect -887 -70 -625 -58
rect -887 -467 -881 -70
rect -631 -467 -625 -70
rect -887 -479 -625 -467
rect -509 -70 -247 -58
rect -509 -467 -503 -70
rect -253 -467 -247 -70
rect -509 -479 -247 -467
rect -131 -70 131 -58
rect -131 -467 -125 -70
rect 125 -467 131 -70
rect -131 -479 131 -467
rect 247 -70 509 -58
rect 247 -467 253 -70
rect 503 -467 509 -70
rect 247 -479 509 -467
rect 625 -70 887 -58
rect 625 -467 631 -70
rect 881 -467 887 -70
rect 625 -479 887 -467
rect -887 -901 -625 -889
rect -887 -1298 -881 -901
rect -631 -1298 -625 -901
rect -887 -1310 -625 -1298
rect -509 -901 -247 -889
rect -509 -1298 -503 -901
rect -253 -1298 -247 -901
rect -509 -1310 -247 -1298
rect -131 -901 131 -889
rect -131 -1298 -125 -901
rect 125 -1298 131 -901
rect -131 -1310 131 -1298
rect 247 -901 509 -889
rect 247 -1298 253 -901
rect 503 -1298 509 -901
rect 247 -1310 509 -1298
rect 625 -901 887 -889
rect 625 -1298 631 -901
rect 881 -1298 887 -901
rect 625 -1310 887 -1298
<< res1p41 >>
rect -899 482 -613 886
rect -521 482 -235 886
rect -143 482 143 886
rect 235 482 521 886
rect 613 482 899 886
rect -899 -886 -613 -482
rect -521 -886 -235 -482
rect -143 -886 143 -482
rect 235 -886 521 -482
rect 613 -886 899 -482
<< properties >>
string FIXED_BBOX -1010 -1429 1010 1429
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 2.0 m 2 nx 5 wmin 1.410 lmin 0.50 rho 2000 val 3.103k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
