magic
tech sky130A
magscale 1 2
timestamp 1689780728
<< error_p >>
rect 36178 1091213 36180 1091297
rect 36262 1091172 36264 1091213
rect 121820 1091172 121822 1091297
rect 136620 1075313 136635 1075328
rect 136540 1075233 136555 1075248
rect 21445 1073352 21460 1073367
rect 21365 1073272 21380 1073287
rect 133187 1068693 133192 1068699
rect 136620 975313 136635 975328
rect 136540 975233 136555 975248
rect 21445 973352 21460 973367
rect 21365 973272 21380 973287
rect 133187 968693 133192 968699
rect 136620 875313 136635 875328
rect 136540 875233 136555 875248
rect 21445 873352 21460 873367
rect 21365 873272 21380 873287
rect 133187 868693 133192 868699
rect 136620 775313 136635 775328
rect 136540 775233 136555 775248
rect 21445 773352 21460 773367
rect 21365 773272 21380 773287
rect 133187 768693 133192 768699
rect 136620 675313 136635 675328
rect 136540 675233 136555 675248
rect 21445 673352 21460 673367
rect 21365 673272 21380 673287
rect 133187 668693 133192 668699
rect 136620 575313 136635 575328
rect 136540 575233 136555 575248
rect 21445 573352 21460 573367
rect 21365 573272 21380 573287
rect 133187 568693 133192 568699
rect 136620 475313 136635 475328
rect 136540 475233 136555 475248
rect 21445 473352 21460 473367
rect 21365 473272 21380 473287
rect 133187 468693 133192 468699
rect 136620 375313 136635 375328
rect 136540 375233 136555 375248
rect 21445 373352 21460 373367
rect 21365 373272 21380 373287
rect 133187 368693 133192 368699
rect 136620 275313 136635 275328
rect 136540 275233 136555 275248
rect 21445 273352 21460 273367
rect 21365 273272 21380 273287
rect 133187 268693 133192 268699
rect 36262 172387 36264 172512
rect 121736 172428 121738 172512
rect 121820 172387 121822 172428
rect 61856 171038 61912 171094
rect 63029 149964 63085 149988
use core3  core3_0
timestamp 1689779843
transform 1 0 6220 0 1 1038962
box 32860 -57400 112380 42940
use core3  core3_1
timestamp 1689779843
transform 1 0 6220 0 1 839000
box 32860 -57400 112380 42940
use core3  core3_3
timestamp 1689779843
transform 1 0 6220 0 1 438800
box 32860 -57400 112380 42940
use core3  core3_4
timestamp 1689779843
transform 1 0 6220 0 1 338800
box 32860 -57400 112380 42940
use core3  core3_5
timestamp 1689779843
transform 1 0 6220 0 1 238800
box 32860 -57400 112380 42940
use core3  core3_6
timestamp 1689779843
transform 1 0 6220 0 1 539000
box 32860 -57400 112380 42940
use core3  core3_7
timestamp 1689779843
transform 1 0 6220 0 1 639000
box 32860 -57400 112380 42940
use core3  core3_8
timestamp 1689779843
transform 1 0 6220 0 1 738800
box 32860 -57400 112380 42940
use core3  core3_9
timestamp 1689779843
transform 1 0 6220 0 1 938800
box 32860 -57400 112380 42940
use frame_modBC  frame_modBC_0 ~/code/hibpm-sky130a-tapeout/mag/frame
timestamp 1689780728
transform 1 0 6000 0 1 1038800
box -6000 -897800 152000 83800
<< end >>
