magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< locali >>
rect 980 3500 1080 3580
rect 1740 3420 2160 3500
rect 3960 3400 4340 3500
rect 6140 3360 6520 3460
rect 8320 3380 8720 3480
rect 880 1400 980 1500
rect 2540 1400 2640 1500
rect 4680 1400 4780 1500
rect 6680 1400 6780 1500
rect 8840 1400 8940 1500
rect 40 -2320 200 -2120
rect 1760 -2320 1920 -2120
rect 3600 -4800 3780 -4580
rect 3280 -6140 3600 -5980
<< viali >>
rect 980 3580 1080 3680
rect 1580 -6140 1760 -5980
<< metal1 >>
rect 968 3680 1092 3686
rect 968 3580 980 3680
rect 1080 3580 1092 3680
rect 968 3574 1092 3580
rect 1668 1340 10472 1564
rect 1686 456 1696 680
rect 1868 456 1878 680
rect 800 -2360 2528 -2200
rect 3564 -3920 4292 -3912
rect 3564 -3988 3728 -3920
rect 3800 -3988 4292 -3920
rect 3564 -4000 4292 -3988
rect 3564 -4460 3660 -4000
rect 3782 -4208 3792 -4028
rect 3852 -4208 3862 -4028
rect 3974 -4208 3984 -4028
rect 4044 -4208 4054 -4028
rect 4166 -4208 4176 -4028
rect 4236 -4208 4246 -4028
rect 4358 -4208 4368 -4028
rect 4428 -4208 4438 -4028
rect 3690 -4432 3700 -4252
rect 3760 -4432 3770 -4252
rect 3878 -4432 3888 -4252
rect 3948 -4432 3958 -4252
rect 4070 -4432 4080 -4252
rect 4140 -4432 4150 -4252
rect 4262 -4432 4272 -4252
rect 4332 -4432 4342 -4252
rect 3564 -4540 4384 -4460
rect 3564 -4920 4584 -4832
rect 3564 -5384 3660 -4920
rect 3782 -5132 3792 -4952
rect 3852 -5132 3862 -4952
rect 3974 -5132 3984 -4952
rect 4044 -5132 4054 -4952
rect 4166 -5132 4176 -4952
rect 4236 -5132 4246 -4952
rect 4358 -5132 4368 -4952
rect 4428 -5132 4438 -4952
rect 4550 -5132 4560 -4952
rect 4620 -5132 4630 -4952
rect 3690 -5352 3700 -5172
rect 3760 -5352 3770 -5172
rect 3878 -5352 3888 -5172
rect 3948 -5352 3958 -5172
rect 4070 -5352 4080 -5172
rect 4140 -5352 4150 -5172
rect 4262 -5352 4272 -5172
rect 4332 -5352 4342 -5172
rect 4454 -5352 4464 -5172
rect 4524 -5352 4534 -5172
rect 4646 -5352 4656 -5172
rect 4716 -5352 4726 -5172
rect 3564 -5540 4680 -5384
rect 1568 -5980 1772 -5974
rect 1568 -6140 1580 -5980
rect 1760 -6140 1772 -5980
rect 3564 -6000 3660 -5540
rect 3782 -5748 3792 -5568
rect 3852 -5748 3862 -5568
rect 3974 -5748 3984 -5568
rect 4044 -5748 4054 -5568
rect 4166 -5748 4176 -5568
rect 4236 -5748 4246 -5568
rect 4358 -5748 4368 -5568
rect 4428 -5748 4438 -5568
rect 4550 -5748 4560 -5568
rect 4620 -5748 4630 -5568
rect 3690 -5972 3700 -5792
rect 3760 -5972 3770 -5792
rect 3878 -5972 3888 -5792
rect 3948 -5972 3958 -5792
rect 4070 -5972 4080 -5792
rect 4140 -5972 4150 -5792
rect 4262 -5972 4272 -5792
rect 4332 -5972 4342 -5792
rect 4454 -5972 4464 -5792
rect 4524 -5972 4534 -5792
rect 4646 -5972 4656 -5792
rect 4716 -5972 4726 -5792
rect 3564 -6104 4584 -6000
rect 1568 -6146 1772 -6140
<< via1 >>
rect 980 3580 1080 3680
rect 1696 456 1868 680
rect 3728 -3988 3800 -3920
rect 3792 -4208 3852 -4028
rect 3984 -4208 4044 -4028
rect 4176 -4208 4236 -4028
rect 4368 -4208 4428 -4028
rect 3700 -4432 3760 -4252
rect 3888 -4432 3948 -4252
rect 4080 -4432 4140 -4252
rect 4272 -4432 4332 -4252
rect 3792 -5132 3852 -4952
rect 3984 -5132 4044 -4952
rect 4176 -5132 4236 -4952
rect 4368 -5132 4428 -4952
rect 4560 -5132 4620 -4952
rect 3700 -5352 3760 -5172
rect 3888 -5352 3948 -5172
rect 4080 -5352 4140 -5172
rect 4272 -5352 4332 -5172
rect 4464 -5352 4524 -5172
rect 4656 -5352 4716 -5172
rect 1580 -6140 1760 -5980
rect 3792 -5748 3852 -5568
rect 3984 -5748 4044 -5568
rect 4176 -5748 4236 -5568
rect 4368 -5748 4428 -5568
rect 4560 -5748 4620 -5568
rect 3700 -5972 3760 -5792
rect 3888 -5972 3948 -5792
rect 4080 -5972 4140 -5792
rect 4272 -5972 4332 -5792
rect 4464 -5972 4524 -5792
rect 4656 -5972 4716 -5792
<< metal2 >>
rect 980 3680 1080 3690
rect 980 3570 1080 3580
rect 3640 1060 10300 1384
rect 1696 680 1868 690
rect 1696 446 1868 456
rect 228 -76 3216 -52
rect 228 -484 948 -76
rect 1776 -484 3216 -76
rect 228 -512 3216 -484
rect 1152 -2660 1924 -2468
rect 3792 -3888 4440 -3864
rect 3792 -3910 3816 -3888
rect 3728 -3920 3816 -3910
rect 3800 -3988 3816 -3920
rect 3728 -3998 3816 -3988
rect 3792 -4028 3816 -3998
rect 4416 -4028 4440 -3888
rect 3852 -4200 3984 -4176
rect 3792 -4218 3852 -4208
rect 4044 -4200 4176 -4176
rect 3984 -4218 4044 -4208
rect 4236 -4200 4368 -4176
rect 4176 -4218 4236 -4208
rect 4428 -4200 4440 -4028
rect 4368 -4218 4428 -4208
rect 3700 -4252 3760 -4242
rect 3580 -4278 3700 -4258
rect 3564 -4288 3700 -4278
rect 3888 -4252 3948 -4242
rect 3760 -4288 3888 -4258
rect 4080 -4252 4140 -4242
rect 3948 -4288 4080 -4258
rect 4272 -4252 4332 -4242
rect 4140 -4260 4164 -4258
rect 4140 -4288 4272 -4260
rect 4180 -4432 4272 -4288
rect 4180 -4472 4332 -4432
rect 3564 -4594 4180 -4584
rect 3792 -4870 4620 -4868
rect 3580 -4880 4620 -4870
rect 4164 -4952 4620 -4880
rect 4164 -5112 4176 -4952
rect 3580 -5122 3792 -5112
rect 3852 -5124 3984 -5112
rect 3792 -5142 3852 -5132
rect 4044 -5124 4176 -5112
rect 3984 -5142 4044 -5132
rect 4236 -5124 4368 -4952
rect 4176 -5142 4236 -5132
rect 4428 -5124 4560 -4952
rect 4368 -5142 4428 -5132
rect 4560 -5142 4620 -5132
rect 3700 -5172 3760 -5162
rect 3888 -5172 3948 -5162
rect 3760 -5352 3888 -5180
rect 4080 -5172 4140 -5162
rect 3948 -5352 4080 -5180
rect 4272 -5172 4332 -5162
rect 4140 -5352 4272 -5180
rect 4464 -5172 4524 -5162
rect 4332 -5196 4464 -5180
rect 4656 -5172 4716 -5162
rect 4524 -5196 4656 -5180
rect 4716 -5196 4836 -5186
rect 3700 -5420 4308 -5352
rect 3700 -5430 4836 -5420
rect 3700 -5436 4716 -5430
rect 3792 -5490 4620 -5484
rect 3580 -5500 4620 -5490
rect 4164 -5568 4620 -5500
rect 4164 -5724 4176 -5568
rect 3580 -5734 3792 -5724
rect 3852 -5740 3984 -5724
rect 3792 -5758 3852 -5748
rect 4044 -5740 4176 -5724
rect 3984 -5758 4044 -5748
rect 4236 -5740 4368 -5568
rect 4176 -5758 4236 -5748
rect 4428 -5740 4560 -5568
rect 4368 -5758 4428 -5748
rect 4560 -5758 4620 -5748
rect 3700 -5792 3760 -5782
rect 1580 -5980 1760 -5970
rect 3888 -5792 3948 -5782
rect 3760 -5972 3888 -5800
rect 4080 -5792 4140 -5782
rect 3948 -5972 4080 -5800
rect 4272 -5792 4332 -5782
rect 4140 -5972 4272 -5800
rect 4464 -5792 4524 -5782
rect 4332 -5816 4464 -5800
rect 4656 -5792 4716 -5782
rect 4524 -5816 4656 -5800
rect 4716 -5816 4832 -5806
rect 3700 -6040 4304 -5972
rect 3700 -6050 4832 -6040
rect 3700 -6056 4716 -6050
rect 1580 -6150 1760 -6140
<< via2 >>
rect 980 3580 1080 3680
rect 1696 456 1868 680
rect 948 -484 1776 -76
rect 3816 -4028 4416 -3888
rect 3816 -4176 3852 -4028
rect 3852 -4176 3984 -4028
rect 3984 -4176 4044 -4028
rect 4044 -4176 4176 -4028
rect 4176 -4176 4236 -4028
rect 4236 -4176 4368 -4028
rect 4368 -4176 4416 -4028
rect 3564 -4432 3700 -4288
rect 3700 -4432 3760 -4288
rect 3760 -4432 3888 -4288
rect 3888 -4432 3948 -4288
rect 3948 -4432 4080 -4288
rect 4080 -4432 4140 -4288
rect 4140 -4432 4180 -4288
rect 3564 -4584 4180 -4432
rect 3580 -4952 4164 -4880
rect 3580 -5112 3792 -4952
rect 3792 -5112 3852 -4952
rect 3852 -5112 3984 -4952
rect 3984 -5112 4044 -4952
rect 4044 -5112 4164 -4952
rect 4308 -5352 4332 -5196
rect 4332 -5352 4464 -5196
rect 4464 -5352 4524 -5196
rect 4524 -5352 4656 -5196
rect 4656 -5352 4716 -5196
rect 4716 -5352 4836 -5196
rect 4308 -5420 4836 -5352
rect 3580 -5568 4164 -5500
rect 3580 -5724 3792 -5568
rect 3792 -5724 3852 -5568
rect 3852 -5724 3984 -5568
rect 3984 -5724 4044 -5568
rect 4044 -5724 4164 -5568
rect 1580 -6140 1760 -5980
rect 4304 -5972 4332 -5816
rect 4332 -5972 4464 -5816
rect 4464 -5972 4524 -5816
rect 4524 -5972 4656 -5816
rect 4656 -5972 4716 -5816
rect 4716 -5972 4832 -5816
rect 4304 -6040 4832 -5972
<< metal3 >>
rect -8 3680 10576 4104
rect -8 3604 980 3680
rect 912 3580 980 3604
rect 1080 3604 10576 3680
rect 1080 3580 1796 3604
rect 912 3468 1796 3580
rect 3132 3472 4016 3604
rect 5312 3504 6196 3604
rect 7492 3520 8376 3604
rect 9692 3532 10576 3604
rect 1686 680 1878 685
rect 1686 456 1696 680
rect 1868 456 1878 680
rect 1686 451 1878 456
rect 932 -76 1796 408
rect 932 -380 948 -76
rect 938 -484 948 -380
rect 1776 -380 1796 -76
rect 3144 -168 10564 304
rect 1776 -484 1786 -380
rect 938 -489 1786 -484
rect 3808 -3883 4448 -168
rect 3806 -3888 4448 -3883
rect 3806 -4176 3816 -3888
rect 4416 -4176 4448 -3888
rect 3806 -4180 4448 -4176
rect 3806 -4181 4426 -4180
rect 3564 -4283 4180 -4272
rect 3554 -4288 4190 -4283
rect 3554 -4584 3564 -4288
rect 4180 -4584 4190 -4288
rect 3554 -4589 4190 -4584
rect 3564 -4880 4180 -4589
rect 3564 -5112 3580 -4880
rect 4164 -5112 4180 -4880
rect 3564 -5500 4180 -5112
rect 886 -5972 896 -5536
rect 1428 -5972 1438 -5536
rect 1570 -5980 1770 -5975
rect 1570 -6140 1580 -5980
rect 1760 -6140 1770 -5980
rect 2606 -5992 2616 -5556
rect 3148 -5992 3158 -5556
rect 3564 -5724 3580 -5500
rect 4164 -5724 4180 -5500
rect 3564 -5740 4180 -5724
rect 4288 -5196 4856 -5180
rect 4288 -5420 4308 -5196
rect 4836 -5420 4856 -5196
rect 4288 -5624 4856 -5420
rect 1570 -6145 1770 -6140
rect 4288 -6164 4304 -5624
rect 4840 -6164 4856 -5624
rect 4288 -6180 4856 -6164
<< via3 >>
rect 896 -5972 1428 -5536
rect 1580 -6140 1760 -5980
rect 2616 -5992 3148 -5556
rect 4304 -5816 4840 -5624
rect 4304 -6040 4832 -5816
rect 4832 -6040 4840 -5816
rect 4304 -6164 4840 -6040
<< metal4 >>
rect 884 -5536 1436 -5520
rect 884 -5972 896 -5536
rect 1428 -5920 1436 -5536
rect 2604 -5556 3156 -5544
rect 1428 -5972 1800 -5920
rect 884 -5980 1800 -5972
rect 884 -6140 1580 -5980
rect 1760 -6140 1800 -5980
rect 884 -6220 1800 -6140
rect 2604 -5992 2616 -5556
rect 3148 -5992 3156 -5556
rect 2604 -6220 3156 -5992
rect 4296 -5624 4848 -5612
rect 4296 -6164 4304 -5624
rect 4840 -6164 4848 -5624
rect 4296 -6220 4848 -6164
rect 192 -6836 5048 -6220
use curr_m  curr_m_0
timestamp 1686659968
transform 1 0 1720 0 1 -1780
box 0 -4400 1624 1656
use curr_m  curr_m_1
timestamp 1686659968
transform 1 0 0 0 1 -1780
box 0 -4400 1624 1656
use currm_p  currm_p_0
timestamp 1686659968
transform 1 0 7460 0 1 -220
box 1200 200 3224 3776
use currm_p  currm_p_1
timestamp 1686659968
transform 1 0 -1320 0 1 -220
box 1200 200 3224 3776
use currm_p  currm_p_2
timestamp 1686659968
transform 1 0 900 0 1 -220
box 1200 200 3224 3776
use currm_p  currm_p_3
timestamp 1686659968
transform 1 0 3080 0 1 -220
box 1200 200 3224 3776
use currm_p  currm_p_4
timestamp 1686659968
transform 1 0 5260 0 1 -220
box 1200 200 3224 3776
use sky130_fd_pr__nfet_01v8_lvt_9B2JGQ  sky130_fd_pr__nfet_01v8_lvt_9B2JGQ_0
timestamp 1686659968
transform 1 0 4063 0 1 -4230
box -503 -410 503 410
use sky130_fd_pr__nfet_01v8_lvt_9U3MKJ  sky130_fd_pr__nfet_01v8_lvt_9U3MKJ_0
timestamp 1686659968
transform 1 0 4207 0 1 -5461
box -647 -719 647 719
<< end >>
