magic
tech sky130A
magscale 1 2
timestamp 1689773955
<< metal1 >>
rect 74 3208 84 3636
rect 1500 3208 1510 3636
rect 74 2376 84 2808
rect 1504 2376 1514 2808
rect 78 1840 88 2268
rect 1504 1840 1514 2268
rect 74 1004 84 1440
rect 1504 1004 1514 1440
rect 336 660 1364 776
rect 286 448 296 628
rect 348 448 358 628
rect 478 448 488 628
rect 540 448 550 628
rect 670 448 680 628
rect 732 448 742 628
rect 862 448 872 628
rect 924 448 934 628
rect 1054 448 1064 628
rect 1116 448 1126 628
rect 1246 448 1256 628
rect 1308 448 1318 628
rect 190 232 200 412
rect 252 232 262 412
rect 382 232 392 412
rect 444 232 454 412
rect 574 232 584 412
rect 636 232 646 412
rect 766 232 776 412
rect 828 232 838 412
rect 958 232 968 412
rect 1020 232 1030 412
rect 1150 232 1160 412
rect 1212 232 1222 412
rect 1342 232 1352 412
rect 1404 232 1414 412
rect 244 84 1268 200
<< via1 >>
rect 84 3208 1500 3636
rect 84 2376 1504 2808
rect 88 1840 1504 2268
rect 84 1004 1504 1440
rect 296 448 348 628
rect 488 448 540 628
rect 680 448 732 628
rect 872 448 924 628
rect 1064 448 1116 628
rect 1256 448 1308 628
rect 200 232 252 412
rect 392 232 444 412
rect 584 232 636 412
rect 776 232 828 412
rect 968 232 1020 412
rect 1160 232 1212 412
rect 1352 232 1404 412
<< metal2 >>
rect 80 3644 1508 3654
rect 80 3198 1508 3208
rect 84 2808 1504 2818
rect 84 2368 464 2376
rect 1128 2368 1504 2376
rect 84 2366 1504 2368
rect 464 2358 1128 2366
rect 84 2278 368 2286
rect 1220 2278 1504 2286
rect 84 2276 1504 2278
rect 368 2268 1220 2276
rect 84 1830 1504 1840
rect 84 1440 1504 1450
rect 84 996 88 1004
rect 1500 996 1504 1004
rect 84 994 1504 996
rect 88 986 1500 994
rect 296 628 1308 986
rect 348 520 488 628
rect 348 464 388 520
rect 452 464 488 520
rect 296 438 348 448
rect 540 520 680 628
rect 540 464 580 520
rect 644 464 680 520
rect 488 438 540 448
rect 732 520 872 628
rect 732 464 772 520
rect 836 464 872 520
rect 680 438 732 448
rect 924 520 1064 628
rect 924 464 964 520
rect 1028 464 1064 520
rect 872 438 924 448
rect 1116 520 1256 628
rect 1116 464 1156 520
rect 1220 464 1256 520
rect 1064 438 1116 448
rect 1256 438 1308 448
rect 200 412 252 422
rect 392 412 444 422
rect 252 340 292 396
rect 356 340 392 396
rect 252 232 392 340
rect 584 412 636 422
rect 444 340 484 396
rect 548 340 584 396
rect 444 232 584 340
rect 776 412 828 422
rect 636 340 672 396
rect 736 340 776 396
rect 636 232 776 340
rect 968 412 1020 422
rect 828 340 868 396
rect 932 340 968 396
rect 828 232 968 340
rect 1160 412 1212 422
rect 1020 340 1060 396
rect 1124 340 1160 396
rect 1020 232 1160 340
rect 1352 412 1404 422
rect 1212 340 1252 396
rect 1316 340 1352 396
rect 1212 232 1352 340
rect 200 60 1404 232
<< via2 >>
rect 80 3636 1508 3644
rect 80 3208 84 3636
rect 84 3208 1500 3636
rect 1500 3208 1508 3636
rect 464 2376 1128 2808
rect 464 2368 1128 2376
rect 84 2268 368 2276
rect 1220 2268 1504 2276
rect 84 1840 88 2268
rect 88 1840 368 2268
rect 1220 1840 1504 2268
rect 88 1004 1500 1440
rect 88 996 1500 1004
<< metal3 >>
rect 70 3644 1518 3649
rect 70 3208 80 3644
rect 1508 3208 1518 3644
rect 70 3203 1518 3208
rect 84 2281 368 3203
rect 454 2808 1138 2813
rect 454 2368 464 2808
rect 1128 2368 1138 2808
rect 454 2363 1138 2368
rect 74 2276 378 2281
rect 74 1840 84 2276
rect 368 1840 378 2276
rect 74 1835 378 1840
rect 464 1445 748 2363
rect 840 1445 1124 2363
rect 1220 2281 1504 3203
rect 1210 2276 1514 2281
rect 1210 1840 1220 2276
rect 1504 1840 1514 2276
rect 1210 1835 1514 1840
rect 78 1440 1510 1445
rect 78 996 88 1440
rect 1500 996 1510 1440
rect 78 991 1510 996
use sky130_fd_pr__nfet_01v8_lvt_F8VELN  sky130_fd_pr__nfet_01v8_lvt_F8VELN_0
timestamp 1684830260
transform 1 0 803 0 1 430
box -743 -410 743 410
use sky130_fd_pr__res_xhigh_po_1p41_FUYU7G  sky130_fd_pr__res_xhigh_po_1p41_FUYU7G_0
timestamp 1689672086
transform 1 0 794 0 1 2322
box -874 -1482 874 1482
<< end >>
