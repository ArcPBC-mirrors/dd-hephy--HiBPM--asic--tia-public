magic
tech sky130A
timestamp 1699354420
<< via4 >>
rect 12341 18139 12619 18259
rect 12341 18019 12979 18139
rect 12341 17899 13219 18019
rect 12341 17779 13459 17899
rect 12341 17659 13699 17779
rect 12341 17539 13939 17659
rect 12341 17419 14179 17539
rect 12341 17141 14299 17419
rect 4061 16699 4339 16819
rect 3461 16219 3739 16339
rect 2981 15739 3139 15859
rect 2861 15341 3139 15739
rect 3341 14861 3739 16219
rect 3461 14741 3739 14861
rect 3941 14261 4339 16699
rect 4541 16579 4699 16699
rect 4061 14141 4339 14261
rect 4421 16339 4819 16579
rect 12341 16421 14179 17141
rect 4181 13459 4339 13579
rect 4061 13339 4339 13459
rect 3581 12739 3739 12859
rect 3461 12619 3739 12739
rect 3341 12341 3739 12619
rect 3461 12221 3739 12341
rect 3941 11981 4339 13339
rect 4061 11861 4339 11981
rect 4421 11621 4939 16339
rect 5141 15739 5299 15859
rect 4541 11501 4939 11621
rect 4661 11381 4939 11501
rect 5021 15499 5419 15739
rect 12341 15581 14059 16421
rect 5021 11261 5539 15499
rect 5141 11021 5539 11261
rect 5621 14899 5899 15019
rect 5621 10781 6019 14899
rect 12341 14861 13939 15581
rect 5741 10661 6019 10781
rect 5861 10541 6019 10661
rect 6221 14179 6379 14299
rect 6221 14059 6499 14179
rect 12341 14141 13819 14861
rect 15221 14779 15499 14899
rect 15221 14659 15859 14779
rect 15101 14539 16099 14659
rect 15101 14419 16459 14539
rect 15101 14299 16699 14419
rect 14981 14141 16699 14299
rect 6221 10301 6619 14059
rect 6341 10181 6619 10301
rect 6821 13339 6979 13459
rect 12341 13421 13699 14141
rect 14981 13939 16579 14141
rect 14861 13901 16579 13939
rect 14861 13661 16459 13901
rect 14861 13459 16339 13661
rect 14741 13421 16339 13459
rect 6821 13219 7099 13339
rect 4061 9979 4459 10099
rect 4061 9859 4699 9979
rect 3941 9739 4939 9859
rect 6821 9821 7219 13219
rect 11141 12619 11299 12739
rect 3941 9619 5179 9739
rect 6941 9701 7219 9821
rect 7421 12379 7699 12619
rect 10661 12499 11419 12619
rect 3821 9499 5419 9619
rect 3821 9379 5659 9499
rect 7421 9461 7819 12379
rect 10301 12139 11419 12499
rect 12341 12581 13579 13421
rect 14741 13219 16219 13421
rect 14621 13181 16219 13219
rect 14621 12941 16099 13181
rect 14621 12739 15979 12941
rect 14501 12701 15979 12739
rect 10301 11981 11539 12139
rect 3821 9259 5899 9379
rect 7541 9341 7819 9461
rect 8021 11779 8179 11899
rect 8021 11539 8299 11779
rect 10421 11621 11539 11981
rect 3701 9139 6139 9259
rect 3701 9019 6379 9139
rect 3581 8899 6619 9019
rect 8021 8981 8419 11539
rect 10541 11419 11539 11621
rect 12341 11741 13459 12581
rect 14501 12461 15859 12701
rect 14501 12379 15739 12461
rect 14381 12221 15739 12379
rect 14381 12019 15619 12221
rect 14261 11981 15619 12019
rect 14261 11741 15499 11981
rect 10541 11179 11659 11419
rect 10301 11059 11659 11179
rect 3581 8779 6859 8899
rect 8141 8861 8419 8981
rect 8621 10939 8779 11059
rect 10061 10939 11659 11059
rect 8621 10699 8899 10939
rect 3581 8741 7099 8779
rect 3701 8659 7099 8741
rect 3701 8621 7219 8659
rect 4061 8539 7219 8621
rect 4061 8501 7579 8539
rect 8621 8501 9019 10699
rect 9821 10661 11659 10939
rect 9941 10579 11659 10661
rect 12341 11021 13339 11741
rect 14261 11659 15379 11741
rect 14141 11501 15379 11659
rect 14141 11299 15259 11501
rect 14021 11261 15259 11299
rect 14021 11021 15139 11261
rect 9941 10421 11779 10579
rect 9101 10099 9379 10219
rect 10061 10181 11779 10421
rect 9101 9859 9499 10099
rect 10181 10061 11779 10181
rect 10301 9859 11779 10061
rect 12341 10301 13219 11021
rect 14021 10939 15019 11021
rect 13901 10781 15019 10939
rect 13901 10579 14899 10781
rect 13781 10541 14899 10579
rect 13781 10301 14779 10541
rect 4421 8419 7579 8501
rect 4421 8381 7699 8419
rect 4781 8299 7699 8381
rect 4781 8261 7939 8299
rect 9101 8261 9619 9859
rect 10301 9821 11899 9859
rect 10421 9581 11899 9821
rect 5141 8179 7939 8261
rect 5141 8141 8179 8179
rect 9221 8141 9619 8261
rect 9701 9379 9859 9499
rect 9701 9259 9979 9379
rect 10541 9341 11899 9581
rect 5501 8059 8179 8141
rect 5501 8021 8419 8059
rect 9341 8021 9499 8141
rect 5861 7939 8419 8021
rect 5861 7901 8659 7939
rect 6221 7819 8659 7901
rect 6221 7781 8899 7819
rect 9701 7781 10099 9259
rect 10661 9139 11899 9341
rect 12341 9581 13099 10301
rect 13781 10219 14659 10301
rect 13661 10061 14659 10219
rect 13661 9859 14539 10061
rect 13541 9821 14539 9859
rect 13541 9581 14419 9821
rect 10661 9101 12019 9139
rect 10781 8861 12019 9101
rect 6701 7699 8899 7781
rect 6701 7661 9139 7699
rect 9821 7661 10099 7781
rect 6941 7579 9139 7661
rect 6941 7541 9379 7579
rect 9941 7541 10099 7661
rect 10301 8419 10579 8659
rect 10901 8621 12019 8861
rect 7421 7459 9379 7541
rect 7421 7421 9619 7459
rect 7781 7339 9619 7421
rect 7781 7301 9859 7339
rect 10301 7301 10699 8419
rect 11021 8381 12019 8621
rect 11141 8299 12019 8381
rect 12341 8741 12979 9581
rect 13541 9499 14299 9581
rect 13421 9341 14299 9499
rect 13421 9101 14179 9341
rect 13421 9019 14059 9101
rect 13301 8861 14059 9019
rect 13301 8741 13939 8861
rect 11141 8141 12139 8299
rect 11261 7901 12139 8141
rect 8141 7219 9859 7301
rect 8141 7181 10099 7219
rect 10421 7181 10699 7301
rect 10901 7579 11179 7819
rect 11381 7781 12139 7901
rect 12341 8021 12859 8741
rect 13301 8659 13819 8741
rect 13181 8501 13819 8659
rect 13181 8419 13699 8501
rect 13061 8261 13699 8419
rect 13061 8059 13579 8261
rect 12941 8021 13579 8059
rect 12341 7781 12739 8021
rect 12941 7781 13459 8021
rect 11381 7661 11899 7781
rect 12941 7661 13339 7781
rect 10901 7421 11299 7579
rect 11501 7541 11659 7661
rect 10901 7301 11179 7421
rect 10901 7181 11059 7301
rect 8501 7099 10099 7181
rect 8501 7061 10339 7099
rect 8861 6979 10339 7061
rect 11981 6979 12739 7099
rect 8861 6941 10579 6979
rect 9221 6859 10579 6941
rect 11741 6859 12979 6979
rect 9221 6821 10699 6859
rect 9581 6701 10699 6821
rect 11621 6739 13219 6859
rect 9941 6581 10699 6701
rect 11501 6619 13339 6739
rect 10300 6460 10580 6581
rect 11381 6499 13339 6619
rect 11381 6379 13459 6499
rect 11261 6259 13459 6379
rect 1541 6139 13579 6259
rect 1421 5741 13579 6139
rect 1541 5621 13579 5741
rect 11261 5501 13459 5621
rect 10421 5299 10579 5419
rect 11381 5381 13459 5501
rect 10061 5179 10699 5299
rect 11381 5261 13339 5381
rect 9701 5059 10699 5179
rect 11501 5141 13339 5261
rect 9341 4939 10699 5059
rect 11621 5021 13219 5141
rect 8981 4901 10699 4939
rect 11741 4901 13099 5021
rect 8981 4819 10459 4901
rect 8621 4781 10459 4819
rect 8621 4699 10219 4781
rect 10660 4699 10940 4820
rect 11981 4781 12859 4901
rect 8261 4661 10219 4699
rect 8261 4579 9979 4661
rect 10541 4579 11059 4699
rect 7781 4541 9979 4579
rect 7781 4459 9739 4541
rect 10301 4459 11059 4579
rect 7421 4421 9739 4459
rect 10181 4421 11059 4459
rect 7421 4339 9499 4421
rect 10181 4339 10939 4421
rect 7061 4301 9499 4339
rect 10061 4301 10939 4339
rect 7061 4219 9259 4301
rect 10061 4219 10819 4301
rect 11141 4219 11539 4339
rect 6701 4181 9259 4219
rect 9821 4181 10819 4219
rect 6701 4099 9019 4181
rect 9821 4099 10699 4181
rect 11021 4099 11779 4219
rect 6341 4061 9019 4099
rect 9701 4061 10699 4099
rect 6341 3979 8779 4061
rect 9701 3979 10579 4061
rect 5981 3941 8779 3979
rect 9461 3941 10579 3979
rect 10901 3941 11899 4099
rect 12101 3979 12379 4099
rect 15701 3979 16699 5899
rect 18941 3979 19939 5899
rect 5981 3859 8539 3941
rect 9461 3859 10459 3941
rect 10901 3859 11779 3941
rect 5621 3821 8539 3859
rect 9341 3821 10459 3859
rect 5621 3739 8299 3821
rect 9341 3739 10339 3821
rect 10781 3739 11779 3859
rect 5261 3701 8299 3739
rect 9221 3701 10339 3739
rect 10661 3701 11779 3739
rect 5261 3619 8059 3701
rect 9221 3619 10219 3701
rect 10661 3619 11659 3701
rect 4901 3581 8059 3619
rect 8981 3581 10219 3619
rect 4901 3499 7819 3581
rect 8981 3499 10099 3581
rect 4421 3461 7819 3499
rect 8861 3461 10099 3499
rect 4421 3379 7579 3461
rect 8861 3379 9979 3461
rect 10541 3379 11659 3619
rect 11981 3379 12499 3979
rect 4181 3341 7579 3379
rect 8621 3341 9979 3379
rect 4181 3259 7339 3341
rect 8621 3259 9859 3341
rect 10421 3259 11659 3379
rect 3821 3221 7339 3259
rect 8501 3221 9859 3259
rect 10301 3221 11659 3259
rect 3821 3139 7099 3221
rect 8501 3139 9739 3221
rect 3701 3101 7099 3139
rect 8381 3101 9739 3139
rect 3701 2981 6859 3101
rect 8381 3019 9619 3101
rect 10301 3019 11539 3221
rect 8141 2981 9619 3019
rect 3821 2861 6619 2981
rect 8141 2899 9499 2981
rect 10181 2899 11539 3019
rect 8021 2861 9499 2899
rect 10061 2861 11539 2899
rect 3941 2741 6379 2861
rect 8021 2779 9379 2861
rect 10061 2779 11419 2861
rect 7901 2741 9379 2779
rect 4181 2621 6139 2741
rect 7901 2659 9259 2741
rect 7661 2621 9259 2659
rect 9941 2621 11419 2779
rect 11861 2659 12499 3379
rect 4301 2501 5899 2621
rect 7661 2539 9139 2621
rect 9941 2539 10699 2621
rect 7541 2501 9139 2539
rect 4421 2381 5659 2501
rect 7541 2419 9019 2501
rect 9821 2419 10699 2539
rect 10901 2501 11419 2621
rect 7301 2381 9019 2419
rect 9701 2381 10699 2419
rect 11141 2381 11299 2501
rect 4661 2261 5419 2381
rect 7301 2299 8899 2381
rect 9701 2299 10579 2381
rect 7181 2261 8899 2299
rect 4781 2141 5179 2261
rect 7181 2179 8779 2261
rect 7061 2141 8779 2179
rect 9581 2141 10579 2299
rect 7061 2059 8659 2141
rect 9581 2059 10459 2141
rect 6821 2021 8659 2059
rect 6821 1939 8539 2021
rect 9461 1939 10459 2059
rect 11741 1939 12499 2659
rect 6701 1901 8539 1939
rect 9341 1901 10459 1939
rect 6701 1819 8419 1901
rect 6581 1781 8419 1819
rect 6581 1699 8299 1781
rect 9341 1699 10339 1901
rect 6341 1661 8299 1699
rect 9221 1661 10339 1699
rect 6341 1541 8179 1661
rect 9221 1579 10219 1661
rect 6341 1421 8059 1541
rect 9101 1459 10219 1579
rect 8981 1421 10219 1459
rect 6581 1301 7939 1421
rect 6941 1181 7819 1301
rect 8981 1219 10099 1421
rect 8861 1181 10099 1219
rect 11621 1301 12499 1939
rect 15701 2981 19939 3979
rect 11621 1181 12379 1301
rect 7301 1061 7699 1181
rect 8861 1099 9979 1181
rect 8741 941 9979 1099
rect 11621 1061 11899 1181
rect 8741 821 9859 941
rect 15701 821 16699 2981
rect 18941 821 19939 2981
rect 20741 5779 23899 5899
rect 24701 5779 27139 5899
rect 20741 5021 24019 5779
rect 24701 5659 27379 5779
rect 24701 5539 27619 5659
rect 24701 5419 27739 5539
rect 24701 5299 27859 5419
rect 24701 5059 27979 5299
rect 20741 4901 23779 5021
rect 24701 4901 28099 5059
rect 20741 3979 21739 4901
rect 20741 3859 23419 3979
rect 20741 2981 23659 3859
rect 24701 3619 25699 4901
rect 26861 4819 28099 4901
rect 26861 4781 28219 4819
rect 26981 4661 28219 4781
rect 27101 4421 28219 4661
rect 27221 4099 28219 4421
rect 27101 3859 28219 4099
rect 26981 3821 28219 3859
rect 29021 3979 30019 5899
rect 32261 3979 33259 5899
rect 34061 5779 35059 5899
rect 37301 5779 38299 5899
rect 34061 5659 35179 5779
rect 37181 5659 38299 5779
rect 34061 5501 35299 5659
rect 34181 5419 35299 5501
rect 37061 5501 38299 5659
rect 37061 5419 38179 5501
rect 34181 5299 35419 5419
rect 36941 5299 38179 5419
rect 34181 5261 35539 5299
rect 34301 5141 35539 5261
rect 36821 5261 38179 5299
rect 36821 5179 38059 5261
rect 34421 5059 35539 5141
rect 36701 5141 38059 5179
rect 34421 5021 35659 5059
rect 34541 4939 35659 5021
rect 36701 5021 37939 5141
rect 36701 4939 37819 5021
rect 34541 4819 35779 4939
rect 36581 4819 37819 4939
rect 34541 4781 35899 4819
rect 34661 4661 35899 4781
rect 34781 4579 35899 4661
rect 36461 4781 37819 4819
rect 36461 4661 37699 4781
rect 36461 4579 37579 4661
rect 34781 4459 36019 4579
rect 36341 4459 37579 4579
rect 34781 4421 36139 4459
rect 34901 4339 36139 4421
rect 36221 4421 37579 4459
rect 36221 4339 37459 4421
rect 34901 4301 37459 4339
rect 35021 4061 37339 4301
rect 26981 3739 28099 3821
rect 26741 3619 28099 3739
rect 24701 3461 28099 3619
rect 24701 3341 27979 3461
rect 24701 3221 27859 3341
rect 24701 3101 27739 3221
rect 24701 2981 27619 3101
rect 29021 2981 33259 3979
rect 35141 3941 37219 4061
rect 35261 3821 37099 3941
rect 35261 3701 36979 3821
rect 35381 3581 36979 3701
rect 35501 3461 36859 3581
rect 35501 3341 36739 3461
rect 20741 1819 21739 2981
rect 24701 2861 27499 2981
rect 24701 2741 27259 2861
rect 24701 2621 27019 2741
rect 20741 1699 23899 1819
rect 20741 941 24019 1699
rect 24701 941 25699 2621
rect 20741 821 23899 941
rect 24821 821 25699 941
rect 29021 941 30019 2981
rect 32261 941 33259 2981
rect 35621 941 36739 3341
rect 29021 821 29899 941
rect 32261 821 33139 941
rect 35741 821 36619 941
<< metal5 >>
rect 12260 18259 12700 18340
rect 3980 16819 4420 16900
rect 3980 16780 4061 16819
rect 3860 16699 4061 16780
rect 4339 16780 4420 16819
rect 4339 16699 4780 16780
rect 3860 16420 3941 16699
rect 3380 16339 3941 16420
rect 3380 16300 3461 16339
rect 3260 16219 3461 16300
rect 3260 15940 3341 16219
rect 2900 15859 3341 15940
rect 2900 15820 2981 15859
rect 2780 15739 2981 15820
rect 2780 15341 2861 15739
rect 3139 15341 3341 15859
rect 2780 15260 3341 15341
rect 3260 14861 3341 15260
rect 3260 14780 3461 14861
rect 3380 14741 3461 14780
rect 3739 14741 3941 16339
rect 3380 14660 3941 14741
rect 3860 14261 3941 14660
rect 4339 16579 4541 16699
rect 4699 16660 4780 16699
rect 4699 16579 4900 16660
rect 3860 14180 4061 14261
rect 3980 14141 4061 14180
rect 4339 14141 4421 16579
rect 4819 16420 4900 16579
rect 4819 16339 5020 16420
rect 3980 14060 4421 14141
rect 4340 13660 4421 14060
rect 4100 13579 4421 13660
rect 4100 13540 4181 13579
rect 3980 13459 4181 13540
rect 3980 13420 4061 13459
rect 3860 13339 4061 13420
rect 3860 12940 3941 13339
rect 3500 12859 3941 12940
rect 3500 12820 3581 12859
rect 3380 12739 3581 12820
rect 3380 12700 3461 12739
rect 3260 12619 3461 12700
rect 3260 12341 3341 12619
rect 3260 12260 3461 12341
rect 3380 12221 3461 12260
rect 3739 12221 3941 12859
rect 3380 12140 3941 12221
rect 3860 11981 3941 12140
rect 3860 11900 4061 11981
rect 3980 11861 4061 11900
rect 4339 11861 4421 13579
rect 3980 11780 4421 11861
rect 4340 11621 4421 11780
rect 4939 15940 5020 16339
rect 4939 15859 5380 15940
rect 4939 15739 5141 15859
rect 5299 15820 5380 15859
rect 5299 15739 5500 15820
rect 4340 11540 4541 11621
rect 4460 11501 4541 11540
rect 4460 11420 4661 11501
rect 4580 11381 4661 11420
rect 4939 11381 5021 15739
rect 5419 15580 5500 15739
rect 5419 15499 5620 15580
rect 4580 11300 5021 11381
rect 4940 11261 5021 11300
rect 5539 15100 5620 15499
rect 5539 15019 5980 15100
rect 4940 11180 5141 11261
rect 5060 11021 5141 11180
rect 5539 11021 5621 15019
rect 5899 14980 5980 15019
rect 5899 14899 6100 14980
rect 5060 10940 5621 11021
rect 5540 10781 5621 10940
rect 6019 14380 6100 14899
rect 6019 14299 6460 14380
rect 5540 10700 5741 10781
rect 5660 10661 5741 10700
rect 5660 10580 5861 10661
rect 5780 10541 5861 10580
rect 6019 10541 6221 14299
rect 6379 14260 6460 14299
rect 6379 14179 6580 14260
rect 6499 14140 6580 14179
rect 6499 14059 6700 14140
rect 5780 10460 6221 10541
rect 6140 10301 6221 10460
rect 6619 13540 6700 14059
rect 6619 13459 7060 13540
rect 6140 10220 6341 10301
rect 6260 10181 6341 10220
rect 6619 10181 6821 13459
rect 6979 13420 7060 13459
rect 6979 13339 7180 13420
rect 7099 13300 7180 13339
rect 7099 13219 7300 13300
rect 3980 10099 4540 10180
rect 6260 10100 6821 10181
rect 3980 9940 4061 10099
rect 4459 10060 4540 10099
rect 4459 9979 4780 10060
rect 3860 9859 4061 9940
rect 4699 9940 4780 9979
rect 4699 9859 5020 9940
rect 3860 9700 3941 9859
rect 4939 9820 5020 9859
rect 6740 9821 6821 10100
rect 7219 12700 7300 13219
rect 11060 12739 11380 12820
rect 11060 12700 11141 12739
rect 7219 12619 7780 12700
rect 4939 9739 5260 9820
rect 6740 9740 6941 9821
rect 3740 9619 3941 9700
rect 5179 9700 5260 9739
rect 6860 9701 6941 9740
rect 7219 9701 7421 12619
rect 7699 12460 7780 12619
rect 10580 12619 11141 12700
rect 11299 12700 11380 12739
rect 11299 12619 11500 12700
rect 10580 12580 10661 12619
rect 10220 12499 10661 12580
rect 7699 12379 7900 12460
rect 5179 9619 5500 9700
rect 6860 9620 7421 9701
rect 3740 9340 3821 9619
rect 5419 9580 5500 9619
rect 5419 9499 5740 9580
rect 5659 9460 5740 9499
rect 7340 9461 7421 9620
rect 7819 11980 7900 12379
rect 10220 11981 10301 12499
rect 11419 12220 11500 12619
rect 11419 12139 11620 12220
rect 7819 11899 8260 11980
rect 10220 11900 10421 11981
rect 5659 9379 5980 9460
rect 7340 9380 7541 9461
rect 3620 9259 3821 9340
rect 5899 9340 5980 9379
rect 7460 9341 7541 9380
rect 7819 9341 8021 11899
rect 8179 11860 8260 11899
rect 8179 11779 8380 11860
rect 8299 11620 8380 11779
rect 10340 11621 10421 11900
rect 8299 11539 8500 11620
rect 10340 11540 10541 11621
rect 5899 9259 6220 9340
rect 7460 9260 8021 9341
rect 3620 9100 3701 9259
rect 6139 9220 6220 9259
rect 6139 9139 6460 9220
rect 3500 9019 3701 9100
rect 6379 9100 6460 9139
rect 6379 9019 6700 9100
rect 3500 8741 3581 9019
rect 6619 8980 6700 9019
rect 7940 8981 8021 9260
rect 8419 11140 8500 11539
rect 10460 11260 10541 11540
rect 11539 11500 11620 12139
rect 11539 11419 11740 11500
rect 10220 11179 10541 11260
rect 10220 11140 10301 11179
rect 8419 11059 8860 11140
rect 6619 8899 6940 8980
rect 7940 8900 8141 8981
rect 6859 8860 6940 8899
rect 8060 8861 8141 8900
rect 8419 8861 8621 11059
rect 8779 11020 8860 11059
rect 9980 11059 10301 11140
rect 9980 11020 10061 11059
rect 8779 10939 8980 11020
rect 8899 10780 8980 10939
rect 9740 10939 10061 11020
rect 8899 10699 9100 10780
rect 6859 8779 7180 8860
rect 8060 8780 8621 8861
rect 3500 8660 3701 8741
rect 3620 8621 3701 8660
rect 7099 8740 7180 8779
rect 7099 8659 7300 8740
rect 3620 8540 4061 8621
rect 3980 8501 4061 8540
rect 7219 8620 7300 8659
rect 7219 8539 7660 8620
rect 3980 8420 4421 8501
rect 4340 8381 4421 8420
rect 7579 8500 7660 8539
rect 8540 8501 8621 8780
rect 9019 10300 9100 10699
rect 9740 10661 9821 10939
rect 9740 10580 9941 10661
rect 9860 10421 9941 10580
rect 11659 10660 11740 11419
rect 11659 10579 11860 10660
rect 9860 10340 10061 10421
rect 9019 10219 9460 10300
rect 9019 8501 9101 10219
rect 9379 10180 9460 10219
rect 9980 10181 10061 10340
rect 9379 10099 9580 10180
rect 9980 10100 10181 10181
rect 9499 9940 9580 10099
rect 10100 10061 10181 10100
rect 10100 9980 10301 10061
rect 9499 9859 9700 9940
rect 7579 8419 7780 8500
rect 8540 8420 9101 8501
rect 4340 8300 4781 8381
rect 4700 8261 4781 8300
rect 7699 8380 7780 8419
rect 7699 8299 8020 8380
rect 4700 8180 5141 8261
rect 5060 8141 5141 8180
rect 7939 8260 8020 8299
rect 9020 8261 9101 8420
rect 9619 9580 9700 9859
rect 10220 9821 10301 9980
rect 11779 9940 11860 10579
rect 11779 9859 11980 9940
rect 10220 9740 10421 9821
rect 10340 9581 10421 9740
rect 9619 9499 9940 9580
rect 10340 9500 10541 9581
rect 7939 8179 8260 8260
rect 9020 8180 9221 8261
rect 5060 8060 5501 8141
rect 5420 8021 5501 8060
rect 8179 8140 8260 8179
rect 9140 8141 9221 8180
rect 9619 8141 9701 9499
rect 9859 9460 9940 9499
rect 9859 9379 10060 9460
rect 9979 9340 10060 9379
rect 10460 9341 10541 9500
rect 9979 9259 10180 9340
rect 10460 9260 10661 9341
rect 8179 8059 8500 8140
rect 9140 8060 9341 8141
rect 5420 7940 5861 8021
rect 5780 7901 5861 7940
rect 8419 8020 8500 8059
rect 9260 8021 9341 8060
rect 9499 8021 9701 8141
rect 8419 7939 8740 8020
rect 9260 7940 9701 8021
rect 5780 7820 6221 7901
rect 6140 7781 6221 7820
rect 8659 7900 8740 7939
rect 8659 7819 8980 7900
rect 6140 7700 6701 7781
rect 6620 7661 6701 7700
rect 8899 7780 8980 7819
rect 9620 7781 9701 7940
rect 10099 8740 10180 9259
rect 10580 9101 10661 9260
rect 11899 9220 11980 9859
rect 11899 9139 12100 9220
rect 10580 9020 10781 9101
rect 10700 8861 10781 9020
rect 10700 8740 10901 8861
rect 10099 8659 10901 8740
rect 8899 7699 9220 7780
rect 9620 7700 9821 7781
rect 6620 7580 6941 7661
rect 6860 7541 6941 7580
rect 9139 7660 9220 7699
rect 9740 7661 9821 7700
rect 9139 7579 9460 7660
rect 6860 7460 7421 7541
rect 7340 7421 7421 7460
rect 9379 7540 9460 7579
rect 9740 7541 9941 7661
rect 10099 7541 10301 8659
rect 10579 8621 10901 8659
rect 10579 8450 11021 8621
rect 10579 8419 10780 8450
rect 9740 7540 10301 7541
rect 9379 7460 10301 7540
rect 9379 7459 9940 7460
rect 7340 7340 7781 7421
rect 7700 7301 7781 7340
rect 9619 7339 9940 7459
rect 7700 7220 8141 7301
rect 8060 7181 8141 7220
rect 9859 7300 9940 7339
rect 10220 7301 10301 7460
rect 10699 7900 10780 8419
rect 10940 8381 11021 8450
rect 10940 8300 11141 8381
rect 11060 8141 11141 8300
rect 12019 8380 12100 9139
rect 12260 8380 12341 18259
rect 12619 18220 12700 18259
rect 12619 18139 13060 18220
rect 12979 18100 13060 18139
rect 12979 18019 13300 18100
rect 13219 17980 13300 18019
rect 13219 17899 13540 17980
rect 13459 17860 13540 17899
rect 13459 17779 13780 17860
rect 13699 17740 13780 17779
rect 13699 17659 14020 17740
rect 13939 17620 14020 17659
rect 13939 17539 14260 17620
rect 14179 17500 14260 17539
rect 14179 17419 14380 17500
rect 14299 17141 14380 17419
rect 14179 17060 14380 17141
rect 14179 16421 14260 17060
rect 14059 16340 14260 16421
rect 14059 15581 14140 16340
rect 13939 15500 14140 15581
rect 13939 14861 14020 15500
rect 13819 14780 14020 14861
rect 15140 14899 15580 14980
rect 13819 14141 13900 14780
rect 15140 14740 15221 14899
rect 15499 14860 15580 14899
rect 15499 14779 15940 14860
rect 15020 14659 15221 14740
rect 15859 14740 15940 14779
rect 15859 14659 16180 14740
rect 15020 14380 15101 14659
rect 16099 14620 16180 14659
rect 16099 14539 16540 14620
rect 16459 14500 16540 14539
rect 16459 14419 16780 14500
rect 13699 14060 13900 14141
rect 14900 14299 15101 14380
rect 13699 13421 13780 14060
rect 14900 14020 14981 14299
rect 16699 14141 16780 14419
rect 14780 13939 14981 14020
rect 16579 14060 16780 14141
rect 14780 13540 14861 13939
rect 16579 13901 16660 14060
rect 16459 13820 16660 13901
rect 16459 13661 16540 13820
rect 13579 13340 13780 13421
rect 14660 13459 14861 13540
rect 16339 13580 16540 13661
rect 13579 12581 13660 13340
rect 14660 13300 14741 13459
rect 16339 13421 16420 13580
rect 14540 13219 14741 13300
rect 16219 13340 16420 13421
rect 14540 12820 14621 13219
rect 16219 13181 16300 13340
rect 16099 13100 16300 13181
rect 16099 12941 16180 13100
rect 13459 12500 13660 12581
rect 14420 12739 14621 12820
rect 15979 12860 16180 12941
rect 13459 11741 13540 12500
rect 14420 12460 14501 12739
rect 15979 12701 16060 12860
rect 15859 12620 16060 12701
rect 15859 12461 15940 12620
rect 14300 12379 14501 12460
rect 15739 12380 15940 12461
rect 14300 12100 14381 12379
rect 15739 12221 15820 12380
rect 13339 11660 13540 11741
rect 14180 12019 14381 12100
rect 15619 12140 15820 12221
rect 14180 11740 14261 12019
rect 15619 11981 15700 12140
rect 15499 11900 15700 11981
rect 15499 11741 15580 11900
rect 13339 11021 13420 11660
rect 14060 11659 14261 11740
rect 15379 11660 15580 11741
rect 14060 11380 14141 11659
rect 15379 11501 15460 11660
rect 13219 10940 13420 11021
rect 13940 11299 14141 11380
rect 15259 11420 15460 11501
rect 13940 11020 14021 11299
rect 15259 11261 15340 11420
rect 15139 11180 15340 11261
rect 15139 11021 15220 11180
rect 13219 10301 13300 10940
rect 13820 10939 14021 11020
rect 15019 10940 15220 11021
rect 13820 10660 13901 10939
rect 15019 10781 15100 10940
rect 13099 10220 13300 10301
rect 13700 10579 13901 10660
rect 14899 10700 15100 10781
rect 13700 10300 13781 10579
rect 14899 10541 14980 10700
rect 14779 10460 14980 10541
rect 14779 10301 14860 10460
rect 13099 9581 13180 10220
rect 13580 10219 13781 10300
rect 14659 10220 14860 10301
rect 13580 9940 13661 10219
rect 14659 10061 14740 10220
rect 12979 9500 13180 9581
rect 13460 9859 13661 9940
rect 14539 9980 14740 10061
rect 13460 9580 13541 9859
rect 14539 9821 14620 9980
rect 14419 9740 14620 9821
rect 14419 9581 14500 9740
rect 12979 8741 13060 9500
rect 13340 9499 13541 9580
rect 14299 9500 14500 9581
rect 13340 9100 13421 9499
rect 14299 9341 14380 9500
rect 14179 9260 14380 9341
rect 14179 9101 14260 9260
rect 12019 8299 12341 8380
rect 11060 8060 11261 8141
rect 11180 7901 11261 8060
rect 11180 7900 11381 7901
rect 10699 7819 11381 7900
rect 10220 7300 10421 7301
rect 9859 7219 10421 7300
rect 10099 7181 10421 7219
rect 10699 7181 10901 7819
rect 11179 7661 11381 7819
rect 12139 7781 12341 8299
rect 12859 8740 13060 8741
rect 13220 9019 13421 9100
rect 14059 9020 14260 9101
rect 13220 8740 13301 9019
rect 14059 8861 14140 9020
rect 13939 8780 14140 8861
rect 13939 8741 14020 8780
rect 12859 8659 13301 8740
rect 13819 8660 14020 8741
rect 12859 8419 13181 8659
rect 13819 8501 13900 8660
rect 13699 8420 13900 8501
rect 12859 8059 13061 8419
rect 13699 8261 13780 8420
rect 13579 8180 13780 8261
rect 12859 8021 12941 8059
rect 13579 8021 13660 8180
rect 12739 7781 12941 8021
rect 13459 7940 13660 8021
rect 13459 7781 13540 7940
rect 11899 7700 12941 7781
rect 11899 7661 11980 7700
rect 11179 7579 11501 7661
rect 11299 7541 11501 7579
rect 11659 7580 11980 7661
rect 12860 7661 12941 7700
rect 13339 7700 13540 7781
rect 13339 7661 13420 7700
rect 12860 7580 13420 7661
rect 11659 7541 11740 7580
rect 11299 7460 11740 7541
rect 11299 7421 11380 7460
rect 11179 7340 11380 7421
rect 11179 7301 11260 7340
rect 11059 7220 11260 7301
rect 11059 7181 11140 7220
rect 8060 7100 8501 7181
rect 8420 7061 8501 7100
rect 10099 7100 11140 7181
rect 10099 7099 10660 7100
rect 8420 6980 8861 7061
rect 8780 6941 8861 6980
rect 10339 6979 10660 7099
rect 11900 7099 12820 7180
rect 11900 7060 11981 7099
rect 8780 6860 9221 6941
rect 9140 6821 9221 6860
rect 10579 6940 10660 6979
rect 11660 6979 11981 7060
rect 12739 7060 12820 7099
rect 12739 6979 13060 7060
rect 11660 6940 11741 6979
rect 10579 6859 10780 6940
rect 9140 6740 9581 6821
rect 9500 6701 9581 6740
rect 9500 6620 9941 6701
rect 9860 6581 9941 6620
rect 10699 6581 10780 6859
rect 11540 6859 11741 6940
rect 12979 6940 13060 6979
rect 12979 6859 13300 6940
rect 11540 6820 11621 6859
rect 11420 6739 11621 6820
rect 13219 6820 13300 6859
rect 13219 6739 13420 6820
rect 11420 6700 11501 6739
rect 9860 6500 10300 6581
rect 10220 6460 10300 6500
rect 10580 6500 10780 6581
rect 11300 6619 11501 6700
rect 10580 6460 10660 6500
rect 11300 6460 11381 6619
rect 13339 6580 13420 6739
rect 13339 6499 13540 6580
rect 10220 6340 10660 6460
rect 11180 6379 11381 6460
rect 11180 6340 11261 6379
rect 1460 6259 11261 6340
rect 13459 6340 13540 6499
rect 13459 6259 13660 6340
rect 1460 6220 1541 6259
rect 1340 6139 1541 6220
rect 1340 5741 1421 6139
rect 1340 5660 1541 5741
rect 1460 5621 1541 5660
rect 13579 5621 13660 6259
rect 1460 5540 11261 5621
rect 10340 5419 10660 5540
rect 11180 5501 11261 5540
rect 13459 5540 13660 5621
rect 15620 5899 16780 5980
rect 11180 5420 11381 5501
rect 10340 5380 10421 5419
rect 9980 5299 10421 5380
rect 10579 5380 10660 5419
rect 10579 5299 10780 5380
rect 9980 5260 10061 5299
rect 9620 5179 10061 5260
rect 9620 5140 9701 5179
rect 9260 5059 9701 5140
rect 9260 5020 9341 5059
rect 8900 4939 9341 5020
rect 8900 4900 8981 4939
rect 10699 4901 10780 5299
rect 11300 5261 11381 5420
rect 13459 5381 13540 5540
rect 13339 5300 13540 5381
rect 11300 5180 11501 5261
rect 11420 5141 11501 5180
rect 13339 5141 13420 5300
rect 11420 5060 11621 5141
rect 11540 5021 11621 5060
rect 13219 5060 13420 5141
rect 13219 5021 13300 5060
rect 11540 4940 11741 5021
rect 8540 4819 8981 4900
rect 10459 4900 10780 4901
rect 11660 4901 11741 4940
rect 13099 4940 13300 5021
rect 13099 4901 13180 4940
rect 10459 4820 11020 4900
rect 11660 4820 11981 4901
rect 8540 4780 8621 4819
rect 10459 4781 10660 4820
rect 8180 4699 8621 4780
rect 10219 4699 10660 4781
rect 10940 4780 11020 4820
rect 11900 4781 11981 4820
rect 12859 4820 13180 4901
rect 12859 4781 12940 4820
rect 10940 4699 11140 4780
rect 11900 4700 12940 4781
rect 8180 4660 8261 4699
rect 10219 4661 10541 4699
rect 7700 4579 8261 4660
rect 9979 4579 10541 4661
rect 7700 4540 7781 4579
rect 9979 4541 10301 4579
rect 7340 4459 7781 4540
rect 9739 4459 10301 4541
rect 7340 4420 7421 4459
rect 9739 4421 10181 4459
rect 11059 4421 11140 4699
rect 6980 4339 7421 4420
rect 9499 4340 10181 4421
rect 6980 4300 7061 4339
rect 9499 4301 9580 4340
rect 6620 4219 7061 4300
rect 6620 4180 6701 4219
rect 9259 4181 9580 4301
rect 6260 4099 6701 4180
rect 9019 4180 9580 4181
rect 9740 4339 10181 4340
rect 10939 4420 11140 4421
rect 10939 4339 11620 4420
rect 9740 4219 10061 4339
rect 10939 4301 11141 4339
rect 10819 4219 11141 4301
rect 11539 4300 11620 4339
rect 11539 4219 11860 4300
rect 9740 4180 9821 4219
rect 10819 4181 11021 4219
rect 9019 4099 9821 4180
rect 10699 4099 11021 4181
rect 11779 4180 11860 4219
rect 11779 4099 12460 4180
rect 6260 4060 6341 4099
rect 9019 4061 9701 4099
rect 10699 4061 10901 4099
rect 5900 3979 6341 4060
rect 8779 3980 9701 4061
rect 5900 3940 5981 3979
rect 8779 3941 8860 3980
rect 5540 3859 5981 3940
rect 8539 3860 8860 3941
rect 9260 3979 9701 3980
rect 5540 3820 5621 3859
rect 8539 3821 8620 3860
rect 5180 3739 5621 3820
rect 8299 3740 8620 3821
rect 9260 3859 9461 3979
rect 10579 3941 10901 4061
rect 11899 3979 12101 4099
rect 12379 4060 12460 4099
rect 12379 3979 12580 4060
rect 11899 3941 11981 3979
rect 10459 3859 10901 3941
rect 9260 3820 9341 3859
rect 10459 3821 10781 3859
rect 5180 3700 5261 3739
rect 8299 3701 8380 3740
rect 4820 3619 5261 3700
rect 8059 3620 8380 3701
rect 9140 3739 9341 3820
rect 10339 3739 10781 3821
rect 9140 3700 9221 3739
rect 10339 3701 10661 3739
rect 11779 3701 11981 3941
rect 4820 3580 4901 3619
rect 8059 3581 8140 3620
rect 4340 3499 4901 3580
rect 7819 3500 8140 3581
rect 8900 3619 9221 3700
rect 10219 3620 10661 3701
rect 8900 3580 8981 3619
rect 10219 3581 10300 3620
rect 4340 3460 4421 3499
rect 7819 3461 7900 3500
rect 4100 3379 4421 3460
rect 7579 3380 7900 3461
rect 8780 3499 8981 3580
rect 8780 3460 8861 3499
rect 10099 3461 10300 3581
rect 4100 3340 4181 3379
rect 7579 3341 7660 3380
rect 3740 3259 4181 3340
rect 7339 3260 7660 3341
rect 8540 3379 8861 3460
rect 9979 3460 10300 3461
rect 10460 3619 10661 3620
rect 10460 3460 10541 3619
rect 9979 3379 10541 3460
rect 11659 3379 11981 3701
rect 8540 3340 8621 3379
rect 9979 3341 10421 3379
rect 3740 3220 3821 3259
rect 7339 3221 7420 3260
rect 3620 3139 3821 3220
rect 7099 3140 7420 3221
rect 8420 3259 8621 3340
rect 9859 3310 10421 3341
rect 9859 3260 10060 3310
rect 8420 3220 8501 3259
rect 9859 3221 9940 3260
rect 3620 2981 3701 3139
rect 7099 3101 7180 3140
rect 6859 3020 7180 3101
rect 8300 3139 8501 3220
rect 9739 3140 9940 3221
rect 10220 3259 10421 3310
rect 8300 3100 8381 3139
rect 9739 3101 9820 3140
rect 6859 2981 6940 3020
rect 3620 2900 3821 2981
rect 3740 2861 3821 2900
rect 6619 2900 6940 2981
rect 8060 3019 8381 3100
rect 9619 3020 9820 3101
rect 10220 3100 10301 3259
rect 11659 3221 11861 3379
rect 8060 2980 8141 3019
rect 9619 2981 9700 3020
rect 6619 2861 6700 2900
rect 3740 2780 3941 2861
rect 3860 2741 3941 2780
rect 6379 2780 6700 2861
rect 7940 2899 8141 2980
rect 9499 2900 9700 2981
rect 10100 3019 10301 3100
rect 11539 3140 11861 3221
rect 10100 2980 10181 3019
rect 7940 2860 8021 2899
rect 9499 2861 9580 2900
rect 6379 2741 6460 2780
rect 3860 2660 4181 2741
rect 4100 2621 4181 2660
rect 6139 2660 6460 2741
rect 7820 2779 8021 2860
rect 9379 2780 9580 2861
rect 9980 2899 10181 2980
rect 9980 2860 10061 2899
rect 11539 2861 11620 3140
rect 7820 2740 7901 2779
rect 9379 2741 9460 2780
rect 6139 2621 6220 2660
rect 4100 2540 4301 2621
rect 4220 2501 4301 2540
rect 5899 2540 6220 2621
rect 7580 2659 7901 2740
rect 9259 2660 9460 2741
rect 9860 2779 10061 2860
rect 7580 2620 7661 2659
rect 9259 2621 9340 2660
rect 5899 2501 5980 2540
rect 4220 2420 4421 2501
rect 4340 2381 4421 2420
rect 5659 2420 5980 2501
rect 7460 2539 7661 2620
rect 9139 2540 9340 2621
rect 9860 2620 9941 2779
rect 11419 2740 11620 2861
rect 11780 2740 11861 3140
rect 11419 2659 11861 2740
rect 7460 2500 7541 2539
rect 9139 2501 9220 2540
rect 5659 2381 5740 2420
rect 4340 2300 4661 2381
rect 4580 2261 4661 2300
rect 5419 2300 5740 2381
rect 7220 2419 7541 2500
rect 9019 2420 9220 2501
rect 9740 2539 9941 2620
rect 9740 2500 9821 2539
rect 7220 2380 7301 2419
rect 9019 2381 9100 2420
rect 5419 2261 5500 2300
rect 4580 2180 4781 2261
rect 4700 2141 4781 2180
rect 5179 2180 5500 2261
rect 7100 2299 7301 2380
rect 8899 2300 9100 2381
rect 9620 2419 9821 2500
rect 10699 2501 10901 2621
rect 11419 2580 11741 2659
rect 11419 2501 11500 2580
rect 10699 2420 11141 2501
rect 9620 2380 9701 2419
rect 10699 2381 10780 2420
rect 7100 2260 7181 2299
rect 8899 2261 8980 2300
rect 5179 2141 5260 2180
rect 4700 2060 5260 2141
rect 6980 2179 7181 2260
rect 8779 2180 8980 2261
rect 9500 2299 9701 2380
rect 10579 2300 10780 2381
rect 11060 2381 11141 2420
rect 11299 2420 11500 2501
rect 11299 2381 11380 2420
rect 11060 2300 11380 2381
rect 6980 2140 7061 2179
rect 8779 2141 8860 2180
rect 6740 2059 7061 2140
rect 8659 2060 8860 2141
rect 9500 2140 9581 2299
rect 10579 2141 10660 2300
rect 6740 2020 6821 2059
rect 8659 2021 8740 2060
rect 6620 1939 6821 2020
rect 8539 1940 8740 2021
rect 9380 2059 9581 2140
rect 10459 2060 10660 2141
rect 9380 2020 9461 2059
rect 6620 1900 6701 1939
rect 8539 1901 8620 1940
rect 6500 1819 6701 1900
rect 8419 1820 8620 1901
rect 9260 1939 9461 2020
rect 6500 1780 6581 1819
rect 8419 1781 8500 1820
rect 6260 1699 6581 1780
rect 8299 1700 8500 1781
rect 9260 1780 9341 1939
rect 10459 1901 10540 2060
rect 11660 2020 11741 2580
rect 6260 1421 6341 1699
rect 8299 1661 8380 1700
rect 8179 1580 8380 1661
rect 9140 1699 9341 1780
rect 10339 1820 10540 1901
rect 11540 1939 11741 2020
rect 9140 1660 9221 1699
rect 10339 1661 10420 1820
rect 8179 1541 8260 1580
rect 8059 1460 8260 1541
rect 9020 1579 9221 1660
rect 10219 1580 10420 1661
rect 9020 1540 9101 1579
rect 8059 1421 8140 1460
rect 6260 1340 6581 1421
rect 6500 1301 6581 1340
rect 7939 1340 8140 1421
rect 8900 1459 9101 1540
rect 7939 1301 8020 1340
rect 6500 1220 6941 1301
rect 6860 1181 6941 1220
rect 7819 1220 8020 1301
rect 8900 1300 8981 1459
rect 10219 1421 10300 1580
rect 7819 1181 7900 1220
rect 6860 1100 7301 1181
rect 7220 1061 7301 1100
rect 7699 1100 7900 1181
rect 8780 1219 8981 1300
rect 10099 1340 10300 1421
rect 8780 1180 8861 1219
rect 10099 1181 10180 1340
rect 7699 1061 7780 1100
rect 7220 980 7780 1061
rect 8660 1099 8861 1180
rect 9979 1100 10180 1181
rect 8660 821 8741 1099
rect 9979 941 10060 1100
rect 11540 1061 11621 1939
rect 12499 1301 12580 3979
rect 12379 1220 12580 1301
rect 12379 1181 12460 1220
rect 11899 1100 12460 1181
rect 11899 1061 11980 1100
rect 11540 980 11980 1061
rect 9859 860 10060 941
rect 9859 821 9940 860
rect 8660 740 9940 821
rect 15620 821 15701 5899
rect 16699 4060 16780 5899
rect 18860 5899 20020 5980
rect 18860 4060 18941 5899
rect 16699 3979 18941 4060
rect 16699 2900 18941 2981
rect 16699 821 16780 2900
rect 15620 740 16780 821
rect 18860 821 18941 2900
rect 19939 821 20020 5899
rect 18860 740 20020 821
rect 20660 5899 23980 5980
rect 20660 821 20741 5899
rect 23899 5860 23980 5899
rect 24620 5899 27220 5980
rect 23899 5779 24100 5860
rect 24019 5021 24100 5779
rect 23779 4940 24100 5021
rect 23779 4901 23860 4940
rect 21739 4820 23860 4901
rect 21739 4060 21820 4820
rect 21739 3979 23500 4060
rect 23419 3940 23500 3979
rect 23419 3859 23740 3940
rect 23659 2981 23740 3859
rect 21739 2900 23740 2981
rect 21739 1900 21820 2900
rect 21739 1819 23980 1900
rect 23899 1780 23980 1819
rect 23899 1699 24100 1780
rect 24019 941 24100 1699
rect 23899 860 24100 941
rect 24620 941 24701 5899
rect 27139 5860 27220 5899
rect 28940 5899 30100 5980
rect 27139 5779 27460 5860
rect 27379 5740 27460 5779
rect 27379 5659 27700 5740
rect 27619 5620 27700 5659
rect 27619 5539 27820 5620
rect 27739 5500 27820 5539
rect 27739 5419 27940 5500
rect 27859 5380 27940 5419
rect 27859 5299 28060 5380
rect 27979 5140 28060 5299
rect 27979 5059 28180 5140
rect 25699 4820 26861 4901
rect 25699 3700 25780 4820
rect 26780 4781 26861 4820
rect 28099 4900 28180 5059
rect 28099 4819 28300 4900
rect 26780 4700 26981 4781
rect 26900 4661 26981 4700
rect 26900 4580 27101 4661
rect 27020 4421 27101 4580
rect 27020 4340 27221 4421
rect 27140 4180 27221 4340
rect 27020 4099 27221 4180
rect 27020 3940 27101 4099
rect 26900 3859 27101 3940
rect 26900 3820 26981 3859
rect 28219 3821 28300 4819
rect 26660 3739 26981 3820
rect 28099 3740 28300 3821
rect 26660 3700 26741 3739
rect 25699 3619 26741 3700
rect 28099 3461 28180 3740
rect 27979 3380 28180 3461
rect 27979 3341 28060 3380
rect 27859 3260 28060 3341
rect 27859 3221 27940 3260
rect 27739 3140 27940 3221
rect 27739 3101 27820 3140
rect 27619 3020 27820 3101
rect 27619 2981 27700 3020
rect 27499 2900 27700 2981
rect 27499 2861 27580 2900
rect 27259 2780 27580 2861
rect 27259 2741 27340 2780
rect 27019 2660 27340 2741
rect 27019 2621 27100 2660
rect 25699 2540 27100 2621
rect 24620 860 24821 941
rect 23899 821 23980 860
rect 20660 740 23980 821
rect 24740 821 24821 860
rect 25699 821 25780 2540
rect 24740 740 25780 821
rect 28940 821 29021 5899
rect 30019 4060 30100 5899
rect 32180 5899 33340 5980
rect 32180 4060 32261 5899
rect 30019 3979 32261 4060
rect 30019 2900 32261 2981
rect 30019 941 30100 2900
rect 29899 860 30100 941
rect 29899 821 29980 860
rect 28940 740 29980 821
rect 32180 821 32261 2900
rect 33259 941 33340 5899
rect 33980 5899 35140 5980
rect 33980 5501 34061 5899
rect 35059 5860 35140 5899
rect 37220 5899 38380 5980
rect 37220 5860 37301 5899
rect 35059 5779 35260 5860
rect 35179 5740 35260 5779
rect 37100 5779 37301 5860
rect 37100 5740 37181 5779
rect 35179 5659 35380 5740
rect 33980 5420 34181 5501
rect 34100 5261 34181 5420
rect 35299 5500 35380 5659
rect 36980 5659 37181 5740
rect 36980 5500 37061 5659
rect 38299 5501 38380 5899
rect 35299 5419 35500 5500
rect 35419 5380 35500 5419
rect 36860 5419 37061 5500
rect 38179 5420 38380 5501
rect 36860 5380 36941 5419
rect 35419 5299 35620 5380
rect 34100 5180 34301 5261
rect 34220 5141 34301 5180
rect 34220 5060 34421 5141
rect 34340 5021 34421 5060
rect 35539 5140 35620 5299
rect 36740 5299 36941 5380
rect 36740 5260 36821 5299
rect 38179 5261 38260 5420
rect 36620 5179 36821 5260
rect 38059 5180 38260 5261
rect 35539 5059 35740 5140
rect 34340 4940 34541 5021
rect 34460 4781 34541 4940
rect 35659 5020 35740 5059
rect 36620 5020 36701 5179
rect 38059 5141 38140 5180
rect 37939 5060 38140 5141
rect 37939 5021 38020 5060
rect 35659 4939 35860 5020
rect 35779 4900 35860 4939
rect 36500 4939 36701 5020
rect 37819 4940 38020 5021
rect 36500 4900 36581 4939
rect 35779 4819 35980 4900
rect 34460 4700 34661 4781
rect 34580 4661 34661 4700
rect 34580 4580 34781 4661
rect 34700 4421 34781 4580
rect 35899 4660 35980 4819
rect 36380 4819 36581 4900
rect 36380 4660 36461 4819
rect 37819 4781 37900 4940
rect 37699 4700 37900 4781
rect 37699 4661 37780 4700
rect 35899 4579 36100 4660
rect 36019 4540 36100 4579
rect 36260 4579 36461 4660
rect 37579 4580 37780 4661
rect 36260 4540 36341 4579
rect 36019 4459 36341 4540
rect 34700 4340 34901 4421
rect 34820 4301 34901 4340
rect 36139 4339 36221 4459
rect 37579 4421 37660 4580
rect 37459 4340 37660 4421
rect 37459 4301 37540 4340
rect 34820 4220 35021 4301
rect 34940 4061 35021 4220
rect 37339 4220 37540 4301
rect 37339 4061 37420 4220
rect 34940 3980 35141 4061
rect 35060 3941 35141 3980
rect 37219 3980 37420 4061
rect 37219 3941 37300 3980
rect 35060 3860 35261 3941
rect 35180 3701 35261 3860
rect 37099 3860 37300 3941
rect 37099 3821 37180 3860
rect 36979 3740 37180 3821
rect 35180 3620 35381 3701
rect 35300 3581 35381 3620
rect 36979 3581 37060 3740
rect 35300 3500 35501 3581
rect 35420 3341 35501 3500
rect 36859 3500 37060 3581
rect 36859 3461 36940 3500
rect 36739 3380 36940 3461
rect 35420 3260 35621 3341
rect 33139 860 33340 941
rect 35540 941 35621 3260
rect 36739 941 36820 3380
rect 35540 860 35741 941
rect 33139 821 33220 860
rect 32180 740 33220 821
rect 35660 821 35741 860
rect 36619 860 36820 941
rect 36619 821 36700 860
rect 35660 740 36700 821
<< end >>
