magic
tech sky130A
magscale 1 2
timestamp 1685096196
<< metal3 >>
rect -1386 2512 1386 2540
rect -1386 -2512 1302 2512
rect 1366 -2512 1386 2512
rect -1386 -2540 1386 -2512
<< via3 >>
rect 1302 -2512 1366 2512
<< mimcap >>
rect -1346 2460 1054 2500
rect -1346 -2460 -1306 2460
rect 1014 -2460 1054 2460
rect -1346 -2500 1054 -2460
<< mimcapcontact >>
rect -1306 -2460 1014 2460
<< metal4 >>
rect 1286 2512 1382 2528
rect -1307 2460 1015 2461
rect -1307 -2460 -1306 2460
rect 1014 -2460 1015 2460
rect -1307 -2461 1015 -2460
rect 1286 -2512 1302 2512
rect 1366 -2512 1382 2512
rect 1286 -2528 1382 -2512
<< properties >>
string FIXED_BBOX -1386 -2540 1094 2540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12 l 25 val 614.06 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
