magic
tech sky130A
magscale 1 2
timestamp 1683627527
<< metal1 >>
rect 1348 3588 3224 3696
rect 1482 3376 1492 3556
rect 1556 3376 1566 3556
rect 1798 3376 1808 3556
rect 1872 3376 1882 3556
rect 2114 3376 2124 3556
rect 2188 3376 2198 3556
rect 2430 3376 2440 3556
rect 2504 3376 2514 3556
rect 2746 3376 2756 3556
rect 2820 3376 2830 3556
rect 1326 3152 1336 3332
rect 1400 3152 1410 3332
rect 1642 3152 1652 3332
rect 1716 3152 1726 3332
rect 1958 3152 1968 3332
rect 2032 3152 2042 3332
rect 2274 3152 2284 3332
rect 2348 3152 2358 3332
rect 2590 3152 2600 3332
rect 2664 3152 2674 3332
rect 2906 3152 2916 3332
rect 2980 3152 2990 3332
rect 3020 3120 3224 3588
rect 1348 2952 3224 3120
rect 1482 2740 1492 2920
rect 1556 2740 1566 2920
rect 1798 2740 1808 2920
rect 1872 2740 1882 2920
rect 2114 2740 2124 2920
rect 2188 2740 2198 2920
rect 2430 2740 2440 2920
rect 2504 2740 2514 2920
rect 2746 2740 2756 2920
rect 2820 2740 2830 2920
rect 1326 2516 1336 2696
rect 1400 2516 1410 2696
rect 1642 2516 1652 2696
rect 1716 2516 1726 2696
rect 1958 2516 1968 2696
rect 2032 2516 2042 2696
rect 2274 2516 2284 2696
rect 2348 2516 2358 2696
rect 2590 2516 2600 2696
rect 2664 2516 2674 2696
rect 2906 2516 2916 2696
rect 2980 2516 2990 2696
rect 3020 2480 3224 2952
rect 1348 2312 3224 2480
rect 1482 2100 1492 2280
rect 1556 2100 1566 2280
rect 1798 2100 1808 2280
rect 1872 2100 1882 2280
rect 2114 2100 2124 2280
rect 2188 2100 2198 2280
rect 2430 2100 2440 2280
rect 2504 2100 2514 2280
rect 2746 2100 2756 2280
rect 2820 2100 2830 2280
rect 1326 1876 1336 2056
rect 1400 1876 1410 2056
rect 1642 1876 1652 2056
rect 1716 1876 1726 2056
rect 1958 1876 1968 2056
rect 2032 1876 2042 2056
rect 2274 1876 2284 2056
rect 2348 1876 2358 2056
rect 2590 1876 2600 2056
rect 2664 1876 2674 2056
rect 2906 1876 2916 2056
rect 2980 1876 2990 2056
rect 3020 1840 3224 2312
rect 1348 1736 3224 1840
rect 2880 1580 3084 1736
rect 1380 1496 3084 1580
rect 1422 1276 1432 1456
rect 1496 1276 1506 1456
rect 1614 1276 1624 1456
rect 1688 1276 1698 1456
rect 1806 1276 1816 1456
rect 1880 1276 1890 1456
rect 1998 1276 2008 1456
rect 2072 1276 2082 1456
rect 2190 1276 2200 1456
rect 2264 1276 2274 1456
rect 2382 1276 2392 1456
rect 2456 1276 2466 1456
rect 2574 1276 2584 1456
rect 2648 1276 2658 1456
rect 2766 1276 2776 1456
rect 2840 1276 2850 1456
rect 1326 1052 1336 1232
rect 1400 1052 1410 1232
rect 1514 1052 1524 1232
rect 1588 1052 1598 1232
rect 1706 1052 1716 1232
rect 1780 1052 1790 1232
rect 1902 1052 1912 1232
rect 1976 1052 1986 1232
rect 2094 1052 2104 1232
rect 2168 1052 2178 1232
rect 2286 1052 2296 1232
rect 2360 1052 2370 1232
rect 2478 1052 2488 1232
rect 2552 1052 2562 1232
rect 2670 1052 2680 1232
rect 2744 1052 2754 1232
rect 2880 1016 3084 1496
rect 1476 860 3084 1016
rect 1422 640 1432 820
rect 1496 640 1506 820
rect 1614 640 1624 820
rect 1688 640 1698 820
rect 1806 640 1816 820
rect 1880 640 1890 820
rect 1998 640 2008 820
rect 2072 640 2082 820
rect 2190 640 2200 820
rect 2264 640 2274 820
rect 2382 640 2392 820
rect 2456 640 2466 820
rect 2574 640 2584 820
rect 2648 640 2658 820
rect 2766 640 2776 820
rect 2840 640 2850 820
rect 1326 416 1336 596
rect 1400 416 1410 596
rect 1514 416 1524 596
rect 1588 416 1598 596
rect 1706 416 1716 596
rect 1780 416 1790 596
rect 1902 416 1912 596
rect 1976 416 1986 596
rect 2094 416 2104 596
rect 2168 416 2178 596
rect 2286 416 2296 596
rect 2360 416 2370 596
rect 2478 416 2488 596
rect 2552 416 2562 596
rect 2670 416 2680 596
rect 2744 416 2754 596
rect 2880 380 3084 860
rect 1380 284 3084 380
<< via1 >>
rect 1492 3376 1556 3556
rect 1808 3376 1872 3556
rect 2124 3376 2188 3556
rect 2440 3376 2504 3556
rect 2756 3376 2820 3556
rect 1336 3152 1400 3332
rect 1652 3152 1716 3332
rect 1968 3152 2032 3332
rect 2284 3152 2348 3332
rect 2600 3152 2664 3332
rect 2916 3152 2980 3332
rect 1492 2740 1556 2920
rect 1808 2740 1872 2920
rect 2124 2740 2188 2920
rect 2440 2740 2504 2920
rect 2756 2740 2820 2920
rect 1336 2516 1400 2696
rect 1652 2516 1716 2696
rect 1968 2516 2032 2696
rect 2284 2516 2348 2696
rect 2600 2516 2664 2696
rect 2916 2516 2980 2696
rect 1492 2100 1556 2280
rect 1808 2100 1872 2280
rect 2124 2100 2188 2280
rect 2440 2100 2504 2280
rect 2756 2100 2820 2280
rect 1336 1876 1400 2056
rect 1652 1876 1716 2056
rect 1968 1876 2032 2056
rect 2284 1876 2348 2056
rect 2600 1876 2664 2056
rect 2916 1876 2980 2056
rect 1432 1276 1496 1456
rect 1624 1276 1688 1456
rect 1816 1276 1880 1456
rect 2008 1276 2072 1456
rect 2200 1276 2264 1456
rect 2392 1276 2456 1456
rect 2584 1276 2648 1456
rect 2776 1276 2840 1456
rect 1336 1052 1400 1232
rect 1524 1052 1588 1232
rect 1716 1052 1780 1232
rect 1912 1052 1976 1232
rect 2104 1052 2168 1232
rect 2296 1052 2360 1232
rect 2488 1052 2552 1232
rect 2680 1052 2744 1232
rect 1432 640 1496 820
rect 1624 640 1688 820
rect 1816 640 1880 820
rect 2008 640 2072 820
rect 2200 640 2264 820
rect 2392 640 2456 820
rect 2584 640 2648 820
rect 2776 640 2840 820
rect 1336 416 1400 596
rect 1524 416 1588 596
rect 1716 416 1780 596
rect 1912 416 1976 596
rect 2104 416 2168 596
rect 2296 416 2360 596
rect 2488 416 2552 596
rect 2680 416 2744 596
<< metal2 >>
rect 1492 3646 2820 3648
rect 1492 3636 3100 3646
rect 1492 3556 2244 3636
rect 1556 3380 1808 3556
rect 1492 3366 1556 3376
rect 1872 3380 2124 3556
rect 1808 3366 1872 3376
rect 2188 3392 2244 3556
rect 2188 3380 2440 3392
rect 2124 3366 2188 3376
rect 2504 3380 2756 3392
rect 2440 3366 2504 3376
rect 2820 3382 3100 3392
rect 2756 3366 2820 3376
rect 1336 3332 1400 3342
rect 1652 3332 1716 3342
rect 1400 3316 1652 3326
rect 1968 3332 2032 3342
rect 1716 3316 1968 3326
rect 2284 3332 2348 3342
rect 2032 3324 2128 3326
rect 2032 3316 2284 3324
rect 2128 3152 2284 3316
rect 2600 3332 2664 3342
rect 2348 3152 2600 3324
rect 2916 3332 2980 3342
rect 2664 3152 2916 3324
rect 1336 3072 1348 3152
rect 2128 3072 2980 3152
rect 1336 3056 2980 3072
rect 2244 3012 3100 3014
rect 1492 3004 3100 3012
rect 1492 2920 2244 3004
rect 1556 2744 1808 2920
rect 1492 2730 1556 2740
rect 1872 2744 2124 2920
rect 1808 2730 1872 2740
rect 2188 2760 2244 2920
rect 2188 2744 2440 2760
rect 2124 2730 2188 2740
rect 2504 2744 2756 2760
rect 2440 2730 2504 2740
rect 2820 2750 3100 2760
rect 2756 2730 2820 2740
rect 1336 2696 1400 2706
rect 1652 2696 1716 2706
rect 1400 2680 1652 2690
rect 1968 2696 2032 2706
rect 1716 2680 1968 2690
rect 2284 2696 2348 2706
rect 2032 2688 2128 2690
rect 2032 2680 2284 2688
rect 2128 2516 2284 2680
rect 2600 2696 2664 2706
rect 2348 2516 2600 2688
rect 2916 2696 2980 2706
rect 2664 2516 2916 2688
rect 1336 2436 1348 2516
rect 2128 2436 2980 2516
rect 1336 2420 2980 2436
rect 2244 2372 3100 2378
rect 1492 2368 3100 2372
rect 1492 2280 2244 2368
rect 1556 2104 1808 2280
rect 1492 2090 1556 2100
rect 1872 2104 2124 2280
rect 1808 2090 1872 2100
rect 2188 2124 2244 2280
rect 2188 2104 2440 2124
rect 2124 2090 2188 2100
rect 2504 2104 2756 2124
rect 2440 2090 2504 2100
rect 2820 2114 3100 2124
rect 2756 2090 2820 2100
rect 1336 2056 1400 2066
rect 1652 2056 1716 2066
rect 1400 2040 1652 2052
rect 1968 2056 2032 2066
rect 1716 2040 1968 2052
rect 2284 2056 2348 2066
rect 2032 2040 2284 2052
rect 2128 1876 2284 2040
rect 2600 2056 2664 2066
rect 2348 1876 2600 2052
rect 2916 2056 2980 2066
rect 2664 1876 2916 2052
rect 1336 1796 1348 1876
rect 2128 1796 2980 1876
rect 1336 1784 2980 1796
rect 1352 1548 2136 1550
rect 1352 1540 2840 1548
rect 2136 1456 2840 1540
rect 2136 1292 2200 1456
rect 1352 1282 1432 1292
rect 1496 1280 1624 1292
rect 1432 1266 1496 1276
rect 1688 1280 1816 1292
rect 1624 1266 1688 1276
rect 1880 1280 2008 1292
rect 1816 1266 1880 1276
rect 2072 1280 2200 1292
rect 2008 1266 2072 1276
rect 2264 1280 2392 1456
rect 2200 1266 2264 1276
rect 2456 1280 2584 1456
rect 2392 1266 2456 1276
rect 2648 1280 2776 1456
rect 2584 1266 2648 1276
rect 2776 1266 2840 1276
rect 1336 1232 1400 1242
rect 1524 1232 1588 1242
rect 1400 1052 1524 1228
rect 1716 1232 1780 1242
rect 1588 1052 1716 1228
rect 1912 1232 1976 1242
rect 1780 1052 1912 1228
rect 2104 1232 2168 1242
rect 1976 1052 2104 1228
rect 2296 1232 2360 1242
rect 2168 1212 2296 1228
rect 2488 1232 2552 1242
rect 2360 1212 2488 1228
rect 2680 1232 2744 1242
rect 2552 1212 2680 1228
rect 2744 1212 3100 1222
rect 2168 1052 2248 1212
rect 1336 972 2248 1052
rect 1336 962 3100 972
rect 1336 960 2744 962
rect 1432 910 2840 912
rect 1352 900 2840 910
rect 2136 820 2840 900
rect 2136 652 2200 820
rect 1352 642 1432 652
rect 1496 642 1624 652
rect 1432 630 1496 640
rect 1688 642 1816 652
rect 1624 630 1688 640
rect 1880 642 2008 652
rect 1816 630 1880 640
rect 2072 644 2200 652
rect 2072 642 2136 644
rect 2008 630 2072 640
rect 2264 644 2392 820
rect 2200 630 2264 640
rect 2456 644 2584 820
rect 2392 630 2456 640
rect 2648 644 2776 820
rect 2584 630 2648 640
rect 2776 630 2840 640
rect 1336 596 1400 606
rect 1524 596 1588 606
rect 1400 416 1524 592
rect 1716 596 1780 606
rect 1588 416 1716 592
rect 1912 596 1976 606
rect 1780 416 1912 592
rect 2104 596 2168 606
rect 1976 416 2104 592
rect 2296 596 2360 606
rect 2168 580 2296 592
rect 2488 596 2552 606
rect 2360 580 2488 592
rect 2680 596 2744 606
rect 2552 580 2680 592
rect 2744 580 3100 590
rect 2168 416 2248 580
rect 1336 340 2248 416
rect 1336 330 3100 340
rect 1336 324 2744 330
<< via2 >>
rect 2244 3556 3100 3636
rect 2244 3392 2440 3556
rect 2440 3392 2504 3556
rect 2504 3392 2756 3556
rect 2756 3392 2820 3556
rect 2820 3392 3100 3556
rect 1348 3152 1400 3316
rect 1400 3152 1652 3316
rect 1652 3152 1716 3316
rect 1716 3152 1968 3316
rect 1968 3152 2032 3316
rect 2032 3152 2128 3316
rect 1348 3072 2128 3152
rect 2244 2920 3100 3004
rect 2244 2760 2440 2920
rect 2440 2760 2504 2920
rect 2504 2760 2756 2920
rect 2756 2760 2820 2920
rect 2820 2760 3100 2920
rect 1348 2516 1400 2680
rect 1400 2516 1652 2680
rect 1652 2516 1716 2680
rect 1716 2516 1968 2680
rect 1968 2516 2032 2680
rect 2032 2516 2128 2680
rect 1348 2436 2128 2516
rect 2244 2280 3100 2368
rect 2244 2124 2440 2280
rect 2440 2124 2504 2280
rect 2504 2124 2756 2280
rect 2756 2124 2820 2280
rect 2820 2124 3100 2280
rect 1348 1876 1400 2040
rect 1400 1876 1652 2040
rect 1652 1876 1716 2040
rect 1716 1876 1968 2040
rect 1968 1876 2032 2040
rect 2032 1876 2128 2040
rect 1348 1796 2128 1876
rect 1352 1456 2136 1540
rect 1352 1292 1432 1456
rect 1432 1292 1496 1456
rect 1496 1292 1624 1456
rect 1624 1292 1688 1456
rect 1688 1292 1816 1456
rect 1816 1292 1880 1456
rect 1880 1292 2008 1456
rect 2008 1292 2072 1456
rect 2072 1292 2136 1456
rect 2248 1052 2296 1212
rect 2296 1052 2360 1212
rect 2360 1052 2488 1212
rect 2488 1052 2552 1212
rect 2552 1052 2680 1212
rect 2680 1052 2744 1212
rect 2744 1052 3100 1212
rect 2248 972 3100 1052
rect 1352 820 2136 900
rect 1352 652 1432 820
rect 1432 652 1496 820
rect 1496 652 1624 820
rect 1624 652 1688 820
rect 1688 652 1816 820
rect 1816 652 1880 820
rect 1880 652 2008 820
rect 2008 652 2072 820
rect 2072 652 2136 820
rect 2248 416 2296 580
rect 2296 416 2360 580
rect 2360 416 2488 580
rect 2488 416 2552 580
rect 2552 416 2680 580
rect 2680 416 2744 580
rect 2744 416 3100 580
rect 2248 340 3100 416
<< metal3 >>
rect 2232 3636 3116 3776
rect 2232 3392 2244 3636
rect 3100 3392 3116 3636
rect 1336 3316 2148 3332
rect 1336 3072 1348 3316
rect 2128 3072 2148 3316
rect 1336 2680 2148 3072
rect 1336 2436 1348 2680
rect 2128 2436 2148 2680
rect 1336 2040 2148 2436
rect 2232 3004 3116 3392
rect 2232 2760 2244 3004
rect 3100 2760 3116 3004
rect 2232 2368 3116 2760
rect 2232 2124 2244 2368
rect 3100 2124 3116 2368
rect 2232 2108 3116 2124
rect 1336 1796 1348 2040
rect 2128 1796 2148 2040
rect 1336 1540 2148 1796
rect 1336 1292 1352 1540
rect 2136 1292 2148 1540
rect 1336 900 2148 1292
rect 1336 652 1352 900
rect 2136 652 2148 900
rect 1336 624 2148 652
rect 2232 1212 3116 1228
rect 2232 972 2248 1212
rect 3100 972 3116 1212
rect 2232 580 3116 972
rect 2232 340 2248 580
rect 3100 340 3116 580
rect 2232 208 3116 340
use sky130_fd_pr__pfet_01v8_QZVKPD  sky130_fd_pr__pfet_01v8_QZVKPD_1
timestamp 1683553987
transform 1 0 2157 0 1 2715
box -957 -1055 957 1055
use sky130_fd_pr__pfet_01v8_VC7ZFX  sky130_fd_pr__pfet_01v8_VC7ZFX_1
timestamp 1683553987
transform 1 0 2087 0 1 937
box -887 -737 887 737
<< end >>
