magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< metal1 >>
rect 4048 2200 4622 2208
rect 2480 2096 4622 2200
rect 2526 1876 2536 2056
rect 2592 1876 2602 2056
rect 2718 1876 2728 2056
rect 2784 1876 2794 2056
rect 2910 1876 2920 2056
rect 2976 1876 2986 2056
rect 3102 1876 3112 2056
rect 3168 1876 3178 2056
rect 3294 1876 3304 2056
rect 3360 1876 3370 2056
rect 3486 1876 3496 2056
rect 3552 1876 3562 2056
rect 3678 1876 3688 2056
rect 3744 1876 3754 2056
rect 3870 1876 3880 2056
rect 3936 1876 3946 2056
rect 4062 1876 4072 2056
rect 4128 1876 4138 2056
rect 4254 1876 4264 2056
rect 4320 1876 4330 2056
rect 2430 1652 2440 1832
rect 2496 1652 2506 1832
rect 2622 1652 2632 1832
rect 2688 1652 2698 1832
rect 2814 1652 2824 1832
rect 2880 1652 2890 1832
rect 3006 1652 3016 1832
rect 3072 1652 3082 1832
rect 3198 1652 3208 1832
rect 3264 1652 3274 1832
rect 3390 1652 3400 1832
rect 3456 1652 3466 1832
rect 3582 1652 3592 1832
rect 3648 1652 3658 1832
rect 3774 1652 3784 1832
rect 3840 1652 3850 1832
rect 3966 1652 3976 1832
rect 4032 1652 4042 1832
rect 4158 1652 4168 1832
rect 4224 1652 4234 1832
rect 4350 1652 4360 1832
rect 4416 1652 4426 1832
rect 4480 1616 4622 2096
rect 2576 1460 4622 1616
rect 2526 1244 2536 1424
rect 2592 1244 2602 1424
rect 2718 1244 2728 1424
rect 2784 1244 2794 1424
rect 2910 1244 2920 1424
rect 2976 1244 2986 1424
rect 3102 1244 3112 1424
rect 3168 1244 3178 1424
rect 3294 1244 3304 1424
rect 3360 1244 3370 1424
rect 3486 1244 3496 1424
rect 3552 1244 3562 1424
rect 3678 1244 3688 1424
rect 3744 1244 3754 1424
rect 3870 1244 3880 1424
rect 3936 1244 3946 1424
rect 4062 1244 4072 1424
rect 4128 1244 4138 1424
rect 4254 1244 4264 1424
rect 4320 1244 4330 1424
rect 2430 1020 2440 1200
rect 2496 1020 2506 1200
rect 2622 1020 2632 1200
rect 2688 1020 2698 1200
rect 2814 1020 2824 1200
rect 2880 1020 2890 1200
rect 3006 1020 3016 1200
rect 3072 1020 3082 1200
rect 3198 1020 3208 1200
rect 3264 1020 3274 1200
rect 3390 1020 3400 1200
rect 3456 1020 3466 1200
rect 3582 1020 3592 1200
rect 3648 1020 3658 1200
rect 3774 1020 3784 1200
rect 3840 1020 3850 1200
rect 3966 1020 3976 1200
rect 4032 1020 4042 1200
rect 4158 1020 4168 1200
rect 4224 1020 4234 1200
rect 4350 1020 4360 1200
rect 4416 1020 4426 1200
rect 4480 980 4622 1460
rect 2480 876 4622 980
rect 2476 500 4276 588
rect 2526 292 2536 472
rect 2592 292 2602 472
rect 2718 292 2728 472
rect 2784 292 2794 472
rect 2910 292 2920 472
rect 2976 292 2986 472
rect 3102 292 3112 472
rect 3168 292 3178 472
rect 3294 292 3304 472
rect 3360 292 3370 472
rect 3486 292 3496 472
rect 3552 292 3562 472
rect 3678 292 3688 472
rect 3744 292 3754 472
rect 3870 292 3880 472
rect 3936 292 3946 472
rect 4062 292 4072 472
rect 4128 292 4138 472
rect 4254 292 4264 472
rect 4320 292 4330 472
rect 2430 68 2440 248
rect 2496 68 2506 248
rect 2622 68 2632 248
rect 2688 68 2698 248
rect 2814 68 2824 248
rect 2880 68 2890 248
rect 3006 68 3016 248
rect 3072 68 3082 248
rect 3198 68 3208 248
rect 3264 68 3274 248
rect 3390 68 3400 248
rect 3456 68 3466 248
rect 3582 68 3592 248
rect 3648 68 3658 248
rect 3774 68 3784 248
rect 3840 68 3850 248
rect 3966 68 3976 248
rect 4032 68 4042 248
rect 4158 68 4168 248
rect 4224 68 4234 248
rect 4350 68 4360 248
rect 4412 68 4422 248
rect 2576 -120 4372 36
rect 2526 -328 2536 -148
rect 2592 -328 2602 -148
rect 2718 -328 2728 -148
rect 2784 -328 2794 -148
rect 2910 -328 2920 -148
rect 2976 -328 2986 -148
rect 3102 -328 3112 -148
rect 3168 -328 3178 -148
rect 3294 -328 3304 -148
rect 3360 -328 3370 -148
rect 3486 -328 3496 -148
rect 3552 -328 3562 -148
rect 3678 -328 3688 -148
rect 3744 -328 3754 -148
rect 3870 -328 3880 -148
rect 3936 -328 3946 -148
rect 4062 -328 4072 -148
rect 4128 -328 4138 -148
rect 4254 -328 4264 -148
rect 4320 -328 4330 -148
rect 2430 -552 2440 -372
rect 2496 -552 2506 -372
rect 2622 -552 2632 -372
rect 2688 -552 2698 -372
rect 2814 -552 2824 -372
rect 2880 -552 2890 -372
rect 3006 -552 3016 -372
rect 3072 -552 3082 -372
rect 3198 -552 3208 -372
rect 3264 -552 3274 -372
rect 3390 -552 3400 -372
rect 3456 -552 3466 -372
rect 3582 -552 3592 -372
rect 3648 -552 3658 -372
rect 3774 -552 3784 -372
rect 3840 -552 3850 -372
rect 3966 -552 3976 -372
rect 4032 -552 4042 -372
rect 4158 -552 4168 -372
rect 4224 -552 4234 -372
rect 4350 -552 4360 -372
rect 4412 -552 4422 -372
rect 2480 -656 4276 -580
rect 2716 -674 4276 -656
<< via1 >>
rect 2536 1876 2592 2056
rect 2728 1876 2784 2056
rect 2920 1876 2976 2056
rect 3112 1876 3168 2056
rect 3304 1876 3360 2056
rect 3496 1876 3552 2056
rect 3688 1876 3744 2056
rect 3880 1876 3936 2056
rect 4072 1876 4128 2056
rect 4264 1876 4320 2056
rect 2440 1652 2496 1832
rect 2632 1652 2688 1832
rect 2824 1652 2880 1832
rect 3016 1652 3072 1832
rect 3208 1652 3264 1832
rect 3400 1652 3456 1832
rect 3592 1652 3648 1832
rect 3784 1652 3840 1832
rect 3976 1652 4032 1832
rect 4168 1652 4224 1832
rect 4360 1652 4416 1832
rect 2536 1244 2592 1424
rect 2728 1244 2784 1424
rect 2920 1244 2976 1424
rect 3112 1244 3168 1424
rect 3304 1244 3360 1424
rect 3496 1244 3552 1424
rect 3688 1244 3744 1424
rect 3880 1244 3936 1424
rect 4072 1244 4128 1424
rect 4264 1244 4320 1424
rect 2440 1020 2496 1200
rect 2632 1020 2688 1200
rect 2824 1020 2880 1200
rect 3016 1020 3072 1200
rect 3208 1020 3264 1200
rect 3400 1020 3456 1200
rect 3592 1020 3648 1200
rect 3784 1020 3840 1200
rect 3976 1020 4032 1200
rect 4168 1020 4224 1200
rect 4360 1020 4416 1200
rect 2536 292 2592 472
rect 2728 292 2784 472
rect 2920 292 2976 472
rect 3112 292 3168 472
rect 3304 292 3360 472
rect 3496 292 3552 472
rect 3688 292 3744 472
rect 3880 292 3936 472
rect 4072 292 4128 472
rect 4264 292 4320 472
rect 2440 68 2496 248
rect 2632 68 2688 248
rect 2824 68 2880 248
rect 3016 68 3072 248
rect 3208 68 3264 248
rect 3400 68 3456 248
rect 3592 68 3648 248
rect 3784 68 3840 248
rect 3976 68 4032 248
rect 4168 68 4224 248
rect 4360 68 4412 248
rect 2536 -328 2592 -148
rect 2728 -328 2784 -148
rect 2920 -328 2976 -148
rect 3112 -328 3168 -148
rect 3304 -328 3360 -148
rect 3496 -328 3552 -148
rect 3688 -328 3744 -148
rect 3880 -328 3936 -148
rect 4072 -328 4128 -148
rect 4264 -328 4320 -148
rect 2440 -552 2496 -372
rect 2632 -552 2688 -372
rect 2824 -552 2880 -372
rect 3016 -552 3072 -372
rect 3208 -552 3264 -372
rect 3400 -552 3456 -372
rect 3592 -552 3648 -372
rect 3784 -552 3840 -372
rect 3976 -552 4032 -372
rect 4168 -552 4224 -372
rect 4360 -552 4412 -372
<< metal2 >>
rect 2532 2056 4524 2152
rect 2532 1880 2536 2056
rect 2592 1880 2728 2056
rect 2536 1866 2592 1876
rect 2784 1880 2920 2056
rect 2728 1866 2784 1876
rect 2976 1880 3112 2056
rect 2920 1866 2976 1876
rect 3168 1880 3304 2056
rect 3112 1866 3168 1876
rect 3360 1880 3496 2056
rect 3304 1866 3360 1876
rect 3552 1880 3688 2056
rect 3496 1866 3552 1876
rect 3744 1880 3880 2056
rect 3688 1866 3744 1876
rect 3936 1880 4072 2056
rect 3880 1866 3936 1876
rect 4128 1880 4264 2056
rect 4072 1866 4128 1876
rect 4320 1880 4524 2056
rect 4264 1866 4320 1876
rect 2440 1834 2496 1842
rect 2632 1834 2688 1842
rect 2824 1834 2880 1842
rect 3016 1834 3072 1842
rect 3208 1834 3264 1842
rect 3400 1834 3456 1842
rect 2436 1832 3456 1834
rect 2436 1652 2440 1832
rect 2496 1652 2632 1832
rect 2688 1652 2824 1832
rect 2880 1652 3016 1832
rect 3072 1652 3208 1832
rect 3264 1652 3400 1832
rect 3592 1832 3648 1842
rect 3456 1652 3592 1828
rect 3784 1832 3840 1842
rect 3648 1652 3784 1828
rect 3976 1832 4032 1842
rect 3840 1652 3976 1828
rect 4168 1832 4224 1842
rect 4032 1652 4168 1828
rect 4360 1832 4416 1842
rect 4224 1652 4360 1828
rect 4416 1652 4428 1828
rect 2436 1556 4428 1652
rect 2524 1424 4516 1520
rect 2524 1248 2536 1424
rect 2592 1248 2728 1424
rect 2536 1234 2592 1244
rect 2784 1248 2920 1424
rect 2728 1234 2784 1244
rect 2976 1248 3112 1424
rect 2920 1234 2976 1244
rect 3168 1248 3304 1424
rect 3112 1234 3168 1244
rect 3360 1248 3496 1424
rect 3304 1234 3360 1244
rect 3552 1248 3688 1424
rect 3496 1234 3552 1244
rect 3744 1248 3880 1424
rect 3688 1234 3744 1244
rect 3936 1248 4072 1424
rect 3880 1234 3936 1244
rect 4128 1248 4264 1424
rect 4072 1234 4128 1244
rect 4320 1248 4516 1424
rect 4264 1234 4320 1244
rect 2440 1202 2496 1210
rect 2632 1202 2688 1210
rect 2824 1202 2880 1210
rect 3016 1202 3072 1210
rect 3208 1202 3264 1210
rect 3400 1202 3456 1210
rect 2436 1200 3456 1202
rect 2436 1020 2440 1200
rect 2496 1020 2632 1200
rect 2688 1020 2824 1200
rect 2880 1020 3016 1200
rect 3072 1020 3208 1200
rect 3264 1020 3400 1200
rect 3592 1200 3648 1210
rect 3456 1020 3592 1196
rect 3784 1200 3840 1210
rect 3648 1020 3784 1196
rect 3976 1200 4032 1210
rect 3840 1020 3976 1196
rect 4168 1200 4224 1210
rect 4032 1020 4168 1196
rect 4360 1200 4416 1210
rect 4224 1020 4360 1196
rect 4416 1020 4428 1196
rect 2436 924 4428 1020
rect 2436 922 3412 924
rect 2532 472 4524 568
rect 2532 296 2536 472
rect 2592 296 2728 472
rect 2536 282 2592 292
rect 2784 296 2920 472
rect 2728 282 2784 292
rect 2976 296 3112 472
rect 2920 282 2976 292
rect 3168 296 3304 472
rect 3112 282 3168 292
rect 3360 296 3496 472
rect 3304 282 3360 292
rect 3552 296 3688 472
rect 3496 282 3552 292
rect 3744 296 3880 472
rect 3688 282 3744 292
rect 3936 296 4072 472
rect 3880 282 3936 292
rect 4128 296 4264 472
rect 4072 282 4128 292
rect 4320 296 4524 472
rect 4264 282 4320 292
rect 2440 254 2496 258
rect 2632 254 2688 258
rect 2824 254 2880 258
rect 3016 254 3072 258
rect 3208 254 3264 258
rect 3400 254 3456 258
rect 2428 248 3456 254
rect 2428 244 2440 248
rect 2400 68 2440 244
rect 2496 68 2632 248
rect 2688 68 2824 248
rect 2880 68 3016 248
rect 3072 68 3208 248
rect 3264 68 3400 248
rect 3592 248 3648 258
rect 3456 68 3592 244
rect 3784 248 3840 258
rect 3648 68 3784 244
rect 3976 248 4032 258
rect 3840 68 3976 244
rect 4168 248 4224 258
rect 4032 68 4168 244
rect 4360 248 4416 258
rect 4224 68 4360 244
rect 4412 68 4416 248
rect 2400 -16 4416 68
rect 2400 -370 2500 -16
rect 2532 -148 4524 -52
rect 2532 -324 2536 -148
rect 2592 -324 2728 -148
rect 2536 -338 2592 -328
rect 2784 -324 2920 -148
rect 2728 -338 2784 -328
rect 2976 -324 3112 -148
rect 2920 -338 2976 -328
rect 3168 -324 3304 -148
rect 3112 -338 3168 -328
rect 3360 -324 3496 -148
rect 3304 -338 3360 -328
rect 3552 -324 3688 -148
rect 3496 -338 3552 -328
rect 3744 -324 3880 -148
rect 3688 -338 3744 -328
rect 3936 -324 4072 -148
rect 3880 -338 3936 -328
rect 4128 -324 4264 -148
rect 4072 -338 4128 -328
rect 4320 -324 4524 -148
rect 4264 -338 4320 -328
rect 2632 -370 2688 -362
rect 2824 -370 2880 -362
rect 3016 -370 3072 -362
rect 3208 -370 3264 -362
rect 3400 -370 3456 -362
rect 2400 -372 3456 -370
rect 3592 -372 3648 -362
rect 3784 -372 3840 -362
rect 3976 -372 4032 -362
rect 4168 -372 4224 -362
rect 4360 -372 4416 -362
rect 2400 -552 2440 -372
rect 2496 -552 2632 -372
rect 2688 -552 2824 -372
rect 2880 -552 3016 -372
rect 3072 -552 3208 -372
rect 3264 -552 3400 -372
rect 3456 -552 3592 -372
rect 3648 -552 3784 -372
rect 3840 -552 3976 -372
rect 4032 -552 4168 -372
rect 4224 -552 4360 -372
rect 4412 -552 4420 -372
rect 2400 -644 4420 -552
rect 2460 -656 2688 -644
use sky130_fd_pr__nfet_01v8_lvt_A46MKJ  sky130_fd_pr__nfet_01v8_lvt_A46MKJ_0
timestamp 1686659968
transform 1 0 3427 0 1 -41
box -1127 -719 1127 719
use sky130_fd_pr__pfet_01v8_8DBWZL  sky130_fd_pr__pfet_01v8_8DBWZL_0
timestamp 1686659968
transform 1 0 3427 0 1 1537
box -1127 -737 1127 737
<< end >>
