magic
tech sky130A
magscale 1 2
timestamp 1689775068
<< error_p >>
rect 13418 29256 13434 29260
rect 145578 29256 145594 29260
rect 13198 29253 13418 29256
rect 145358 29253 145578 29256
rect 675 28987 691 29215
rect 132835 28996 132842 29220
rect 691 28984 702 28987
rect 132842 28984 132862 28996
rect 13138 22004 13158 22016
rect 145298 22013 145309 22016
rect 13158 21780 13165 22004
rect 145309 21785 145325 22013
rect 422 21744 642 21747
rect 132582 21744 132802 21747
rect 406 21740 422 21744
rect 132566 21740 132582 21744
rect 13418 9256 13434 9260
rect 145578 9256 145594 9260
rect 13198 9253 13418 9256
rect 145358 9253 145578 9256
rect 675 8987 691 9215
rect 132835 8996 132842 9220
rect 691 8984 702 8987
rect 132842 8984 132862 8996
rect 13138 2004 13158 2016
rect 145298 2013 145309 2016
rect 13158 1780 13165 2004
rect 145309 1785 145325 2013
rect 422 1744 642 1747
rect 132582 1744 132802 1747
rect 406 1740 422 1744
rect 132566 1740 132582 1744
rect 13418 -10744 13434 -10740
rect 145578 -10744 145594 -10740
rect 13198 -10747 13418 -10744
rect 145358 -10747 145578 -10744
rect 675 -11013 691 -10785
rect 132835 -11004 132842 -10780
rect 691 -11016 702 -11013
rect 132842 -11016 132862 -11004
rect 13138 -17996 13158 -17984
rect 145298 -17987 145309 -17984
rect 13158 -18220 13165 -17996
rect 145309 -18215 145325 -17987
rect 422 -18256 642 -18253
rect 132582 -18256 132802 -18253
rect 406 -18260 422 -18256
rect 132566 -18260 132582 -18256
rect 13418 -30744 13434 -30740
rect 145578 -30744 145594 -30740
rect 13198 -30747 13418 -30744
rect 145358 -30747 145578 -30744
rect 675 -31013 691 -30785
rect 132835 -31004 132842 -30780
rect 691 -31016 702 -31013
rect 132842 -31016 132862 -31004
rect 13138 -37996 13158 -37984
rect 145298 -37987 145309 -37984
rect 13158 -38220 13165 -37996
rect 145309 -38215 145325 -37987
rect 422 -38256 642 -38253
rect 132582 -38256 132802 -38253
rect 406 -38260 422 -38256
rect 132566 -38260 132582 -38256
rect 13418 -50744 13434 -50740
rect 145578 -50744 145594 -50740
rect 13198 -50747 13418 -50744
rect 145358 -50747 145578 -50744
rect 675 -51013 691 -50785
rect 132835 -51004 132842 -50780
rect 691 -51016 702 -51013
rect 132842 -51016 132862 -51004
rect 13418 -70744 13434 -70740
rect 145578 -70744 145594 -70740
rect 13198 -70747 13418 -70744
rect 145358 -70747 145578 -70744
rect 675 -71013 691 -70785
rect 132835 -71004 132842 -70780
rect 691 -71016 702 -71013
rect 132842 -71016 132862 -71004
rect 13138 -77996 13158 -77984
rect 145298 -77987 145309 -77984
rect 13158 -78220 13165 -77996
rect 145309 -78215 145325 -77987
rect 422 -78256 642 -78253
rect 132582 -78256 132802 -78253
rect 406 -78260 422 -78256
rect 132566 -78260 132582 -78256
rect 13418 -90744 13434 -90740
rect 145578 -90744 145594 -90740
rect 13198 -90747 13418 -90744
rect 145358 -90747 145578 -90744
rect 675 -91013 691 -90785
rect 132835 -91004 132842 -90780
rect 691 -91016 702 -91013
rect 132842 -91016 132862 -91004
rect 13138 -97996 13158 -97984
rect 145298 -97987 145309 -97984
rect 13158 -98220 13165 -97996
rect 145309 -98215 145325 -97987
rect 422 -98256 642 -98253
rect 132582 -98256 132802 -98253
rect 406 -98260 422 -98256
rect 132566 -98260 132582 -98256
rect 13418 -110744 13434 -110740
rect 145578 -110744 145594 -110740
rect 13198 -110747 13418 -110744
rect 145358 -110747 145578 -110744
rect 675 -111013 691 -110785
rect 132835 -111004 132842 -110780
rect 691 -111016 702 -111013
rect 132842 -111016 132862 -111004
rect 13138 -117996 13158 -117984
rect 145298 -117987 145309 -117984
rect 13158 -118220 13165 -117996
rect 145309 -118215 145325 -117987
rect 422 -118256 642 -118253
rect 132582 -118256 132802 -118253
rect 406 -118260 422 -118256
rect 132566 -118260 132582 -118256
rect 13418 -130744 13434 -130740
rect 145578 -130744 145594 -130740
rect 13198 -130747 13418 -130744
rect 145358 -130747 145578 -130744
rect 675 -131013 691 -130785
rect 132835 -131004 132842 -130780
rect 691 -131016 702 -131013
rect 132842 -131016 132862 -131004
rect 13138 -137996 13158 -137984
rect 145298 -137987 145309 -137984
rect 13158 -138220 13165 -137996
rect 145309 -138215 145325 -137987
rect 422 -138256 642 -138253
rect 132582 -138256 132802 -138253
rect 406 -138260 422 -138256
rect 132566 -138260 132582 -138256
rect 13418 -150744 13434 -150740
rect 145578 -150744 145594 -150740
rect 13198 -150747 13418 -150744
rect 145358 -150747 145578 -150744
rect 675 -151013 691 -150785
rect 132835 -151004 132842 -150780
rect 691 -151016 702 -151013
rect 132842 -151016 132862 -151004
rect 13418 -170744 13434 -170740
rect 145578 -170744 145594 -170740
rect 13198 -170747 13418 -170744
rect 145358 -170747 145578 -170744
rect 675 -171013 691 -170785
rect 132835 -171004 132842 -170780
rect 691 -171016 702 -171013
rect 132842 -171016 132862 -171004
rect 13138 -177996 13158 -177984
rect 145298 -177987 145309 -177984
rect 13158 -178220 13165 -177996
rect 145309 -178215 145325 -177987
rect 422 -178256 642 -178253
rect 132582 -178256 132802 -178253
rect 406 -178260 422 -178256
rect 132566 -178260 132582 -178256
rect 13418 -190744 13434 -190740
rect 145578 -190744 145594 -190740
rect 13198 -190747 13418 -190744
rect 145358 -190747 145578 -190744
rect 675 -191013 691 -190785
rect 132835 -191004 132842 -190780
rect 691 -191016 702 -191013
rect 132842 -191016 132862 -191004
rect 13138 -197996 13158 -197984
rect 145298 -197987 145309 -197984
rect 13158 -198220 13165 -197996
rect 145309 -198215 145325 -197987
rect 422 -198256 642 -198253
rect 132582 -198256 132802 -198253
rect 406 -198260 422 -198256
rect 132566 -198260 132582 -198256
rect 13418 -210744 13434 -210740
rect 145578 -210744 145594 -210740
rect 13198 -210747 13418 -210744
rect 145358 -210747 145578 -210744
rect 675 -211013 691 -210785
rect 132835 -211004 132842 -210780
rect 691 -211016 702 -211013
rect 132842 -211016 132862 -211004
rect 13138 -217996 13158 -217984
rect 145298 -217987 145309 -217984
rect 13158 -218220 13165 -217996
rect 145309 -218215 145325 -217987
rect 422 -218256 642 -218253
rect 132582 -218256 132802 -218253
rect 406 -218260 422 -218256
rect 132566 -218260 132582 -218256
rect 13418 -230744 13434 -230740
rect 145578 -230744 145594 -230740
rect 13198 -230747 13418 -230744
rect 145358 -230747 145578 -230744
rect 675 -231013 691 -230785
rect 132835 -231004 132842 -230780
rect 691 -231016 702 -231013
rect 132842 -231016 132862 -231004
rect 13138 -237996 13158 -237984
rect 145298 -237987 145309 -237984
rect 13158 -238220 13165 -237996
rect 145309 -238215 145325 -237987
rect 422 -238256 642 -238253
rect 132582 -238256 132802 -238253
rect 406 -238260 422 -238256
rect 132566 -238260 132582 -238256
rect 13418 -250744 13434 -250740
rect 145578 -250744 145594 -250740
rect 13198 -250747 13418 -250744
rect 145358 -250747 145578 -250744
rect 675 -251013 691 -250785
rect 132835 -251004 132842 -250780
rect 691 -251016 702 -251013
rect 132842 -251016 132862 -251004
rect 13418 -270744 13434 -270740
rect 145578 -270744 145594 -270740
rect 13198 -270747 13418 -270744
rect 145358 -270747 145578 -270744
rect 675 -271013 691 -270785
rect 132835 -271004 132842 -270780
rect 691 -271016 702 -271013
rect 132842 -271016 132862 -271004
rect 13138 -277996 13158 -277984
rect 145298 -277987 145309 -277984
rect 13158 -278220 13165 -277996
rect 145309 -278215 145325 -277987
rect 422 -278256 642 -278253
rect 132582 -278256 132802 -278253
rect 406 -278260 422 -278256
rect 132566 -278260 132582 -278256
rect 13418 -290744 13434 -290740
rect 145578 -290744 145594 -290740
rect 13198 -290747 13418 -290744
rect 145358 -290747 145578 -290744
rect 675 -291013 691 -290785
rect 132835 -291004 132842 -290780
rect 691 -291016 702 -291013
rect 132842 -291016 132862 -291004
rect 13138 -297996 13158 -297984
rect 145298 -297987 145309 -297984
rect 13158 -298220 13165 -297996
rect 145309 -298215 145325 -297987
rect 422 -298256 642 -298253
rect 132582 -298256 132802 -298253
rect 406 -298260 422 -298256
rect 132566 -298260 132582 -298256
rect 13418 -310744 13434 -310740
rect 145578 -310744 145594 -310740
rect 13198 -310747 13418 -310744
rect 145358 -310747 145578 -310744
rect 675 -311013 691 -310785
rect 132835 -311004 132842 -310780
rect 691 -311016 702 -311013
rect 132842 -311016 132862 -311004
rect 13138 -317996 13158 -317984
rect 145298 -317987 145309 -317984
rect 13158 -318220 13165 -317996
rect 145309 -318215 145325 -317987
rect 422 -318256 642 -318253
rect 132582 -318256 132802 -318253
rect 406 -318260 422 -318256
rect 132566 -318260 132582 -318256
rect 13418 -330744 13434 -330740
rect 145578 -330744 145594 -330740
rect 13198 -330747 13418 -330744
rect 145358 -330747 145578 -330744
rect 675 -331013 691 -330785
rect 132835 -331004 132842 -330780
rect 691 -331016 702 -331013
rect 132842 -331016 132862 -331004
rect 13138 -337996 13158 -337984
rect 145298 -337987 145309 -337984
rect 13158 -338220 13165 -337996
rect 145309 -338215 145325 -337987
rect 422 -338256 642 -338253
rect 132582 -338256 132802 -338253
rect 406 -338260 422 -338256
rect 132566 -338260 132582 -338256
rect 13418 -350744 13434 -350740
rect 145578 -350744 145594 -350740
rect 13198 -350747 13418 -350744
rect 145358 -350747 145578 -350744
rect 675 -351013 691 -350785
rect 132835 -351004 132842 -350780
rect 691 -351016 702 -351013
rect 132842 -351016 132862 -351004
rect 13418 -370744 13434 -370740
rect 145578 -370744 145594 -370740
rect 13198 -370747 13418 -370744
rect 145358 -370747 145578 -370744
rect 675 -371013 691 -370785
rect 132835 -371004 132842 -370780
rect 691 -371016 702 -371013
rect 132842 -371016 132862 -371004
rect 13138 -377996 13158 -377984
rect 145298 -377987 145309 -377984
rect 13158 -378220 13165 -377996
rect 145309 -378215 145325 -377987
rect 422 -378256 642 -378253
rect 132582 -378256 132802 -378253
rect 406 -378260 422 -378256
rect 132566 -378260 132582 -378256
rect 13418 -390744 13434 -390740
rect 145578 -390744 145594 -390740
rect 13198 -390747 13418 -390744
rect 145358 -390747 145578 -390744
rect 675 -391013 691 -390785
rect 132835 -391004 132842 -390780
rect 691 -391016 702 -391013
rect 132842 -391016 132862 -391004
rect 13138 -397996 13158 -397984
rect 145298 -397987 145309 -397984
rect 13158 -398220 13165 -397996
rect 145309 -398215 145325 -397987
rect 422 -398256 642 -398253
rect 132582 -398256 132802 -398253
rect 406 -398260 422 -398256
rect 132566 -398260 132582 -398256
rect 13418 -410744 13434 -410740
rect 145578 -410744 145594 -410740
rect 13198 -410747 13418 -410744
rect 145358 -410747 145578 -410744
rect 675 -411013 691 -410785
rect 132835 -411004 132842 -410780
rect 691 -411016 702 -411013
rect 132842 -411016 132862 -411004
rect 13138 -417996 13158 -417984
rect 145298 -417987 145309 -417984
rect 13158 -418220 13165 -417996
rect 145309 -418215 145325 -417987
rect 422 -418256 642 -418253
rect 132582 -418256 132802 -418253
rect 406 -418260 422 -418256
rect 132566 -418260 132582 -418256
rect 13418 -430744 13434 -430740
rect 145578 -430744 145594 -430740
rect 13198 -430747 13418 -430744
rect 145358 -430747 145578 -430744
rect 675 -431013 691 -430785
rect 132835 -431004 132842 -430780
rect 691 -431016 702 -431013
rect 132842 -431016 132862 -431004
rect 13138 -437996 13158 -437984
rect 145298 -437987 145309 -437984
rect 13158 -438220 13165 -437996
rect 145309 -438215 145325 -437987
rect 422 -438256 642 -438253
rect 132582 -438256 132802 -438253
rect 406 -438260 422 -438256
rect 132566 -438260 132582 -438256
rect 13418 -450744 13434 -450740
rect 145578 -450744 145594 -450740
rect 13198 -450747 13418 -450744
rect 145358 -450747 145578 -450744
rect 675 -451013 691 -450785
rect 132835 -451004 132842 -450780
rect 691 -451016 702 -451013
rect 132842 -451016 132862 -451004
rect 13418 -470744 13434 -470740
rect 145578 -470744 145594 -470740
rect 13198 -470747 13418 -470744
rect 145358 -470747 145578 -470744
rect 675 -471013 691 -470785
rect 132835 -471004 132842 -470780
rect 691 -471016 702 -471013
rect 132842 -471016 132862 -471004
rect 13138 -477996 13158 -477984
rect 145298 -477987 145309 -477984
rect 13158 -478220 13165 -477996
rect 145309 -478215 145325 -477987
rect 422 -478256 642 -478253
rect 132582 -478256 132802 -478253
rect 406 -478260 422 -478256
rect 132566 -478260 132582 -478256
rect 13418 -490744 13434 -490740
rect 145578 -490744 145594 -490740
rect 13198 -490747 13418 -490744
rect 145358 -490747 145578 -490744
rect 675 -491013 691 -490785
rect 132835 -491004 132842 -490780
rect 691 -491016 702 -491013
rect 132842 -491016 132862 -491004
rect 13138 -497996 13158 -497984
rect 145298 -497987 145309 -497984
rect 13158 -498220 13165 -497996
rect 145309 -498215 145325 -497987
rect 422 -498256 642 -498253
rect 132582 -498256 132802 -498253
rect 406 -498260 422 -498256
rect 132566 -498260 132582 -498256
rect 13418 -510744 13434 -510740
rect 145578 -510744 145594 -510740
rect 13198 -510747 13418 -510744
rect 145358 -510747 145578 -510744
rect 675 -511013 691 -510785
rect 132835 -511004 132842 -510780
rect 691 -511016 702 -511013
rect 132842 -511016 132862 -511004
rect 13138 -517996 13158 -517984
rect 145298 -517987 145309 -517984
rect 13158 -518220 13165 -517996
rect 145309 -518215 145325 -517987
rect 422 -518256 642 -518253
rect 132582 -518256 132802 -518253
rect 406 -518260 422 -518256
rect 132566 -518260 132582 -518256
rect 13418 -530744 13434 -530740
rect 145578 -530744 145594 -530740
rect 13198 -530747 13418 -530744
rect 145358 -530747 145578 -530744
rect 675 -531013 691 -530785
rect 132835 -531004 132842 -530780
rect 691 -531016 702 -531013
rect 132842 -531016 132862 -531004
rect 13138 -537996 13158 -537984
rect 145298 -537987 145309 -537984
rect 13158 -538220 13165 -537996
rect 145309 -538215 145325 -537987
rect 422 -538256 642 -538253
rect 132582 -538256 132802 -538253
rect 406 -538260 422 -538256
rect 132566 -538260 132582 -538256
rect 13418 -550744 13434 -550740
rect 145578 -550744 145594 -550740
rect 13198 -550747 13418 -550744
rect 145358 -550747 145578 -550744
rect 675 -551013 691 -550785
rect 132835 -551004 132842 -550780
rect 691 -551016 702 -551013
rect 132842 -551016 132862 -551004
rect 13418 -570744 13434 -570740
rect 145578 -570744 145594 -570740
rect 13198 -570747 13418 -570744
rect 145358 -570747 145578 -570744
rect 675 -571013 691 -570785
rect 132835 -571004 132842 -570780
rect 691 -571016 702 -571013
rect 132842 -571016 132862 -571004
rect 13138 -577996 13158 -577984
rect 145298 -577987 145309 -577984
rect 13158 -578220 13165 -577996
rect 145309 -578215 145325 -577987
rect 422 -578256 642 -578253
rect 132582 -578256 132802 -578253
rect 406 -578260 422 -578256
rect 132566 -578260 132582 -578256
rect 13418 -590744 13434 -590740
rect 145578 -590744 145594 -590740
rect 13198 -590747 13418 -590744
rect 145358 -590747 145578 -590744
rect 675 -591013 691 -590785
rect 132835 -591004 132842 -590780
rect 691 -591016 702 -591013
rect 132842 -591016 132862 -591004
rect 13138 -597996 13158 -597984
rect 145298 -597987 145309 -597984
rect 13158 -598220 13165 -597996
rect 145309 -598215 145325 -597987
rect 422 -598256 642 -598253
rect 132582 -598256 132802 -598253
rect 406 -598260 422 -598256
rect 132566 -598260 132582 -598256
rect 13418 -610744 13434 -610740
rect 145578 -610744 145594 -610740
rect 13198 -610747 13418 -610744
rect 145358 -610747 145578 -610744
rect 675 -611013 691 -610785
rect 132835 -611004 132842 -610780
rect 691 -611016 702 -611013
rect 132842 -611016 132862 -611004
rect 13138 -617996 13158 -617984
rect 145298 -617987 145309 -617984
rect 13158 -618220 13165 -617996
rect 145309 -618215 145325 -617987
rect 422 -618256 642 -618253
rect 132582 -618256 132802 -618253
rect 406 -618260 422 -618256
rect 132566 -618260 132582 -618256
rect 13418 -630744 13434 -630740
rect 145578 -630744 145594 -630740
rect 13198 -630747 13418 -630744
rect 145358 -630747 145578 -630744
rect 675 -631013 691 -630785
rect 132835 -631004 132842 -630780
rect 691 -631016 702 -631013
rect 132842 -631016 132862 -631004
rect 13138 -637996 13158 -637984
rect 145298 -637987 145309 -637984
rect 13158 -638220 13165 -637996
rect 145309 -638215 145325 -637987
rect 422 -638256 642 -638253
rect 132582 -638256 132802 -638253
rect 406 -638260 422 -638256
rect 132566 -638260 132582 -638256
rect 13418 -650744 13434 -650740
rect 145578 -650744 145594 -650740
rect 13198 -650747 13418 -650744
rect 145358 -650747 145578 -650744
rect 675 -651013 691 -650785
rect 132835 -651004 132842 -650780
rect 691 -651016 702 -651013
rect 132842 -651016 132862 -651004
rect 13418 -670744 13434 -670740
rect 145578 -670744 145594 -670740
rect 13198 -670747 13418 -670744
rect 145358 -670747 145578 -670744
rect 675 -671013 691 -670785
rect 132835 -671004 132842 -670780
rect 691 -671016 702 -671013
rect 132842 -671016 132862 -671004
rect 13138 -677996 13158 -677984
rect 145298 -677987 145309 -677984
rect 13158 -678220 13165 -677996
rect 145309 -678215 145325 -677987
rect 422 -678256 642 -678253
rect 132582 -678256 132802 -678253
rect 406 -678260 422 -678256
rect 132566 -678260 132582 -678256
rect 13418 -690744 13434 -690740
rect 145578 -690744 145594 -690740
rect 13198 -690747 13418 -690744
rect 145358 -690747 145578 -690744
rect 675 -691013 691 -690785
rect 132835 -691004 132842 -690780
rect 691 -691016 702 -691013
rect 132842 -691016 132862 -691004
rect 13138 -697996 13158 -697984
rect 145298 -697987 145309 -697984
rect 13158 -698220 13165 -697996
rect 145309 -698215 145325 -697987
rect 422 -698256 642 -698253
rect 132582 -698256 132802 -698253
rect 406 -698260 422 -698256
rect 132566 -698260 132582 -698256
rect 13418 -710744 13434 -710740
rect 145578 -710744 145594 -710740
rect 13198 -710747 13418 -710744
rect 145358 -710747 145578 -710744
rect 675 -711013 691 -710785
rect 132835 -711004 132842 -710780
rect 691 -711016 702 -711013
rect 132842 -711016 132862 -711004
rect 13138 -717996 13158 -717984
rect 145298 -717987 145309 -717984
rect 13158 -718220 13165 -717996
rect 145309 -718215 145325 -717987
rect 422 -718256 642 -718253
rect 132582 -718256 132802 -718253
rect 406 -718260 422 -718256
rect 132566 -718260 132582 -718256
rect 13418 -730744 13434 -730740
rect 145578 -730744 145594 -730740
rect 13198 -730747 13418 -730744
rect 145358 -730747 145578 -730744
rect 675 -731013 691 -730785
rect 132835 -731004 132842 -730780
rect 691 -731016 702 -731013
rect 132842 -731016 132862 -731004
rect 13138 -737996 13158 -737984
rect 145298 -737987 145309 -737984
rect 13158 -738220 13165 -737996
rect 145309 -738215 145325 -737987
rect 422 -738256 642 -738253
rect 132582 -738256 132802 -738253
rect 406 -738260 422 -738256
rect 132566 -738260 132582 -738256
rect 13418 -750744 13434 -750740
rect 145578 -750744 145594 -750740
rect 13198 -750747 13418 -750744
rect 145358 -750747 145578 -750744
rect 675 -751013 691 -750785
rect 132835 -751004 132842 -750780
rect 691 -751016 702 -751013
rect 132842 -751016 132862 -751004
rect 13418 -770744 13434 -770740
rect 145578 -770744 145594 -770740
rect 13198 -770747 13418 -770744
rect 145358 -770747 145578 -770744
rect 675 -771013 691 -770785
rect 132835 -771004 132842 -770780
rect 691 -771016 702 -771013
rect 132842 -771016 132862 -771004
rect 13138 -777996 13158 -777984
rect 145298 -777987 145309 -777984
rect 13158 -778220 13165 -777996
rect 145309 -778215 145325 -777987
rect 422 -778256 642 -778253
rect 132582 -778256 132802 -778253
rect 406 -778260 422 -778256
rect 132566 -778260 132582 -778256
rect 13418 -790744 13434 -790740
rect 145578 -790744 145594 -790740
rect 13198 -790747 13418 -790744
rect 145358 -790747 145578 -790744
rect 675 -791013 691 -790785
rect 132835 -791004 132842 -790780
rect 691 -791016 702 -791013
rect 132842 -791016 132862 -791004
rect 13138 -797996 13158 -797984
rect 145298 -797987 145309 -797984
rect 13158 -798220 13165 -797996
rect 145309 -798215 145325 -797987
rect 422 -798256 642 -798253
rect 132582 -798256 132802 -798253
rect 406 -798260 422 -798256
rect 132566 -798260 132582 -798256
rect 13418 -810744 13434 -810740
rect 145578 -810744 145594 -810740
rect 13198 -810747 13418 -810744
rect 145358 -810747 145578 -810744
rect 675 -811013 691 -810785
rect 132835 -811004 132842 -810780
rect 691 -811016 702 -811013
rect 132842 -811016 132862 -811004
rect 13138 -817996 13158 -817984
rect 145298 -817987 145309 -817984
rect 13158 -818220 13165 -817996
rect 145309 -818215 145325 -817987
rect 422 -818256 642 -818253
rect 132582 -818256 132802 -818253
rect 406 -818260 422 -818256
rect 132566 -818260 132582 -818256
rect 13418 -830744 13434 -830740
rect 145578 -830744 145594 -830740
rect 13198 -830747 13418 -830744
rect 145358 -830747 145578 -830744
rect 675 -831013 691 -830785
rect 132835 -831004 132842 -830780
rect 691 -831016 702 -831013
rect 132842 -831016 132862 -831004
rect 13138 -837996 13158 -837984
rect 145298 -837987 145309 -837984
rect 13158 -838220 13165 -837996
rect 145309 -838215 145325 -837987
rect 422 -838256 642 -838253
rect 132582 -838256 132802 -838253
rect 406 -838260 422 -838256
rect 132566 -838260 132582 -838256
rect 13418 -850744 13434 -850740
rect 145578 -850744 145594 -850740
rect 13198 -850747 13418 -850744
rect 145358 -850747 145578 -850744
rect 675 -851013 691 -850785
rect 132835 -851004 132842 -850780
rect 691 -851016 702 -851013
rect 132842 -851016 132862 -851004
<< error_s >>
rect 47740 77378 47744 77394
rect 68740 77378 68744 77394
rect 89740 77380 89742 77394
rect 89742 77378 89744 77380
rect 110740 77378 110744 77394
rect 47744 77158 47747 77378
rect 68744 77158 68747 77378
rect 89744 77337 89747 77378
rect 110744 77158 110747 77378
rect 34987 77109 35215 77125
rect 55987 77109 56215 77125
rect 76987 77109 77215 77125
rect 97987 77109 98215 77125
rect 34984 77098 34987 77109
rect 55984 77098 55987 77109
rect 76984 77098 76987 77109
rect 97984 77098 97987 77109
rect 48004 64642 48016 64662
rect 69004 64642 69016 64662
rect 90004 64642 90016 64662
rect 111004 64642 111016 64662
rect 47780 64635 48004 64642
rect 68780 64635 69004 64642
rect 89780 64635 90004 64642
rect 110780 64635 111004 64642
rect 35253 64382 35256 64390
rect 56253 64382 56256 64390
rect 77253 64382 77256 64390
rect 98253 64382 98256 64390
rect 35256 64366 35260 64382
rect 56256 64366 56260 64382
rect 77256 64366 77260 64382
rect 98256 64366 98260 64382
rect 30178 52413 30180 52497
rect 30262 52372 30264 52413
rect 115820 52372 115822 52497
rect 13138 42004 13158 42016
rect 145298 42013 145309 42016
rect 13158 41780 13165 42004
rect 145309 41785 145325 42013
rect 422 41744 642 41747
rect 132582 41744 132802 41747
rect 406 41740 422 41744
rect 132566 41740 132582 41744
rect 13138 -57996 13158 -57984
rect 145298 -57987 145309 -57984
rect 13158 -58220 13165 -57996
rect 145309 -58215 145325 -57987
rect 422 -58256 642 -58253
rect 132582 -58256 132802 -58253
rect 406 -58260 422 -58256
rect 132566 -58260 132582 -58256
rect 13138 -157996 13158 -157984
rect 145298 -157987 145309 -157984
rect 13158 -158220 13165 -157996
rect 145309 -158215 145325 -157987
rect 422 -158256 642 -158253
rect 132582 -158256 132802 -158253
rect 406 -158260 422 -158256
rect 132566 -158260 132582 -158256
rect 13138 -257996 13158 -257984
rect 145298 -257987 145309 -257984
rect 13158 -258220 13165 -257996
rect 145309 -258215 145325 -257987
rect 422 -258256 642 -258253
rect 132582 -258256 132802 -258253
rect 406 -258260 422 -258256
rect 132566 -258260 132582 -258256
rect 13138 -357996 13158 -357984
rect 145298 -357987 145309 -357984
rect 13158 -358220 13165 -357996
rect 145309 -358215 145325 -357987
rect 422 -358256 642 -358253
rect 132582 -358256 132802 -358253
rect 406 -358260 422 -358256
rect 132566 -358260 132582 -358256
rect 13138 -457996 13158 -457984
rect 145298 -457987 145309 -457984
rect 13158 -458220 13165 -457996
rect 145309 -458215 145325 -457987
rect 422 -458256 642 -458253
rect 132582 -458256 132802 -458253
rect 406 -458260 422 -458256
rect 132566 -458260 132582 -458256
rect 13138 -557996 13158 -557984
rect 145298 -557987 145309 -557984
rect 13158 -558220 13165 -557996
rect 145309 -558215 145325 -557987
rect 422 -558256 642 -558253
rect 132582 -558256 132802 -558253
rect 406 -558260 422 -558256
rect 132566 -558260 132582 -558256
rect 13138 -657996 13158 -657984
rect 145298 -657987 145309 -657984
rect 13158 -658220 13165 -657996
rect 145309 -658215 145325 -657987
rect 422 -658256 642 -658253
rect 132582 -658256 132802 -658253
rect 406 -658260 422 -658256
rect 132566 -658260 132582 -658256
rect 13138 -757996 13158 -757984
rect 145298 -757987 145309 -757984
rect 13158 -758220 13165 -757996
rect 145309 -758215 145325 -757987
rect 422 -758256 642 -758253
rect 132582 -758256 132802 -758253
rect 406 -758260 422 -758256
rect 132566 -758260 132582 -758256
rect 30262 -866413 30264 -866288
rect 115736 -866372 115738 -866288
rect 115820 -866413 115822 -866372
rect 47740 -878382 47744 -878366
rect 68740 -878382 68744 -878366
rect 89740 -878382 89744 -878366
rect 110740 -878382 110744 -878366
rect 47744 -878390 47747 -878382
rect 68744 -878390 68747 -878382
rect 89744 -878390 89747 -878382
rect 110744 -878390 110747 -878382
rect 34996 -878642 35220 -878635
rect 55996 -878642 56220 -878635
rect 76996 -878642 77220 -878635
rect 97996 -878642 98220 -878635
rect 34984 -878662 34996 -878642
rect 55984 -878662 55996 -878642
rect 76984 -878662 76996 -878642
rect 97984 -878662 97996 -878642
rect 48013 -891109 48016 -891098
rect 69013 -891109 69016 -891098
rect 90013 -891109 90016 -891098
rect 111013 -891109 111016 -891098
rect 47785 -891125 48013 -891109
rect 68785 -891125 69013 -891109
rect 89785 -891125 90013 -891109
rect 110785 -891125 111013 -891109
rect 35253 -891378 35256 -891158
rect 56253 -891378 56256 -891337
rect 77253 -891378 77256 -891337
rect 98253 -891378 98256 -891158
rect 35256 -891394 35260 -891378
rect 56256 -891380 56258 -891378
rect 77256 -891380 77258 -891378
rect 56258 -891394 56260 -891380
rect 77258 -891394 77260 -891380
rect 98256 -891394 98260 -891378
use frameBC_unit  frameBC_unit_0
timestamp 1689774372
transform 1 0 0 0 1 -300000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_1
timestamp 1689774372
transform 1 0 0 0 1 -800000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_2
timestamp 1689774372
transform 1 0 0 0 1 -400000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_3
timestamp 1689774372
transform 1 0 0 0 1 -700000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_4
timestamp 1689774372
transform 1 0 0 0 1 -600000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_5
timestamp 1689774372
transform 1 0 0 0 1 -500000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_6
timestamp 1689774372
transform 1 0 0 0 1 -200000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_7
timestamp 1689774372
transform 1 0 0 0 1 -100000
box -6000 -57000 152000 43000
use frameBC_unit  frameBC_unit_8
timestamp 1689774372
transform 1 0 0 0 1 0
box -6000 -57000 152000 43000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683767628
transform -1 0 112000 0 -1 -857800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_1
timestamp 1683767628
transform -1 0 91000 0 -1 -857800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_2
timestamp 1683767628
transform 1 0 97000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_3
timestamp 1683767628
transform -1 0 70000 0 -1 -857800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_6
timestamp 1683767628
transform 1 0 55000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_7
timestamp 1683767628
transform 1 0 76000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_9
timestamp 1683767628
transform 1 0 34000 0 1 43800
box 0 0 15000 40000
use sky130_ef_io__analog_pad  sky130_ef_io__analog_pad_10
timestamp 1683767628
transform -1 0 49000 0 -1 -857800
box 0 0 15000 40000
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_4 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683767628
transform 1 0 74000 0 1 44207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_5
timestamp 1683767628
transform -1 0 76000 0 -1 -858207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_7
timestamp 1683767628
transform 1 0 95000 0 1 44207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_9
timestamp 1683767628
transform 1 0 53000 0 1 44207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_10
timestamp 1683767628
transform -1 0 55000 0 -1 -858207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_11
timestamp 1683767628
transform -1 0 97000 0 -1 -858207
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_4 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683767628
transform 1 0 70000 0 1 44207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_5
timestamp 1683767628
transform -1 0 74000 0 -1 -858207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_7
timestamp 1683767628
transform 1 0 91000 0 1 44207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_9
timestamp 1683767628
transform 1 0 49000 0 1 44207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_10
timestamp 1683767628
transform -1 0 53000 0 -1 -858207
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_14
timestamp 1683767628
transform -1 0 95000 0 -1 -858207
box 0 0 4000 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683767628
transform 1 0 112000 0 1 43000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_1
timestamp 1683767628
transform 1 0 112000 0 -1 -857000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_3
timestamp 1683767628
transform -1 0 34000 0 -1 -857000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_4
timestamp 1683767628
transform -1 0 34000 0 1 43000
box 0 0 40000 40800
<< end >>
