magic
tech sky130A
magscale 1 2
timestamp 1684833579
<< metal3 >>
rect -1786 1012 1786 1040
rect -1786 -1012 1702 1012
rect 1766 -1012 1786 1012
rect -1786 -1040 1786 -1012
<< via3 >>
rect 1702 -1012 1766 1012
<< mimcap >>
rect -1746 960 1454 1000
rect -1746 -960 -1706 960
rect 1414 -960 1454 960
rect -1746 -1000 1454 -960
<< mimcapcontact >>
rect -1706 -960 1414 960
<< metal4 >>
rect 1686 1012 1782 1028
rect -1707 960 1415 961
rect -1707 -960 -1706 960
rect 1414 -960 1415 960
rect -1707 -961 1415 -960
rect 1686 -1012 1702 1012
rect 1766 -1012 1782 1012
rect 1686 -1028 1782 -1012
<< properties >>
string FIXED_BBOX -1786 -1040 1494 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16 l 10 val 329.88 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
