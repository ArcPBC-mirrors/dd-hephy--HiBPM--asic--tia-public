magic
tech sky130A
magscale 1 2
timestamp 1684167095
<< locali >>
rect 1320 1520 1400 4160
rect 2680 1520 2760 4160
rect 4040 1520 4120 4160
rect 5400 1520 5480 4160
rect 6760 1520 6840 4160
rect 8120 1520 8200 4160
rect 9480 1520 9560 4160
rect 40 1420 10840 1520
rect 1320 40 1400 1420
rect 2680 40 2760 1420
rect 4040 40 4120 1420
rect 5400 40 5480 1420
rect 6760 40 6840 1420
rect 8120 40 8200 1420
rect 9480 40 9560 1420
<< metal1 >>
rect 180 1360 10880 1580
<< metal2 >>
rect 236 1076 10232 1344
<< metal3 >>
rect 74 3764 646 4076
rect 74 2892 84 3764
rect 636 2892 646 3764
rect 1434 3764 2006 4076
rect 2794 3764 3366 4076
rect 1434 2892 1444 3764
rect 1996 2892 2006 3764
rect 2790 2892 2800 3764
rect 3352 3188 3366 3764
rect 4154 3764 4726 4076
rect 3352 2892 3362 3188
rect 4154 2892 4164 3764
rect 4716 2892 4726 3764
rect 5514 3764 6086 4076
rect 5514 2892 5524 3764
rect 6076 2892 6086 3764
rect 6874 3764 7446 4076
rect 6874 2892 6884 3764
rect 7436 2892 7446 3764
rect 8234 3764 8806 4076
rect 8234 2892 8244 3764
rect 8796 2892 8806 3764
rect 9594 3764 10166 4076
rect 9594 2892 9604 3764
rect 10156 2892 10166 3764
rect 38 16 48 660
rect 568 16 578 660
rect 1398 16 1408 660
rect 1928 16 1938 660
rect 2758 16 2768 660
rect 3288 16 3298 660
rect 4118 20 4128 664
rect 4648 20 4658 664
rect 5478 16 5488 660
rect 6008 16 6018 660
rect 6838 16 6848 660
rect 7368 16 7378 660
rect 8198 16 8208 660
rect 8728 16 8738 660
rect 9558 16 9568 660
rect 10088 16 10098 660
<< via3 >>
rect 84 2892 636 3764
rect 1444 2892 1996 3764
rect 2800 2892 3352 3764
rect 4164 2892 4716 3764
rect 5524 2892 6076 3764
rect 6884 2892 7436 3764
rect 8244 2892 8796 3764
rect 9604 2892 10156 3764
rect 48 16 568 660
rect 1408 16 1928 660
rect 2768 16 3288 660
rect 4128 20 4648 664
rect 5488 16 6008 660
rect 6848 16 7368 660
rect 8208 16 8728 660
rect 9568 16 10088 660
<< metal4 >>
rect 83 3764 637 3765
rect 1443 3764 1997 3765
rect 2799 3764 3353 3765
rect 4163 3764 4717 3765
rect 5523 3764 6077 3765
rect 6883 3764 7437 3765
rect 8243 3764 8797 3765
rect 9603 3764 10157 3765
rect 83 2892 84 3764
rect 636 2892 1444 3764
rect 1996 2892 2800 3764
rect 3352 2892 4164 3764
rect 4716 2892 5524 3764
rect 6076 2892 6884 3764
rect 7436 2892 8244 3764
rect 8796 2892 9604 3764
rect 10156 2892 10157 3764
rect 83 2891 637 2892
rect 1443 2891 1997 2892
rect 2799 2891 3353 2892
rect 4163 2891 4717 2892
rect 5523 2891 6077 2892
rect 6883 2891 7437 2892
rect 8243 2891 8797 2892
rect 9603 2891 10157 2892
rect 32 664 10828 960
rect 32 660 4128 664
rect 32 16 48 660
rect 568 16 1408 660
rect 1928 16 2768 660
rect 3288 20 4128 660
rect 4648 660 10828 664
rect 4648 20 5488 660
rect 3288 16 5488 20
rect 6008 16 6848 660
rect 7368 16 8208 660
rect 8728 16 9568 660
rect 10088 16 10828 660
rect 32 -4 10828 16
use bias2_currm  bias2_currm_0
timestamp 1684167095
transform 1 0 9480 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_1
timestamp 1684167095
transform 1 0 -40 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_2
timestamp 1684167095
transform 1 0 1320 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_3
timestamp 1684167095
transform 1 0 2680 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_4
timestamp 1684167095
transform 1 0 4040 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_5
timestamp 1684167095
transform 1 0 5400 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_6
timestamp 1684167095
transform 1 0 6760 0 1 1620
box 40 -1620 1408 2586
use bias2_currm  bias2_currm_7
timestamp 1684167095
transform 1 0 8120 0 1 1620
box 40 -1620 1408 2586
<< end >>
