magic
tech sky130A
magscale 1 2
timestamp 1689778135
<< error_p >>
rect 53740 174178 53744 174194
rect 74740 174178 74744 174194
rect 95740 174178 95744 174194
rect 116740 174178 116744 174194
rect 53744 173958 53747 174178
rect 74744 173958 74747 174178
rect 95744 173958 95747 174178
rect 116744 173958 116747 174178
rect 40987 173909 41215 173925
rect 61987 173909 62215 173925
rect 82987 173909 83215 173925
rect 103987 173909 104215 173925
rect 40984 173898 40987 173909
rect 61984 173898 61987 173909
rect 82984 173898 82987 173909
rect 103984 173898 103987 173909
rect 54004 161442 54016 161462
rect 75004 161442 75016 161462
rect 96004 161442 96016 161462
rect 117004 161442 117016 161462
rect 53780 161435 54004 161442
rect 74780 161435 75004 161442
rect 95780 161435 96004 161442
rect 116780 161435 117004 161442
rect 41253 161182 41256 161190
rect 62253 161182 62256 161190
rect 83253 161182 83256 161402
rect 104253 161182 104256 161190
rect 41256 161166 41260 161182
rect 62256 161166 62260 161182
rect 83256 161166 83260 161182
rect 104256 161166 104260 161182
rect 36178 149213 36180 149297
rect 36262 149172 36264 149213
rect 121820 149172 121822 149297
rect 19138 138804 19158 138816
rect 151298 138813 151309 138816
rect 19158 138580 19165 138804
rect 151309 138585 151325 138813
rect 6422 138544 6642 138547
rect 138582 138544 138802 138547
rect 6406 138540 6422 138544
rect 138566 138540 138582 138544
rect 19418 126056 19434 126060
rect 151578 126056 151594 126060
rect 19198 126053 19418 126056
rect 151358 126053 151578 126056
rect 6675 125787 6691 126015
rect 138835 125796 138842 126020
rect 6691 125784 6702 125787
rect 138842 125784 138862 125796
rect 19138 117804 19158 117816
rect 151298 117813 151309 117816
rect 19158 117580 19165 117804
rect 151309 117585 151325 117813
rect 6422 117544 6642 117547
rect 138582 117544 138802 117547
rect 6406 117540 6422 117544
rect 138566 117540 138582 117544
rect 19418 105056 19434 105060
rect 151578 105056 151594 105060
rect 19198 105053 19418 105056
rect 151358 105053 151578 105056
rect 6675 104787 6691 105015
rect 138835 104796 138842 105020
rect 6691 104784 6702 104787
rect 138842 104784 138862 104796
rect 7583 96800 8483 97115
rect 19138 96804 19158 96816
rect 151298 96813 151309 96816
rect 19158 96580 19165 96804
rect 151309 96585 151325 96813
rect 6422 96544 6642 96547
rect 138582 96544 138802 96547
rect 6406 96311 6422 96544
rect 19252 96490 19472 96493
rect 19472 96257 19488 96490
rect 138566 96311 138582 96544
rect 151537 96490 151632 96493
rect 151632 96257 151648 96490
rect 6102 96224 6322 96227
rect 6086 95991 6102 96224
rect 138256 96218 138482 96227
rect 19572 96160 19802 96173
rect 19802 95937 19808 96160
rect 138246 95991 138256 96218
rect 151732 96170 151952 96173
rect 151952 96053 151968 96170
rect 5782 95904 6002 95907
rect 137942 95904 138162 95907
rect 5766 95774 5782 95904
rect 19892 95850 20112 95853
rect 20112 95617 20128 95850
rect 137926 95671 137942 95904
rect 152069 95850 152272 95853
rect 152272 95784 152288 95850
rect 5420 95542 5640 95545
rect 137580 95542 137800 95545
rect 5404 95518 5420 95542
rect 20200 95518 20436 95531
rect 137564 95518 137580 95542
rect 152360 95518 152596 95531
rect 9275 95323 9309 95357
rect 12297 95323 12331 95357
rect 145669 95323 145703 95357
rect 148691 95323 148725 95357
rect 9275 95285 9347 95321
rect 12259 95285 12331 95321
rect 145669 95285 145741 95321
rect 148653 95285 148725 95321
rect 9275 85279 9347 85315
rect 12259 85279 12331 85315
rect 145669 85279 145741 85315
rect 148653 85279 148725 85315
rect 9275 85243 9309 85277
rect 12297 85243 12331 85277
rect 145669 85243 145703 85277
rect 148691 85243 148725 85277
rect 5404 85069 5640 85082
rect 20420 85058 20436 85082
rect 137564 85069 137800 85082
rect 152580 85058 152596 85082
rect 20200 85055 20420 85058
rect 152360 85055 152580 85058
rect 5712 84750 5728 84816
rect 5728 84747 5931 84750
rect 20058 84696 20074 84929
rect 137872 84750 137888 84983
rect 137888 84747 138108 84750
rect 152218 84696 152234 84826
rect 19838 84693 20058 84696
rect 151998 84693 152218 84696
rect 6032 84430 6048 84547
rect 6048 84427 6268 84430
rect 19744 84382 19754 84609
rect 138192 84440 138198 84663
rect 138198 84427 138428 84440
rect 19518 84373 19744 84382
rect 151898 84376 151914 84609
rect 151678 84373 151898 84376
rect 6352 84110 6368 84343
rect 6368 84107 6463 84110
rect 19418 84056 19434 84289
rect 138512 84110 138528 84343
rect 138528 84107 138748 84110
rect 151578 84056 151594 84289
rect 19198 84053 19418 84056
rect 151358 84053 151578 84056
rect 6675 83787 6691 84015
rect 138835 83796 138842 84020
rect 6691 83784 6702 83787
rect 138842 83784 138862 83796
rect 19138 75804 19158 75816
rect 151298 75813 151309 75816
rect 19158 75580 19165 75804
rect 151309 75585 151325 75813
rect 6422 75544 6642 75547
rect 138582 75544 138802 75547
rect 6406 75311 6422 75544
rect 19252 75490 19472 75493
rect 19472 75257 19488 75490
rect 138566 75311 138582 75544
rect 151537 75490 151632 75493
rect 151632 75257 151648 75490
rect 6102 75224 6322 75227
rect 6086 74991 6102 75224
rect 138256 75218 138482 75227
rect 19572 75160 19802 75173
rect 19802 74937 19808 75160
rect 138246 74991 138256 75218
rect 151732 75170 151952 75173
rect 151952 75053 151968 75170
rect 5782 74904 6002 74907
rect 137942 74904 138162 74907
rect 5766 74774 5782 74904
rect 19892 74850 20112 74853
rect 20112 74617 20128 74850
rect 137926 74671 137942 74904
rect 152069 74850 152272 74853
rect 152272 74617 152288 74850
rect 5420 74542 5640 74545
rect 137580 74542 137800 74545
rect 5404 74518 5420 74542
rect 20200 74518 20436 74531
rect 137564 74518 137580 74542
rect 152360 74518 152596 74531
rect 9275 74323 9309 74357
rect 12297 74323 12331 74357
rect 9275 74285 9347 74321
rect 12259 74285 12331 74321
rect 9275 64279 9347 64315
rect 12259 64279 12331 64315
rect 9275 64243 9309 64277
rect 12297 64243 12331 64277
rect 5404 64069 5640 64082
rect 20420 64058 20436 64082
rect 137564 64069 137800 64082
rect 152580 64058 152596 64082
rect 20200 64055 20420 64058
rect 152360 64055 152580 64058
rect 5712 63750 5728 63816
rect 5728 63747 5931 63750
rect 20058 63696 20074 63929
rect 137872 63750 137888 63983
rect 137888 63747 138108 63750
rect 152218 63696 152234 63929
rect 19838 63693 20058 63696
rect 151998 63693 152218 63696
rect 6032 63430 6048 63547
rect 6048 63427 6268 63430
rect 19744 63382 19754 63609
rect 138192 63440 138198 63663
rect 138198 63427 138428 63440
rect 19518 63373 19744 63382
rect 151898 63376 151914 63609
rect 151678 63373 151898 63376
rect 6352 63110 6368 63343
rect 6368 63107 6463 63110
rect 19418 63056 19434 63289
rect 138512 63110 138528 63343
rect 138528 63107 138748 63110
rect 151578 63056 151594 63289
rect 19198 63053 19418 63056
rect 151358 63053 151578 63056
rect 6675 62787 6691 63015
rect 138835 62796 138842 63020
rect 6691 62784 6702 62787
rect 138842 62784 138862 62796
rect 19138 54804 19158 54816
rect 151298 54813 151309 54816
rect 19158 54580 19165 54804
rect 151309 54585 151325 54813
rect 6422 54544 6642 54547
rect 138582 54544 138802 54547
rect 6406 54311 6422 54544
rect 19252 54490 19472 54493
rect 19472 54257 19488 54490
rect 138566 54311 138582 54544
rect 151537 54490 151632 54493
rect 151632 54257 151648 54490
rect 6102 54224 6322 54227
rect 6086 53991 6102 54224
rect 138256 54218 138482 54227
rect 19572 54160 19802 54173
rect 19802 53937 19808 54160
rect 138246 53991 138256 54218
rect 151732 54170 151952 54173
rect 151952 54053 151968 54170
rect 5782 53904 6002 53907
rect 137942 53904 138162 53907
rect 5766 53671 5782 53904
rect 19892 53850 20112 53853
rect 20112 53617 20128 53850
rect 137926 53671 137942 53904
rect 152069 53850 152272 53853
rect 152272 53784 152288 53850
rect 5420 53542 5640 53545
rect 137580 53542 137800 53545
rect 5404 53518 5420 53542
rect 20200 53518 20436 53531
rect 137564 53518 137580 53542
rect 152360 53518 152596 53531
rect 145669 53323 145703 53357
rect 148691 53323 148725 53357
rect 145669 53285 145741 53321
rect 148653 53285 148725 53321
rect 145669 43279 145741 43315
rect 148653 43279 148725 43315
rect 145669 43243 145703 43277
rect 148691 43243 148725 43277
rect 5404 43069 5640 43082
rect 20420 43058 20436 43082
rect 137564 43069 137800 43082
rect 152580 43058 152596 43082
rect 20200 43055 20420 43058
rect 152360 43055 152580 43058
rect 5712 42750 5728 42983
rect 5728 42747 5931 42750
rect 20058 42696 20074 42929
rect 137872 42750 137888 42983
rect 137888 42747 138108 42750
rect 152218 42696 152234 42826
rect 19838 42693 20058 42696
rect 151998 42693 152218 42696
rect 6032 42430 6048 42547
rect 6048 42427 6268 42430
rect 19744 42382 19754 42609
rect 138192 42440 138198 42663
rect 138198 42427 138428 42440
rect 19518 42373 19744 42382
rect 151898 42376 151914 42609
rect 151678 42373 151898 42376
rect 6352 42110 6368 42343
rect 6368 42107 6463 42110
rect 19418 42056 19434 42289
rect 138512 42110 138528 42343
rect 138528 42107 138748 42110
rect 151578 42056 151594 42289
rect 19198 42053 19418 42056
rect 151358 42053 151578 42056
rect 6675 41787 6691 42015
rect 138835 41796 138842 42020
rect 6691 41784 6702 41787
rect 138842 41784 138862 41796
rect 53740 19418 53744 19434
rect 74740 19418 74744 19434
rect 95540 19418 95744 19434
rect 116740 19418 116744 19434
rect 53744 19410 53747 19418
rect 74744 19410 74747 19418
rect 95744 19198 95747 19418
rect 116744 19410 116747 19418
rect 40996 19158 41220 19165
rect 61996 19158 62220 19165
rect 82996 19158 83220 19165
rect 103996 19158 104220 19165
rect 40984 19138 40996 19158
rect 61984 19138 61996 19158
rect 82984 19138 82996 19158
rect 103984 19138 103996 19158
rect 54013 6691 54016 6702
rect 75013 6691 75016 6702
rect 96013 6691 96016 6702
rect 117013 6691 117016 6702
rect 53785 6675 54013 6691
rect 74785 6675 75013 6691
rect 95785 6675 96013 6691
rect 116785 6675 117013 6691
rect 41253 6422 41256 6642
rect 62253 6422 62256 6463
rect 83253 6422 83256 6642
rect 41256 6406 41260 6422
rect 62256 6420 62258 6422
rect 62258 6406 62260 6420
rect 83256 6406 83260 6422
rect 95690 6368 95693 6463
rect 104253 6422 104256 6642
rect 104256 6406 104260 6422
rect 95540 6352 95690 6368
<< metal3 >>
rect 82100 140100 86900 141400
rect 92100 140000 97000 141700
rect 39400 135000 40300 139700
rect 39100 124900 40400 129700
rect 117900 113900 119600 118700
rect 117900 103900 119600 108600
rect 118100 71900 118900 76700
rect 117900 61800 118700 66700
rect 38700 50900 41500 55800
rect 38700 40800 41500 45700
rect 82000 39400 86800 40000
rect 92100 39500 96900 40100
use core1B  core1B_0
timestamp 1689778135
transform 1 0 -34 0 1 14
box 39460 39580 118400 141020
use frame  frame_1 ~/code/hibpm-sky130a-tapeout/mag/frame
timestamp 1687287864
transform 1 0 6000 0 1 96800
box -6000 -96800 152000 83800
<< end >>
