magic
tech sky130A
magscale 1 2
timestamp 1686659968
<< metal1 >>
rect 5076 2064 6872 2160
rect 5026 1852 5036 2036
rect 5092 1852 5102 2036
rect 5218 1852 5228 2036
rect 5284 1852 5294 2036
rect 5410 1852 5420 2036
rect 5476 1852 5486 2036
rect 5602 1852 5612 2036
rect 5668 1852 5678 2036
rect 5794 1852 5804 2036
rect 5860 1852 5870 2036
rect 5986 1852 5996 2036
rect 6052 1852 6062 2036
rect 6178 1852 6188 2036
rect 6244 1852 6254 2036
rect 6370 1852 6380 2036
rect 6436 1852 6446 2036
rect 6562 1852 6572 2036
rect 6628 1852 6638 2036
rect 6754 1852 6764 2036
rect 6820 1852 6830 2036
rect 4930 1632 4940 1816
rect 4996 1632 5006 1816
rect 5122 1632 5132 1816
rect 5188 1632 5198 1816
rect 5314 1632 5324 1816
rect 5380 1632 5390 1816
rect 5506 1632 5516 1816
rect 5572 1632 5582 1816
rect 5698 1632 5708 1816
rect 5764 1632 5774 1816
rect 5890 1632 5900 1816
rect 5956 1632 5966 1816
rect 6082 1632 6092 1816
rect 6148 1632 6158 1816
rect 6274 1632 6284 1816
rect 6340 1632 6350 1816
rect 6466 1632 6476 1816
rect 6532 1632 6542 1816
rect 6658 1632 6668 1816
rect 6724 1632 6734 1816
rect 6850 1632 6860 1816
rect 6916 1632 6926 1816
rect 4980 1448 6776 1604
rect 5026 1236 5036 1420
rect 5092 1236 5102 1420
rect 5218 1236 5228 1420
rect 5284 1236 5294 1420
rect 5410 1236 5420 1420
rect 5476 1236 5486 1420
rect 5602 1236 5612 1420
rect 5668 1236 5678 1420
rect 5794 1236 5804 1420
rect 5860 1236 5870 1420
rect 5986 1236 5996 1420
rect 6052 1236 6062 1420
rect 6178 1236 6188 1420
rect 6244 1236 6254 1420
rect 6370 1236 6380 1420
rect 6436 1236 6446 1420
rect 6562 1236 6572 1420
rect 6628 1236 6638 1420
rect 6754 1236 6764 1420
rect 6820 1236 6830 1420
rect 4930 1016 4940 1200
rect 4996 1016 5006 1200
rect 5122 1016 5132 1200
rect 5188 1016 5198 1200
rect 5314 1016 5324 1200
rect 5380 1016 5390 1200
rect 5506 1016 5516 1200
rect 5572 1016 5582 1200
rect 5698 1016 5708 1200
rect 5764 1016 5774 1200
rect 5890 1016 5900 1200
rect 5956 1016 5966 1200
rect 6082 1016 6092 1200
rect 6148 1016 6158 1200
rect 6274 1016 6284 1200
rect 6340 1016 6350 1200
rect 6466 1016 6476 1200
rect 6532 1016 6542 1200
rect 6658 1016 6668 1200
rect 6724 1016 6734 1200
rect 6850 1016 6860 1200
rect 6916 1016 6926 1200
rect 5076 828 6872 984
rect 5026 616 5036 800
rect 5092 616 5102 800
rect 5218 616 5228 800
rect 5284 616 5294 800
rect 5410 616 5420 800
rect 5476 616 5486 800
rect 5602 616 5612 800
rect 5668 616 5678 800
rect 5794 616 5804 800
rect 5860 616 5870 800
rect 5986 616 5996 800
rect 6052 616 6062 800
rect 6178 616 6188 800
rect 6244 616 6254 800
rect 6370 616 6380 800
rect 6436 616 6446 800
rect 6562 616 6572 800
rect 6628 616 6638 800
rect 6754 616 6764 800
rect 6820 616 6830 800
rect 4930 396 4940 580
rect 4996 396 5006 580
rect 5122 396 5132 580
rect 5188 396 5198 580
rect 5314 396 5324 580
rect 5380 396 5390 580
rect 5506 396 5516 580
rect 5572 396 5582 580
rect 5698 396 5708 580
rect 5764 396 5774 580
rect 5890 396 5900 580
rect 5956 396 5966 580
rect 6082 396 6092 580
rect 6148 396 6158 580
rect 6274 396 6284 580
rect 6340 396 6350 580
rect 6466 396 6476 580
rect 6532 396 6542 580
rect 6658 396 6668 580
rect 6724 396 6734 580
rect 6850 396 6860 580
rect 6916 396 6926 580
rect 4980 212 6776 368
rect 5026 0 5036 184
rect 5092 0 5102 184
rect 5218 0 5228 184
rect 5284 0 5294 184
rect 5410 0 5420 184
rect 5476 0 5486 184
rect 5602 0 5612 184
rect 5668 0 5678 184
rect 5794 0 5804 184
rect 5860 0 5870 184
rect 5986 0 5996 184
rect 6052 0 6062 184
rect 6178 0 6188 184
rect 6244 0 6254 184
rect 6370 0 6380 184
rect 6436 0 6446 184
rect 6562 0 6572 184
rect 6628 0 6638 184
rect 6754 0 6764 184
rect 6820 0 6830 184
rect 4930 -220 4940 -36
rect 4996 -220 5006 -36
rect 5122 -220 5132 -36
rect 5188 -220 5198 -36
rect 5314 -220 5324 -36
rect 5380 -220 5390 -36
rect 5506 -220 5516 -36
rect 5572 -220 5582 -36
rect 5698 -220 5708 -36
rect 5764 -220 5774 -36
rect 5890 -220 5900 -36
rect 5956 -220 5966 -36
rect 6082 -220 6092 -36
rect 6148 -220 6158 -36
rect 6274 -220 6284 -36
rect 6340 -220 6350 -36
rect 6466 -220 6476 -36
rect 6532 -220 6542 -36
rect 6658 -220 6668 -36
rect 6724 -220 6734 -36
rect 6850 -220 6860 -36
rect 6916 -220 6926 -36
rect 5076 -408 6872 -252
rect 5026 -620 5036 -436
rect 5092 -620 5102 -436
rect 5218 -620 5228 -436
rect 5284 -620 5294 -436
rect 5410 -620 5420 -436
rect 5476 -620 5486 -436
rect 5602 -620 5612 -436
rect 5668 -620 5678 -436
rect 5794 -620 5804 -436
rect 5860 -620 5870 -436
rect 5986 -620 5996 -436
rect 6052 -620 6062 -436
rect 6178 -620 6188 -436
rect 6244 -620 6254 -436
rect 6370 -620 6380 -436
rect 6436 -620 6446 -436
rect 6562 -620 6572 -436
rect 6628 -620 6638 -436
rect 6754 -620 6764 -436
rect 6820 -620 6830 -436
rect 4930 -840 4940 -656
rect 4996 -840 5006 -656
rect 5122 -840 5132 -656
rect 5188 -840 5198 -656
rect 5314 -840 5324 -656
rect 5380 -840 5390 -656
rect 5506 -840 5516 -656
rect 5572 -840 5582 -656
rect 5698 -840 5708 -656
rect 5764 -840 5774 -656
rect 5890 -840 5900 -656
rect 5956 -840 5966 -656
rect 6082 -840 6092 -656
rect 6148 -840 6158 -656
rect 6274 -840 6284 -656
rect 6340 -840 6350 -656
rect 6466 -840 6476 -656
rect 6532 -840 6542 -656
rect 6658 -840 6668 -656
rect 6724 -840 6734 -656
rect 6850 -840 6860 -656
rect 6916 -840 6926 -656
rect 4980 -1024 6776 -868
rect 5026 -1236 5036 -1052
rect 5092 -1236 5102 -1052
rect 5218 -1236 5228 -1052
rect 5284 -1236 5294 -1052
rect 5410 -1236 5420 -1052
rect 5476 -1236 5486 -1052
rect 5602 -1236 5612 -1052
rect 5668 -1236 5678 -1052
rect 5794 -1236 5804 -1052
rect 5860 -1236 5870 -1052
rect 5986 -1236 5996 -1052
rect 6052 -1236 6062 -1052
rect 6178 -1236 6188 -1052
rect 6244 -1236 6254 -1052
rect 6370 -1236 6380 -1052
rect 6436 -1236 6446 -1052
rect 6562 -1236 6572 -1052
rect 6628 -1236 6638 -1052
rect 6754 -1236 6764 -1052
rect 6820 -1236 6830 -1052
rect 4930 -1456 4940 -1272
rect 4996 -1456 5006 -1272
rect 5122 -1456 5132 -1272
rect 5188 -1456 5198 -1272
rect 5314 -1456 5324 -1272
rect 5380 -1456 5390 -1272
rect 5506 -1456 5516 -1272
rect 5572 -1456 5582 -1272
rect 5698 -1456 5708 -1272
rect 5764 -1456 5774 -1272
rect 5890 -1456 5900 -1272
rect 5956 -1456 5966 -1272
rect 6082 -1456 6092 -1272
rect 6148 -1456 6158 -1272
rect 6274 -1456 6284 -1272
rect 6340 -1456 6350 -1272
rect 6466 -1456 6476 -1272
rect 6532 -1456 6542 -1272
rect 6658 -1456 6668 -1272
rect 6724 -1456 6734 -1272
rect 6850 -1456 6860 -1272
rect 6916 -1456 6926 -1272
rect 5076 -1644 6872 -1488
rect 5026 -1856 5036 -1672
rect 5092 -1856 5102 -1672
rect 5218 -1856 5228 -1672
rect 5284 -1856 5294 -1672
rect 5410 -1856 5420 -1672
rect 5476 -1856 5486 -1672
rect 5602 -1856 5612 -1672
rect 5668 -1856 5678 -1672
rect 5794 -1856 5804 -1672
rect 5860 -1856 5870 -1672
rect 5986 -1856 5996 -1672
rect 6052 -1856 6062 -1672
rect 6178 -1856 6188 -1672
rect 6244 -1856 6254 -1672
rect 6370 -1856 6380 -1672
rect 6436 -1856 6446 -1672
rect 6562 -1856 6572 -1672
rect 6628 -1856 6638 -1672
rect 6754 -1856 6764 -1672
rect 6820 -1856 6830 -1672
rect 4930 -2076 4940 -1892
rect 4996 -2076 5006 -1892
rect 5122 -2076 5132 -1892
rect 5188 -2076 5198 -1892
rect 5314 -2076 5324 -1892
rect 5380 -2076 5390 -1892
rect 5506 -2076 5516 -1892
rect 5572 -2076 5582 -1892
rect 5698 -2076 5708 -1892
rect 5764 -2076 5774 -1892
rect 5890 -2076 5900 -1892
rect 5956 -2076 5966 -1892
rect 6082 -2076 6092 -1892
rect 6148 -2076 6158 -1892
rect 6274 -2076 6284 -1892
rect 6340 -2076 6350 -1892
rect 6466 -2076 6476 -1892
rect 6532 -2076 6542 -1892
rect 6658 -2076 6668 -1892
rect 6724 -2076 6734 -1892
rect 6850 -2076 6860 -1892
rect 6916 -2076 6926 -1892
rect 4980 -2260 6776 -2104
rect 5026 -2472 5036 -2288
rect 5092 -2472 5102 -2288
rect 5218 -2472 5228 -2288
rect 5284 -2472 5294 -2288
rect 5410 -2472 5420 -2288
rect 5476 -2472 5486 -2288
rect 5602 -2472 5612 -2288
rect 5668 -2472 5678 -2288
rect 5794 -2472 5804 -2288
rect 5860 -2472 5870 -2288
rect 5986 -2472 5996 -2288
rect 6052 -2472 6062 -2288
rect 6178 -2472 6188 -2288
rect 6244 -2472 6254 -2288
rect 6370 -2472 6380 -2288
rect 6436 -2472 6446 -2288
rect 6562 -2472 6572 -2288
rect 6628 -2472 6638 -2288
rect 6754 -2472 6764 -2288
rect 6820 -2472 6830 -2288
rect 4930 -2692 4940 -2508
rect 4996 -2692 5006 -2508
rect 5122 -2692 5132 -2508
rect 5188 -2692 5198 -2508
rect 5314 -2692 5324 -2508
rect 5380 -2692 5390 -2508
rect 5506 -2692 5516 -2508
rect 5572 -2692 5582 -2508
rect 5698 -2692 5708 -2508
rect 5764 -2692 5774 -2508
rect 5890 -2692 5900 -2508
rect 5956 -2692 5966 -2508
rect 6082 -2692 6092 -2508
rect 6148 -2692 6158 -2508
rect 6274 -2692 6284 -2508
rect 6340 -2692 6350 -2508
rect 6466 -2692 6476 -2508
rect 6532 -2692 6542 -2508
rect 6658 -2692 6668 -2508
rect 6724 -2692 6734 -2508
rect 6850 -2692 6860 -2508
rect 6916 -2692 6926 -2508
rect 5076 -2880 6872 -2724
rect 5026 -3092 5036 -2908
rect 5092 -3092 5102 -2908
rect 5218 -3092 5228 -2908
rect 5284 -3092 5294 -2908
rect 5410 -3092 5420 -2908
rect 5476 -3092 5486 -2908
rect 5602 -3092 5612 -2908
rect 5668 -3092 5678 -2908
rect 5794 -3092 5804 -2908
rect 5860 -3092 5870 -2908
rect 5986 -3092 5996 -2908
rect 6052 -3092 6062 -2908
rect 6178 -3092 6188 -2908
rect 6244 -3092 6254 -2908
rect 6370 -3092 6380 -2908
rect 6436 -3092 6446 -2908
rect 6562 -3092 6572 -2908
rect 6628 -3092 6638 -2908
rect 6754 -3092 6764 -2908
rect 6820 -3092 6830 -2908
rect 4930 -3312 4940 -3128
rect 4996 -3312 5006 -3128
rect 5122 -3312 5132 -3128
rect 5188 -3312 5198 -3128
rect 5314 -3312 5324 -3128
rect 5380 -3312 5390 -3128
rect 5506 -3312 5516 -3128
rect 5572 -3312 5582 -3128
rect 5698 -3312 5708 -3128
rect 5764 -3312 5774 -3128
rect 5890 -3312 5900 -3128
rect 5956 -3312 5966 -3128
rect 6082 -3312 6092 -3128
rect 6148 -3312 6158 -3128
rect 6274 -3312 6284 -3128
rect 6340 -3312 6350 -3128
rect 6466 -3312 6476 -3128
rect 6532 -3312 6542 -3128
rect 6658 -3312 6668 -3128
rect 6724 -3312 6734 -3128
rect 6850 -3312 6860 -3128
rect 6916 -3312 6926 -3128
rect 4980 -3436 6776 -3340
<< via1 >>
rect 5036 1852 5092 2036
rect 5228 1852 5284 2036
rect 5420 1852 5476 2036
rect 5612 1852 5668 2036
rect 5804 1852 5860 2036
rect 5996 1852 6052 2036
rect 6188 1852 6244 2036
rect 6380 1852 6436 2036
rect 6572 1852 6628 2036
rect 6764 1852 6820 2036
rect 4940 1632 4996 1816
rect 5132 1632 5188 1816
rect 5324 1632 5380 1816
rect 5516 1632 5572 1816
rect 5708 1632 5764 1816
rect 5900 1632 5956 1816
rect 6092 1632 6148 1816
rect 6284 1632 6340 1816
rect 6476 1632 6532 1816
rect 6668 1632 6724 1816
rect 6860 1632 6916 1816
rect 5036 1236 5092 1420
rect 5228 1236 5284 1420
rect 5420 1236 5476 1420
rect 5612 1236 5668 1420
rect 5804 1236 5860 1420
rect 5996 1236 6052 1420
rect 6188 1236 6244 1420
rect 6380 1236 6436 1420
rect 6572 1236 6628 1420
rect 6764 1236 6820 1420
rect 4940 1016 4996 1200
rect 5132 1016 5188 1200
rect 5324 1016 5380 1200
rect 5516 1016 5572 1200
rect 5708 1016 5764 1200
rect 5900 1016 5956 1200
rect 6092 1016 6148 1200
rect 6284 1016 6340 1200
rect 6476 1016 6532 1200
rect 6668 1016 6724 1200
rect 6860 1016 6916 1200
rect 5036 616 5092 800
rect 5228 616 5284 800
rect 5420 616 5476 800
rect 5612 616 5668 800
rect 5804 616 5860 800
rect 5996 616 6052 800
rect 6188 616 6244 800
rect 6380 616 6436 800
rect 6572 616 6628 800
rect 6764 616 6820 800
rect 4940 396 4996 580
rect 5132 396 5188 580
rect 5324 396 5380 580
rect 5516 396 5572 580
rect 5708 396 5764 580
rect 5900 396 5956 580
rect 6092 396 6148 580
rect 6284 396 6340 580
rect 6476 396 6532 580
rect 6668 396 6724 580
rect 6860 396 6916 580
rect 5036 0 5092 184
rect 5228 0 5284 184
rect 5420 0 5476 184
rect 5612 0 5668 184
rect 5804 0 5860 184
rect 5996 0 6052 184
rect 6188 0 6244 184
rect 6380 0 6436 184
rect 6572 0 6628 184
rect 6764 0 6820 184
rect 4940 -220 4996 -36
rect 5132 -220 5188 -36
rect 5324 -220 5380 -36
rect 5516 -220 5572 -36
rect 5708 -220 5764 -36
rect 5900 -220 5956 -36
rect 6092 -220 6148 -36
rect 6284 -220 6340 -36
rect 6476 -220 6532 -36
rect 6668 -220 6724 -36
rect 6860 -220 6916 -36
rect 5036 -620 5092 -436
rect 5228 -620 5284 -436
rect 5420 -620 5476 -436
rect 5612 -620 5668 -436
rect 5804 -620 5860 -436
rect 5996 -620 6052 -436
rect 6188 -620 6244 -436
rect 6380 -620 6436 -436
rect 6572 -620 6628 -436
rect 6764 -620 6820 -436
rect 4940 -840 4996 -656
rect 5132 -840 5188 -656
rect 5324 -840 5380 -656
rect 5516 -840 5572 -656
rect 5708 -840 5764 -656
rect 5900 -840 5956 -656
rect 6092 -840 6148 -656
rect 6284 -840 6340 -656
rect 6476 -840 6532 -656
rect 6668 -840 6724 -656
rect 6860 -840 6916 -656
rect 5036 -1236 5092 -1052
rect 5228 -1236 5284 -1052
rect 5420 -1236 5476 -1052
rect 5612 -1236 5668 -1052
rect 5804 -1236 5860 -1052
rect 5996 -1236 6052 -1052
rect 6188 -1236 6244 -1052
rect 6380 -1236 6436 -1052
rect 6572 -1236 6628 -1052
rect 6764 -1236 6820 -1052
rect 4940 -1456 4996 -1272
rect 5132 -1456 5188 -1272
rect 5324 -1456 5380 -1272
rect 5516 -1456 5572 -1272
rect 5708 -1456 5764 -1272
rect 5900 -1456 5956 -1272
rect 6092 -1456 6148 -1272
rect 6284 -1456 6340 -1272
rect 6476 -1456 6532 -1272
rect 6668 -1456 6724 -1272
rect 6860 -1456 6916 -1272
rect 5036 -1856 5092 -1672
rect 5228 -1856 5284 -1672
rect 5420 -1856 5476 -1672
rect 5612 -1856 5668 -1672
rect 5804 -1856 5860 -1672
rect 5996 -1856 6052 -1672
rect 6188 -1856 6244 -1672
rect 6380 -1856 6436 -1672
rect 6572 -1856 6628 -1672
rect 6764 -1856 6820 -1672
rect 4940 -2076 4996 -1892
rect 5132 -2076 5188 -1892
rect 5324 -2076 5380 -1892
rect 5516 -2076 5572 -1892
rect 5708 -2076 5764 -1892
rect 5900 -2076 5956 -1892
rect 6092 -2076 6148 -1892
rect 6284 -2076 6340 -1892
rect 6476 -2076 6532 -1892
rect 6668 -2076 6724 -1892
rect 6860 -2076 6916 -1892
rect 5036 -2472 5092 -2288
rect 5228 -2472 5284 -2288
rect 5420 -2472 5476 -2288
rect 5612 -2472 5668 -2288
rect 5804 -2472 5860 -2288
rect 5996 -2472 6052 -2288
rect 6188 -2472 6244 -2288
rect 6380 -2472 6436 -2288
rect 6572 -2472 6628 -2288
rect 6764 -2472 6820 -2288
rect 4940 -2692 4996 -2508
rect 5132 -2692 5188 -2508
rect 5324 -2692 5380 -2508
rect 5516 -2692 5572 -2508
rect 5708 -2692 5764 -2508
rect 5900 -2692 5956 -2508
rect 6092 -2692 6148 -2508
rect 6284 -2692 6340 -2508
rect 6476 -2692 6532 -2508
rect 6668 -2692 6724 -2508
rect 6860 -2692 6916 -2508
rect 5036 -3092 5092 -2908
rect 5228 -3092 5284 -2908
rect 5420 -3092 5476 -2908
rect 5612 -3092 5668 -2908
rect 5804 -3092 5860 -2908
rect 5996 -3092 6052 -2908
rect 6188 -3092 6244 -2908
rect 6380 -3092 6436 -2908
rect 6572 -3092 6628 -2908
rect 6764 -3092 6820 -2908
rect 4940 -3312 4996 -3128
rect 5132 -3312 5188 -3128
rect 5324 -3312 5380 -3128
rect 5516 -3312 5572 -3128
rect 5708 -3312 5764 -3128
rect 5900 -3312 5956 -3128
rect 6092 -3312 6148 -3128
rect 6284 -3312 6340 -3128
rect 6476 -3312 6532 -3128
rect 6668 -3312 6724 -3128
rect 6860 -3312 6916 -3128
<< metal2 >>
rect 6084 2064 6956 2074
rect 5032 2036 6084 2048
rect 5032 1856 5036 2036
rect 5092 1856 5228 2036
rect 5036 1842 5092 1852
rect 5284 1856 5420 2036
rect 5228 1842 5284 1852
rect 5476 1856 5612 2036
rect 5420 1842 5476 1852
rect 5668 1856 5804 2036
rect 5612 1842 5668 1852
rect 5860 1856 5996 2036
rect 5804 1842 5860 1852
rect 6052 1864 6084 2036
rect 6052 1856 6188 1864
rect 6084 1854 6188 1856
rect 5996 1842 6052 1852
rect 6244 1854 6380 1864
rect 6188 1842 6244 1852
rect 6436 1854 6572 1864
rect 6380 1842 6436 1852
rect 6628 1854 6764 1864
rect 6572 1842 6628 1852
rect 6820 1854 6956 1864
rect 6764 1842 6820 1852
rect 4940 1816 4996 1826
rect 4932 1804 4940 1814
rect 5132 1816 5188 1826
rect 4996 1804 5132 1814
rect 5324 1816 5380 1826
rect 5188 1804 5324 1814
rect 5516 1816 5572 1826
rect 5380 1804 5516 1814
rect 5708 1816 5764 1826
rect 5572 1804 5708 1814
rect 5900 1816 5956 1826
rect 5764 1804 5900 1814
rect 6092 1816 6148 1826
rect 5956 1632 6092 1812
rect 6284 1816 6340 1826
rect 6148 1632 6284 1812
rect 6476 1816 6532 1826
rect 6340 1632 6476 1812
rect 6668 1816 6724 1826
rect 6532 1632 6668 1812
rect 6860 1816 6916 1826
rect 6724 1632 6860 1812
rect 5916 1620 6916 1632
rect 4932 1606 5916 1616
rect 6088 1448 6960 1458
rect 5032 1420 6088 1432
rect 5032 1240 5036 1420
rect 5092 1240 5228 1420
rect 5036 1226 5092 1236
rect 5284 1240 5420 1420
rect 5228 1226 5284 1236
rect 5476 1240 5612 1420
rect 5420 1226 5476 1236
rect 5668 1240 5804 1420
rect 5612 1226 5668 1236
rect 5860 1240 5996 1420
rect 5804 1226 5860 1236
rect 6052 1248 6088 1420
rect 6052 1240 6188 1248
rect 6088 1238 6188 1240
rect 5996 1226 6052 1236
rect 6244 1238 6380 1248
rect 6188 1226 6244 1236
rect 6436 1238 6572 1248
rect 6380 1226 6436 1236
rect 6628 1238 6764 1248
rect 6572 1226 6628 1236
rect 6820 1238 6960 1248
rect 6764 1226 6820 1236
rect 4940 1200 4996 1210
rect 4936 1184 4940 1196
rect 5132 1200 5188 1210
rect 4996 1184 5132 1196
rect 5324 1200 5380 1210
rect 5188 1184 5324 1196
rect 5516 1200 5572 1210
rect 5380 1184 5516 1196
rect 5708 1200 5764 1210
rect 5572 1184 5708 1196
rect 5900 1200 5956 1210
rect 5764 1184 5900 1196
rect 6092 1200 6148 1210
rect 5956 1016 6092 1196
rect 6284 1200 6340 1210
rect 6148 1016 6284 1196
rect 6476 1200 6532 1210
rect 6340 1016 6476 1196
rect 6668 1200 6724 1210
rect 6532 1016 6668 1196
rect 6860 1200 6916 1210
rect 6724 1016 6860 1196
rect 5920 1004 6916 1016
rect 4936 986 5920 996
rect 6088 832 6960 842
rect 5032 800 6088 812
rect 5032 620 5036 800
rect 5092 620 5228 800
rect 5036 606 5092 616
rect 5284 620 5420 800
rect 5228 606 5284 616
rect 5476 620 5612 800
rect 5420 606 5476 616
rect 5668 620 5804 800
rect 5612 606 5668 616
rect 5860 620 5996 800
rect 5804 606 5860 616
rect 6052 632 6088 800
rect 6052 620 6188 632
rect 5996 606 6052 616
rect 6244 620 6380 632
rect 6188 606 6244 616
rect 6436 620 6572 632
rect 6380 606 6436 616
rect 6628 620 6764 632
rect 6572 606 6628 616
rect 6820 622 6960 632
rect 6820 620 6824 622
rect 6764 606 6820 616
rect 4940 580 4996 590
rect 4932 568 4940 578
rect 5132 580 5188 590
rect 4996 568 5132 578
rect 5324 580 5380 590
rect 5188 568 5324 578
rect 5516 580 5572 590
rect 5380 568 5516 578
rect 5708 580 5764 590
rect 5572 568 5708 578
rect 5900 580 5956 590
rect 5764 568 5900 578
rect 6092 580 6148 590
rect 5956 396 6092 576
rect 6284 580 6340 590
rect 6148 396 6284 576
rect 6476 580 6532 590
rect 6340 396 6476 576
rect 6668 580 6724 590
rect 6532 396 6668 576
rect 6860 580 6916 590
rect 6724 396 6860 576
rect 5916 384 6916 396
rect 4932 370 5916 380
rect 6088 212 6960 222
rect 5032 184 6088 196
rect 5032 4 5036 184
rect 5092 4 5228 184
rect 5036 -10 5092 0
rect 5284 4 5420 184
rect 5228 -10 5284 0
rect 5476 4 5612 184
rect 5420 -10 5476 0
rect 5668 4 5804 184
rect 5612 -10 5668 0
rect 5860 4 5996 184
rect 5804 -10 5860 0
rect 6052 12 6088 184
rect 6052 4 6188 12
rect 6088 2 6188 4
rect 5996 -10 6052 0
rect 6244 2 6380 12
rect 6188 -10 6244 0
rect 6436 2 6572 12
rect 6380 -10 6436 0
rect 6628 2 6764 12
rect 6572 -10 6628 0
rect 6820 2 6960 12
rect 6764 -10 6820 0
rect 4940 -36 4996 -26
rect 4928 -48 4940 -38
rect 5132 -36 5188 -26
rect 4996 -48 5132 -38
rect 5324 -36 5380 -26
rect 5188 -48 5324 -38
rect 5516 -36 5572 -26
rect 5380 -48 5516 -38
rect 5708 -36 5764 -26
rect 5572 -48 5708 -38
rect 5900 -36 5956 -26
rect 5764 -48 5900 -38
rect 6092 -36 6148 -26
rect 5956 -220 6092 -40
rect 6284 -36 6340 -26
rect 6148 -220 6284 -40
rect 6476 -36 6532 -26
rect 6340 -220 6476 -40
rect 6668 -36 6724 -26
rect 6532 -220 6668 -40
rect 6860 -36 6916 -26
rect 6724 -220 6860 -40
rect 5912 -232 6916 -220
rect 4928 -246 5912 -236
rect 6088 -408 6960 -398
rect 5032 -436 6088 -424
rect 5032 -616 5036 -436
rect 5092 -616 5228 -436
rect 5036 -630 5092 -620
rect 5284 -616 5420 -436
rect 5228 -630 5284 -620
rect 5476 -616 5612 -436
rect 5420 -630 5476 -620
rect 5668 -616 5804 -436
rect 5612 -630 5668 -620
rect 5860 -616 5996 -436
rect 5804 -630 5860 -620
rect 6052 -608 6088 -436
rect 6052 -616 6188 -608
rect 6088 -618 6188 -616
rect 5996 -630 6052 -620
rect 6244 -618 6380 -608
rect 6188 -630 6244 -620
rect 6436 -618 6572 -608
rect 6380 -630 6436 -620
rect 6628 -618 6764 -608
rect 6572 -630 6628 -620
rect 6820 -618 6960 -608
rect 6764 -630 6820 -620
rect 4940 -656 4996 -646
rect 4936 -662 4940 -660
rect 4932 -672 4940 -662
rect 5132 -656 5188 -646
rect 4996 -672 5132 -660
rect 5324 -656 5380 -646
rect 5188 -672 5324 -660
rect 5516 -656 5572 -646
rect 5380 -672 5516 -660
rect 5708 -656 5764 -646
rect 5572 -672 5708 -660
rect 5900 -656 5956 -646
rect 5764 -672 5900 -660
rect 6092 -656 6148 -646
rect 5956 -840 6092 -660
rect 6284 -656 6340 -646
rect 6148 -840 6284 -660
rect 6476 -656 6532 -646
rect 6340 -840 6476 -660
rect 6668 -656 6724 -646
rect 6532 -840 6668 -660
rect 6860 -656 6916 -646
rect 6724 -840 6860 -660
rect 5916 -852 6916 -840
rect 4932 -870 5916 -860
rect 6088 -1024 6960 -1014
rect 5032 -1052 6088 -1040
rect 5032 -1232 5036 -1052
rect 5092 -1232 5228 -1052
rect 5036 -1246 5092 -1236
rect 5284 -1232 5420 -1052
rect 5228 -1246 5284 -1236
rect 5476 -1232 5612 -1052
rect 5420 -1246 5476 -1236
rect 5668 -1232 5804 -1052
rect 5612 -1246 5668 -1236
rect 5860 -1232 5996 -1052
rect 5804 -1246 5860 -1236
rect 6052 -1224 6088 -1052
rect 6052 -1232 6188 -1224
rect 6088 -1234 6188 -1232
rect 5996 -1246 6052 -1236
rect 6244 -1234 6380 -1224
rect 6188 -1246 6244 -1236
rect 6436 -1234 6572 -1224
rect 6380 -1246 6436 -1236
rect 6628 -1234 6764 -1224
rect 6572 -1246 6628 -1236
rect 6820 -1234 6960 -1224
rect 6764 -1246 6820 -1236
rect 4940 -1272 4996 -1262
rect 4932 -1284 4940 -1274
rect 5132 -1272 5188 -1262
rect 4996 -1284 5132 -1274
rect 5324 -1272 5380 -1262
rect 5188 -1284 5324 -1274
rect 5516 -1272 5572 -1262
rect 5380 -1284 5516 -1274
rect 5708 -1272 5764 -1262
rect 5572 -1284 5708 -1274
rect 5900 -1272 5956 -1262
rect 5764 -1284 5900 -1274
rect 6092 -1272 6148 -1262
rect 5956 -1456 6092 -1276
rect 6284 -1272 6340 -1262
rect 6148 -1456 6284 -1276
rect 6476 -1272 6532 -1262
rect 6340 -1456 6476 -1276
rect 6668 -1272 6724 -1262
rect 6532 -1456 6668 -1276
rect 6860 -1272 6916 -1262
rect 6724 -1456 6860 -1276
rect 5916 -1468 6916 -1456
rect 4932 -1482 5916 -1472
rect 6088 -1640 6960 -1630
rect 5032 -1672 6088 -1660
rect 5032 -1852 5036 -1672
rect 5092 -1852 5228 -1672
rect 5036 -1866 5092 -1856
rect 5284 -1852 5420 -1672
rect 5228 -1866 5284 -1856
rect 5476 -1852 5612 -1672
rect 5420 -1866 5476 -1856
rect 5668 -1852 5804 -1672
rect 5612 -1866 5668 -1856
rect 5860 -1852 5996 -1672
rect 5804 -1866 5860 -1856
rect 6052 -1840 6088 -1672
rect 6052 -1852 6188 -1840
rect 5996 -1866 6052 -1856
rect 6244 -1852 6380 -1840
rect 6188 -1866 6244 -1856
rect 6436 -1852 6572 -1840
rect 6380 -1866 6436 -1856
rect 6628 -1852 6764 -1840
rect 6572 -1866 6628 -1856
rect 6820 -1850 6960 -1840
rect 6820 -1852 6824 -1850
rect 6764 -1866 6820 -1856
rect 4940 -1892 4996 -1882
rect 4936 -1898 4940 -1896
rect 4928 -1908 4940 -1898
rect 5132 -1892 5188 -1882
rect 4996 -1908 5132 -1896
rect 5324 -1892 5380 -1882
rect 5188 -1908 5324 -1896
rect 5516 -1892 5572 -1882
rect 5380 -1908 5516 -1896
rect 5708 -1892 5764 -1882
rect 5572 -1908 5708 -1896
rect 5900 -1892 5956 -1882
rect 5764 -1908 5900 -1896
rect 6092 -1892 6148 -1882
rect 5956 -2076 6092 -1896
rect 6284 -1892 6340 -1882
rect 6148 -2076 6284 -1896
rect 6476 -1892 6532 -1882
rect 6340 -2076 6476 -1896
rect 6668 -1892 6724 -1882
rect 6532 -2076 6668 -1896
rect 6860 -1892 6916 -1882
rect 6724 -2076 6860 -1896
rect 5912 -2088 6916 -2076
rect 4928 -2106 5912 -2096
rect 6084 -2260 6956 -2250
rect 5032 -2288 6084 -2276
rect 5032 -2468 5036 -2288
rect 5092 -2468 5228 -2288
rect 5036 -2482 5092 -2472
rect 5284 -2468 5420 -2288
rect 5228 -2482 5284 -2472
rect 5476 -2468 5612 -2288
rect 5420 -2482 5476 -2472
rect 5668 -2468 5804 -2288
rect 5612 -2482 5668 -2472
rect 5860 -2468 5996 -2288
rect 5804 -2482 5860 -2472
rect 6052 -2460 6084 -2288
rect 6052 -2468 6188 -2460
rect 6084 -2470 6188 -2468
rect 5996 -2482 6052 -2472
rect 6244 -2470 6380 -2460
rect 6188 -2482 6244 -2472
rect 6436 -2470 6572 -2460
rect 6380 -2482 6436 -2472
rect 6628 -2470 6764 -2460
rect 6572 -2482 6628 -2472
rect 6820 -2470 6956 -2460
rect 6764 -2482 6820 -2472
rect 4940 -2508 4996 -2498
rect 4928 -2520 4940 -2510
rect 5132 -2508 5188 -2498
rect 4996 -2520 5132 -2510
rect 5324 -2508 5380 -2498
rect 5188 -2520 5324 -2510
rect 5516 -2508 5572 -2498
rect 5380 -2520 5516 -2510
rect 5708 -2508 5764 -2498
rect 5572 -2520 5708 -2510
rect 5900 -2508 5956 -2498
rect 5764 -2520 5900 -2510
rect 6092 -2508 6148 -2498
rect 5956 -2692 6092 -2512
rect 6284 -2508 6340 -2498
rect 6148 -2692 6284 -2512
rect 6476 -2508 6532 -2498
rect 6340 -2692 6476 -2512
rect 6668 -2508 6724 -2498
rect 6532 -2692 6668 -2512
rect 6860 -2508 6916 -2498
rect 6724 -2692 6860 -2512
rect 5912 -2704 6916 -2692
rect 4928 -2718 5912 -2708
rect 6084 -2880 6956 -2870
rect 5032 -2908 6084 -2896
rect 5032 -3088 5036 -2908
rect 5092 -3088 5228 -2908
rect 5036 -3102 5092 -3092
rect 5284 -3088 5420 -2908
rect 5228 -3102 5284 -3092
rect 5476 -3088 5612 -2908
rect 5420 -3102 5476 -3092
rect 5668 -3088 5804 -2908
rect 5612 -3102 5668 -3092
rect 5860 -3088 5996 -2908
rect 5804 -3102 5860 -3092
rect 6052 -3080 6084 -2908
rect 6052 -3088 6188 -3080
rect 6084 -3090 6188 -3088
rect 5996 -3102 6052 -3092
rect 6244 -3090 6380 -3080
rect 6188 -3102 6244 -3092
rect 6436 -3090 6572 -3080
rect 6380 -3102 6436 -3092
rect 6628 -3090 6764 -3080
rect 6572 -3102 6628 -3092
rect 6820 -3090 6956 -3080
rect 6764 -3102 6820 -3092
rect 4940 -3128 4996 -3118
rect 4936 -3134 4940 -3132
rect 4928 -3144 4940 -3134
rect 5132 -3128 5188 -3118
rect 4996 -3144 5132 -3132
rect 5324 -3128 5380 -3118
rect 5188 -3144 5324 -3132
rect 5516 -3128 5572 -3118
rect 5380 -3144 5516 -3132
rect 5708 -3128 5764 -3118
rect 5572 -3144 5708 -3132
rect 5900 -3128 5956 -3118
rect 5764 -3144 5900 -3132
rect 6092 -3128 6148 -3118
rect 5956 -3312 6092 -3132
rect 6284 -3128 6340 -3118
rect 6148 -3312 6284 -3132
rect 6476 -3128 6532 -3118
rect 6340 -3312 6476 -3132
rect 6668 -3128 6724 -3118
rect 6532 -3312 6668 -3132
rect 6860 -3128 6916 -3118
rect 6724 -3312 6860 -3132
rect 5912 -3324 6916 -3312
rect 4928 -3342 5912 -3332
<< via2 >>
rect 6084 2036 6956 2064
rect 6084 1864 6188 2036
rect 6188 1864 6244 2036
rect 6244 1864 6380 2036
rect 6380 1864 6436 2036
rect 6436 1864 6572 2036
rect 6572 1864 6628 2036
rect 6628 1864 6764 2036
rect 6764 1864 6820 2036
rect 6820 1864 6956 2036
rect 4932 1632 4940 1804
rect 4940 1632 4996 1804
rect 4996 1632 5132 1804
rect 5132 1632 5188 1804
rect 5188 1632 5324 1804
rect 5324 1632 5380 1804
rect 5380 1632 5516 1804
rect 5516 1632 5572 1804
rect 5572 1632 5708 1804
rect 5708 1632 5764 1804
rect 5764 1632 5900 1804
rect 5900 1632 5916 1804
rect 4932 1616 5916 1632
rect 6088 1420 6960 1448
rect 6088 1248 6188 1420
rect 6188 1248 6244 1420
rect 6244 1248 6380 1420
rect 6380 1248 6436 1420
rect 6436 1248 6572 1420
rect 6572 1248 6628 1420
rect 6628 1248 6764 1420
rect 6764 1248 6820 1420
rect 6820 1248 6960 1420
rect 4936 1016 4940 1184
rect 4940 1016 4996 1184
rect 4996 1016 5132 1184
rect 5132 1016 5188 1184
rect 5188 1016 5324 1184
rect 5324 1016 5380 1184
rect 5380 1016 5516 1184
rect 5516 1016 5572 1184
rect 5572 1016 5708 1184
rect 5708 1016 5764 1184
rect 5764 1016 5900 1184
rect 5900 1016 5920 1184
rect 4936 996 5920 1016
rect 6088 800 6960 832
rect 6088 632 6188 800
rect 6188 632 6244 800
rect 6244 632 6380 800
rect 6380 632 6436 800
rect 6436 632 6572 800
rect 6572 632 6628 800
rect 6628 632 6764 800
rect 6764 632 6820 800
rect 6820 632 6960 800
rect 4932 396 4940 568
rect 4940 396 4996 568
rect 4996 396 5132 568
rect 5132 396 5188 568
rect 5188 396 5324 568
rect 5324 396 5380 568
rect 5380 396 5516 568
rect 5516 396 5572 568
rect 5572 396 5708 568
rect 5708 396 5764 568
rect 5764 396 5900 568
rect 5900 396 5916 568
rect 4932 380 5916 396
rect 6088 184 6960 212
rect 6088 12 6188 184
rect 6188 12 6244 184
rect 6244 12 6380 184
rect 6380 12 6436 184
rect 6436 12 6572 184
rect 6572 12 6628 184
rect 6628 12 6764 184
rect 6764 12 6820 184
rect 6820 12 6960 184
rect 4928 -220 4940 -48
rect 4940 -220 4996 -48
rect 4996 -220 5132 -48
rect 5132 -220 5188 -48
rect 5188 -220 5324 -48
rect 5324 -220 5380 -48
rect 5380 -220 5516 -48
rect 5516 -220 5572 -48
rect 5572 -220 5708 -48
rect 5708 -220 5764 -48
rect 5764 -220 5900 -48
rect 5900 -220 5912 -48
rect 4928 -236 5912 -220
rect 6088 -436 6960 -408
rect 6088 -608 6188 -436
rect 6188 -608 6244 -436
rect 6244 -608 6380 -436
rect 6380 -608 6436 -436
rect 6436 -608 6572 -436
rect 6572 -608 6628 -436
rect 6628 -608 6764 -436
rect 6764 -608 6820 -436
rect 6820 -608 6960 -436
rect 4932 -840 4940 -672
rect 4940 -840 4996 -672
rect 4996 -840 5132 -672
rect 5132 -840 5188 -672
rect 5188 -840 5324 -672
rect 5324 -840 5380 -672
rect 5380 -840 5516 -672
rect 5516 -840 5572 -672
rect 5572 -840 5708 -672
rect 5708 -840 5764 -672
rect 5764 -840 5900 -672
rect 5900 -840 5916 -672
rect 4932 -860 5916 -840
rect 6088 -1052 6960 -1024
rect 6088 -1224 6188 -1052
rect 6188 -1224 6244 -1052
rect 6244 -1224 6380 -1052
rect 6380 -1224 6436 -1052
rect 6436 -1224 6572 -1052
rect 6572 -1224 6628 -1052
rect 6628 -1224 6764 -1052
rect 6764 -1224 6820 -1052
rect 6820 -1224 6960 -1052
rect 4932 -1456 4940 -1284
rect 4940 -1456 4996 -1284
rect 4996 -1456 5132 -1284
rect 5132 -1456 5188 -1284
rect 5188 -1456 5324 -1284
rect 5324 -1456 5380 -1284
rect 5380 -1456 5516 -1284
rect 5516 -1456 5572 -1284
rect 5572 -1456 5708 -1284
rect 5708 -1456 5764 -1284
rect 5764 -1456 5900 -1284
rect 5900 -1456 5916 -1284
rect 4932 -1472 5916 -1456
rect 6088 -1672 6960 -1640
rect 6088 -1840 6188 -1672
rect 6188 -1840 6244 -1672
rect 6244 -1840 6380 -1672
rect 6380 -1840 6436 -1672
rect 6436 -1840 6572 -1672
rect 6572 -1840 6628 -1672
rect 6628 -1840 6764 -1672
rect 6764 -1840 6820 -1672
rect 6820 -1840 6960 -1672
rect 4928 -2076 4940 -1908
rect 4940 -2076 4996 -1908
rect 4996 -2076 5132 -1908
rect 5132 -2076 5188 -1908
rect 5188 -2076 5324 -1908
rect 5324 -2076 5380 -1908
rect 5380 -2076 5516 -1908
rect 5516 -2076 5572 -1908
rect 5572 -2076 5708 -1908
rect 5708 -2076 5764 -1908
rect 5764 -2076 5900 -1908
rect 5900 -2076 5912 -1908
rect 4928 -2096 5912 -2076
rect 6084 -2288 6956 -2260
rect 6084 -2460 6188 -2288
rect 6188 -2460 6244 -2288
rect 6244 -2460 6380 -2288
rect 6380 -2460 6436 -2288
rect 6436 -2460 6572 -2288
rect 6572 -2460 6628 -2288
rect 6628 -2460 6764 -2288
rect 6764 -2460 6820 -2288
rect 6820 -2460 6956 -2288
rect 4928 -2692 4940 -2520
rect 4940 -2692 4996 -2520
rect 4996 -2692 5132 -2520
rect 5132 -2692 5188 -2520
rect 5188 -2692 5324 -2520
rect 5324 -2692 5380 -2520
rect 5380 -2692 5516 -2520
rect 5516 -2692 5572 -2520
rect 5572 -2692 5708 -2520
rect 5708 -2692 5764 -2520
rect 5764 -2692 5900 -2520
rect 5900 -2692 5912 -2520
rect 4928 -2708 5912 -2692
rect 6084 -2908 6956 -2880
rect 6084 -3080 6188 -2908
rect 6188 -3080 6244 -2908
rect 6244 -3080 6380 -2908
rect 6380 -3080 6436 -2908
rect 6436 -3080 6572 -2908
rect 6572 -3080 6628 -2908
rect 6628 -3080 6764 -2908
rect 6764 -3080 6820 -2908
rect 6820 -3080 6956 -2908
rect 4928 -3312 4940 -3144
rect 4940 -3312 4996 -3144
rect 4996 -3312 5132 -3144
rect 5132 -3312 5188 -3144
rect 5188 -3312 5324 -3144
rect 5324 -3312 5380 -3144
rect 5380 -3312 5516 -3144
rect 5516 -3312 5572 -3144
rect 5572 -3312 5708 -3144
rect 5708 -3312 5764 -3144
rect 5764 -3312 5900 -3144
rect 5900 -3312 5912 -3144
rect 4928 -3332 5912 -3312
<< metal3 >>
rect 6074 2064 6966 2069
rect 6074 1864 6084 2064
rect 6956 1864 6966 2064
rect 6074 1859 6966 1864
rect 4924 1809 5924 1812
rect 4922 1804 5926 1809
rect 4922 1616 4932 1804
rect 5916 1616 5926 1804
rect 4922 1611 5926 1616
rect 4924 1189 5924 1611
rect 6084 1453 6960 1859
rect 6078 1448 6970 1453
rect 6078 1248 6088 1448
rect 6960 1248 6970 1448
rect 6078 1243 6970 1248
rect 4924 1184 5930 1189
rect 4924 996 4936 1184
rect 5920 996 5930 1184
rect 4924 991 5930 996
rect 4924 573 5924 991
rect 6084 837 6960 1243
rect 6078 832 6970 837
rect 6078 632 6088 832
rect 6960 632 6970 832
rect 6078 627 6970 632
rect 4922 568 5926 573
rect 4922 380 4932 568
rect 5916 380 5926 568
rect 4922 375 5926 380
rect 4922 -48 5924 375
rect 6084 217 6960 627
rect 6078 212 6970 217
rect 6078 12 6088 212
rect 6960 12 6970 212
rect 6078 7 6970 12
rect 4922 -236 4928 -48
rect 5912 -236 5924 -48
rect 4922 -324 5924 -236
rect 4924 -667 5924 -324
rect 6084 -403 6960 7
rect 6078 -408 6970 -403
rect 6078 -608 6088 -408
rect 6960 -608 6970 -408
rect 6078 -613 6970 -608
rect 4922 -672 5926 -667
rect 4922 -860 4932 -672
rect 5916 -860 5926 -672
rect 4922 -865 5926 -860
rect 4924 -1279 5924 -865
rect 6084 -1019 6960 -613
rect 6078 -1024 6970 -1019
rect 6078 -1224 6088 -1024
rect 6960 -1224 6970 -1024
rect 6078 -1229 6970 -1224
rect 4922 -1284 5926 -1279
rect 4922 -1472 4932 -1284
rect 5916 -1472 5926 -1284
rect 4922 -1477 5926 -1472
rect 4924 -1903 5924 -1477
rect 6084 -1635 6960 -1229
rect 6078 -1640 6970 -1635
rect 6078 -1840 6088 -1640
rect 6960 -1840 6970 -1640
rect 6078 -1845 6970 -1840
rect 4918 -1908 5924 -1903
rect 4918 -2096 4928 -1908
rect 5912 -2096 5924 -1908
rect 4918 -2101 5924 -2096
rect 4924 -2515 5924 -2101
rect 6084 -2255 6960 -1845
rect 6074 -2260 6966 -2255
rect 6074 -2460 6084 -2260
rect 6956 -2460 6966 -2260
rect 6074 -2465 6966 -2460
rect 4918 -2520 5924 -2515
rect 4918 -2708 4928 -2520
rect 5912 -2708 5924 -2520
rect 4918 -2713 5924 -2708
rect 4924 -3139 5924 -2713
rect 6084 -2875 6960 -2465
rect 6074 -2880 6966 -2875
rect 6074 -3080 6084 -2880
rect 6956 -3080 6966 -2880
rect 6074 -3085 6966 -3080
rect 6084 -3088 6960 -3085
rect 4918 -3144 5924 -3139
rect 4918 -3332 4928 -3144
rect 5912 -3324 5924 -3144
rect 5912 -3332 5922 -3324
rect 4918 -3337 5922 -3332
use sky130_fd_pr__nfet_01v8_lvt_S9AFLJ  sky130_fd_pr__nfet_01v8_lvt_S9AFLJ_1
timestamp 1686659968
transform 1 0 5927 0 1 -638
box -1127 -2882 1127 2882
<< end >>
