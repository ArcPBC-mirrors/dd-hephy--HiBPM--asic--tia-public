magic
tech sky130A
magscale 1 2
timestamp 1683553776
<< nwell >>
rect -562 -1373 562 1373
<< pmos >>
rect -366 754 -266 1154
rect -208 754 -108 1154
rect -50 754 50 1154
rect 108 754 208 1154
rect 266 754 366 1154
rect -366 118 -266 518
rect -208 118 -108 518
rect -50 118 50 518
rect 108 118 208 518
rect 266 118 366 518
rect -366 -518 -266 -118
rect -208 -518 -108 -118
rect -50 -518 50 -118
rect 108 -518 208 -118
rect 266 -518 366 -118
rect -366 -1154 -266 -754
rect -208 -1154 -108 -754
rect -50 -1154 50 -754
rect 108 -1154 208 -754
rect 266 -1154 366 -754
<< pdiff >>
rect -424 1142 -366 1154
rect -424 766 -412 1142
rect -378 766 -366 1142
rect -424 754 -366 766
rect -266 1142 -208 1154
rect -266 766 -254 1142
rect -220 766 -208 1142
rect -266 754 -208 766
rect -108 1142 -50 1154
rect -108 766 -96 1142
rect -62 766 -50 1142
rect -108 754 -50 766
rect 50 1142 108 1154
rect 50 766 62 1142
rect 96 766 108 1142
rect 50 754 108 766
rect 208 1142 266 1154
rect 208 766 220 1142
rect 254 766 266 1142
rect 208 754 266 766
rect 366 1142 424 1154
rect 366 766 378 1142
rect 412 766 424 1142
rect 366 754 424 766
rect -424 506 -366 518
rect -424 130 -412 506
rect -378 130 -366 506
rect -424 118 -366 130
rect -266 506 -208 518
rect -266 130 -254 506
rect -220 130 -208 506
rect -266 118 -208 130
rect -108 506 -50 518
rect -108 130 -96 506
rect -62 130 -50 506
rect -108 118 -50 130
rect 50 506 108 518
rect 50 130 62 506
rect 96 130 108 506
rect 50 118 108 130
rect 208 506 266 518
rect 208 130 220 506
rect 254 130 266 506
rect 208 118 266 130
rect 366 506 424 518
rect 366 130 378 506
rect 412 130 424 506
rect 366 118 424 130
rect -424 -130 -366 -118
rect -424 -506 -412 -130
rect -378 -506 -366 -130
rect -424 -518 -366 -506
rect -266 -130 -208 -118
rect -266 -506 -254 -130
rect -220 -506 -208 -130
rect -266 -518 -208 -506
rect -108 -130 -50 -118
rect -108 -506 -96 -130
rect -62 -506 -50 -130
rect -108 -518 -50 -506
rect 50 -130 108 -118
rect 50 -506 62 -130
rect 96 -506 108 -130
rect 50 -518 108 -506
rect 208 -130 266 -118
rect 208 -506 220 -130
rect 254 -506 266 -130
rect 208 -518 266 -506
rect 366 -130 424 -118
rect 366 -506 378 -130
rect 412 -506 424 -130
rect 366 -518 424 -506
rect -424 -766 -366 -754
rect -424 -1142 -412 -766
rect -378 -1142 -366 -766
rect -424 -1154 -366 -1142
rect -266 -766 -208 -754
rect -266 -1142 -254 -766
rect -220 -1142 -208 -766
rect -266 -1154 -208 -1142
rect -108 -766 -50 -754
rect -108 -1142 -96 -766
rect -62 -1142 -50 -766
rect -108 -1154 -50 -1142
rect 50 -766 108 -754
rect 50 -1142 62 -766
rect 96 -1142 108 -766
rect 50 -1154 108 -1142
rect 208 -766 266 -754
rect 208 -1142 220 -766
rect 254 -1142 266 -766
rect 208 -1154 266 -1142
rect 366 -766 424 -754
rect 366 -1142 378 -766
rect 412 -1142 424 -766
rect 366 -1154 424 -1142
<< pdiffc >>
rect -412 766 -378 1142
rect -254 766 -220 1142
rect -96 766 -62 1142
rect 62 766 96 1142
rect 220 766 254 1142
rect 378 766 412 1142
rect -412 130 -378 506
rect -254 130 -220 506
rect -96 130 -62 506
rect 62 130 96 506
rect 220 130 254 506
rect 378 130 412 506
rect -412 -506 -378 -130
rect -254 -506 -220 -130
rect -96 -506 -62 -130
rect 62 -506 96 -130
rect 220 -506 254 -130
rect 378 -506 412 -130
rect -412 -1142 -378 -766
rect -254 -1142 -220 -766
rect -96 -1142 -62 -766
rect 62 -1142 96 -766
rect 220 -1142 254 -766
rect 378 -1142 412 -766
<< nsubdiff >>
rect -526 1303 -430 1337
rect 430 1303 526 1337
rect -526 1241 -492 1303
rect 492 1241 526 1303
rect -526 -1303 -492 -1241
rect 492 -1303 526 -1241
rect -526 -1337 -430 -1303
rect 430 -1337 526 -1303
<< nsubdiffcont >>
rect -430 1303 430 1337
rect -526 -1241 -492 1241
rect 492 -1241 526 1241
rect -430 -1337 430 -1303
<< poly >>
rect -366 1235 -266 1251
rect -366 1201 -350 1235
rect -282 1201 -266 1235
rect -366 1154 -266 1201
rect -208 1235 -108 1251
rect -208 1201 -192 1235
rect -124 1201 -108 1235
rect -208 1154 -108 1201
rect -50 1235 50 1251
rect -50 1201 -34 1235
rect 34 1201 50 1235
rect -50 1154 50 1201
rect 108 1235 208 1251
rect 108 1201 124 1235
rect 192 1201 208 1235
rect 108 1154 208 1201
rect 266 1235 366 1251
rect 266 1201 282 1235
rect 350 1201 366 1235
rect 266 1154 366 1201
rect -366 707 -266 754
rect -366 673 -350 707
rect -282 673 -266 707
rect -366 657 -266 673
rect -208 707 -108 754
rect -208 673 -192 707
rect -124 673 -108 707
rect -208 657 -108 673
rect -50 707 50 754
rect -50 673 -34 707
rect 34 673 50 707
rect -50 657 50 673
rect 108 707 208 754
rect 108 673 124 707
rect 192 673 208 707
rect 108 657 208 673
rect 266 707 366 754
rect 266 673 282 707
rect 350 673 366 707
rect 266 657 366 673
rect -366 599 -266 615
rect -366 565 -350 599
rect -282 565 -266 599
rect -366 518 -266 565
rect -208 599 -108 615
rect -208 565 -192 599
rect -124 565 -108 599
rect -208 518 -108 565
rect -50 599 50 615
rect -50 565 -34 599
rect 34 565 50 599
rect -50 518 50 565
rect 108 599 208 615
rect 108 565 124 599
rect 192 565 208 599
rect 108 518 208 565
rect 266 599 366 615
rect 266 565 282 599
rect 350 565 366 599
rect 266 518 366 565
rect -366 71 -266 118
rect -366 37 -350 71
rect -282 37 -266 71
rect -366 21 -266 37
rect -208 71 -108 118
rect -208 37 -192 71
rect -124 37 -108 71
rect -208 21 -108 37
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect 108 71 208 118
rect 108 37 124 71
rect 192 37 208 71
rect 108 21 208 37
rect 266 71 366 118
rect 266 37 282 71
rect 350 37 366 71
rect 266 21 366 37
rect -366 -37 -266 -21
rect -366 -71 -350 -37
rect -282 -71 -266 -37
rect -366 -118 -266 -71
rect -208 -37 -108 -21
rect -208 -71 -192 -37
rect -124 -71 -108 -37
rect -208 -118 -108 -71
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect 108 -37 208 -21
rect 108 -71 124 -37
rect 192 -71 208 -37
rect 108 -118 208 -71
rect 266 -37 366 -21
rect 266 -71 282 -37
rect 350 -71 366 -37
rect 266 -118 366 -71
rect -366 -565 -266 -518
rect -366 -599 -350 -565
rect -282 -599 -266 -565
rect -366 -615 -266 -599
rect -208 -565 -108 -518
rect -208 -599 -192 -565
rect -124 -599 -108 -565
rect -208 -615 -108 -599
rect -50 -565 50 -518
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -50 -615 50 -599
rect 108 -565 208 -518
rect 108 -599 124 -565
rect 192 -599 208 -565
rect 108 -615 208 -599
rect 266 -565 366 -518
rect 266 -599 282 -565
rect 350 -599 366 -565
rect 266 -615 366 -599
rect -366 -673 -266 -657
rect -366 -707 -350 -673
rect -282 -707 -266 -673
rect -366 -754 -266 -707
rect -208 -673 -108 -657
rect -208 -707 -192 -673
rect -124 -707 -108 -673
rect -208 -754 -108 -707
rect -50 -673 50 -657
rect -50 -707 -34 -673
rect 34 -707 50 -673
rect -50 -754 50 -707
rect 108 -673 208 -657
rect 108 -707 124 -673
rect 192 -707 208 -673
rect 108 -754 208 -707
rect 266 -673 366 -657
rect 266 -707 282 -673
rect 350 -707 366 -673
rect 266 -754 366 -707
rect -366 -1201 -266 -1154
rect -366 -1235 -350 -1201
rect -282 -1235 -266 -1201
rect -366 -1251 -266 -1235
rect -208 -1201 -108 -1154
rect -208 -1235 -192 -1201
rect -124 -1235 -108 -1201
rect -208 -1251 -108 -1235
rect -50 -1201 50 -1154
rect -50 -1235 -34 -1201
rect 34 -1235 50 -1201
rect -50 -1251 50 -1235
rect 108 -1201 208 -1154
rect 108 -1235 124 -1201
rect 192 -1235 208 -1201
rect 108 -1251 208 -1235
rect 266 -1201 366 -1154
rect 266 -1235 282 -1201
rect 350 -1235 366 -1201
rect 266 -1251 366 -1235
<< polycont >>
rect -350 1201 -282 1235
rect -192 1201 -124 1235
rect -34 1201 34 1235
rect 124 1201 192 1235
rect 282 1201 350 1235
rect -350 673 -282 707
rect -192 673 -124 707
rect -34 673 34 707
rect 124 673 192 707
rect 282 673 350 707
rect -350 565 -282 599
rect -192 565 -124 599
rect -34 565 34 599
rect 124 565 192 599
rect 282 565 350 599
rect -350 37 -282 71
rect -192 37 -124 71
rect -34 37 34 71
rect 124 37 192 71
rect 282 37 350 71
rect -350 -71 -282 -37
rect -192 -71 -124 -37
rect -34 -71 34 -37
rect 124 -71 192 -37
rect 282 -71 350 -37
rect -350 -599 -282 -565
rect -192 -599 -124 -565
rect -34 -599 34 -565
rect 124 -599 192 -565
rect 282 -599 350 -565
rect -350 -707 -282 -673
rect -192 -707 -124 -673
rect -34 -707 34 -673
rect 124 -707 192 -673
rect 282 -707 350 -673
rect -350 -1235 -282 -1201
rect -192 -1235 -124 -1201
rect -34 -1235 34 -1201
rect 124 -1235 192 -1201
rect 282 -1235 350 -1201
<< locali >>
rect -526 1303 -430 1337
rect 430 1303 526 1337
rect -526 1241 -492 1303
rect 492 1241 526 1303
rect -366 1201 -350 1235
rect -282 1201 -266 1235
rect -208 1201 -192 1235
rect -124 1201 -108 1235
rect -50 1201 -34 1235
rect 34 1201 50 1235
rect 108 1201 124 1235
rect 192 1201 208 1235
rect 266 1201 282 1235
rect 350 1201 366 1235
rect -412 1142 -378 1158
rect -412 750 -378 766
rect -254 1142 -220 1158
rect -254 750 -220 766
rect -96 1142 -62 1158
rect -96 750 -62 766
rect 62 1142 96 1158
rect 62 750 96 766
rect 220 1142 254 1158
rect 220 750 254 766
rect 378 1142 412 1158
rect 378 750 412 766
rect -366 673 -350 707
rect -282 673 -266 707
rect -208 673 -192 707
rect -124 673 -108 707
rect -50 673 -34 707
rect 34 673 50 707
rect 108 673 124 707
rect 192 673 208 707
rect 266 673 282 707
rect 350 673 366 707
rect -366 565 -350 599
rect -282 565 -266 599
rect -208 565 -192 599
rect -124 565 -108 599
rect -50 565 -34 599
rect 34 565 50 599
rect 108 565 124 599
rect 192 565 208 599
rect 266 565 282 599
rect 350 565 366 599
rect -412 506 -378 522
rect -412 114 -378 130
rect -254 506 -220 522
rect -254 114 -220 130
rect -96 506 -62 522
rect -96 114 -62 130
rect 62 506 96 522
rect 62 114 96 130
rect 220 506 254 522
rect 220 114 254 130
rect 378 506 412 522
rect 378 114 412 130
rect -366 37 -350 71
rect -282 37 -266 71
rect -208 37 -192 71
rect -124 37 -108 71
rect -50 37 -34 71
rect 34 37 50 71
rect 108 37 124 71
rect 192 37 208 71
rect 266 37 282 71
rect 350 37 366 71
rect -366 -71 -350 -37
rect -282 -71 -266 -37
rect -208 -71 -192 -37
rect -124 -71 -108 -37
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect 108 -71 124 -37
rect 192 -71 208 -37
rect 266 -71 282 -37
rect 350 -71 366 -37
rect -412 -130 -378 -114
rect -412 -522 -378 -506
rect -254 -130 -220 -114
rect -254 -522 -220 -506
rect -96 -130 -62 -114
rect -96 -522 -62 -506
rect 62 -130 96 -114
rect 62 -522 96 -506
rect 220 -130 254 -114
rect 220 -522 254 -506
rect 378 -130 412 -114
rect 378 -522 412 -506
rect -366 -599 -350 -565
rect -282 -599 -266 -565
rect -208 -599 -192 -565
rect -124 -599 -108 -565
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect 108 -599 124 -565
rect 192 -599 208 -565
rect 266 -599 282 -565
rect 350 -599 366 -565
rect -366 -707 -350 -673
rect -282 -707 -266 -673
rect -208 -707 -192 -673
rect -124 -707 -108 -673
rect -50 -707 -34 -673
rect 34 -707 50 -673
rect 108 -707 124 -673
rect 192 -707 208 -673
rect 266 -707 282 -673
rect 350 -707 366 -673
rect -412 -766 -378 -750
rect -412 -1158 -378 -1142
rect -254 -766 -220 -750
rect -254 -1158 -220 -1142
rect -96 -766 -62 -750
rect -96 -1158 -62 -1142
rect 62 -766 96 -750
rect 62 -1158 96 -1142
rect 220 -766 254 -750
rect 220 -1158 254 -1142
rect 378 -766 412 -750
rect 378 -1158 412 -1142
rect -366 -1235 -350 -1201
rect -282 -1235 -266 -1201
rect -208 -1235 -192 -1201
rect -124 -1235 -108 -1201
rect -50 -1235 -34 -1201
rect 34 -1235 50 -1201
rect 108 -1235 124 -1201
rect 192 -1235 208 -1201
rect 266 -1235 282 -1201
rect 350 -1235 366 -1201
rect -526 -1303 -492 -1241
rect 492 -1303 526 -1241
rect -526 -1337 -430 -1303
rect 430 -1337 526 -1303
<< viali >>
rect -350 1201 -282 1235
rect -192 1201 -124 1235
rect -34 1201 34 1235
rect 124 1201 192 1235
rect 282 1201 350 1235
rect -412 766 -378 1142
rect -254 766 -220 1142
rect -96 766 -62 1142
rect 62 766 96 1142
rect 220 766 254 1142
rect 378 766 412 1142
rect -350 673 -282 707
rect -192 673 -124 707
rect -34 673 34 707
rect 124 673 192 707
rect 282 673 350 707
rect -350 565 -282 599
rect -192 565 -124 599
rect -34 565 34 599
rect 124 565 192 599
rect 282 565 350 599
rect -412 130 -378 506
rect -254 130 -220 506
rect -96 130 -62 506
rect 62 130 96 506
rect 220 130 254 506
rect 378 130 412 506
rect -350 37 -282 71
rect -192 37 -124 71
rect -34 37 34 71
rect 124 37 192 71
rect 282 37 350 71
rect -350 -71 -282 -37
rect -192 -71 -124 -37
rect -34 -71 34 -37
rect 124 -71 192 -37
rect 282 -71 350 -37
rect -412 -506 -378 -130
rect -254 -506 -220 -130
rect -96 -506 -62 -130
rect 62 -506 96 -130
rect 220 -506 254 -130
rect 378 -506 412 -130
rect -350 -599 -282 -565
rect -192 -599 -124 -565
rect -34 -599 34 -565
rect 124 -599 192 -565
rect 282 -599 350 -565
rect -350 -707 -282 -673
rect -192 -707 -124 -673
rect -34 -707 34 -673
rect 124 -707 192 -673
rect 282 -707 350 -673
rect -412 -1142 -378 -766
rect -254 -1142 -220 -766
rect -96 -1142 -62 -766
rect 62 -1142 96 -766
rect 220 -1142 254 -766
rect 378 -1142 412 -766
rect -350 -1235 -282 -1201
rect -192 -1235 -124 -1201
rect -34 -1235 34 -1201
rect 124 -1235 192 -1201
rect 282 -1235 350 -1201
<< metal1 >>
rect -362 1235 -270 1241
rect -362 1201 -350 1235
rect -282 1201 -270 1235
rect -362 1195 -270 1201
rect -204 1235 -112 1241
rect -204 1201 -192 1235
rect -124 1201 -112 1235
rect -204 1195 -112 1201
rect -46 1235 46 1241
rect -46 1201 -34 1235
rect 34 1201 46 1235
rect -46 1195 46 1201
rect 112 1235 204 1241
rect 112 1201 124 1235
rect 192 1201 204 1235
rect 112 1195 204 1201
rect 270 1235 362 1241
rect 270 1201 282 1235
rect 350 1201 362 1235
rect 270 1195 362 1201
rect -418 1142 -372 1154
rect -418 766 -412 1142
rect -378 766 -372 1142
rect -418 754 -372 766
rect -260 1142 -214 1154
rect -260 766 -254 1142
rect -220 766 -214 1142
rect -260 754 -214 766
rect -102 1142 -56 1154
rect -102 766 -96 1142
rect -62 766 -56 1142
rect -102 754 -56 766
rect 56 1142 102 1154
rect 56 766 62 1142
rect 96 766 102 1142
rect 56 754 102 766
rect 214 1142 260 1154
rect 214 766 220 1142
rect 254 766 260 1142
rect 214 754 260 766
rect 372 1142 418 1154
rect 372 766 378 1142
rect 412 766 418 1142
rect 372 754 418 766
rect -362 707 -270 713
rect -362 673 -350 707
rect -282 673 -270 707
rect -362 667 -270 673
rect -204 707 -112 713
rect -204 673 -192 707
rect -124 673 -112 707
rect -204 667 -112 673
rect -46 707 46 713
rect -46 673 -34 707
rect 34 673 46 707
rect -46 667 46 673
rect 112 707 204 713
rect 112 673 124 707
rect 192 673 204 707
rect 112 667 204 673
rect 270 707 362 713
rect 270 673 282 707
rect 350 673 362 707
rect 270 667 362 673
rect -362 599 -270 605
rect -362 565 -350 599
rect -282 565 -270 599
rect -362 559 -270 565
rect -204 599 -112 605
rect -204 565 -192 599
rect -124 565 -112 599
rect -204 559 -112 565
rect -46 599 46 605
rect -46 565 -34 599
rect 34 565 46 599
rect -46 559 46 565
rect 112 599 204 605
rect 112 565 124 599
rect 192 565 204 599
rect 112 559 204 565
rect 270 599 362 605
rect 270 565 282 599
rect 350 565 362 599
rect 270 559 362 565
rect -418 506 -372 518
rect -418 130 -412 506
rect -378 130 -372 506
rect -418 118 -372 130
rect -260 506 -214 518
rect -260 130 -254 506
rect -220 130 -214 506
rect -260 118 -214 130
rect -102 506 -56 518
rect -102 130 -96 506
rect -62 130 -56 506
rect -102 118 -56 130
rect 56 506 102 518
rect 56 130 62 506
rect 96 130 102 506
rect 56 118 102 130
rect 214 506 260 518
rect 214 130 220 506
rect 254 130 260 506
rect 214 118 260 130
rect 372 506 418 518
rect 372 130 378 506
rect 412 130 418 506
rect 372 118 418 130
rect -362 71 -270 77
rect -362 37 -350 71
rect -282 37 -270 71
rect -362 31 -270 37
rect -204 71 -112 77
rect -204 37 -192 71
rect -124 37 -112 71
rect -204 31 -112 37
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect 112 71 204 77
rect 112 37 124 71
rect 192 37 204 71
rect 112 31 204 37
rect 270 71 362 77
rect 270 37 282 71
rect 350 37 362 71
rect 270 31 362 37
rect -362 -37 -270 -31
rect -362 -71 -350 -37
rect -282 -71 -270 -37
rect -362 -77 -270 -71
rect -204 -37 -112 -31
rect -204 -71 -192 -37
rect -124 -71 -112 -37
rect -204 -77 -112 -71
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect 112 -37 204 -31
rect 112 -71 124 -37
rect 192 -71 204 -37
rect 112 -77 204 -71
rect 270 -37 362 -31
rect 270 -71 282 -37
rect 350 -71 362 -37
rect 270 -77 362 -71
rect -418 -130 -372 -118
rect -418 -506 -412 -130
rect -378 -506 -372 -130
rect -418 -518 -372 -506
rect -260 -130 -214 -118
rect -260 -506 -254 -130
rect -220 -506 -214 -130
rect -260 -518 -214 -506
rect -102 -130 -56 -118
rect -102 -506 -96 -130
rect -62 -506 -56 -130
rect -102 -518 -56 -506
rect 56 -130 102 -118
rect 56 -506 62 -130
rect 96 -506 102 -130
rect 56 -518 102 -506
rect 214 -130 260 -118
rect 214 -506 220 -130
rect 254 -506 260 -130
rect 214 -518 260 -506
rect 372 -130 418 -118
rect 372 -506 378 -130
rect 412 -506 418 -130
rect 372 -518 418 -506
rect -362 -565 -270 -559
rect -362 -599 -350 -565
rect -282 -599 -270 -565
rect -362 -605 -270 -599
rect -204 -565 -112 -559
rect -204 -599 -192 -565
rect -124 -599 -112 -565
rect -204 -605 -112 -599
rect -46 -565 46 -559
rect -46 -599 -34 -565
rect 34 -599 46 -565
rect -46 -605 46 -599
rect 112 -565 204 -559
rect 112 -599 124 -565
rect 192 -599 204 -565
rect 112 -605 204 -599
rect 270 -565 362 -559
rect 270 -599 282 -565
rect 350 -599 362 -565
rect 270 -605 362 -599
rect -362 -673 -270 -667
rect -362 -707 -350 -673
rect -282 -707 -270 -673
rect -362 -713 -270 -707
rect -204 -673 -112 -667
rect -204 -707 -192 -673
rect -124 -707 -112 -673
rect -204 -713 -112 -707
rect -46 -673 46 -667
rect -46 -707 -34 -673
rect 34 -707 46 -673
rect -46 -713 46 -707
rect 112 -673 204 -667
rect 112 -707 124 -673
rect 192 -707 204 -673
rect 112 -713 204 -707
rect 270 -673 362 -667
rect 270 -707 282 -673
rect 350 -707 362 -673
rect 270 -713 362 -707
rect -418 -766 -372 -754
rect -418 -1142 -412 -766
rect -378 -1142 -372 -766
rect -418 -1154 -372 -1142
rect -260 -766 -214 -754
rect -260 -1142 -254 -766
rect -220 -1142 -214 -766
rect -260 -1154 -214 -1142
rect -102 -766 -56 -754
rect -102 -1142 -96 -766
rect -62 -1142 -56 -766
rect -102 -1154 -56 -1142
rect 56 -766 102 -754
rect 56 -1142 62 -766
rect 96 -1142 102 -766
rect 56 -1154 102 -1142
rect 214 -766 260 -754
rect 214 -1142 220 -766
rect 254 -1142 260 -766
rect 214 -1154 260 -1142
rect 372 -766 418 -754
rect 372 -1142 378 -766
rect 412 -1142 418 -766
rect 372 -1154 418 -1142
rect -362 -1201 -270 -1195
rect -362 -1235 -350 -1201
rect -282 -1235 -270 -1201
rect -362 -1241 -270 -1235
rect -204 -1201 -112 -1195
rect -204 -1235 -192 -1201
rect -124 -1235 -112 -1201
rect -204 -1241 -112 -1235
rect -46 -1201 46 -1195
rect -46 -1235 -34 -1201
rect 34 -1235 46 -1201
rect -46 -1241 46 -1235
rect 112 -1201 204 -1195
rect 112 -1235 124 -1201
rect 192 -1235 204 -1201
rect 112 -1241 204 -1235
rect 270 -1201 362 -1195
rect 270 -1235 282 -1201
rect 350 -1235 362 -1201
rect 270 -1241 362 -1235
<< properties >>
string FIXED_BBOX -509 -1320 509 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.5 m 4 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
