magic
tech sky130A
magscale 1 2
timestamp 1683557511
<< nwell >>
rect -2913 1381 -1647 1963
rect -1393 1381 -127 1963
rect 127 1381 1393 1963
rect 1647 1381 2913 1963
rect -2913 545 -1647 1127
rect -1393 545 -127 1127
rect 127 545 1393 1127
rect 1647 545 2913 1127
rect -2913 -291 -1647 291
rect -1393 -291 -127 291
rect 127 -291 1393 291
rect 1647 -291 2913 291
rect -2913 -1127 -1647 -545
rect -1393 -1127 -127 -545
rect 127 -1127 1393 -545
rect 1647 -1127 2913 -545
rect -2913 -1963 -1647 -1381
rect -1393 -1963 -127 -1381
rect 127 -1963 1393 -1381
rect 1647 -1963 2913 -1381
<< pwell >>
rect -3023 1963 3023 2073
rect -3023 1381 -2913 1963
rect -1647 1381 -1393 1963
rect -127 1381 127 1963
rect 1393 1381 1647 1963
rect 2913 1381 3023 1963
rect -3023 1127 3023 1381
rect -3023 545 -2913 1127
rect -1647 545 -1393 1127
rect -127 545 127 1127
rect 1393 545 1647 1127
rect 2913 545 3023 1127
rect -3023 291 3023 545
rect -3023 -291 -2913 291
rect -1647 -291 -1393 291
rect -127 -291 127 291
rect 1393 -291 1647 291
rect 2913 -291 3023 291
rect -3023 -545 3023 -291
rect -3023 -1127 -2913 -545
rect -1647 -1127 -1393 -545
rect -127 -1127 127 -545
rect 1393 -1127 1647 -545
rect 2913 -1127 3023 -545
rect -3023 -1381 3023 -1127
rect -3023 -1963 -2913 -1381
rect -1647 -1963 -1393 -1381
rect -127 -1963 127 -1381
rect 1393 -1963 1647 -1381
rect 2913 -1963 3023 -1381
rect -3023 -2073 3023 -1963
<< varactor >>
rect -2780 1472 -1780 1872
rect -1260 1472 -260 1872
rect 260 1472 1260 1872
rect 1780 1472 2780 1872
rect -2780 636 -1780 1036
rect -1260 636 -260 1036
rect 260 636 1260 1036
rect 1780 636 2780 1036
rect -2780 -200 -1780 200
rect -1260 -200 -260 200
rect 260 -200 1260 200
rect 1780 -200 2780 200
rect -2780 -1036 -1780 -636
rect -1260 -1036 -260 -636
rect 260 -1036 1260 -636
rect 1780 -1036 2780 -636
rect -2780 -1872 -1780 -1472
rect -1260 -1872 -260 -1472
rect 260 -1872 1260 -1472
rect 1780 -1872 2780 -1472
<< psubdiff >>
rect -2987 2003 -2891 2037
rect 2891 2003 2987 2037
rect -2987 1941 -2953 2003
rect 2953 1941 2987 2003
rect -2987 -2003 -2953 -1941
rect 2953 -2003 2987 -1941
rect -2987 -2037 -2891 -2003
rect 2891 -2037 2987 -2003
<< nsubdiff >>
rect -2877 1848 -2780 1872
rect -2877 1496 -2865 1848
rect -2831 1496 -2780 1848
rect -2877 1472 -2780 1496
rect -1780 1848 -1683 1872
rect -1780 1496 -1729 1848
rect -1695 1496 -1683 1848
rect -1780 1472 -1683 1496
rect -1357 1848 -1260 1872
rect -1357 1496 -1345 1848
rect -1311 1496 -1260 1848
rect -1357 1472 -1260 1496
rect -260 1848 -163 1872
rect -260 1496 -209 1848
rect -175 1496 -163 1848
rect -260 1472 -163 1496
rect 163 1848 260 1872
rect 163 1496 175 1848
rect 209 1496 260 1848
rect 163 1472 260 1496
rect 1260 1848 1357 1872
rect 1260 1496 1311 1848
rect 1345 1496 1357 1848
rect 1260 1472 1357 1496
rect 1683 1848 1780 1872
rect 1683 1496 1695 1848
rect 1729 1496 1780 1848
rect 1683 1472 1780 1496
rect 2780 1848 2877 1872
rect 2780 1496 2831 1848
rect 2865 1496 2877 1848
rect 2780 1472 2877 1496
rect -2877 1012 -2780 1036
rect -2877 660 -2865 1012
rect -2831 660 -2780 1012
rect -2877 636 -2780 660
rect -1780 1012 -1683 1036
rect -1780 660 -1729 1012
rect -1695 660 -1683 1012
rect -1780 636 -1683 660
rect -1357 1012 -1260 1036
rect -1357 660 -1345 1012
rect -1311 660 -1260 1012
rect -1357 636 -1260 660
rect -260 1012 -163 1036
rect -260 660 -209 1012
rect -175 660 -163 1012
rect -260 636 -163 660
rect 163 1012 260 1036
rect 163 660 175 1012
rect 209 660 260 1012
rect 163 636 260 660
rect 1260 1012 1357 1036
rect 1260 660 1311 1012
rect 1345 660 1357 1012
rect 1260 636 1357 660
rect 1683 1012 1780 1036
rect 1683 660 1695 1012
rect 1729 660 1780 1012
rect 1683 636 1780 660
rect 2780 1012 2877 1036
rect 2780 660 2831 1012
rect 2865 660 2877 1012
rect 2780 636 2877 660
rect -2877 176 -2780 200
rect -2877 -176 -2865 176
rect -2831 -176 -2780 176
rect -2877 -200 -2780 -176
rect -1780 176 -1683 200
rect -1780 -176 -1729 176
rect -1695 -176 -1683 176
rect -1780 -200 -1683 -176
rect -1357 176 -1260 200
rect -1357 -176 -1345 176
rect -1311 -176 -1260 176
rect -1357 -200 -1260 -176
rect -260 176 -163 200
rect -260 -176 -209 176
rect -175 -176 -163 176
rect -260 -200 -163 -176
rect 163 176 260 200
rect 163 -176 175 176
rect 209 -176 260 176
rect 163 -200 260 -176
rect 1260 176 1357 200
rect 1260 -176 1311 176
rect 1345 -176 1357 176
rect 1260 -200 1357 -176
rect 1683 176 1780 200
rect 1683 -176 1695 176
rect 1729 -176 1780 176
rect 1683 -200 1780 -176
rect 2780 176 2877 200
rect 2780 -176 2831 176
rect 2865 -176 2877 176
rect 2780 -200 2877 -176
rect -2877 -660 -2780 -636
rect -2877 -1012 -2865 -660
rect -2831 -1012 -2780 -660
rect -2877 -1036 -2780 -1012
rect -1780 -660 -1683 -636
rect -1780 -1012 -1729 -660
rect -1695 -1012 -1683 -660
rect -1780 -1036 -1683 -1012
rect -1357 -660 -1260 -636
rect -1357 -1012 -1345 -660
rect -1311 -1012 -1260 -660
rect -1357 -1036 -1260 -1012
rect -260 -660 -163 -636
rect -260 -1012 -209 -660
rect -175 -1012 -163 -660
rect -260 -1036 -163 -1012
rect 163 -660 260 -636
rect 163 -1012 175 -660
rect 209 -1012 260 -660
rect 163 -1036 260 -1012
rect 1260 -660 1357 -636
rect 1260 -1012 1311 -660
rect 1345 -1012 1357 -660
rect 1260 -1036 1357 -1012
rect 1683 -660 1780 -636
rect 1683 -1012 1695 -660
rect 1729 -1012 1780 -660
rect 1683 -1036 1780 -1012
rect 2780 -660 2877 -636
rect 2780 -1012 2831 -660
rect 2865 -1012 2877 -660
rect 2780 -1036 2877 -1012
rect -2877 -1496 -2780 -1472
rect -2877 -1848 -2865 -1496
rect -2831 -1848 -2780 -1496
rect -2877 -1872 -2780 -1848
rect -1780 -1496 -1683 -1472
rect -1780 -1848 -1729 -1496
rect -1695 -1848 -1683 -1496
rect -1780 -1872 -1683 -1848
rect -1357 -1496 -1260 -1472
rect -1357 -1848 -1345 -1496
rect -1311 -1848 -1260 -1496
rect -1357 -1872 -1260 -1848
rect -260 -1496 -163 -1472
rect -260 -1848 -209 -1496
rect -175 -1848 -163 -1496
rect -260 -1872 -163 -1848
rect 163 -1496 260 -1472
rect 163 -1848 175 -1496
rect 209 -1848 260 -1496
rect 163 -1872 260 -1848
rect 1260 -1496 1357 -1472
rect 1260 -1848 1311 -1496
rect 1345 -1848 1357 -1496
rect 1260 -1872 1357 -1848
rect 1683 -1496 1780 -1472
rect 1683 -1848 1695 -1496
rect 1729 -1848 1780 -1496
rect 1683 -1872 1780 -1848
rect 2780 -1496 2877 -1472
rect 2780 -1848 2831 -1496
rect 2865 -1848 2877 -1496
rect 2780 -1872 2877 -1848
<< psubdiffcont >>
rect -2891 2003 2891 2037
rect -2987 -1941 -2953 1941
rect 2953 -1941 2987 1941
rect -2891 -2037 2891 -2003
<< nsubdiffcont >>
rect -2865 1496 -2831 1848
rect -1729 1496 -1695 1848
rect -1345 1496 -1311 1848
rect -209 1496 -175 1848
rect 175 1496 209 1848
rect 1311 1496 1345 1848
rect 1695 1496 1729 1848
rect 2831 1496 2865 1848
rect -2865 660 -2831 1012
rect -1729 660 -1695 1012
rect -1345 660 -1311 1012
rect -209 660 -175 1012
rect 175 660 209 1012
rect 1311 660 1345 1012
rect 1695 660 1729 1012
rect 2831 660 2865 1012
rect -2865 -176 -2831 176
rect -1729 -176 -1695 176
rect -1345 -176 -1311 176
rect -209 -176 -175 176
rect 175 -176 209 176
rect 1311 -176 1345 176
rect 1695 -176 1729 176
rect 2831 -176 2865 176
rect -2865 -1012 -2831 -660
rect -1729 -1012 -1695 -660
rect -1345 -1012 -1311 -660
rect -209 -1012 -175 -660
rect 175 -1012 209 -660
rect 1311 -1012 1345 -660
rect 1695 -1012 1729 -660
rect 2831 -1012 2865 -660
rect -2865 -1848 -2831 -1496
rect -1729 -1848 -1695 -1496
rect -1345 -1848 -1311 -1496
rect -209 -1848 -175 -1496
rect 175 -1848 209 -1496
rect 1311 -1848 1345 -1496
rect 1695 -1848 1729 -1496
rect 2831 -1848 2865 -1496
<< poly >>
rect -2780 1944 -1780 1960
rect -2780 1910 -2764 1944
rect -1796 1910 -1780 1944
rect -2780 1872 -1780 1910
rect -1260 1944 -260 1960
rect -1260 1910 -1244 1944
rect -276 1910 -260 1944
rect -1260 1872 -260 1910
rect 260 1944 1260 1960
rect 260 1910 276 1944
rect 1244 1910 1260 1944
rect 260 1872 1260 1910
rect 1780 1944 2780 1960
rect 1780 1910 1796 1944
rect 2764 1910 2780 1944
rect 1780 1872 2780 1910
rect -2780 1434 -1780 1472
rect -2780 1400 -2764 1434
rect -1796 1400 -1780 1434
rect -2780 1384 -1780 1400
rect -1260 1434 -260 1472
rect -1260 1400 -1244 1434
rect -276 1400 -260 1434
rect -1260 1384 -260 1400
rect 260 1434 1260 1472
rect 260 1400 276 1434
rect 1244 1400 1260 1434
rect 260 1384 1260 1400
rect 1780 1434 2780 1472
rect 1780 1400 1796 1434
rect 2764 1400 2780 1434
rect 1780 1384 2780 1400
rect -2780 1108 -1780 1124
rect -2780 1074 -2764 1108
rect -1796 1074 -1780 1108
rect -2780 1036 -1780 1074
rect -1260 1108 -260 1124
rect -1260 1074 -1244 1108
rect -276 1074 -260 1108
rect -1260 1036 -260 1074
rect 260 1108 1260 1124
rect 260 1074 276 1108
rect 1244 1074 1260 1108
rect 260 1036 1260 1074
rect 1780 1108 2780 1124
rect 1780 1074 1796 1108
rect 2764 1074 2780 1108
rect 1780 1036 2780 1074
rect -2780 598 -1780 636
rect -2780 564 -2764 598
rect -1796 564 -1780 598
rect -2780 548 -1780 564
rect -1260 598 -260 636
rect -1260 564 -1244 598
rect -276 564 -260 598
rect -1260 548 -260 564
rect 260 598 1260 636
rect 260 564 276 598
rect 1244 564 1260 598
rect 260 548 1260 564
rect 1780 598 2780 636
rect 1780 564 1796 598
rect 2764 564 2780 598
rect 1780 548 2780 564
rect -2780 272 -1780 288
rect -2780 238 -2764 272
rect -1796 238 -1780 272
rect -2780 200 -1780 238
rect -1260 272 -260 288
rect -1260 238 -1244 272
rect -276 238 -260 272
rect -1260 200 -260 238
rect 260 272 1260 288
rect 260 238 276 272
rect 1244 238 1260 272
rect 260 200 1260 238
rect 1780 272 2780 288
rect 1780 238 1796 272
rect 2764 238 2780 272
rect 1780 200 2780 238
rect -2780 -238 -1780 -200
rect -2780 -272 -2764 -238
rect -1796 -272 -1780 -238
rect -2780 -288 -1780 -272
rect -1260 -238 -260 -200
rect -1260 -272 -1244 -238
rect -276 -272 -260 -238
rect -1260 -288 -260 -272
rect 260 -238 1260 -200
rect 260 -272 276 -238
rect 1244 -272 1260 -238
rect 260 -288 1260 -272
rect 1780 -238 2780 -200
rect 1780 -272 1796 -238
rect 2764 -272 2780 -238
rect 1780 -288 2780 -272
rect -2780 -564 -1780 -548
rect -2780 -598 -2764 -564
rect -1796 -598 -1780 -564
rect -2780 -636 -1780 -598
rect -1260 -564 -260 -548
rect -1260 -598 -1244 -564
rect -276 -598 -260 -564
rect -1260 -636 -260 -598
rect 260 -564 1260 -548
rect 260 -598 276 -564
rect 1244 -598 1260 -564
rect 260 -636 1260 -598
rect 1780 -564 2780 -548
rect 1780 -598 1796 -564
rect 2764 -598 2780 -564
rect 1780 -636 2780 -598
rect -2780 -1074 -1780 -1036
rect -2780 -1108 -2764 -1074
rect -1796 -1108 -1780 -1074
rect -2780 -1124 -1780 -1108
rect -1260 -1074 -260 -1036
rect -1260 -1108 -1244 -1074
rect -276 -1108 -260 -1074
rect -1260 -1124 -260 -1108
rect 260 -1074 1260 -1036
rect 260 -1108 276 -1074
rect 1244 -1108 1260 -1074
rect 260 -1124 1260 -1108
rect 1780 -1074 2780 -1036
rect 1780 -1108 1796 -1074
rect 2764 -1108 2780 -1074
rect 1780 -1124 2780 -1108
rect -2780 -1400 -1780 -1384
rect -2780 -1434 -2764 -1400
rect -1796 -1434 -1780 -1400
rect -2780 -1472 -1780 -1434
rect -1260 -1400 -260 -1384
rect -1260 -1434 -1244 -1400
rect -276 -1434 -260 -1400
rect -1260 -1472 -260 -1434
rect 260 -1400 1260 -1384
rect 260 -1434 276 -1400
rect 1244 -1434 1260 -1400
rect 260 -1472 1260 -1434
rect 1780 -1400 2780 -1384
rect 1780 -1434 1796 -1400
rect 2764 -1434 2780 -1400
rect 1780 -1472 2780 -1434
rect -2780 -1910 -1780 -1872
rect -2780 -1944 -2764 -1910
rect -1796 -1944 -1780 -1910
rect -2780 -1960 -1780 -1944
rect -1260 -1910 -260 -1872
rect -1260 -1944 -1244 -1910
rect -276 -1944 -260 -1910
rect -1260 -1960 -260 -1944
rect 260 -1910 1260 -1872
rect 260 -1944 276 -1910
rect 1244 -1944 1260 -1910
rect 260 -1960 1260 -1944
rect 1780 -1910 2780 -1872
rect 1780 -1944 1796 -1910
rect 2764 -1944 2780 -1910
rect 1780 -1960 2780 -1944
<< polycont >>
rect -2764 1910 -1796 1944
rect -1244 1910 -276 1944
rect 276 1910 1244 1944
rect 1796 1910 2764 1944
rect -2764 1400 -1796 1434
rect -1244 1400 -276 1434
rect 276 1400 1244 1434
rect 1796 1400 2764 1434
rect -2764 1074 -1796 1108
rect -1244 1074 -276 1108
rect 276 1074 1244 1108
rect 1796 1074 2764 1108
rect -2764 564 -1796 598
rect -1244 564 -276 598
rect 276 564 1244 598
rect 1796 564 2764 598
rect -2764 238 -1796 272
rect -1244 238 -276 272
rect 276 238 1244 272
rect 1796 238 2764 272
rect -2764 -272 -1796 -238
rect -1244 -272 -276 -238
rect 276 -272 1244 -238
rect 1796 -272 2764 -238
rect -2764 -598 -1796 -564
rect -1244 -598 -276 -564
rect 276 -598 1244 -564
rect 1796 -598 2764 -564
rect -2764 -1108 -1796 -1074
rect -1244 -1108 -276 -1074
rect 276 -1108 1244 -1074
rect 1796 -1108 2764 -1074
rect -2764 -1434 -1796 -1400
rect -1244 -1434 -276 -1400
rect 276 -1434 1244 -1400
rect 1796 -1434 2764 -1400
rect -2764 -1944 -1796 -1910
rect -1244 -1944 -276 -1910
rect 276 -1944 1244 -1910
rect 1796 -1944 2764 -1910
<< locali >>
rect -2987 2003 -2891 2037
rect 2891 2003 2987 2037
rect -2987 1941 -2953 2003
rect -2780 1910 -2764 1944
rect -1796 1910 -1780 1944
rect -1260 1910 -1244 1944
rect -276 1910 -260 1944
rect 260 1910 276 1944
rect 1244 1910 1260 1944
rect 1780 1910 1796 1944
rect 2764 1910 2780 1944
rect 2953 1941 2987 2003
rect -2865 1848 -2831 1864
rect -2865 1480 -2831 1496
rect -1729 1848 -1695 1864
rect -1729 1480 -1695 1496
rect -1345 1848 -1311 1864
rect -1345 1480 -1311 1496
rect -209 1848 -175 1864
rect -209 1480 -175 1496
rect 175 1848 209 1864
rect 175 1480 209 1496
rect 1311 1848 1345 1864
rect 1311 1480 1345 1496
rect 1695 1848 1729 1864
rect 1695 1480 1729 1496
rect 2831 1848 2865 1864
rect 2831 1480 2865 1496
rect -2780 1400 -2764 1434
rect -1796 1400 -1780 1434
rect -1260 1400 -1244 1434
rect -276 1400 -260 1434
rect 260 1400 276 1434
rect 1244 1400 1260 1434
rect 1780 1400 1796 1434
rect 2764 1400 2780 1434
rect -2780 1074 -2764 1108
rect -1796 1074 -1780 1108
rect -1260 1074 -1244 1108
rect -276 1074 -260 1108
rect 260 1074 276 1108
rect 1244 1074 1260 1108
rect 1780 1074 1796 1108
rect 2764 1074 2780 1108
rect -2865 1012 -2831 1028
rect -2865 644 -2831 660
rect -1729 1012 -1695 1028
rect -1729 644 -1695 660
rect -1345 1012 -1311 1028
rect -1345 644 -1311 660
rect -209 1012 -175 1028
rect -209 644 -175 660
rect 175 1012 209 1028
rect 175 644 209 660
rect 1311 1012 1345 1028
rect 1311 644 1345 660
rect 1695 1012 1729 1028
rect 1695 644 1729 660
rect 2831 1012 2865 1028
rect 2831 644 2865 660
rect -2780 564 -2764 598
rect -1796 564 -1780 598
rect -1260 564 -1244 598
rect -276 564 -260 598
rect 260 564 276 598
rect 1244 564 1260 598
rect 1780 564 1796 598
rect 2764 564 2780 598
rect -2780 238 -2764 272
rect -1796 238 -1780 272
rect -1260 238 -1244 272
rect -276 238 -260 272
rect 260 238 276 272
rect 1244 238 1260 272
rect 1780 238 1796 272
rect 2764 238 2780 272
rect -2865 176 -2831 192
rect -2865 -192 -2831 -176
rect -1729 176 -1695 192
rect -1729 -192 -1695 -176
rect -1345 176 -1311 192
rect -1345 -192 -1311 -176
rect -209 176 -175 192
rect -209 -192 -175 -176
rect 175 176 209 192
rect 175 -192 209 -176
rect 1311 176 1345 192
rect 1311 -192 1345 -176
rect 1695 176 1729 192
rect 1695 -192 1729 -176
rect 2831 176 2865 192
rect 2831 -192 2865 -176
rect -2780 -272 -2764 -238
rect -1796 -272 -1780 -238
rect -1260 -272 -1244 -238
rect -276 -272 -260 -238
rect 260 -272 276 -238
rect 1244 -272 1260 -238
rect 1780 -272 1796 -238
rect 2764 -272 2780 -238
rect -2780 -598 -2764 -564
rect -1796 -598 -1780 -564
rect -1260 -598 -1244 -564
rect -276 -598 -260 -564
rect 260 -598 276 -564
rect 1244 -598 1260 -564
rect 1780 -598 1796 -564
rect 2764 -598 2780 -564
rect -2865 -660 -2831 -644
rect -2865 -1028 -2831 -1012
rect -1729 -660 -1695 -644
rect -1729 -1028 -1695 -1012
rect -1345 -660 -1311 -644
rect -1345 -1028 -1311 -1012
rect -209 -660 -175 -644
rect -209 -1028 -175 -1012
rect 175 -660 209 -644
rect 175 -1028 209 -1012
rect 1311 -660 1345 -644
rect 1311 -1028 1345 -1012
rect 1695 -660 1729 -644
rect 1695 -1028 1729 -1012
rect 2831 -660 2865 -644
rect 2831 -1028 2865 -1012
rect -2780 -1108 -2764 -1074
rect -1796 -1108 -1780 -1074
rect -1260 -1108 -1244 -1074
rect -276 -1108 -260 -1074
rect 260 -1108 276 -1074
rect 1244 -1108 1260 -1074
rect 1780 -1108 1796 -1074
rect 2764 -1108 2780 -1074
rect -2780 -1434 -2764 -1400
rect -1796 -1434 -1780 -1400
rect -1260 -1434 -1244 -1400
rect -276 -1434 -260 -1400
rect 260 -1434 276 -1400
rect 1244 -1434 1260 -1400
rect 1780 -1434 1796 -1400
rect 2764 -1434 2780 -1400
rect -2865 -1496 -2831 -1480
rect -2865 -1864 -2831 -1848
rect -1729 -1496 -1695 -1480
rect -1729 -1864 -1695 -1848
rect -1345 -1496 -1311 -1480
rect -1345 -1864 -1311 -1848
rect -209 -1496 -175 -1480
rect -209 -1864 -175 -1848
rect 175 -1496 209 -1480
rect 175 -1864 209 -1848
rect 1311 -1496 1345 -1480
rect 1311 -1864 1345 -1848
rect 1695 -1496 1729 -1480
rect 1695 -1864 1729 -1848
rect 2831 -1496 2865 -1480
rect 2831 -1864 2865 -1848
rect -2987 -2003 -2953 -1941
rect -2780 -1944 -2764 -1910
rect -1796 -1944 -1780 -1910
rect -1260 -1944 -1244 -1910
rect -276 -1944 -260 -1910
rect 260 -1944 276 -1910
rect 1244 -1944 1260 -1910
rect 1780 -1944 1796 -1910
rect 2764 -1944 2780 -1910
rect 2953 -2003 2987 -1941
rect -2987 -2037 -2891 -2003
rect 2891 -2037 2987 -2003
<< viali >>
rect -2764 1910 -1796 1944
rect -1244 1910 -276 1944
rect 276 1910 1244 1944
rect 1796 1910 2764 1944
rect -2865 1496 -2831 1848
rect -1729 1496 -1695 1848
rect -1345 1496 -1311 1848
rect -209 1496 -175 1848
rect 175 1496 209 1848
rect 1311 1496 1345 1848
rect 1695 1496 1729 1848
rect 2831 1496 2865 1848
rect -2764 1400 -1796 1434
rect -1244 1400 -276 1434
rect 276 1400 1244 1434
rect 1796 1400 2764 1434
rect -2764 1074 -1796 1108
rect -1244 1074 -276 1108
rect 276 1074 1244 1108
rect 1796 1074 2764 1108
rect -2865 660 -2831 1012
rect -1729 660 -1695 1012
rect -1345 660 -1311 1012
rect -209 660 -175 1012
rect 175 660 209 1012
rect 1311 660 1345 1012
rect 1695 660 1729 1012
rect 2831 660 2865 1012
rect -2764 564 -1796 598
rect -1244 564 -276 598
rect 276 564 1244 598
rect 1796 564 2764 598
rect -2764 238 -1796 272
rect -1244 238 -276 272
rect 276 238 1244 272
rect 1796 238 2764 272
rect -2865 -176 -2831 176
rect -1729 -176 -1695 176
rect -1345 -176 -1311 176
rect -209 -176 -175 176
rect 175 -176 209 176
rect 1311 -176 1345 176
rect 1695 -176 1729 176
rect 2831 -176 2865 176
rect -2764 -272 -1796 -238
rect -1244 -272 -276 -238
rect 276 -272 1244 -238
rect 1796 -272 2764 -238
rect -2764 -598 -1796 -564
rect -1244 -598 -276 -564
rect 276 -598 1244 -564
rect 1796 -598 2764 -564
rect -2865 -1012 -2831 -660
rect -1729 -1012 -1695 -660
rect -1345 -1012 -1311 -660
rect -209 -1012 -175 -660
rect 175 -1012 209 -660
rect 1311 -1012 1345 -660
rect 1695 -1012 1729 -660
rect 2831 -1012 2865 -660
rect -2764 -1108 -1796 -1074
rect -1244 -1108 -276 -1074
rect 276 -1108 1244 -1074
rect 1796 -1108 2764 -1074
rect -2764 -1434 -1796 -1400
rect -1244 -1434 -276 -1400
rect 276 -1434 1244 -1400
rect 1796 -1434 2764 -1400
rect -2865 -1848 -2831 -1496
rect -1729 -1848 -1695 -1496
rect -1345 -1848 -1311 -1496
rect -209 -1848 -175 -1496
rect 175 -1848 209 -1496
rect 1311 -1848 1345 -1496
rect 1695 -1848 1729 -1496
rect 2831 -1848 2865 -1496
rect -2764 -1944 -1796 -1910
rect -1244 -1944 -276 -1910
rect 276 -1944 1244 -1910
rect 1796 -1944 2764 -1910
<< metal1 >>
rect -2776 1944 -1784 1950
rect -2776 1910 -2764 1944
rect -1796 1910 -1784 1944
rect -2776 1904 -1784 1910
rect -1256 1944 -264 1950
rect -1256 1910 -1244 1944
rect -276 1910 -264 1944
rect -1256 1904 -264 1910
rect 264 1944 1256 1950
rect 264 1910 276 1944
rect 1244 1910 1256 1944
rect 264 1904 1256 1910
rect 1784 1944 2776 1950
rect 1784 1910 1796 1944
rect 2764 1910 2776 1944
rect 1784 1904 2776 1910
rect -2871 1848 -2825 1860
rect -1735 1848 -1689 1860
rect -2871 1496 -2865 1848
rect -2831 1496 -1729 1848
rect -1695 1496 -1689 1848
rect -2871 1484 -2825 1496
rect -1735 1484 -1689 1496
rect -1351 1848 -1305 1860
rect -215 1848 -169 1860
rect -1351 1496 -1345 1848
rect -1311 1496 -209 1848
rect -175 1496 -169 1848
rect -1351 1484 -1305 1496
rect -215 1484 -169 1496
rect 169 1848 215 1860
rect 1305 1848 1351 1860
rect 169 1496 175 1848
rect 209 1496 1311 1848
rect 1345 1496 1351 1848
rect 169 1484 215 1496
rect 1305 1484 1351 1496
rect 1689 1848 1735 1860
rect 2825 1848 2871 1860
rect 1689 1496 1695 1848
rect 1729 1496 2831 1848
rect 2865 1496 2871 1848
rect 1689 1484 1735 1496
rect 2825 1484 2871 1496
rect -2776 1434 -1784 1440
rect -2776 1400 -2764 1434
rect -1796 1400 -1784 1434
rect -2776 1394 -1784 1400
rect -1256 1434 -264 1440
rect -1256 1400 -1244 1434
rect -276 1400 -264 1434
rect -1256 1394 -264 1400
rect 264 1434 1256 1440
rect 264 1400 276 1434
rect 1244 1400 1256 1434
rect 264 1394 1256 1400
rect 1784 1434 2776 1440
rect 1784 1400 1796 1434
rect 2764 1400 2776 1434
rect 1784 1394 2776 1400
rect -2776 1108 -1784 1114
rect -2776 1074 -2764 1108
rect -1796 1074 -1784 1108
rect -2776 1068 -1784 1074
rect -1256 1108 -264 1114
rect -1256 1074 -1244 1108
rect -276 1074 -264 1108
rect -1256 1068 -264 1074
rect 264 1108 1256 1114
rect 264 1074 276 1108
rect 1244 1074 1256 1108
rect 264 1068 1256 1074
rect 1784 1108 2776 1114
rect 1784 1074 1796 1108
rect 2764 1074 2776 1108
rect 1784 1068 2776 1074
rect -2871 1012 -2825 1024
rect -1735 1012 -1689 1024
rect -2871 660 -2865 1012
rect -2831 660 -1729 1012
rect -1695 660 -1689 1012
rect -2871 648 -2825 660
rect -1735 648 -1689 660
rect -1351 1012 -1305 1024
rect -215 1012 -169 1024
rect -1351 660 -1345 1012
rect -1311 660 -209 1012
rect -175 660 -169 1012
rect -1351 648 -1305 660
rect -215 648 -169 660
rect 169 1012 215 1024
rect 1305 1012 1351 1024
rect 169 660 175 1012
rect 209 660 1311 1012
rect 1345 660 1351 1012
rect 169 648 215 660
rect 1305 648 1351 660
rect 1689 1012 1735 1024
rect 2825 1012 2871 1024
rect 1689 660 1695 1012
rect 1729 660 2831 1012
rect 2865 660 2871 1012
rect 1689 648 1735 660
rect 2825 648 2871 660
rect -2776 598 -1784 604
rect -2776 564 -2764 598
rect -1796 564 -1784 598
rect -2776 558 -1784 564
rect -1256 598 -264 604
rect -1256 564 -1244 598
rect -276 564 -264 598
rect -1256 558 -264 564
rect 264 598 1256 604
rect 264 564 276 598
rect 1244 564 1256 598
rect 264 558 1256 564
rect 1784 598 2776 604
rect 1784 564 1796 598
rect 2764 564 2776 598
rect 1784 558 2776 564
rect -2776 272 -1784 278
rect -2776 238 -2764 272
rect -1796 238 -1784 272
rect -2776 232 -1784 238
rect -1256 272 -264 278
rect -1256 238 -1244 272
rect -276 238 -264 272
rect -1256 232 -264 238
rect 264 272 1256 278
rect 264 238 276 272
rect 1244 238 1256 272
rect 264 232 1256 238
rect 1784 272 2776 278
rect 1784 238 1796 272
rect 2764 238 2776 272
rect 1784 232 2776 238
rect -2871 176 -2825 188
rect -1735 176 -1689 188
rect -2871 -176 -2865 176
rect -2831 -176 -1729 176
rect -1695 -176 -1689 176
rect -2871 -188 -2825 -176
rect -1735 -188 -1689 -176
rect -1351 176 -1305 188
rect -215 176 -169 188
rect -1351 -176 -1345 176
rect -1311 -176 -209 176
rect -175 -176 -169 176
rect -1351 -188 -1305 -176
rect -215 -188 -169 -176
rect 169 176 215 188
rect 1305 176 1351 188
rect 169 -176 175 176
rect 209 -176 1311 176
rect 1345 -176 1351 176
rect 169 -188 215 -176
rect 1305 -188 1351 -176
rect 1689 176 1735 188
rect 2825 176 2871 188
rect 1689 -176 1695 176
rect 1729 -176 2831 176
rect 2865 -176 2871 176
rect 1689 -188 1735 -176
rect 2825 -188 2871 -176
rect -2776 -238 -1784 -232
rect -2776 -272 -2764 -238
rect -1796 -272 -1784 -238
rect -2776 -278 -1784 -272
rect -1256 -238 -264 -232
rect -1256 -272 -1244 -238
rect -276 -272 -264 -238
rect -1256 -278 -264 -272
rect 264 -238 1256 -232
rect 264 -272 276 -238
rect 1244 -272 1256 -238
rect 264 -278 1256 -272
rect 1784 -238 2776 -232
rect 1784 -272 1796 -238
rect 2764 -272 2776 -238
rect 1784 -278 2776 -272
rect -2776 -564 -1784 -558
rect -2776 -598 -2764 -564
rect -1796 -598 -1784 -564
rect -2776 -604 -1784 -598
rect -1256 -564 -264 -558
rect -1256 -598 -1244 -564
rect -276 -598 -264 -564
rect -1256 -604 -264 -598
rect 264 -564 1256 -558
rect 264 -598 276 -564
rect 1244 -598 1256 -564
rect 264 -604 1256 -598
rect 1784 -564 2776 -558
rect 1784 -598 1796 -564
rect 2764 -598 2776 -564
rect 1784 -604 2776 -598
rect -2871 -660 -2825 -648
rect -1735 -660 -1689 -648
rect -2871 -1012 -2865 -660
rect -2831 -1012 -1729 -660
rect -1695 -1012 -1689 -660
rect -2871 -1024 -2825 -1012
rect -1735 -1024 -1689 -1012
rect -1351 -660 -1305 -648
rect -215 -660 -169 -648
rect -1351 -1012 -1345 -660
rect -1311 -1012 -209 -660
rect -175 -1012 -169 -660
rect -1351 -1024 -1305 -1012
rect -215 -1024 -169 -1012
rect 169 -660 215 -648
rect 1305 -660 1351 -648
rect 169 -1012 175 -660
rect 209 -1012 1311 -660
rect 1345 -1012 1351 -660
rect 169 -1024 215 -1012
rect 1305 -1024 1351 -1012
rect 1689 -660 1735 -648
rect 2825 -660 2871 -648
rect 1689 -1012 1695 -660
rect 1729 -1012 2831 -660
rect 2865 -1012 2871 -660
rect 1689 -1024 1735 -1012
rect 2825 -1024 2871 -1012
rect -2776 -1074 -1784 -1068
rect -2776 -1108 -2764 -1074
rect -1796 -1108 -1784 -1074
rect -2776 -1114 -1784 -1108
rect -1256 -1074 -264 -1068
rect -1256 -1108 -1244 -1074
rect -276 -1108 -264 -1074
rect -1256 -1114 -264 -1108
rect 264 -1074 1256 -1068
rect 264 -1108 276 -1074
rect 1244 -1108 1256 -1074
rect 264 -1114 1256 -1108
rect 1784 -1074 2776 -1068
rect 1784 -1108 1796 -1074
rect 2764 -1108 2776 -1074
rect 1784 -1114 2776 -1108
rect -2776 -1400 -1784 -1394
rect -2776 -1434 -2764 -1400
rect -1796 -1434 -1784 -1400
rect -2776 -1440 -1784 -1434
rect -1256 -1400 -264 -1394
rect -1256 -1434 -1244 -1400
rect -276 -1434 -264 -1400
rect -1256 -1440 -264 -1434
rect 264 -1400 1256 -1394
rect 264 -1434 276 -1400
rect 1244 -1434 1256 -1400
rect 264 -1440 1256 -1434
rect 1784 -1400 2776 -1394
rect 1784 -1434 1796 -1400
rect 2764 -1434 2776 -1400
rect 1784 -1440 2776 -1434
rect -2871 -1496 -2825 -1484
rect -1735 -1496 -1689 -1484
rect -2871 -1848 -2865 -1496
rect -2831 -1848 -1729 -1496
rect -1695 -1848 -1689 -1496
rect -2871 -1860 -2825 -1848
rect -1735 -1860 -1689 -1848
rect -1351 -1496 -1305 -1484
rect -215 -1496 -169 -1484
rect -1351 -1848 -1345 -1496
rect -1311 -1848 -209 -1496
rect -175 -1848 -169 -1496
rect -1351 -1860 -1305 -1848
rect -215 -1860 -169 -1848
rect 169 -1496 215 -1484
rect 1305 -1496 1351 -1484
rect 169 -1848 175 -1496
rect 209 -1848 1311 -1496
rect 1345 -1848 1351 -1496
rect 169 -1860 215 -1848
rect 1305 -1860 1351 -1848
rect 1689 -1496 1735 -1484
rect 2825 -1496 2871 -1484
rect 1689 -1848 1695 -1496
rect 1729 -1848 2831 -1496
rect 2865 -1848 2871 -1496
rect 1689 -1860 1735 -1848
rect 2825 -1860 2871 -1848
rect -2776 -1910 -1784 -1904
rect -2776 -1944 -2764 -1910
rect -1796 -1944 -1784 -1910
rect -2776 -1950 -1784 -1944
rect -1256 -1910 -264 -1904
rect -1256 -1944 -1244 -1910
rect -276 -1944 -264 -1910
rect -1256 -1950 -264 -1944
rect 264 -1910 1256 -1904
rect 264 -1944 276 -1910
rect 1244 -1944 1256 -1910
rect 264 -1950 1256 -1944
rect 1784 -1910 2776 -1904
rect 1784 -1944 1796 -1910
rect 2764 -1944 2776 -1910
rect 1784 -1950 2776 -1944
<< properties >>
string FIXED_BBOX -2970 -2020 2970 2020
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 2 l 5 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 gshield 1
<< end >>
