magic
tech sky130A
magscale 1 2
timestamp 1683809155
<< error_p >>
rect -1421 1199 -1363 1205
rect -1229 1199 -1171 1205
rect -1037 1199 -979 1205
rect -845 1199 -787 1205
rect -653 1199 -595 1205
rect -461 1199 -403 1205
rect -269 1199 -211 1205
rect -77 1199 -19 1205
rect 115 1199 173 1205
rect 307 1199 365 1205
rect 499 1199 557 1205
rect 691 1199 749 1205
rect 883 1199 941 1205
rect 1075 1199 1133 1205
rect 1267 1199 1325 1205
rect -1421 1165 -1409 1199
rect -1229 1165 -1217 1199
rect -1037 1165 -1025 1199
rect -845 1165 -833 1199
rect -653 1165 -641 1199
rect -461 1165 -449 1199
rect -269 1165 -257 1199
rect -77 1165 -65 1199
rect 115 1165 127 1199
rect 307 1165 319 1199
rect 499 1165 511 1199
rect 691 1165 703 1199
rect 883 1165 895 1199
rect 1075 1165 1087 1199
rect 1267 1165 1279 1199
rect -1421 1159 -1363 1165
rect -1229 1159 -1171 1165
rect -1037 1159 -979 1165
rect -845 1159 -787 1165
rect -653 1159 -595 1165
rect -461 1159 -403 1165
rect -269 1159 -211 1165
rect -77 1159 -19 1165
rect 115 1159 173 1165
rect 307 1159 365 1165
rect 499 1159 557 1165
rect 691 1159 749 1165
rect 883 1159 941 1165
rect 1075 1159 1133 1165
rect 1267 1159 1325 1165
rect -1325 689 -1267 695
rect -1133 689 -1075 695
rect -941 689 -883 695
rect -749 689 -691 695
rect -557 689 -499 695
rect -365 689 -307 695
rect -173 689 -115 695
rect 19 689 77 695
rect 211 689 269 695
rect 403 689 461 695
rect 595 689 653 695
rect 787 689 845 695
rect 979 689 1037 695
rect 1171 689 1229 695
rect 1363 689 1421 695
rect -1325 655 -1313 689
rect -1133 655 -1121 689
rect -941 655 -929 689
rect -749 655 -737 689
rect -557 655 -545 689
rect -365 655 -353 689
rect -173 655 -161 689
rect 19 655 31 689
rect 211 655 223 689
rect 403 655 415 689
rect 595 655 607 689
rect 787 655 799 689
rect 979 655 991 689
rect 1171 655 1183 689
rect 1363 655 1375 689
rect -1325 649 -1267 655
rect -1133 649 -1075 655
rect -941 649 -883 655
rect -749 649 -691 655
rect -557 649 -499 655
rect -365 649 -307 655
rect -173 649 -115 655
rect 19 649 77 655
rect 211 649 269 655
rect 403 649 461 655
rect 595 649 653 655
rect 787 649 845 655
rect 979 649 1037 655
rect 1171 649 1229 655
rect 1363 649 1421 655
rect -1325 581 -1267 587
rect -1133 581 -1075 587
rect -941 581 -883 587
rect -749 581 -691 587
rect -557 581 -499 587
rect -365 581 -307 587
rect -173 581 -115 587
rect 19 581 77 587
rect 211 581 269 587
rect 403 581 461 587
rect 595 581 653 587
rect 787 581 845 587
rect 979 581 1037 587
rect 1171 581 1229 587
rect 1363 581 1421 587
rect -1325 547 -1313 581
rect -1133 547 -1121 581
rect -941 547 -929 581
rect -749 547 -737 581
rect -557 547 -545 581
rect -365 547 -353 581
rect -173 547 -161 581
rect 19 547 31 581
rect 211 547 223 581
rect 403 547 415 581
rect 595 547 607 581
rect 787 547 799 581
rect 979 547 991 581
rect 1171 547 1183 581
rect 1363 547 1375 581
rect -1325 541 -1267 547
rect -1133 541 -1075 547
rect -941 541 -883 547
rect -749 541 -691 547
rect -557 541 -499 547
rect -365 541 -307 547
rect -173 541 -115 547
rect 19 541 77 547
rect 211 541 269 547
rect 403 541 461 547
rect 595 541 653 547
rect 787 541 845 547
rect 979 541 1037 547
rect 1171 541 1229 547
rect 1363 541 1421 547
rect -1421 71 -1363 77
rect -1229 71 -1171 77
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect 1267 71 1325 77
rect -1421 37 -1409 71
rect -1229 37 -1217 71
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect 1267 37 1279 71
rect -1421 31 -1363 37
rect -1229 31 -1171 37
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect 1267 31 1325 37
rect -1421 -37 -1363 -31
rect -1229 -37 -1171 -31
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect 1267 -37 1325 -31
rect -1421 -71 -1409 -37
rect -1229 -71 -1217 -37
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect 1267 -71 1279 -37
rect -1421 -77 -1363 -71
rect -1229 -77 -1171 -71
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect 1267 -77 1325 -71
rect -1325 -547 -1267 -541
rect -1133 -547 -1075 -541
rect -941 -547 -883 -541
rect -749 -547 -691 -541
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect 595 -547 653 -541
rect 787 -547 845 -541
rect 979 -547 1037 -541
rect 1171 -547 1229 -541
rect 1363 -547 1421 -541
rect -1325 -581 -1313 -547
rect -1133 -581 -1121 -547
rect -941 -581 -929 -547
rect -749 -581 -737 -547
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect 595 -581 607 -547
rect 787 -581 799 -547
rect 979 -581 991 -547
rect 1171 -581 1183 -547
rect 1363 -581 1375 -547
rect -1325 -587 -1267 -581
rect -1133 -587 -1075 -581
rect -941 -587 -883 -581
rect -749 -587 -691 -581
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
rect 595 -587 653 -581
rect 787 -587 845 -581
rect 979 -587 1037 -581
rect 1171 -587 1229 -581
rect 1363 -587 1421 -581
rect -1325 -655 -1267 -649
rect -1133 -655 -1075 -649
rect -941 -655 -883 -649
rect -749 -655 -691 -649
rect -557 -655 -499 -649
rect -365 -655 -307 -649
rect -173 -655 -115 -649
rect 19 -655 77 -649
rect 211 -655 269 -649
rect 403 -655 461 -649
rect 595 -655 653 -649
rect 787 -655 845 -649
rect 979 -655 1037 -649
rect 1171 -655 1229 -649
rect 1363 -655 1421 -649
rect -1325 -689 -1313 -655
rect -1133 -689 -1121 -655
rect -941 -689 -929 -655
rect -749 -689 -737 -655
rect -557 -689 -545 -655
rect -365 -689 -353 -655
rect -173 -689 -161 -655
rect 19 -689 31 -655
rect 211 -689 223 -655
rect 403 -689 415 -655
rect 595 -689 607 -655
rect 787 -689 799 -655
rect 979 -689 991 -655
rect 1171 -689 1183 -655
rect 1363 -689 1375 -655
rect -1325 -695 -1267 -689
rect -1133 -695 -1075 -689
rect -941 -695 -883 -689
rect -749 -695 -691 -689
rect -557 -695 -499 -689
rect -365 -695 -307 -689
rect -173 -695 -115 -689
rect 19 -695 77 -689
rect 211 -695 269 -689
rect 403 -695 461 -689
rect 595 -695 653 -689
rect 787 -695 845 -689
rect 979 -695 1037 -689
rect 1171 -695 1229 -689
rect 1363 -695 1421 -689
rect -1421 -1165 -1363 -1159
rect -1229 -1165 -1171 -1159
rect -1037 -1165 -979 -1159
rect -845 -1165 -787 -1159
rect -653 -1165 -595 -1159
rect -461 -1165 -403 -1159
rect -269 -1165 -211 -1159
rect -77 -1165 -19 -1159
rect 115 -1165 173 -1159
rect 307 -1165 365 -1159
rect 499 -1165 557 -1159
rect 691 -1165 749 -1159
rect 883 -1165 941 -1159
rect 1075 -1165 1133 -1159
rect 1267 -1165 1325 -1159
rect -1421 -1199 -1409 -1165
rect -1229 -1199 -1217 -1165
rect -1037 -1199 -1025 -1165
rect -845 -1199 -833 -1165
rect -653 -1199 -641 -1165
rect -461 -1199 -449 -1165
rect -269 -1199 -257 -1165
rect -77 -1199 -65 -1165
rect 115 -1199 127 -1165
rect 307 -1199 319 -1165
rect 499 -1199 511 -1165
rect 691 -1199 703 -1165
rect 883 -1199 895 -1165
rect 1075 -1199 1087 -1165
rect 1267 -1199 1279 -1165
rect -1421 -1205 -1363 -1199
rect -1229 -1205 -1171 -1199
rect -1037 -1205 -979 -1199
rect -845 -1205 -787 -1199
rect -653 -1205 -595 -1199
rect -461 -1205 -403 -1199
rect -269 -1205 -211 -1199
rect -77 -1205 -19 -1199
rect 115 -1205 173 -1199
rect 307 -1205 365 -1199
rect 499 -1205 557 -1199
rect 691 -1205 749 -1199
rect 883 -1205 941 -1199
rect 1075 -1205 1133 -1199
rect 1267 -1205 1325 -1199
<< pwell >>
rect -1607 -1337 1607 1337
<< nmoslvt >>
rect -1407 727 -1377 1127
rect -1311 727 -1281 1127
rect -1215 727 -1185 1127
rect -1119 727 -1089 1127
rect -1023 727 -993 1127
rect -927 727 -897 1127
rect -831 727 -801 1127
rect -735 727 -705 1127
rect -639 727 -609 1127
rect -543 727 -513 1127
rect -447 727 -417 1127
rect -351 727 -321 1127
rect -255 727 -225 1127
rect -159 727 -129 1127
rect -63 727 -33 1127
rect 33 727 63 1127
rect 129 727 159 1127
rect 225 727 255 1127
rect 321 727 351 1127
rect 417 727 447 1127
rect 513 727 543 1127
rect 609 727 639 1127
rect 705 727 735 1127
rect 801 727 831 1127
rect 897 727 927 1127
rect 993 727 1023 1127
rect 1089 727 1119 1127
rect 1185 727 1215 1127
rect 1281 727 1311 1127
rect 1377 727 1407 1127
rect -1407 109 -1377 509
rect -1311 109 -1281 509
rect -1215 109 -1185 509
rect -1119 109 -1089 509
rect -1023 109 -993 509
rect -927 109 -897 509
rect -831 109 -801 509
rect -735 109 -705 509
rect -639 109 -609 509
rect -543 109 -513 509
rect -447 109 -417 509
rect -351 109 -321 509
rect -255 109 -225 509
rect -159 109 -129 509
rect -63 109 -33 509
rect 33 109 63 509
rect 129 109 159 509
rect 225 109 255 509
rect 321 109 351 509
rect 417 109 447 509
rect 513 109 543 509
rect 609 109 639 509
rect 705 109 735 509
rect 801 109 831 509
rect 897 109 927 509
rect 993 109 1023 509
rect 1089 109 1119 509
rect 1185 109 1215 509
rect 1281 109 1311 509
rect 1377 109 1407 509
rect -1407 -509 -1377 -109
rect -1311 -509 -1281 -109
rect -1215 -509 -1185 -109
rect -1119 -509 -1089 -109
rect -1023 -509 -993 -109
rect -927 -509 -897 -109
rect -831 -509 -801 -109
rect -735 -509 -705 -109
rect -639 -509 -609 -109
rect -543 -509 -513 -109
rect -447 -509 -417 -109
rect -351 -509 -321 -109
rect -255 -509 -225 -109
rect -159 -509 -129 -109
rect -63 -509 -33 -109
rect 33 -509 63 -109
rect 129 -509 159 -109
rect 225 -509 255 -109
rect 321 -509 351 -109
rect 417 -509 447 -109
rect 513 -509 543 -109
rect 609 -509 639 -109
rect 705 -509 735 -109
rect 801 -509 831 -109
rect 897 -509 927 -109
rect 993 -509 1023 -109
rect 1089 -509 1119 -109
rect 1185 -509 1215 -109
rect 1281 -509 1311 -109
rect 1377 -509 1407 -109
rect -1407 -1127 -1377 -727
rect -1311 -1127 -1281 -727
rect -1215 -1127 -1185 -727
rect -1119 -1127 -1089 -727
rect -1023 -1127 -993 -727
rect -927 -1127 -897 -727
rect -831 -1127 -801 -727
rect -735 -1127 -705 -727
rect -639 -1127 -609 -727
rect -543 -1127 -513 -727
rect -447 -1127 -417 -727
rect -351 -1127 -321 -727
rect -255 -1127 -225 -727
rect -159 -1127 -129 -727
rect -63 -1127 -33 -727
rect 33 -1127 63 -727
rect 129 -1127 159 -727
rect 225 -1127 255 -727
rect 321 -1127 351 -727
rect 417 -1127 447 -727
rect 513 -1127 543 -727
rect 609 -1127 639 -727
rect 705 -1127 735 -727
rect 801 -1127 831 -727
rect 897 -1127 927 -727
rect 993 -1127 1023 -727
rect 1089 -1127 1119 -727
rect 1185 -1127 1215 -727
rect 1281 -1127 1311 -727
rect 1377 -1127 1407 -727
<< ndiff >>
rect -1469 1115 -1407 1127
rect -1469 739 -1457 1115
rect -1423 739 -1407 1115
rect -1469 727 -1407 739
rect -1377 1115 -1311 1127
rect -1377 739 -1361 1115
rect -1327 739 -1311 1115
rect -1377 727 -1311 739
rect -1281 1115 -1215 1127
rect -1281 739 -1265 1115
rect -1231 739 -1215 1115
rect -1281 727 -1215 739
rect -1185 1115 -1119 1127
rect -1185 739 -1169 1115
rect -1135 739 -1119 1115
rect -1185 727 -1119 739
rect -1089 1115 -1023 1127
rect -1089 739 -1073 1115
rect -1039 739 -1023 1115
rect -1089 727 -1023 739
rect -993 1115 -927 1127
rect -993 739 -977 1115
rect -943 739 -927 1115
rect -993 727 -927 739
rect -897 1115 -831 1127
rect -897 739 -881 1115
rect -847 739 -831 1115
rect -897 727 -831 739
rect -801 1115 -735 1127
rect -801 739 -785 1115
rect -751 739 -735 1115
rect -801 727 -735 739
rect -705 1115 -639 1127
rect -705 739 -689 1115
rect -655 739 -639 1115
rect -705 727 -639 739
rect -609 1115 -543 1127
rect -609 739 -593 1115
rect -559 739 -543 1115
rect -609 727 -543 739
rect -513 1115 -447 1127
rect -513 739 -497 1115
rect -463 739 -447 1115
rect -513 727 -447 739
rect -417 1115 -351 1127
rect -417 739 -401 1115
rect -367 739 -351 1115
rect -417 727 -351 739
rect -321 1115 -255 1127
rect -321 739 -305 1115
rect -271 739 -255 1115
rect -321 727 -255 739
rect -225 1115 -159 1127
rect -225 739 -209 1115
rect -175 739 -159 1115
rect -225 727 -159 739
rect -129 1115 -63 1127
rect -129 739 -113 1115
rect -79 739 -63 1115
rect -129 727 -63 739
rect -33 1115 33 1127
rect -33 739 -17 1115
rect 17 739 33 1115
rect -33 727 33 739
rect 63 1115 129 1127
rect 63 739 79 1115
rect 113 739 129 1115
rect 63 727 129 739
rect 159 1115 225 1127
rect 159 739 175 1115
rect 209 739 225 1115
rect 159 727 225 739
rect 255 1115 321 1127
rect 255 739 271 1115
rect 305 739 321 1115
rect 255 727 321 739
rect 351 1115 417 1127
rect 351 739 367 1115
rect 401 739 417 1115
rect 351 727 417 739
rect 447 1115 513 1127
rect 447 739 463 1115
rect 497 739 513 1115
rect 447 727 513 739
rect 543 1115 609 1127
rect 543 739 559 1115
rect 593 739 609 1115
rect 543 727 609 739
rect 639 1115 705 1127
rect 639 739 655 1115
rect 689 739 705 1115
rect 639 727 705 739
rect 735 1115 801 1127
rect 735 739 751 1115
rect 785 739 801 1115
rect 735 727 801 739
rect 831 1115 897 1127
rect 831 739 847 1115
rect 881 739 897 1115
rect 831 727 897 739
rect 927 1115 993 1127
rect 927 739 943 1115
rect 977 739 993 1115
rect 927 727 993 739
rect 1023 1115 1089 1127
rect 1023 739 1039 1115
rect 1073 739 1089 1115
rect 1023 727 1089 739
rect 1119 1115 1185 1127
rect 1119 739 1135 1115
rect 1169 739 1185 1115
rect 1119 727 1185 739
rect 1215 1115 1281 1127
rect 1215 739 1231 1115
rect 1265 739 1281 1115
rect 1215 727 1281 739
rect 1311 1115 1377 1127
rect 1311 739 1327 1115
rect 1361 739 1377 1115
rect 1311 727 1377 739
rect 1407 1115 1469 1127
rect 1407 739 1423 1115
rect 1457 739 1469 1115
rect 1407 727 1469 739
rect -1469 497 -1407 509
rect -1469 121 -1457 497
rect -1423 121 -1407 497
rect -1469 109 -1407 121
rect -1377 497 -1311 509
rect -1377 121 -1361 497
rect -1327 121 -1311 497
rect -1377 109 -1311 121
rect -1281 497 -1215 509
rect -1281 121 -1265 497
rect -1231 121 -1215 497
rect -1281 109 -1215 121
rect -1185 497 -1119 509
rect -1185 121 -1169 497
rect -1135 121 -1119 497
rect -1185 109 -1119 121
rect -1089 497 -1023 509
rect -1089 121 -1073 497
rect -1039 121 -1023 497
rect -1089 109 -1023 121
rect -993 497 -927 509
rect -993 121 -977 497
rect -943 121 -927 497
rect -993 109 -927 121
rect -897 497 -831 509
rect -897 121 -881 497
rect -847 121 -831 497
rect -897 109 -831 121
rect -801 497 -735 509
rect -801 121 -785 497
rect -751 121 -735 497
rect -801 109 -735 121
rect -705 497 -639 509
rect -705 121 -689 497
rect -655 121 -639 497
rect -705 109 -639 121
rect -609 497 -543 509
rect -609 121 -593 497
rect -559 121 -543 497
rect -609 109 -543 121
rect -513 497 -447 509
rect -513 121 -497 497
rect -463 121 -447 497
rect -513 109 -447 121
rect -417 497 -351 509
rect -417 121 -401 497
rect -367 121 -351 497
rect -417 109 -351 121
rect -321 497 -255 509
rect -321 121 -305 497
rect -271 121 -255 497
rect -321 109 -255 121
rect -225 497 -159 509
rect -225 121 -209 497
rect -175 121 -159 497
rect -225 109 -159 121
rect -129 497 -63 509
rect -129 121 -113 497
rect -79 121 -63 497
rect -129 109 -63 121
rect -33 497 33 509
rect -33 121 -17 497
rect 17 121 33 497
rect -33 109 33 121
rect 63 497 129 509
rect 63 121 79 497
rect 113 121 129 497
rect 63 109 129 121
rect 159 497 225 509
rect 159 121 175 497
rect 209 121 225 497
rect 159 109 225 121
rect 255 497 321 509
rect 255 121 271 497
rect 305 121 321 497
rect 255 109 321 121
rect 351 497 417 509
rect 351 121 367 497
rect 401 121 417 497
rect 351 109 417 121
rect 447 497 513 509
rect 447 121 463 497
rect 497 121 513 497
rect 447 109 513 121
rect 543 497 609 509
rect 543 121 559 497
rect 593 121 609 497
rect 543 109 609 121
rect 639 497 705 509
rect 639 121 655 497
rect 689 121 705 497
rect 639 109 705 121
rect 735 497 801 509
rect 735 121 751 497
rect 785 121 801 497
rect 735 109 801 121
rect 831 497 897 509
rect 831 121 847 497
rect 881 121 897 497
rect 831 109 897 121
rect 927 497 993 509
rect 927 121 943 497
rect 977 121 993 497
rect 927 109 993 121
rect 1023 497 1089 509
rect 1023 121 1039 497
rect 1073 121 1089 497
rect 1023 109 1089 121
rect 1119 497 1185 509
rect 1119 121 1135 497
rect 1169 121 1185 497
rect 1119 109 1185 121
rect 1215 497 1281 509
rect 1215 121 1231 497
rect 1265 121 1281 497
rect 1215 109 1281 121
rect 1311 497 1377 509
rect 1311 121 1327 497
rect 1361 121 1377 497
rect 1311 109 1377 121
rect 1407 497 1469 509
rect 1407 121 1423 497
rect 1457 121 1469 497
rect 1407 109 1469 121
rect -1469 -121 -1407 -109
rect -1469 -497 -1457 -121
rect -1423 -497 -1407 -121
rect -1469 -509 -1407 -497
rect -1377 -121 -1311 -109
rect -1377 -497 -1361 -121
rect -1327 -497 -1311 -121
rect -1377 -509 -1311 -497
rect -1281 -121 -1215 -109
rect -1281 -497 -1265 -121
rect -1231 -497 -1215 -121
rect -1281 -509 -1215 -497
rect -1185 -121 -1119 -109
rect -1185 -497 -1169 -121
rect -1135 -497 -1119 -121
rect -1185 -509 -1119 -497
rect -1089 -121 -1023 -109
rect -1089 -497 -1073 -121
rect -1039 -497 -1023 -121
rect -1089 -509 -1023 -497
rect -993 -121 -927 -109
rect -993 -497 -977 -121
rect -943 -497 -927 -121
rect -993 -509 -927 -497
rect -897 -121 -831 -109
rect -897 -497 -881 -121
rect -847 -497 -831 -121
rect -897 -509 -831 -497
rect -801 -121 -735 -109
rect -801 -497 -785 -121
rect -751 -497 -735 -121
rect -801 -509 -735 -497
rect -705 -121 -639 -109
rect -705 -497 -689 -121
rect -655 -497 -639 -121
rect -705 -509 -639 -497
rect -609 -121 -543 -109
rect -609 -497 -593 -121
rect -559 -497 -543 -121
rect -609 -509 -543 -497
rect -513 -121 -447 -109
rect -513 -497 -497 -121
rect -463 -497 -447 -121
rect -513 -509 -447 -497
rect -417 -121 -351 -109
rect -417 -497 -401 -121
rect -367 -497 -351 -121
rect -417 -509 -351 -497
rect -321 -121 -255 -109
rect -321 -497 -305 -121
rect -271 -497 -255 -121
rect -321 -509 -255 -497
rect -225 -121 -159 -109
rect -225 -497 -209 -121
rect -175 -497 -159 -121
rect -225 -509 -159 -497
rect -129 -121 -63 -109
rect -129 -497 -113 -121
rect -79 -497 -63 -121
rect -129 -509 -63 -497
rect -33 -121 33 -109
rect -33 -497 -17 -121
rect 17 -497 33 -121
rect -33 -509 33 -497
rect 63 -121 129 -109
rect 63 -497 79 -121
rect 113 -497 129 -121
rect 63 -509 129 -497
rect 159 -121 225 -109
rect 159 -497 175 -121
rect 209 -497 225 -121
rect 159 -509 225 -497
rect 255 -121 321 -109
rect 255 -497 271 -121
rect 305 -497 321 -121
rect 255 -509 321 -497
rect 351 -121 417 -109
rect 351 -497 367 -121
rect 401 -497 417 -121
rect 351 -509 417 -497
rect 447 -121 513 -109
rect 447 -497 463 -121
rect 497 -497 513 -121
rect 447 -509 513 -497
rect 543 -121 609 -109
rect 543 -497 559 -121
rect 593 -497 609 -121
rect 543 -509 609 -497
rect 639 -121 705 -109
rect 639 -497 655 -121
rect 689 -497 705 -121
rect 639 -509 705 -497
rect 735 -121 801 -109
rect 735 -497 751 -121
rect 785 -497 801 -121
rect 735 -509 801 -497
rect 831 -121 897 -109
rect 831 -497 847 -121
rect 881 -497 897 -121
rect 831 -509 897 -497
rect 927 -121 993 -109
rect 927 -497 943 -121
rect 977 -497 993 -121
rect 927 -509 993 -497
rect 1023 -121 1089 -109
rect 1023 -497 1039 -121
rect 1073 -497 1089 -121
rect 1023 -509 1089 -497
rect 1119 -121 1185 -109
rect 1119 -497 1135 -121
rect 1169 -497 1185 -121
rect 1119 -509 1185 -497
rect 1215 -121 1281 -109
rect 1215 -497 1231 -121
rect 1265 -497 1281 -121
rect 1215 -509 1281 -497
rect 1311 -121 1377 -109
rect 1311 -497 1327 -121
rect 1361 -497 1377 -121
rect 1311 -509 1377 -497
rect 1407 -121 1469 -109
rect 1407 -497 1423 -121
rect 1457 -497 1469 -121
rect 1407 -509 1469 -497
rect -1469 -739 -1407 -727
rect -1469 -1115 -1457 -739
rect -1423 -1115 -1407 -739
rect -1469 -1127 -1407 -1115
rect -1377 -739 -1311 -727
rect -1377 -1115 -1361 -739
rect -1327 -1115 -1311 -739
rect -1377 -1127 -1311 -1115
rect -1281 -739 -1215 -727
rect -1281 -1115 -1265 -739
rect -1231 -1115 -1215 -739
rect -1281 -1127 -1215 -1115
rect -1185 -739 -1119 -727
rect -1185 -1115 -1169 -739
rect -1135 -1115 -1119 -739
rect -1185 -1127 -1119 -1115
rect -1089 -739 -1023 -727
rect -1089 -1115 -1073 -739
rect -1039 -1115 -1023 -739
rect -1089 -1127 -1023 -1115
rect -993 -739 -927 -727
rect -993 -1115 -977 -739
rect -943 -1115 -927 -739
rect -993 -1127 -927 -1115
rect -897 -739 -831 -727
rect -897 -1115 -881 -739
rect -847 -1115 -831 -739
rect -897 -1127 -831 -1115
rect -801 -739 -735 -727
rect -801 -1115 -785 -739
rect -751 -1115 -735 -739
rect -801 -1127 -735 -1115
rect -705 -739 -639 -727
rect -705 -1115 -689 -739
rect -655 -1115 -639 -739
rect -705 -1127 -639 -1115
rect -609 -739 -543 -727
rect -609 -1115 -593 -739
rect -559 -1115 -543 -739
rect -609 -1127 -543 -1115
rect -513 -739 -447 -727
rect -513 -1115 -497 -739
rect -463 -1115 -447 -739
rect -513 -1127 -447 -1115
rect -417 -739 -351 -727
rect -417 -1115 -401 -739
rect -367 -1115 -351 -739
rect -417 -1127 -351 -1115
rect -321 -739 -255 -727
rect -321 -1115 -305 -739
rect -271 -1115 -255 -739
rect -321 -1127 -255 -1115
rect -225 -739 -159 -727
rect -225 -1115 -209 -739
rect -175 -1115 -159 -739
rect -225 -1127 -159 -1115
rect -129 -739 -63 -727
rect -129 -1115 -113 -739
rect -79 -1115 -63 -739
rect -129 -1127 -63 -1115
rect -33 -739 33 -727
rect -33 -1115 -17 -739
rect 17 -1115 33 -739
rect -33 -1127 33 -1115
rect 63 -739 129 -727
rect 63 -1115 79 -739
rect 113 -1115 129 -739
rect 63 -1127 129 -1115
rect 159 -739 225 -727
rect 159 -1115 175 -739
rect 209 -1115 225 -739
rect 159 -1127 225 -1115
rect 255 -739 321 -727
rect 255 -1115 271 -739
rect 305 -1115 321 -739
rect 255 -1127 321 -1115
rect 351 -739 417 -727
rect 351 -1115 367 -739
rect 401 -1115 417 -739
rect 351 -1127 417 -1115
rect 447 -739 513 -727
rect 447 -1115 463 -739
rect 497 -1115 513 -739
rect 447 -1127 513 -1115
rect 543 -739 609 -727
rect 543 -1115 559 -739
rect 593 -1115 609 -739
rect 543 -1127 609 -1115
rect 639 -739 705 -727
rect 639 -1115 655 -739
rect 689 -1115 705 -739
rect 639 -1127 705 -1115
rect 735 -739 801 -727
rect 735 -1115 751 -739
rect 785 -1115 801 -739
rect 735 -1127 801 -1115
rect 831 -739 897 -727
rect 831 -1115 847 -739
rect 881 -1115 897 -739
rect 831 -1127 897 -1115
rect 927 -739 993 -727
rect 927 -1115 943 -739
rect 977 -1115 993 -739
rect 927 -1127 993 -1115
rect 1023 -739 1089 -727
rect 1023 -1115 1039 -739
rect 1073 -1115 1089 -739
rect 1023 -1127 1089 -1115
rect 1119 -739 1185 -727
rect 1119 -1115 1135 -739
rect 1169 -1115 1185 -739
rect 1119 -1127 1185 -1115
rect 1215 -739 1281 -727
rect 1215 -1115 1231 -739
rect 1265 -1115 1281 -739
rect 1215 -1127 1281 -1115
rect 1311 -739 1377 -727
rect 1311 -1115 1327 -739
rect 1361 -1115 1377 -739
rect 1311 -1127 1377 -1115
rect 1407 -739 1469 -727
rect 1407 -1115 1423 -739
rect 1457 -1115 1469 -739
rect 1407 -1127 1469 -1115
<< ndiffc >>
rect -1457 739 -1423 1115
rect -1361 739 -1327 1115
rect -1265 739 -1231 1115
rect -1169 739 -1135 1115
rect -1073 739 -1039 1115
rect -977 739 -943 1115
rect -881 739 -847 1115
rect -785 739 -751 1115
rect -689 739 -655 1115
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect 655 739 689 1115
rect 751 739 785 1115
rect 847 739 881 1115
rect 943 739 977 1115
rect 1039 739 1073 1115
rect 1135 739 1169 1115
rect 1231 739 1265 1115
rect 1327 739 1361 1115
rect 1423 739 1457 1115
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect -1457 -1115 -1423 -739
rect -1361 -1115 -1327 -739
rect -1265 -1115 -1231 -739
rect -1169 -1115 -1135 -739
rect -1073 -1115 -1039 -739
rect -977 -1115 -943 -739
rect -881 -1115 -847 -739
rect -785 -1115 -751 -739
rect -689 -1115 -655 -739
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect 655 -1115 689 -739
rect 751 -1115 785 -739
rect 847 -1115 881 -739
rect 943 -1115 977 -739
rect 1039 -1115 1073 -739
rect 1135 -1115 1169 -739
rect 1231 -1115 1265 -739
rect 1327 -1115 1361 -739
rect 1423 -1115 1457 -739
<< psubdiff >>
rect -1571 1267 -1475 1301
rect 1475 1267 1571 1301
rect -1571 1205 -1537 1267
rect 1537 1205 1571 1267
rect -1571 -1267 -1537 -1205
rect 1537 -1267 1571 -1205
rect -1571 -1301 -1475 -1267
rect 1475 -1301 1571 -1267
<< psubdiffcont >>
rect -1475 1267 1475 1301
rect -1571 -1205 -1537 1205
rect 1537 -1205 1571 1205
rect -1475 -1301 1475 -1267
<< poly >>
rect -1425 1199 -1359 1215
rect -1425 1165 -1409 1199
rect -1375 1165 -1359 1199
rect -1425 1149 -1359 1165
rect -1233 1199 -1167 1215
rect -1233 1165 -1217 1199
rect -1183 1165 -1167 1199
rect -1407 1127 -1377 1149
rect -1311 1127 -1281 1153
rect -1233 1149 -1167 1165
rect -1041 1199 -975 1215
rect -1041 1165 -1025 1199
rect -991 1165 -975 1199
rect -1215 1127 -1185 1149
rect -1119 1127 -1089 1153
rect -1041 1149 -975 1165
rect -849 1199 -783 1215
rect -849 1165 -833 1199
rect -799 1165 -783 1199
rect -1023 1127 -993 1149
rect -927 1127 -897 1153
rect -849 1149 -783 1165
rect -657 1199 -591 1215
rect -657 1165 -641 1199
rect -607 1165 -591 1199
rect -831 1127 -801 1149
rect -735 1127 -705 1153
rect -657 1149 -591 1165
rect -465 1199 -399 1215
rect -465 1165 -449 1199
rect -415 1165 -399 1199
rect -639 1127 -609 1149
rect -543 1127 -513 1153
rect -465 1149 -399 1165
rect -273 1199 -207 1215
rect -273 1165 -257 1199
rect -223 1165 -207 1199
rect -447 1127 -417 1149
rect -351 1127 -321 1153
rect -273 1149 -207 1165
rect -81 1199 -15 1215
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect -255 1127 -225 1149
rect -159 1127 -129 1153
rect -81 1149 -15 1165
rect 111 1199 177 1215
rect 111 1165 127 1199
rect 161 1165 177 1199
rect -63 1127 -33 1149
rect 33 1127 63 1153
rect 111 1149 177 1165
rect 303 1199 369 1215
rect 303 1165 319 1199
rect 353 1165 369 1199
rect 129 1127 159 1149
rect 225 1127 255 1153
rect 303 1149 369 1165
rect 495 1199 561 1215
rect 495 1165 511 1199
rect 545 1165 561 1199
rect 321 1127 351 1149
rect 417 1127 447 1153
rect 495 1149 561 1165
rect 687 1199 753 1215
rect 687 1165 703 1199
rect 737 1165 753 1199
rect 513 1127 543 1149
rect 609 1127 639 1153
rect 687 1149 753 1165
rect 879 1199 945 1215
rect 879 1165 895 1199
rect 929 1165 945 1199
rect 705 1127 735 1149
rect 801 1127 831 1153
rect 879 1149 945 1165
rect 1071 1199 1137 1215
rect 1071 1165 1087 1199
rect 1121 1165 1137 1199
rect 897 1127 927 1149
rect 993 1127 1023 1153
rect 1071 1149 1137 1165
rect 1263 1199 1329 1215
rect 1263 1165 1279 1199
rect 1313 1165 1329 1199
rect 1089 1127 1119 1149
rect 1185 1127 1215 1153
rect 1263 1149 1329 1165
rect 1281 1127 1311 1149
rect 1377 1127 1407 1153
rect -1407 701 -1377 727
rect -1311 705 -1281 727
rect -1329 689 -1263 705
rect -1215 701 -1185 727
rect -1119 705 -1089 727
rect -1329 655 -1313 689
rect -1279 655 -1263 689
rect -1329 639 -1263 655
rect -1137 689 -1071 705
rect -1023 701 -993 727
rect -927 705 -897 727
rect -1137 655 -1121 689
rect -1087 655 -1071 689
rect -1137 639 -1071 655
rect -945 689 -879 705
rect -831 701 -801 727
rect -735 705 -705 727
rect -945 655 -929 689
rect -895 655 -879 689
rect -945 639 -879 655
rect -753 689 -687 705
rect -639 701 -609 727
rect -543 705 -513 727
rect -753 655 -737 689
rect -703 655 -687 689
rect -753 639 -687 655
rect -561 689 -495 705
rect -447 701 -417 727
rect -351 705 -321 727
rect -561 655 -545 689
rect -511 655 -495 689
rect -561 639 -495 655
rect -369 689 -303 705
rect -255 701 -225 727
rect -159 705 -129 727
rect -369 655 -353 689
rect -319 655 -303 689
rect -369 639 -303 655
rect -177 689 -111 705
rect -63 701 -33 727
rect 33 705 63 727
rect -177 655 -161 689
rect -127 655 -111 689
rect -177 639 -111 655
rect 15 689 81 705
rect 129 701 159 727
rect 225 705 255 727
rect 15 655 31 689
rect 65 655 81 689
rect 15 639 81 655
rect 207 689 273 705
rect 321 701 351 727
rect 417 705 447 727
rect 207 655 223 689
rect 257 655 273 689
rect 207 639 273 655
rect 399 689 465 705
rect 513 701 543 727
rect 609 705 639 727
rect 399 655 415 689
rect 449 655 465 689
rect 399 639 465 655
rect 591 689 657 705
rect 705 701 735 727
rect 801 705 831 727
rect 591 655 607 689
rect 641 655 657 689
rect 591 639 657 655
rect 783 689 849 705
rect 897 701 927 727
rect 993 705 1023 727
rect 783 655 799 689
rect 833 655 849 689
rect 783 639 849 655
rect 975 689 1041 705
rect 1089 701 1119 727
rect 1185 705 1215 727
rect 975 655 991 689
rect 1025 655 1041 689
rect 975 639 1041 655
rect 1167 689 1233 705
rect 1281 701 1311 727
rect 1377 705 1407 727
rect 1167 655 1183 689
rect 1217 655 1233 689
rect 1167 639 1233 655
rect 1359 689 1425 705
rect 1359 655 1375 689
rect 1409 655 1425 689
rect 1359 639 1425 655
rect -1329 581 -1263 597
rect -1329 547 -1313 581
rect -1279 547 -1263 581
rect -1407 509 -1377 535
rect -1329 531 -1263 547
rect -1137 581 -1071 597
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -1311 509 -1281 531
rect -1215 509 -1185 535
rect -1137 531 -1071 547
rect -945 581 -879 597
rect -945 547 -929 581
rect -895 547 -879 581
rect -1119 509 -1089 531
rect -1023 509 -993 535
rect -945 531 -879 547
rect -753 581 -687 597
rect -753 547 -737 581
rect -703 547 -687 581
rect -927 509 -897 531
rect -831 509 -801 535
rect -753 531 -687 547
rect -561 581 -495 597
rect -561 547 -545 581
rect -511 547 -495 581
rect -735 509 -705 531
rect -639 509 -609 535
rect -561 531 -495 547
rect -369 581 -303 597
rect -369 547 -353 581
rect -319 547 -303 581
rect -543 509 -513 531
rect -447 509 -417 535
rect -369 531 -303 547
rect -177 581 -111 597
rect -177 547 -161 581
rect -127 547 -111 581
rect -351 509 -321 531
rect -255 509 -225 535
rect -177 531 -111 547
rect 15 581 81 597
rect 15 547 31 581
rect 65 547 81 581
rect -159 509 -129 531
rect -63 509 -33 535
rect 15 531 81 547
rect 207 581 273 597
rect 207 547 223 581
rect 257 547 273 581
rect 33 509 63 531
rect 129 509 159 535
rect 207 531 273 547
rect 399 581 465 597
rect 399 547 415 581
rect 449 547 465 581
rect 225 509 255 531
rect 321 509 351 535
rect 399 531 465 547
rect 591 581 657 597
rect 591 547 607 581
rect 641 547 657 581
rect 417 509 447 531
rect 513 509 543 535
rect 591 531 657 547
rect 783 581 849 597
rect 783 547 799 581
rect 833 547 849 581
rect 609 509 639 531
rect 705 509 735 535
rect 783 531 849 547
rect 975 581 1041 597
rect 975 547 991 581
rect 1025 547 1041 581
rect 801 509 831 531
rect 897 509 927 535
rect 975 531 1041 547
rect 1167 581 1233 597
rect 1167 547 1183 581
rect 1217 547 1233 581
rect 993 509 1023 531
rect 1089 509 1119 535
rect 1167 531 1233 547
rect 1359 581 1425 597
rect 1359 547 1375 581
rect 1409 547 1425 581
rect 1185 509 1215 531
rect 1281 509 1311 535
rect 1359 531 1425 547
rect 1377 509 1407 531
rect -1407 87 -1377 109
rect -1425 71 -1359 87
rect -1311 83 -1281 109
rect -1215 87 -1185 109
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1425 21 -1359 37
rect -1233 71 -1167 87
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1233 21 -1167 37
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1185 83 1215 109
rect 1281 87 1311 109
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect 1263 71 1329 87
rect 1377 83 1407 109
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1263 21 1329 37
rect -1425 -37 -1359 -21
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1425 -87 -1359 -71
rect -1233 -37 -1167 -21
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -83
rect -1233 -87 -1167 -71
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1263 -37 1329 -21
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1089 -109 1119 -87
rect 1185 -109 1215 -83
rect 1263 -87 1329 -71
rect 1281 -109 1311 -87
rect 1377 -109 1407 -83
rect -1407 -535 -1377 -509
rect -1311 -531 -1281 -509
rect -1329 -547 -1263 -531
rect -1215 -535 -1185 -509
rect -1119 -531 -1089 -509
rect -1329 -581 -1313 -547
rect -1279 -581 -1263 -547
rect -1329 -597 -1263 -581
rect -1137 -547 -1071 -531
rect -1023 -535 -993 -509
rect -927 -531 -897 -509
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -1137 -597 -1071 -581
rect -945 -547 -879 -531
rect -831 -535 -801 -509
rect -735 -531 -705 -509
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -945 -597 -879 -581
rect -753 -547 -687 -531
rect -639 -535 -609 -509
rect -543 -531 -513 -509
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -753 -597 -687 -581
rect -561 -547 -495 -531
rect -447 -535 -417 -509
rect -351 -531 -321 -509
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -255 -535 -225 -509
rect -159 -531 -129 -509
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -63 -535 -33 -509
rect 33 -531 63 -509
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 129 -535 159 -509
rect 225 -531 255 -509
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 321 -535 351 -509
rect 417 -531 447 -509
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 513 -535 543 -509
rect 609 -531 639 -509
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
rect 591 -547 657 -531
rect 705 -535 735 -509
rect 801 -531 831 -509
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 591 -597 657 -581
rect 783 -547 849 -531
rect 897 -535 927 -509
rect 993 -531 1023 -509
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 783 -597 849 -581
rect 975 -547 1041 -531
rect 1089 -535 1119 -509
rect 1185 -531 1215 -509
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 975 -597 1041 -581
rect 1167 -547 1233 -531
rect 1281 -535 1311 -509
rect 1377 -531 1407 -509
rect 1167 -581 1183 -547
rect 1217 -581 1233 -547
rect 1167 -597 1233 -581
rect 1359 -547 1425 -531
rect 1359 -581 1375 -547
rect 1409 -581 1425 -547
rect 1359 -597 1425 -581
rect -1329 -655 -1263 -639
rect -1329 -689 -1313 -655
rect -1279 -689 -1263 -655
rect -1407 -727 -1377 -701
rect -1329 -705 -1263 -689
rect -1137 -655 -1071 -639
rect -1137 -689 -1121 -655
rect -1087 -689 -1071 -655
rect -1311 -727 -1281 -705
rect -1215 -727 -1185 -701
rect -1137 -705 -1071 -689
rect -945 -655 -879 -639
rect -945 -689 -929 -655
rect -895 -689 -879 -655
rect -1119 -727 -1089 -705
rect -1023 -727 -993 -701
rect -945 -705 -879 -689
rect -753 -655 -687 -639
rect -753 -689 -737 -655
rect -703 -689 -687 -655
rect -927 -727 -897 -705
rect -831 -727 -801 -701
rect -753 -705 -687 -689
rect -561 -655 -495 -639
rect -561 -689 -545 -655
rect -511 -689 -495 -655
rect -735 -727 -705 -705
rect -639 -727 -609 -701
rect -561 -705 -495 -689
rect -369 -655 -303 -639
rect -369 -689 -353 -655
rect -319 -689 -303 -655
rect -543 -727 -513 -705
rect -447 -727 -417 -701
rect -369 -705 -303 -689
rect -177 -655 -111 -639
rect -177 -689 -161 -655
rect -127 -689 -111 -655
rect -351 -727 -321 -705
rect -255 -727 -225 -701
rect -177 -705 -111 -689
rect 15 -655 81 -639
rect 15 -689 31 -655
rect 65 -689 81 -655
rect -159 -727 -129 -705
rect -63 -727 -33 -701
rect 15 -705 81 -689
rect 207 -655 273 -639
rect 207 -689 223 -655
rect 257 -689 273 -655
rect 33 -727 63 -705
rect 129 -727 159 -701
rect 207 -705 273 -689
rect 399 -655 465 -639
rect 399 -689 415 -655
rect 449 -689 465 -655
rect 225 -727 255 -705
rect 321 -727 351 -701
rect 399 -705 465 -689
rect 591 -655 657 -639
rect 591 -689 607 -655
rect 641 -689 657 -655
rect 417 -727 447 -705
rect 513 -727 543 -701
rect 591 -705 657 -689
rect 783 -655 849 -639
rect 783 -689 799 -655
rect 833 -689 849 -655
rect 609 -727 639 -705
rect 705 -727 735 -701
rect 783 -705 849 -689
rect 975 -655 1041 -639
rect 975 -689 991 -655
rect 1025 -689 1041 -655
rect 801 -727 831 -705
rect 897 -727 927 -701
rect 975 -705 1041 -689
rect 1167 -655 1233 -639
rect 1167 -689 1183 -655
rect 1217 -689 1233 -655
rect 993 -727 1023 -705
rect 1089 -727 1119 -701
rect 1167 -705 1233 -689
rect 1359 -655 1425 -639
rect 1359 -689 1375 -655
rect 1409 -689 1425 -655
rect 1185 -727 1215 -705
rect 1281 -727 1311 -701
rect 1359 -705 1425 -689
rect 1377 -727 1407 -705
rect -1407 -1149 -1377 -1127
rect -1425 -1165 -1359 -1149
rect -1311 -1153 -1281 -1127
rect -1215 -1149 -1185 -1127
rect -1425 -1199 -1409 -1165
rect -1375 -1199 -1359 -1165
rect -1425 -1215 -1359 -1199
rect -1233 -1165 -1167 -1149
rect -1119 -1153 -1089 -1127
rect -1023 -1149 -993 -1127
rect -1233 -1199 -1217 -1165
rect -1183 -1199 -1167 -1165
rect -1233 -1215 -1167 -1199
rect -1041 -1165 -975 -1149
rect -927 -1153 -897 -1127
rect -831 -1149 -801 -1127
rect -1041 -1199 -1025 -1165
rect -991 -1199 -975 -1165
rect -1041 -1215 -975 -1199
rect -849 -1165 -783 -1149
rect -735 -1153 -705 -1127
rect -639 -1149 -609 -1127
rect -849 -1199 -833 -1165
rect -799 -1199 -783 -1165
rect -849 -1215 -783 -1199
rect -657 -1165 -591 -1149
rect -543 -1153 -513 -1127
rect -447 -1149 -417 -1127
rect -657 -1199 -641 -1165
rect -607 -1199 -591 -1165
rect -657 -1215 -591 -1199
rect -465 -1165 -399 -1149
rect -351 -1153 -321 -1127
rect -255 -1149 -225 -1127
rect -465 -1199 -449 -1165
rect -415 -1199 -399 -1165
rect -465 -1215 -399 -1199
rect -273 -1165 -207 -1149
rect -159 -1153 -129 -1127
rect -63 -1149 -33 -1127
rect -273 -1199 -257 -1165
rect -223 -1199 -207 -1165
rect -273 -1215 -207 -1199
rect -81 -1165 -15 -1149
rect 33 -1153 63 -1127
rect 129 -1149 159 -1127
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect -81 -1215 -15 -1199
rect 111 -1165 177 -1149
rect 225 -1153 255 -1127
rect 321 -1149 351 -1127
rect 111 -1199 127 -1165
rect 161 -1199 177 -1165
rect 111 -1215 177 -1199
rect 303 -1165 369 -1149
rect 417 -1153 447 -1127
rect 513 -1149 543 -1127
rect 303 -1199 319 -1165
rect 353 -1199 369 -1165
rect 303 -1215 369 -1199
rect 495 -1165 561 -1149
rect 609 -1153 639 -1127
rect 705 -1149 735 -1127
rect 495 -1199 511 -1165
rect 545 -1199 561 -1165
rect 495 -1215 561 -1199
rect 687 -1165 753 -1149
rect 801 -1153 831 -1127
rect 897 -1149 927 -1127
rect 687 -1199 703 -1165
rect 737 -1199 753 -1165
rect 687 -1215 753 -1199
rect 879 -1165 945 -1149
rect 993 -1153 1023 -1127
rect 1089 -1149 1119 -1127
rect 879 -1199 895 -1165
rect 929 -1199 945 -1165
rect 879 -1215 945 -1199
rect 1071 -1165 1137 -1149
rect 1185 -1153 1215 -1127
rect 1281 -1149 1311 -1127
rect 1071 -1199 1087 -1165
rect 1121 -1199 1137 -1165
rect 1071 -1215 1137 -1199
rect 1263 -1165 1329 -1149
rect 1377 -1153 1407 -1127
rect 1263 -1199 1279 -1165
rect 1313 -1199 1329 -1165
rect 1263 -1215 1329 -1199
<< polycont >>
rect -1409 1165 -1375 1199
rect -1217 1165 -1183 1199
rect -1025 1165 -991 1199
rect -833 1165 -799 1199
rect -641 1165 -607 1199
rect -449 1165 -415 1199
rect -257 1165 -223 1199
rect -65 1165 -31 1199
rect 127 1165 161 1199
rect 319 1165 353 1199
rect 511 1165 545 1199
rect 703 1165 737 1199
rect 895 1165 929 1199
rect 1087 1165 1121 1199
rect 1279 1165 1313 1199
rect -1313 655 -1279 689
rect -1121 655 -1087 689
rect -929 655 -895 689
rect -737 655 -703 689
rect -545 655 -511 689
rect -353 655 -319 689
rect -161 655 -127 689
rect 31 655 65 689
rect 223 655 257 689
rect 415 655 449 689
rect 607 655 641 689
rect 799 655 833 689
rect 991 655 1025 689
rect 1183 655 1217 689
rect 1375 655 1409 689
rect -1313 547 -1279 581
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect 1183 547 1217 581
rect 1375 547 1409 581
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect -1313 -581 -1279 -547
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect 1183 -581 1217 -547
rect 1375 -581 1409 -547
rect -1313 -689 -1279 -655
rect -1121 -689 -1087 -655
rect -929 -689 -895 -655
rect -737 -689 -703 -655
rect -545 -689 -511 -655
rect -353 -689 -319 -655
rect -161 -689 -127 -655
rect 31 -689 65 -655
rect 223 -689 257 -655
rect 415 -689 449 -655
rect 607 -689 641 -655
rect 799 -689 833 -655
rect 991 -689 1025 -655
rect 1183 -689 1217 -655
rect 1375 -689 1409 -655
rect -1409 -1199 -1375 -1165
rect -1217 -1199 -1183 -1165
rect -1025 -1199 -991 -1165
rect -833 -1199 -799 -1165
rect -641 -1199 -607 -1165
rect -449 -1199 -415 -1165
rect -257 -1199 -223 -1165
rect -65 -1199 -31 -1165
rect 127 -1199 161 -1165
rect 319 -1199 353 -1165
rect 511 -1199 545 -1165
rect 703 -1199 737 -1165
rect 895 -1199 929 -1165
rect 1087 -1199 1121 -1165
rect 1279 -1199 1313 -1165
<< locali >>
rect -1571 1267 -1475 1301
rect 1475 1267 1571 1301
rect -1571 1205 -1537 1267
rect 1537 1205 1571 1267
rect -1425 1165 -1409 1199
rect -1375 1165 -1359 1199
rect -1233 1165 -1217 1199
rect -1183 1165 -1167 1199
rect -1041 1165 -1025 1199
rect -991 1165 -975 1199
rect -849 1165 -833 1199
rect -799 1165 -783 1199
rect -657 1165 -641 1199
rect -607 1165 -591 1199
rect -465 1165 -449 1199
rect -415 1165 -399 1199
rect -273 1165 -257 1199
rect -223 1165 -207 1199
rect -81 1165 -65 1199
rect -31 1165 -15 1199
rect 111 1165 127 1199
rect 161 1165 177 1199
rect 303 1165 319 1199
rect 353 1165 369 1199
rect 495 1165 511 1199
rect 545 1165 561 1199
rect 687 1165 703 1199
rect 737 1165 753 1199
rect 879 1165 895 1199
rect 929 1165 945 1199
rect 1071 1165 1087 1199
rect 1121 1165 1137 1199
rect 1263 1165 1279 1199
rect 1313 1165 1329 1199
rect -1457 1115 -1423 1131
rect -1457 723 -1423 739
rect -1361 1115 -1327 1131
rect -1361 723 -1327 739
rect -1265 1115 -1231 1131
rect -1265 723 -1231 739
rect -1169 1115 -1135 1131
rect -1169 723 -1135 739
rect -1073 1115 -1039 1131
rect -1073 723 -1039 739
rect -977 1115 -943 1131
rect -977 723 -943 739
rect -881 1115 -847 1131
rect -881 723 -847 739
rect -785 1115 -751 1131
rect -785 723 -751 739
rect -689 1115 -655 1131
rect -689 723 -655 739
rect -593 1115 -559 1131
rect -593 723 -559 739
rect -497 1115 -463 1131
rect -497 723 -463 739
rect -401 1115 -367 1131
rect -401 723 -367 739
rect -305 1115 -271 1131
rect -305 723 -271 739
rect -209 1115 -175 1131
rect -209 723 -175 739
rect -113 1115 -79 1131
rect -113 723 -79 739
rect -17 1115 17 1131
rect -17 723 17 739
rect 79 1115 113 1131
rect 79 723 113 739
rect 175 1115 209 1131
rect 175 723 209 739
rect 271 1115 305 1131
rect 271 723 305 739
rect 367 1115 401 1131
rect 367 723 401 739
rect 463 1115 497 1131
rect 463 723 497 739
rect 559 1115 593 1131
rect 559 723 593 739
rect 655 1115 689 1131
rect 655 723 689 739
rect 751 1115 785 1131
rect 751 723 785 739
rect 847 1115 881 1131
rect 847 723 881 739
rect 943 1115 977 1131
rect 943 723 977 739
rect 1039 1115 1073 1131
rect 1039 723 1073 739
rect 1135 1115 1169 1131
rect 1135 723 1169 739
rect 1231 1115 1265 1131
rect 1231 723 1265 739
rect 1327 1115 1361 1131
rect 1327 723 1361 739
rect 1423 1115 1457 1131
rect 1423 723 1457 739
rect -1329 655 -1313 689
rect -1279 655 -1263 689
rect -1137 655 -1121 689
rect -1087 655 -1071 689
rect -945 655 -929 689
rect -895 655 -879 689
rect -753 655 -737 689
rect -703 655 -687 689
rect -561 655 -545 689
rect -511 655 -495 689
rect -369 655 -353 689
rect -319 655 -303 689
rect -177 655 -161 689
rect -127 655 -111 689
rect 15 655 31 689
rect 65 655 81 689
rect 207 655 223 689
rect 257 655 273 689
rect 399 655 415 689
rect 449 655 465 689
rect 591 655 607 689
rect 641 655 657 689
rect 783 655 799 689
rect 833 655 849 689
rect 975 655 991 689
rect 1025 655 1041 689
rect 1167 655 1183 689
rect 1217 655 1233 689
rect 1359 655 1375 689
rect 1409 655 1425 689
rect -1329 547 -1313 581
rect -1279 547 -1263 581
rect -1137 547 -1121 581
rect -1087 547 -1071 581
rect -945 547 -929 581
rect -895 547 -879 581
rect -753 547 -737 581
rect -703 547 -687 581
rect -561 547 -545 581
rect -511 547 -495 581
rect -369 547 -353 581
rect -319 547 -303 581
rect -177 547 -161 581
rect -127 547 -111 581
rect 15 547 31 581
rect 65 547 81 581
rect 207 547 223 581
rect 257 547 273 581
rect 399 547 415 581
rect 449 547 465 581
rect 591 547 607 581
rect 641 547 657 581
rect 783 547 799 581
rect 833 547 849 581
rect 975 547 991 581
rect 1025 547 1041 581
rect 1167 547 1183 581
rect 1217 547 1233 581
rect 1359 547 1375 581
rect 1409 547 1425 581
rect -1457 497 -1423 513
rect -1457 105 -1423 121
rect -1361 497 -1327 513
rect -1361 105 -1327 121
rect -1265 497 -1231 513
rect -1265 105 -1231 121
rect -1169 497 -1135 513
rect -1169 105 -1135 121
rect -1073 497 -1039 513
rect -1073 105 -1039 121
rect -977 497 -943 513
rect -977 105 -943 121
rect -881 497 -847 513
rect -881 105 -847 121
rect -785 497 -751 513
rect -785 105 -751 121
rect -689 497 -655 513
rect -689 105 -655 121
rect -593 497 -559 513
rect -593 105 -559 121
rect -497 497 -463 513
rect -497 105 -463 121
rect -401 497 -367 513
rect -401 105 -367 121
rect -305 497 -271 513
rect -305 105 -271 121
rect -209 497 -175 513
rect -209 105 -175 121
rect -113 497 -79 513
rect -113 105 -79 121
rect -17 497 17 513
rect -17 105 17 121
rect 79 497 113 513
rect 79 105 113 121
rect 175 497 209 513
rect 175 105 209 121
rect 271 497 305 513
rect 271 105 305 121
rect 367 497 401 513
rect 367 105 401 121
rect 463 497 497 513
rect 463 105 497 121
rect 559 497 593 513
rect 559 105 593 121
rect 655 497 689 513
rect 655 105 689 121
rect 751 497 785 513
rect 751 105 785 121
rect 847 497 881 513
rect 847 105 881 121
rect 943 497 977 513
rect 943 105 977 121
rect 1039 497 1073 513
rect 1039 105 1073 121
rect 1135 497 1169 513
rect 1135 105 1169 121
rect 1231 497 1265 513
rect 1231 105 1265 121
rect 1327 497 1361 513
rect 1327 105 1361 121
rect 1423 497 1457 513
rect 1423 105 1457 121
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1263 37 1279 71
rect 1313 37 1329 71
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect -1457 -121 -1423 -105
rect -1457 -513 -1423 -497
rect -1361 -121 -1327 -105
rect -1361 -513 -1327 -497
rect -1265 -121 -1231 -105
rect -1265 -513 -1231 -497
rect -1169 -121 -1135 -105
rect -1169 -513 -1135 -497
rect -1073 -121 -1039 -105
rect -1073 -513 -1039 -497
rect -977 -121 -943 -105
rect -977 -513 -943 -497
rect -881 -121 -847 -105
rect -881 -513 -847 -497
rect -785 -121 -751 -105
rect -785 -513 -751 -497
rect -689 -121 -655 -105
rect -689 -513 -655 -497
rect -593 -121 -559 -105
rect -593 -513 -559 -497
rect -497 -121 -463 -105
rect -497 -513 -463 -497
rect -401 -121 -367 -105
rect -401 -513 -367 -497
rect -305 -121 -271 -105
rect -305 -513 -271 -497
rect -209 -121 -175 -105
rect -209 -513 -175 -497
rect -113 -121 -79 -105
rect -113 -513 -79 -497
rect -17 -121 17 -105
rect -17 -513 17 -497
rect 79 -121 113 -105
rect 79 -513 113 -497
rect 175 -121 209 -105
rect 175 -513 209 -497
rect 271 -121 305 -105
rect 271 -513 305 -497
rect 367 -121 401 -105
rect 367 -513 401 -497
rect 463 -121 497 -105
rect 463 -513 497 -497
rect 559 -121 593 -105
rect 559 -513 593 -497
rect 655 -121 689 -105
rect 655 -513 689 -497
rect 751 -121 785 -105
rect 751 -513 785 -497
rect 847 -121 881 -105
rect 847 -513 881 -497
rect 943 -121 977 -105
rect 943 -513 977 -497
rect 1039 -121 1073 -105
rect 1039 -513 1073 -497
rect 1135 -121 1169 -105
rect 1135 -513 1169 -497
rect 1231 -121 1265 -105
rect 1231 -513 1265 -497
rect 1327 -121 1361 -105
rect 1327 -513 1361 -497
rect 1423 -121 1457 -105
rect 1423 -513 1457 -497
rect -1329 -581 -1313 -547
rect -1279 -581 -1263 -547
rect -1137 -581 -1121 -547
rect -1087 -581 -1071 -547
rect -945 -581 -929 -547
rect -895 -581 -879 -547
rect -753 -581 -737 -547
rect -703 -581 -687 -547
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 591 -581 607 -547
rect 641 -581 657 -547
rect 783 -581 799 -547
rect 833 -581 849 -547
rect 975 -581 991 -547
rect 1025 -581 1041 -547
rect 1167 -581 1183 -547
rect 1217 -581 1233 -547
rect 1359 -581 1375 -547
rect 1409 -581 1425 -547
rect -1329 -689 -1313 -655
rect -1279 -689 -1263 -655
rect -1137 -689 -1121 -655
rect -1087 -689 -1071 -655
rect -945 -689 -929 -655
rect -895 -689 -879 -655
rect -753 -689 -737 -655
rect -703 -689 -687 -655
rect -561 -689 -545 -655
rect -511 -689 -495 -655
rect -369 -689 -353 -655
rect -319 -689 -303 -655
rect -177 -689 -161 -655
rect -127 -689 -111 -655
rect 15 -689 31 -655
rect 65 -689 81 -655
rect 207 -689 223 -655
rect 257 -689 273 -655
rect 399 -689 415 -655
rect 449 -689 465 -655
rect 591 -689 607 -655
rect 641 -689 657 -655
rect 783 -689 799 -655
rect 833 -689 849 -655
rect 975 -689 991 -655
rect 1025 -689 1041 -655
rect 1167 -689 1183 -655
rect 1217 -689 1233 -655
rect 1359 -689 1375 -655
rect 1409 -689 1425 -655
rect -1457 -739 -1423 -723
rect -1457 -1131 -1423 -1115
rect -1361 -739 -1327 -723
rect -1361 -1131 -1327 -1115
rect -1265 -739 -1231 -723
rect -1265 -1131 -1231 -1115
rect -1169 -739 -1135 -723
rect -1169 -1131 -1135 -1115
rect -1073 -739 -1039 -723
rect -1073 -1131 -1039 -1115
rect -977 -739 -943 -723
rect -977 -1131 -943 -1115
rect -881 -739 -847 -723
rect -881 -1131 -847 -1115
rect -785 -739 -751 -723
rect -785 -1131 -751 -1115
rect -689 -739 -655 -723
rect -689 -1131 -655 -1115
rect -593 -739 -559 -723
rect -593 -1131 -559 -1115
rect -497 -739 -463 -723
rect -497 -1131 -463 -1115
rect -401 -739 -367 -723
rect -401 -1131 -367 -1115
rect -305 -739 -271 -723
rect -305 -1131 -271 -1115
rect -209 -739 -175 -723
rect -209 -1131 -175 -1115
rect -113 -739 -79 -723
rect -113 -1131 -79 -1115
rect -17 -739 17 -723
rect -17 -1131 17 -1115
rect 79 -739 113 -723
rect 79 -1131 113 -1115
rect 175 -739 209 -723
rect 175 -1131 209 -1115
rect 271 -739 305 -723
rect 271 -1131 305 -1115
rect 367 -739 401 -723
rect 367 -1131 401 -1115
rect 463 -739 497 -723
rect 463 -1131 497 -1115
rect 559 -739 593 -723
rect 559 -1131 593 -1115
rect 655 -739 689 -723
rect 655 -1131 689 -1115
rect 751 -739 785 -723
rect 751 -1131 785 -1115
rect 847 -739 881 -723
rect 847 -1131 881 -1115
rect 943 -739 977 -723
rect 943 -1131 977 -1115
rect 1039 -739 1073 -723
rect 1039 -1131 1073 -1115
rect 1135 -739 1169 -723
rect 1135 -1131 1169 -1115
rect 1231 -739 1265 -723
rect 1231 -1131 1265 -1115
rect 1327 -739 1361 -723
rect 1327 -1131 1361 -1115
rect 1423 -739 1457 -723
rect 1423 -1131 1457 -1115
rect -1425 -1199 -1409 -1165
rect -1375 -1199 -1359 -1165
rect -1233 -1199 -1217 -1165
rect -1183 -1199 -1167 -1165
rect -1041 -1199 -1025 -1165
rect -991 -1199 -975 -1165
rect -849 -1199 -833 -1165
rect -799 -1199 -783 -1165
rect -657 -1199 -641 -1165
rect -607 -1199 -591 -1165
rect -465 -1199 -449 -1165
rect -415 -1199 -399 -1165
rect -273 -1199 -257 -1165
rect -223 -1199 -207 -1165
rect -81 -1199 -65 -1165
rect -31 -1199 -15 -1165
rect 111 -1199 127 -1165
rect 161 -1199 177 -1165
rect 303 -1199 319 -1165
rect 353 -1199 369 -1165
rect 495 -1199 511 -1165
rect 545 -1199 561 -1165
rect 687 -1199 703 -1165
rect 737 -1199 753 -1165
rect 879 -1199 895 -1165
rect 929 -1199 945 -1165
rect 1071 -1199 1087 -1165
rect 1121 -1199 1137 -1165
rect 1263 -1199 1279 -1165
rect 1313 -1199 1329 -1165
rect -1571 -1267 -1537 -1205
rect 1537 -1267 1571 -1205
rect -1571 -1301 -1475 -1267
rect 1475 -1301 1571 -1267
<< viali >>
rect -1409 1165 -1375 1199
rect -1217 1165 -1183 1199
rect -1025 1165 -991 1199
rect -833 1165 -799 1199
rect -641 1165 -607 1199
rect -449 1165 -415 1199
rect -257 1165 -223 1199
rect -65 1165 -31 1199
rect 127 1165 161 1199
rect 319 1165 353 1199
rect 511 1165 545 1199
rect 703 1165 737 1199
rect 895 1165 929 1199
rect 1087 1165 1121 1199
rect 1279 1165 1313 1199
rect -1457 739 -1423 1115
rect -1361 739 -1327 1115
rect -1265 739 -1231 1115
rect -1169 739 -1135 1115
rect -1073 739 -1039 1115
rect -977 739 -943 1115
rect -881 739 -847 1115
rect -785 739 -751 1115
rect -689 739 -655 1115
rect -593 739 -559 1115
rect -497 739 -463 1115
rect -401 739 -367 1115
rect -305 739 -271 1115
rect -209 739 -175 1115
rect -113 739 -79 1115
rect -17 739 17 1115
rect 79 739 113 1115
rect 175 739 209 1115
rect 271 739 305 1115
rect 367 739 401 1115
rect 463 739 497 1115
rect 559 739 593 1115
rect 655 739 689 1115
rect 751 739 785 1115
rect 847 739 881 1115
rect 943 739 977 1115
rect 1039 739 1073 1115
rect 1135 739 1169 1115
rect 1231 739 1265 1115
rect 1327 739 1361 1115
rect 1423 739 1457 1115
rect -1313 655 -1279 689
rect -1121 655 -1087 689
rect -929 655 -895 689
rect -737 655 -703 689
rect -545 655 -511 689
rect -353 655 -319 689
rect -161 655 -127 689
rect 31 655 65 689
rect 223 655 257 689
rect 415 655 449 689
rect 607 655 641 689
rect 799 655 833 689
rect 991 655 1025 689
rect 1183 655 1217 689
rect 1375 655 1409 689
rect -1313 547 -1279 581
rect -1121 547 -1087 581
rect -929 547 -895 581
rect -737 547 -703 581
rect -545 547 -511 581
rect -353 547 -319 581
rect -161 547 -127 581
rect 31 547 65 581
rect 223 547 257 581
rect 415 547 449 581
rect 607 547 641 581
rect 799 547 833 581
rect 991 547 1025 581
rect 1183 547 1217 581
rect 1375 547 1409 581
rect -1457 121 -1423 497
rect -1361 121 -1327 497
rect -1265 121 -1231 497
rect -1169 121 -1135 497
rect -1073 121 -1039 497
rect -977 121 -943 497
rect -881 121 -847 497
rect -785 121 -751 497
rect -689 121 -655 497
rect -593 121 -559 497
rect -497 121 -463 497
rect -401 121 -367 497
rect -305 121 -271 497
rect -209 121 -175 497
rect -113 121 -79 497
rect -17 121 17 497
rect 79 121 113 497
rect 175 121 209 497
rect 271 121 305 497
rect 367 121 401 497
rect 463 121 497 497
rect 559 121 593 497
rect 655 121 689 497
rect 751 121 785 497
rect 847 121 881 497
rect 943 121 977 497
rect 1039 121 1073 497
rect 1135 121 1169 497
rect 1231 121 1265 497
rect 1327 121 1361 497
rect 1423 121 1457 497
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect -1457 -497 -1423 -121
rect -1361 -497 -1327 -121
rect -1265 -497 -1231 -121
rect -1169 -497 -1135 -121
rect -1073 -497 -1039 -121
rect -977 -497 -943 -121
rect -881 -497 -847 -121
rect -785 -497 -751 -121
rect -689 -497 -655 -121
rect -593 -497 -559 -121
rect -497 -497 -463 -121
rect -401 -497 -367 -121
rect -305 -497 -271 -121
rect -209 -497 -175 -121
rect -113 -497 -79 -121
rect -17 -497 17 -121
rect 79 -497 113 -121
rect 175 -497 209 -121
rect 271 -497 305 -121
rect 367 -497 401 -121
rect 463 -497 497 -121
rect 559 -497 593 -121
rect 655 -497 689 -121
rect 751 -497 785 -121
rect 847 -497 881 -121
rect 943 -497 977 -121
rect 1039 -497 1073 -121
rect 1135 -497 1169 -121
rect 1231 -497 1265 -121
rect 1327 -497 1361 -121
rect 1423 -497 1457 -121
rect -1313 -581 -1279 -547
rect -1121 -581 -1087 -547
rect -929 -581 -895 -547
rect -737 -581 -703 -547
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
rect 607 -581 641 -547
rect 799 -581 833 -547
rect 991 -581 1025 -547
rect 1183 -581 1217 -547
rect 1375 -581 1409 -547
rect -1313 -689 -1279 -655
rect -1121 -689 -1087 -655
rect -929 -689 -895 -655
rect -737 -689 -703 -655
rect -545 -689 -511 -655
rect -353 -689 -319 -655
rect -161 -689 -127 -655
rect 31 -689 65 -655
rect 223 -689 257 -655
rect 415 -689 449 -655
rect 607 -689 641 -655
rect 799 -689 833 -655
rect 991 -689 1025 -655
rect 1183 -689 1217 -655
rect 1375 -689 1409 -655
rect -1457 -1115 -1423 -739
rect -1361 -1115 -1327 -739
rect -1265 -1115 -1231 -739
rect -1169 -1115 -1135 -739
rect -1073 -1115 -1039 -739
rect -977 -1115 -943 -739
rect -881 -1115 -847 -739
rect -785 -1115 -751 -739
rect -689 -1115 -655 -739
rect -593 -1115 -559 -739
rect -497 -1115 -463 -739
rect -401 -1115 -367 -739
rect -305 -1115 -271 -739
rect -209 -1115 -175 -739
rect -113 -1115 -79 -739
rect -17 -1115 17 -739
rect 79 -1115 113 -739
rect 175 -1115 209 -739
rect 271 -1115 305 -739
rect 367 -1115 401 -739
rect 463 -1115 497 -739
rect 559 -1115 593 -739
rect 655 -1115 689 -739
rect 751 -1115 785 -739
rect 847 -1115 881 -739
rect 943 -1115 977 -739
rect 1039 -1115 1073 -739
rect 1135 -1115 1169 -739
rect 1231 -1115 1265 -739
rect 1327 -1115 1361 -739
rect 1423 -1115 1457 -739
rect -1409 -1199 -1375 -1165
rect -1217 -1199 -1183 -1165
rect -1025 -1199 -991 -1165
rect -833 -1199 -799 -1165
rect -641 -1199 -607 -1165
rect -449 -1199 -415 -1165
rect -257 -1199 -223 -1165
rect -65 -1199 -31 -1165
rect 127 -1199 161 -1165
rect 319 -1199 353 -1165
rect 511 -1199 545 -1165
rect 703 -1199 737 -1165
rect 895 -1199 929 -1165
rect 1087 -1199 1121 -1165
rect 1279 -1199 1313 -1165
<< metal1 >>
rect -1421 1199 -1363 1205
rect -1421 1165 -1409 1199
rect -1375 1165 -1363 1199
rect -1421 1159 -1363 1165
rect -1229 1199 -1171 1205
rect -1229 1165 -1217 1199
rect -1183 1165 -1171 1199
rect -1229 1159 -1171 1165
rect -1037 1199 -979 1205
rect -1037 1165 -1025 1199
rect -991 1165 -979 1199
rect -1037 1159 -979 1165
rect -845 1199 -787 1205
rect -845 1165 -833 1199
rect -799 1165 -787 1199
rect -845 1159 -787 1165
rect -653 1199 -595 1205
rect -653 1165 -641 1199
rect -607 1165 -595 1199
rect -653 1159 -595 1165
rect -461 1199 -403 1205
rect -461 1165 -449 1199
rect -415 1165 -403 1199
rect -461 1159 -403 1165
rect -269 1199 -211 1205
rect -269 1165 -257 1199
rect -223 1165 -211 1199
rect -269 1159 -211 1165
rect -77 1199 -19 1205
rect -77 1165 -65 1199
rect -31 1165 -19 1199
rect -77 1159 -19 1165
rect 115 1199 173 1205
rect 115 1165 127 1199
rect 161 1165 173 1199
rect 115 1159 173 1165
rect 307 1199 365 1205
rect 307 1165 319 1199
rect 353 1165 365 1199
rect 307 1159 365 1165
rect 499 1199 557 1205
rect 499 1165 511 1199
rect 545 1165 557 1199
rect 499 1159 557 1165
rect 691 1199 749 1205
rect 691 1165 703 1199
rect 737 1165 749 1199
rect 691 1159 749 1165
rect 883 1199 941 1205
rect 883 1165 895 1199
rect 929 1165 941 1199
rect 883 1159 941 1165
rect 1075 1199 1133 1205
rect 1075 1165 1087 1199
rect 1121 1165 1133 1199
rect 1075 1159 1133 1165
rect 1267 1199 1325 1205
rect 1267 1165 1279 1199
rect 1313 1165 1325 1199
rect 1267 1159 1325 1165
rect -1463 1115 -1417 1127
rect -1463 739 -1457 1115
rect -1423 739 -1417 1115
rect -1463 727 -1417 739
rect -1367 1115 -1321 1127
rect -1367 739 -1361 1115
rect -1327 739 -1321 1115
rect -1367 727 -1321 739
rect -1271 1115 -1225 1127
rect -1271 739 -1265 1115
rect -1231 739 -1225 1115
rect -1271 727 -1225 739
rect -1175 1115 -1129 1127
rect -1175 739 -1169 1115
rect -1135 739 -1129 1115
rect -1175 727 -1129 739
rect -1079 1115 -1033 1127
rect -1079 739 -1073 1115
rect -1039 739 -1033 1115
rect -1079 727 -1033 739
rect -983 1115 -937 1127
rect -983 739 -977 1115
rect -943 739 -937 1115
rect -983 727 -937 739
rect -887 1115 -841 1127
rect -887 739 -881 1115
rect -847 739 -841 1115
rect -887 727 -841 739
rect -791 1115 -745 1127
rect -791 739 -785 1115
rect -751 739 -745 1115
rect -791 727 -745 739
rect -695 1115 -649 1127
rect -695 739 -689 1115
rect -655 739 -649 1115
rect -695 727 -649 739
rect -599 1115 -553 1127
rect -599 739 -593 1115
rect -559 739 -553 1115
rect -599 727 -553 739
rect -503 1115 -457 1127
rect -503 739 -497 1115
rect -463 739 -457 1115
rect -503 727 -457 739
rect -407 1115 -361 1127
rect -407 739 -401 1115
rect -367 739 -361 1115
rect -407 727 -361 739
rect -311 1115 -265 1127
rect -311 739 -305 1115
rect -271 739 -265 1115
rect -311 727 -265 739
rect -215 1115 -169 1127
rect -215 739 -209 1115
rect -175 739 -169 1115
rect -215 727 -169 739
rect -119 1115 -73 1127
rect -119 739 -113 1115
rect -79 739 -73 1115
rect -119 727 -73 739
rect -23 1115 23 1127
rect -23 739 -17 1115
rect 17 739 23 1115
rect -23 727 23 739
rect 73 1115 119 1127
rect 73 739 79 1115
rect 113 739 119 1115
rect 73 727 119 739
rect 169 1115 215 1127
rect 169 739 175 1115
rect 209 739 215 1115
rect 169 727 215 739
rect 265 1115 311 1127
rect 265 739 271 1115
rect 305 739 311 1115
rect 265 727 311 739
rect 361 1115 407 1127
rect 361 739 367 1115
rect 401 739 407 1115
rect 361 727 407 739
rect 457 1115 503 1127
rect 457 739 463 1115
rect 497 739 503 1115
rect 457 727 503 739
rect 553 1115 599 1127
rect 553 739 559 1115
rect 593 739 599 1115
rect 553 727 599 739
rect 649 1115 695 1127
rect 649 739 655 1115
rect 689 739 695 1115
rect 649 727 695 739
rect 745 1115 791 1127
rect 745 739 751 1115
rect 785 739 791 1115
rect 745 727 791 739
rect 841 1115 887 1127
rect 841 739 847 1115
rect 881 739 887 1115
rect 841 727 887 739
rect 937 1115 983 1127
rect 937 739 943 1115
rect 977 739 983 1115
rect 937 727 983 739
rect 1033 1115 1079 1127
rect 1033 739 1039 1115
rect 1073 739 1079 1115
rect 1033 727 1079 739
rect 1129 1115 1175 1127
rect 1129 739 1135 1115
rect 1169 739 1175 1115
rect 1129 727 1175 739
rect 1225 1115 1271 1127
rect 1225 739 1231 1115
rect 1265 739 1271 1115
rect 1225 727 1271 739
rect 1321 1115 1367 1127
rect 1321 739 1327 1115
rect 1361 739 1367 1115
rect 1321 727 1367 739
rect 1417 1115 1463 1127
rect 1417 739 1423 1115
rect 1457 739 1463 1115
rect 1417 727 1463 739
rect -1325 689 -1267 695
rect -1325 655 -1313 689
rect -1279 655 -1267 689
rect -1325 649 -1267 655
rect -1133 689 -1075 695
rect -1133 655 -1121 689
rect -1087 655 -1075 689
rect -1133 649 -1075 655
rect -941 689 -883 695
rect -941 655 -929 689
rect -895 655 -883 689
rect -941 649 -883 655
rect -749 689 -691 695
rect -749 655 -737 689
rect -703 655 -691 689
rect -749 649 -691 655
rect -557 689 -499 695
rect -557 655 -545 689
rect -511 655 -499 689
rect -557 649 -499 655
rect -365 689 -307 695
rect -365 655 -353 689
rect -319 655 -307 689
rect -365 649 -307 655
rect -173 689 -115 695
rect -173 655 -161 689
rect -127 655 -115 689
rect -173 649 -115 655
rect 19 689 77 695
rect 19 655 31 689
rect 65 655 77 689
rect 19 649 77 655
rect 211 689 269 695
rect 211 655 223 689
rect 257 655 269 689
rect 211 649 269 655
rect 403 689 461 695
rect 403 655 415 689
rect 449 655 461 689
rect 403 649 461 655
rect 595 689 653 695
rect 595 655 607 689
rect 641 655 653 689
rect 595 649 653 655
rect 787 689 845 695
rect 787 655 799 689
rect 833 655 845 689
rect 787 649 845 655
rect 979 689 1037 695
rect 979 655 991 689
rect 1025 655 1037 689
rect 979 649 1037 655
rect 1171 689 1229 695
rect 1171 655 1183 689
rect 1217 655 1229 689
rect 1171 649 1229 655
rect 1363 689 1421 695
rect 1363 655 1375 689
rect 1409 655 1421 689
rect 1363 649 1421 655
rect -1325 581 -1267 587
rect -1325 547 -1313 581
rect -1279 547 -1267 581
rect -1325 541 -1267 547
rect -1133 581 -1075 587
rect -1133 547 -1121 581
rect -1087 547 -1075 581
rect -1133 541 -1075 547
rect -941 581 -883 587
rect -941 547 -929 581
rect -895 547 -883 581
rect -941 541 -883 547
rect -749 581 -691 587
rect -749 547 -737 581
rect -703 547 -691 581
rect -749 541 -691 547
rect -557 581 -499 587
rect -557 547 -545 581
rect -511 547 -499 581
rect -557 541 -499 547
rect -365 581 -307 587
rect -365 547 -353 581
rect -319 547 -307 581
rect -365 541 -307 547
rect -173 581 -115 587
rect -173 547 -161 581
rect -127 547 -115 581
rect -173 541 -115 547
rect 19 581 77 587
rect 19 547 31 581
rect 65 547 77 581
rect 19 541 77 547
rect 211 581 269 587
rect 211 547 223 581
rect 257 547 269 581
rect 211 541 269 547
rect 403 581 461 587
rect 403 547 415 581
rect 449 547 461 581
rect 403 541 461 547
rect 595 581 653 587
rect 595 547 607 581
rect 641 547 653 581
rect 595 541 653 547
rect 787 581 845 587
rect 787 547 799 581
rect 833 547 845 581
rect 787 541 845 547
rect 979 581 1037 587
rect 979 547 991 581
rect 1025 547 1037 581
rect 979 541 1037 547
rect 1171 581 1229 587
rect 1171 547 1183 581
rect 1217 547 1229 581
rect 1171 541 1229 547
rect 1363 581 1421 587
rect 1363 547 1375 581
rect 1409 547 1421 581
rect 1363 541 1421 547
rect -1463 497 -1417 509
rect -1463 121 -1457 497
rect -1423 121 -1417 497
rect -1463 109 -1417 121
rect -1367 497 -1321 509
rect -1367 121 -1361 497
rect -1327 121 -1321 497
rect -1367 109 -1321 121
rect -1271 497 -1225 509
rect -1271 121 -1265 497
rect -1231 121 -1225 497
rect -1271 109 -1225 121
rect -1175 497 -1129 509
rect -1175 121 -1169 497
rect -1135 121 -1129 497
rect -1175 109 -1129 121
rect -1079 497 -1033 509
rect -1079 121 -1073 497
rect -1039 121 -1033 497
rect -1079 109 -1033 121
rect -983 497 -937 509
rect -983 121 -977 497
rect -943 121 -937 497
rect -983 109 -937 121
rect -887 497 -841 509
rect -887 121 -881 497
rect -847 121 -841 497
rect -887 109 -841 121
rect -791 497 -745 509
rect -791 121 -785 497
rect -751 121 -745 497
rect -791 109 -745 121
rect -695 497 -649 509
rect -695 121 -689 497
rect -655 121 -649 497
rect -695 109 -649 121
rect -599 497 -553 509
rect -599 121 -593 497
rect -559 121 -553 497
rect -599 109 -553 121
rect -503 497 -457 509
rect -503 121 -497 497
rect -463 121 -457 497
rect -503 109 -457 121
rect -407 497 -361 509
rect -407 121 -401 497
rect -367 121 -361 497
rect -407 109 -361 121
rect -311 497 -265 509
rect -311 121 -305 497
rect -271 121 -265 497
rect -311 109 -265 121
rect -215 497 -169 509
rect -215 121 -209 497
rect -175 121 -169 497
rect -215 109 -169 121
rect -119 497 -73 509
rect -119 121 -113 497
rect -79 121 -73 497
rect -119 109 -73 121
rect -23 497 23 509
rect -23 121 -17 497
rect 17 121 23 497
rect -23 109 23 121
rect 73 497 119 509
rect 73 121 79 497
rect 113 121 119 497
rect 73 109 119 121
rect 169 497 215 509
rect 169 121 175 497
rect 209 121 215 497
rect 169 109 215 121
rect 265 497 311 509
rect 265 121 271 497
rect 305 121 311 497
rect 265 109 311 121
rect 361 497 407 509
rect 361 121 367 497
rect 401 121 407 497
rect 361 109 407 121
rect 457 497 503 509
rect 457 121 463 497
rect 497 121 503 497
rect 457 109 503 121
rect 553 497 599 509
rect 553 121 559 497
rect 593 121 599 497
rect 553 109 599 121
rect 649 497 695 509
rect 649 121 655 497
rect 689 121 695 497
rect 649 109 695 121
rect 745 497 791 509
rect 745 121 751 497
rect 785 121 791 497
rect 745 109 791 121
rect 841 497 887 509
rect 841 121 847 497
rect 881 121 887 497
rect 841 109 887 121
rect 937 497 983 509
rect 937 121 943 497
rect 977 121 983 497
rect 937 109 983 121
rect 1033 497 1079 509
rect 1033 121 1039 497
rect 1073 121 1079 497
rect 1033 109 1079 121
rect 1129 497 1175 509
rect 1129 121 1135 497
rect 1169 121 1175 497
rect 1129 109 1175 121
rect 1225 497 1271 509
rect 1225 121 1231 497
rect 1265 121 1271 497
rect 1225 109 1271 121
rect 1321 497 1367 509
rect 1321 121 1327 497
rect 1361 121 1367 497
rect 1321 109 1367 121
rect 1417 497 1463 509
rect 1417 121 1423 497
rect 1457 121 1463 497
rect 1417 109 1463 121
rect -1421 71 -1363 77
rect -1421 37 -1409 71
rect -1375 37 -1363 71
rect -1421 31 -1363 37
rect -1229 71 -1171 77
rect -1229 37 -1217 71
rect -1183 37 -1171 71
rect -1229 31 -1171 37
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect 1267 71 1325 77
rect 1267 37 1279 71
rect 1313 37 1325 71
rect 1267 31 1325 37
rect -1421 -37 -1363 -31
rect -1421 -71 -1409 -37
rect -1375 -71 -1363 -37
rect -1421 -77 -1363 -71
rect -1229 -37 -1171 -31
rect -1229 -71 -1217 -37
rect -1183 -71 -1171 -37
rect -1229 -77 -1171 -71
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect 1267 -37 1325 -31
rect 1267 -71 1279 -37
rect 1313 -71 1325 -37
rect 1267 -77 1325 -71
rect -1463 -121 -1417 -109
rect -1463 -497 -1457 -121
rect -1423 -497 -1417 -121
rect -1463 -509 -1417 -497
rect -1367 -121 -1321 -109
rect -1367 -497 -1361 -121
rect -1327 -497 -1321 -121
rect -1367 -509 -1321 -497
rect -1271 -121 -1225 -109
rect -1271 -497 -1265 -121
rect -1231 -497 -1225 -121
rect -1271 -509 -1225 -497
rect -1175 -121 -1129 -109
rect -1175 -497 -1169 -121
rect -1135 -497 -1129 -121
rect -1175 -509 -1129 -497
rect -1079 -121 -1033 -109
rect -1079 -497 -1073 -121
rect -1039 -497 -1033 -121
rect -1079 -509 -1033 -497
rect -983 -121 -937 -109
rect -983 -497 -977 -121
rect -943 -497 -937 -121
rect -983 -509 -937 -497
rect -887 -121 -841 -109
rect -887 -497 -881 -121
rect -847 -497 -841 -121
rect -887 -509 -841 -497
rect -791 -121 -745 -109
rect -791 -497 -785 -121
rect -751 -497 -745 -121
rect -791 -509 -745 -497
rect -695 -121 -649 -109
rect -695 -497 -689 -121
rect -655 -497 -649 -121
rect -695 -509 -649 -497
rect -599 -121 -553 -109
rect -599 -497 -593 -121
rect -559 -497 -553 -121
rect -599 -509 -553 -497
rect -503 -121 -457 -109
rect -503 -497 -497 -121
rect -463 -497 -457 -121
rect -503 -509 -457 -497
rect -407 -121 -361 -109
rect -407 -497 -401 -121
rect -367 -497 -361 -121
rect -407 -509 -361 -497
rect -311 -121 -265 -109
rect -311 -497 -305 -121
rect -271 -497 -265 -121
rect -311 -509 -265 -497
rect -215 -121 -169 -109
rect -215 -497 -209 -121
rect -175 -497 -169 -121
rect -215 -509 -169 -497
rect -119 -121 -73 -109
rect -119 -497 -113 -121
rect -79 -497 -73 -121
rect -119 -509 -73 -497
rect -23 -121 23 -109
rect -23 -497 -17 -121
rect 17 -497 23 -121
rect -23 -509 23 -497
rect 73 -121 119 -109
rect 73 -497 79 -121
rect 113 -497 119 -121
rect 73 -509 119 -497
rect 169 -121 215 -109
rect 169 -497 175 -121
rect 209 -497 215 -121
rect 169 -509 215 -497
rect 265 -121 311 -109
rect 265 -497 271 -121
rect 305 -497 311 -121
rect 265 -509 311 -497
rect 361 -121 407 -109
rect 361 -497 367 -121
rect 401 -497 407 -121
rect 361 -509 407 -497
rect 457 -121 503 -109
rect 457 -497 463 -121
rect 497 -497 503 -121
rect 457 -509 503 -497
rect 553 -121 599 -109
rect 553 -497 559 -121
rect 593 -497 599 -121
rect 553 -509 599 -497
rect 649 -121 695 -109
rect 649 -497 655 -121
rect 689 -497 695 -121
rect 649 -509 695 -497
rect 745 -121 791 -109
rect 745 -497 751 -121
rect 785 -497 791 -121
rect 745 -509 791 -497
rect 841 -121 887 -109
rect 841 -497 847 -121
rect 881 -497 887 -121
rect 841 -509 887 -497
rect 937 -121 983 -109
rect 937 -497 943 -121
rect 977 -497 983 -121
rect 937 -509 983 -497
rect 1033 -121 1079 -109
rect 1033 -497 1039 -121
rect 1073 -497 1079 -121
rect 1033 -509 1079 -497
rect 1129 -121 1175 -109
rect 1129 -497 1135 -121
rect 1169 -497 1175 -121
rect 1129 -509 1175 -497
rect 1225 -121 1271 -109
rect 1225 -497 1231 -121
rect 1265 -497 1271 -121
rect 1225 -509 1271 -497
rect 1321 -121 1367 -109
rect 1321 -497 1327 -121
rect 1361 -497 1367 -121
rect 1321 -509 1367 -497
rect 1417 -121 1463 -109
rect 1417 -497 1423 -121
rect 1457 -497 1463 -121
rect 1417 -509 1463 -497
rect -1325 -547 -1267 -541
rect -1325 -581 -1313 -547
rect -1279 -581 -1267 -547
rect -1325 -587 -1267 -581
rect -1133 -547 -1075 -541
rect -1133 -581 -1121 -547
rect -1087 -581 -1075 -547
rect -1133 -587 -1075 -581
rect -941 -547 -883 -541
rect -941 -581 -929 -547
rect -895 -581 -883 -547
rect -941 -587 -883 -581
rect -749 -547 -691 -541
rect -749 -581 -737 -547
rect -703 -581 -691 -547
rect -749 -587 -691 -581
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
rect 595 -547 653 -541
rect 595 -581 607 -547
rect 641 -581 653 -547
rect 595 -587 653 -581
rect 787 -547 845 -541
rect 787 -581 799 -547
rect 833 -581 845 -547
rect 787 -587 845 -581
rect 979 -547 1037 -541
rect 979 -581 991 -547
rect 1025 -581 1037 -547
rect 979 -587 1037 -581
rect 1171 -547 1229 -541
rect 1171 -581 1183 -547
rect 1217 -581 1229 -547
rect 1171 -587 1229 -581
rect 1363 -547 1421 -541
rect 1363 -581 1375 -547
rect 1409 -581 1421 -547
rect 1363 -587 1421 -581
rect -1325 -655 -1267 -649
rect -1325 -689 -1313 -655
rect -1279 -689 -1267 -655
rect -1325 -695 -1267 -689
rect -1133 -655 -1075 -649
rect -1133 -689 -1121 -655
rect -1087 -689 -1075 -655
rect -1133 -695 -1075 -689
rect -941 -655 -883 -649
rect -941 -689 -929 -655
rect -895 -689 -883 -655
rect -941 -695 -883 -689
rect -749 -655 -691 -649
rect -749 -689 -737 -655
rect -703 -689 -691 -655
rect -749 -695 -691 -689
rect -557 -655 -499 -649
rect -557 -689 -545 -655
rect -511 -689 -499 -655
rect -557 -695 -499 -689
rect -365 -655 -307 -649
rect -365 -689 -353 -655
rect -319 -689 -307 -655
rect -365 -695 -307 -689
rect -173 -655 -115 -649
rect -173 -689 -161 -655
rect -127 -689 -115 -655
rect -173 -695 -115 -689
rect 19 -655 77 -649
rect 19 -689 31 -655
rect 65 -689 77 -655
rect 19 -695 77 -689
rect 211 -655 269 -649
rect 211 -689 223 -655
rect 257 -689 269 -655
rect 211 -695 269 -689
rect 403 -655 461 -649
rect 403 -689 415 -655
rect 449 -689 461 -655
rect 403 -695 461 -689
rect 595 -655 653 -649
rect 595 -689 607 -655
rect 641 -689 653 -655
rect 595 -695 653 -689
rect 787 -655 845 -649
rect 787 -689 799 -655
rect 833 -689 845 -655
rect 787 -695 845 -689
rect 979 -655 1037 -649
rect 979 -689 991 -655
rect 1025 -689 1037 -655
rect 979 -695 1037 -689
rect 1171 -655 1229 -649
rect 1171 -689 1183 -655
rect 1217 -689 1229 -655
rect 1171 -695 1229 -689
rect 1363 -655 1421 -649
rect 1363 -689 1375 -655
rect 1409 -689 1421 -655
rect 1363 -695 1421 -689
rect -1463 -739 -1417 -727
rect -1463 -1115 -1457 -739
rect -1423 -1115 -1417 -739
rect -1463 -1127 -1417 -1115
rect -1367 -739 -1321 -727
rect -1367 -1115 -1361 -739
rect -1327 -1115 -1321 -739
rect -1367 -1127 -1321 -1115
rect -1271 -739 -1225 -727
rect -1271 -1115 -1265 -739
rect -1231 -1115 -1225 -739
rect -1271 -1127 -1225 -1115
rect -1175 -739 -1129 -727
rect -1175 -1115 -1169 -739
rect -1135 -1115 -1129 -739
rect -1175 -1127 -1129 -1115
rect -1079 -739 -1033 -727
rect -1079 -1115 -1073 -739
rect -1039 -1115 -1033 -739
rect -1079 -1127 -1033 -1115
rect -983 -739 -937 -727
rect -983 -1115 -977 -739
rect -943 -1115 -937 -739
rect -983 -1127 -937 -1115
rect -887 -739 -841 -727
rect -887 -1115 -881 -739
rect -847 -1115 -841 -739
rect -887 -1127 -841 -1115
rect -791 -739 -745 -727
rect -791 -1115 -785 -739
rect -751 -1115 -745 -739
rect -791 -1127 -745 -1115
rect -695 -739 -649 -727
rect -695 -1115 -689 -739
rect -655 -1115 -649 -739
rect -695 -1127 -649 -1115
rect -599 -739 -553 -727
rect -599 -1115 -593 -739
rect -559 -1115 -553 -739
rect -599 -1127 -553 -1115
rect -503 -739 -457 -727
rect -503 -1115 -497 -739
rect -463 -1115 -457 -739
rect -503 -1127 -457 -1115
rect -407 -739 -361 -727
rect -407 -1115 -401 -739
rect -367 -1115 -361 -739
rect -407 -1127 -361 -1115
rect -311 -739 -265 -727
rect -311 -1115 -305 -739
rect -271 -1115 -265 -739
rect -311 -1127 -265 -1115
rect -215 -739 -169 -727
rect -215 -1115 -209 -739
rect -175 -1115 -169 -739
rect -215 -1127 -169 -1115
rect -119 -739 -73 -727
rect -119 -1115 -113 -739
rect -79 -1115 -73 -739
rect -119 -1127 -73 -1115
rect -23 -739 23 -727
rect -23 -1115 -17 -739
rect 17 -1115 23 -739
rect -23 -1127 23 -1115
rect 73 -739 119 -727
rect 73 -1115 79 -739
rect 113 -1115 119 -739
rect 73 -1127 119 -1115
rect 169 -739 215 -727
rect 169 -1115 175 -739
rect 209 -1115 215 -739
rect 169 -1127 215 -1115
rect 265 -739 311 -727
rect 265 -1115 271 -739
rect 305 -1115 311 -739
rect 265 -1127 311 -1115
rect 361 -739 407 -727
rect 361 -1115 367 -739
rect 401 -1115 407 -739
rect 361 -1127 407 -1115
rect 457 -739 503 -727
rect 457 -1115 463 -739
rect 497 -1115 503 -739
rect 457 -1127 503 -1115
rect 553 -739 599 -727
rect 553 -1115 559 -739
rect 593 -1115 599 -739
rect 553 -1127 599 -1115
rect 649 -739 695 -727
rect 649 -1115 655 -739
rect 689 -1115 695 -739
rect 649 -1127 695 -1115
rect 745 -739 791 -727
rect 745 -1115 751 -739
rect 785 -1115 791 -739
rect 745 -1127 791 -1115
rect 841 -739 887 -727
rect 841 -1115 847 -739
rect 881 -1115 887 -739
rect 841 -1127 887 -1115
rect 937 -739 983 -727
rect 937 -1115 943 -739
rect 977 -1115 983 -739
rect 937 -1127 983 -1115
rect 1033 -739 1079 -727
rect 1033 -1115 1039 -739
rect 1073 -1115 1079 -739
rect 1033 -1127 1079 -1115
rect 1129 -739 1175 -727
rect 1129 -1115 1135 -739
rect 1169 -1115 1175 -739
rect 1129 -1127 1175 -1115
rect 1225 -739 1271 -727
rect 1225 -1115 1231 -739
rect 1265 -1115 1271 -739
rect 1225 -1127 1271 -1115
rect 1321 -739 1367 -727
rect 1321 -1115 1327 -739
rect 1361 -1115 1367 -739
rect 1321 -1127 1367 -1115
rect 1417 -739 1463 -727
rect 1417 -1115 1423 -739
rect 1457 -1115 1463 -739
rect 1417 -1127 1463 -1115
rect -1421 -1165 -1363 -1159
rect -1421 -1199 -1409 -1165
rect -1375 -1199 -1363 -1165
rect -1421 -1205 -1363 -1199
rect -1229 -1165 -1171 -1159
rect -1229 -1199 -1217 -1165
rect -1183 -1199 -1171 -1165
rect -1229 -1205 -1171 -1199
rect -1037 -1165 -979 -1159
rect -1037 -1199 -1025 -1165
rect -991 -1199 -979 -1165
rect -1037 -1205 -979 -1199
rect -845 -1165 -787 -1159
rect -845 -1199 -833 -1165
rect -799 -1199 -787 -1165
rect -845 -1205 -787 -1199
rect -653 -1165 -595 -1159
rect -653 -1199 -641 -1165
rect -607 -1199 -595 -1165
rect -653 -1205 -595 -1199
rect -461 -1165 -403 -1159
rect -461 -1199 -449 -1165
rect -415 -1199 -403 -1165
rect -461 -1205 -403 -1199
rect -269 -1165 -211 -1159
rect -269 -1199 -257 -1165
rect -223 -1199 -211 -1165
rect -269 -1205 -211 -1199
rect -77 -1165 -19 -1159
rect -77 -1199 -65 -1165
rect -31 -1199 -19 -1165
rect -77 -1205 -19 -1199
rect 115 -1165 173 -1159
rect 115 -1199 127 -1165
rect 161 -1199 173 -1165
rect 115 -1205 173 -1199
rect 307 -1165 365 -1159
rect 307 -1199 319 -1165
rect 353 -1199 365 -1165
rect 307 -1205 365 -1199
rect 499 -1165 557 -1159
rect 499 -1199 511 -1165
rect 545 -1199 557 -1165
rect 499 -1205 557 -1199
rect 691 -1165 749 -1159
rect 691 -1199 703 -1165
rect 737 -1199 749 -1165
rect 691 -1205 749 -1199
rect 883 -1165 941 -1159
rect 883 -1199 895 -1165
rect 929 -1199 941 -1165
rect 883 -1205 941 -1199
rect 1075 -1165 1133 -1159
rect 1075 -1199 1087 -1165
rect 1121 -1199 1133 -1165
rect 1075 -1205 1133 -1199
rect 1267 -1165 1325 -1159
rect 1267 -1199 1279 -1165
rect 1313 -1199 1325 -1165
rect 1267 -1205 1325 -1199
<< properties >>
string FIXED_BBOX -1554 -1284 1554 1284
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 4 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
