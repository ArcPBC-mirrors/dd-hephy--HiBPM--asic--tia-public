magic
tech sky130A
magscale 1 2
timestamp 1683736741
<< pwell >>
rect -554 -719 554 719
<< nmoslvt >>
rect -358 109 -158 509
rect -100 109 100 509
rect 158 109 358 509
rect -358 -509 -158 -109
rect -100 -509 100 -109
rect 158 -509 358 -109
<< ndiff >>
rect -416 497 -358 509
rect -416 121 -404 497
rect -370 121 -358 497
rect -416 109 -358 121
rect -158 497 -100 509
rect -158 121 -146 497
rect -112 121 -100 497
rect -158 109 -100 121
rect 100 497 158 509
rect 100 121 112 497
rect 146 121 158 497
rect 100 109 158 121
rect 358 497 416 509
rect 358 121 370 497
rect 404 121 416 497
rect 358 109 416 121
rect -416 -121 -358 -109
rect -416 -497 -404 -121
rect -370 -497 -358 -121
rect -416 -509 -358 -497
rect -158 -121 -100 -109
rect -158 -497 -146 -121
rect -112 -497 -100 -121
rect -158 -509 -100 -497
rect 100 -121 158 -109
rect 100 -497 112 -121
rect 146 -497 158 -121
rect 100 -509 158 -497
rect 358 -121 416 -109
rect 358 -497 370 -121
rect 404 -497 416 -121
rect 358 -509 416 -497
<< ndiffc >>
rect -404 121 -370 497
rect -146 121 -112 497
rect 112 121 146 497
rect 370 121 404 497
rect -404 -497 -370 -121
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect 370 -497 404 -121
<< psubdiff >>
rect -518 649 -422 683
rect 422 649 518 683
rect -518 587 -484 649
rect 484 587 518 649
rect -518 -649 -484 -587
rect 484 -649 518 -587
rect -518 -683 -422 -649
rect 422 -683 518 -649
<< psubdiffcont >>
rect -422 649 422 683
rect -518 -587 -484 587
rect 484 -587 518 587
rect -422 -683 422 -649
<< poly >>
rect -358 581 -158 597
rect -358 547 -342 581
rect -174 547 -158 581
rect -358 509 -158 547
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 509 100 547
rect 158 581 358 597
rect 158 547 174 581
rect 342 547 358 581
rect 158 509 358 547
rect -358 71 -158 109
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 109
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -109 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -109 358 -71
rect -358 -547 -158 -509
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -358 -597 -158 -581
rect -100 -547 100 -509
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
rect 158 -547 358 -509
rect 158 -581 174 -547
rect 342 -581 358 -547
rect 158 -597 358 -581
<< polycont >>
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
<< locali >>
rect -518 649 -422 683
rect 422 649 518 683
rect -518 587 -484 649
rect 484 587 518 649
rect -358 547 -342 581
rect -174 547 -158 581
rect -100 547 -84 581
rect 84 547 100 581
rect 158 547 174 581
rect 342 547 358 581
rect -404 497 -370 513
rect -404 105 -370 121
rect -146 497 -112 513
rect -146 105 -112 121
rect 112 497 146 513
rect 112 105 146 121
rect 370 497 404 513
rect 370 105 404 121
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect -404 -121 -370 -105
rect -404 -513 -370 -497
rect -146 -121 -112 -105
rect -146 -513 -112 -497
rect 112 -121 146 -105
rect 112 -513 146 -497
rect 370 -121 404 -105
rect 370 -513 404 -497
rect -358 -581 -342 -547
rect -174 -581 -158 -547
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect 158 -581 174 -547
rect 342 -581 358 -547
rect -518 -649 -484 -587
rect 484 -649 518 -587
rect -518 -683 -422 -649
rect 422 -683 518 -649
<< viali >>
rect -342 547 -174 581
rect -84 547 84 581
rect 174 547 342 581
rect -404 121 -370 497
rect -146 121 -112 497
rect 112 121 146 497
rect 370 121 404 497
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect -404 -497 -370 -121
rect -146 -497 -112 -121
rect 112 -497 146 -121
rect 370 -497 404 -121
rect -342 -581 -174 -547
rect -84 -581 84 -547
rect 174 -581 342 -547
<< metal1 >>
rect -354 581 -162 587
rect -354 547 -342 581
rect -174 547 -162 581
rect -354 541 -162 547
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect 162 581 354 587
rect 162 547 174 581
rect 342 547 354 581
rect 162 541 354 547
rect -410 497 -364 509
rect -410 121 -404 497
rect -370 121 -364 497
rect -410 109 -364 121
rect -152 497 -106 509
rect -152 121 -146 497
rect -112 121 -106 497
rect -152 109 -106 121
rect 106 497 152 509
rect 106 121 112 497
rect 146 121 152 497
rect 106 109 152 121
rect 364 497 410 509
rect 364 121 370 497
rect 404 121 410 497
rect 364 109 410 121
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect -410 -121 -364 -109
rect -410 -497 -404 -121
rect -370 -497 -364 -121
rect -410 -509 -364 -497
rect -152 -121 -106 -109
rect -152 -497 -146 -121
rect -112 -497 -106 -121
rect -152 -509 -106 -497
rect 106 -121 152 -109
rect 106 -497 112 -121
rect 146 -497 152 -121
rect 106 -509 152 -497
rect 364 -121 410 -109
rect 364 -497 370 -121
rect 404 -497 410 -121
rect 364 -509 410 -497
rect -354 -547 -162 -541
rect -354 -581 -342 -547
rect -174 -581 -162 -547
rect -354 -587 -162 -581
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
rect 162 -547 354 -541
rect 162 -581 174 -547
rect 342 -581 354 -547
rect 162 -587 354 -581
<< properties >>
string FIXED_BBOX -501 -666 501 666
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 1 m 2 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
