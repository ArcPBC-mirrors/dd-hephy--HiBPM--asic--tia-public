magic
tech sky130A
magscale 1 2
timestamp 1686510802
<< locali >>
rect 1420 16760 11980 16860
rect 1420 12560 11980 12660
rect 1420 8360 11980 8460
rect 900 4480 1420 4500
rect 900 4260 940 4480
rect 1260 4260 1420 4480
rect 900 4160 11980 4260
rect 1340 1520 1440 4160
rect 60 1420 1480 1520
rect 1420 -40 11980 60
<< viali >>
rect 940 4260 1260 4480
<< metal1 >>
rect 3716 16716 3852 16968
rect 3660 12516 3852 12720
rect 3644 8312 3852 8520
rect 928 4480 1272 4486
rect 928 4260 940 4480
rect 1260 4260 1272 4480
rect 928 4254 1272 4260
rect 2356 4116 2492 4332
rect 11980 1020 12860 1380
rect 1440 800 1708 816
rect 1000 680 1708 800
rect 1440 664 1708 680
rect 152 160 220 392
rect 152 68 332 160
rect 344 140 412 392
rect 536 140 604 392
rect 728 140 796 392
rect 920 140 988 392
rect 2364 -76 2492 132
<< via1 >>
rect 940 4260 1260 4480
<< metal2 >>
rect 1040 17900 1680 18140
rect 1040 14440 1200 17900
rect 1040 14140 1700 14440
rect 1040 9720 1200 14140
rect 1040 9500 1700 9720
rect 1040 7940 1200 9500
rect 1040 7700 1820 7940
rect 940 4480 1260 4490
rect 940 4250 1260 4260
<< via2 >>
rect 940 4260 1260 4480
<< metal3 >>
rect 930 4480 1270 4485
rect 930 4260 940 4480
rect 1260 4260 1270 4480
rect 930 4255 1270 4260
rect 90 3180 100 4100
rect 660 3180 670 4100
rect -160 0 300 400
<< via3 >>
rect 940 4260 1260 4480
rect 100 3180 660 4100
<< metal4 >>
rect 100 19680 11540 20580
rect 100 16380 1280 19680
rect 1420 16800 12860 17800
rect 100 15480 11540 16380
rect 100 12180 1280 15480
rect 12020 13600 12860 16800
rect 1420 12600 12860 13600
rect 100 11280 11540 12180
rect 100 7980 1280 11280
rect 12020 9400 12860 12600
rect 1420 8400 12860 9400
rect 100 7080 11540 7980
rect 100 4480 1280 7080
rect 12020 5200 12860 8400
rect 100 4260 940 4480
rect 1260 4260 1280 4480
rect 100 4101 1280 4260
rect 1420 4200 12860 5200
rect 99 4100 1280 4101
rect 99 3180 100 4100
rect 660 3780 1280 4100
rect 660 3180 11540 3780
rect 99 3179 11540 3180
rect 100 2880 11540 3179
rect 100 -420 1280 2880
rect 11800 0 12860 980
rect 100 -1320 11540 -420
rect 11680 -4200 12860 -3220
use bias2_currm  bias2_currm_0
timestamp 1684167095
transform 1 0 -20 0 1 1620
box 40 -1620 1408 2586
use bias2_currm_x8  bias2_currm_x8_0
timestamp 1684167095
transform 1 0 1380 0 1 -4196
box 0 -4 10888 4206
use bias2_currm_x8  bias2_currm_x8_1
timestamp 1684167095
transform 1 0 1380 0 1 16804
box 0 -4 10888 4206
use bias2_currm_x8  bias2_currm_x8_2
timestamp 1684167095
transform 1 0 1380 0 1 4
box 0 -4 10888 4206
use bias2_currm_x8  bias2_currm_x8_3
timestamp 1684167095
transform 1 0 1380 0 1 4204
box 0 -4 10888 4206
use bias2_currm_x8  bias2_currm_x8_4
timestamp 1684167095
transform 1 0 1380 0 1 8404
box 0 -4 10888 4206
use bias2_currm_x8  bias2_currm_x8_5
timestamp 1684167095
transform 1 0 1380 0 1 12604
box 0 -4 10888 4206
<< labels >>
rlabel metal3 -140 40 40 380 1 I_in
port 1 n
rlabel metal4 200 19160 1180 20480 1 VP
port 2 n
rlabel metal4 12300 4400 12760 5000 1 I_Out_Driver
port 3 n
rlabel metal4 12320 140 12780 740 1 I_Out_TIA
port 4 n
rlabel metal4 12300 -4060 12760 -3460 1 I_Out_ref
port 5 n
rlabel metal2 1300 9520 1400 9700 1 vm1d
<< end >>
